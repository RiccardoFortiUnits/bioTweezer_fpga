`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
btFygjM0KQLlXPreW38zB7garVUJSqLx88XlIZ0WrKfDAx3qfS/vVyrPMkC8bgeP
lsaixKha5nHXZwvt6xcv//th1yw4jzYXf8DDY48LB+an8qkWlcIoxrxe0KGGFnav
ABL8ElD+kg0owSaD6KLYQ6NvL4EWdiXrmDBYAwxYTDM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
Jy2U55MMoHZIKXcFnYe6TLDlIR4mga0bLYNii+4dsZXc1+7Gh13z5VuREyEpfAnD
NODKz6ZnjmNOZ66kS3Es3rgarJ5qyD4s4X9nO0oudZaMI5MOsOSvSQeTl9AFRQ8a
wBXz+ifCinR/3ZgNMdQIzi+JZEw6U2Wbl7rR0PZj0O+PCWNVqe4UNw8OFqyDdwUM
9udRTwzWsrS01C1vKMKcIl1srvAUknICfr27/q+D6HYGu3gR1zjt7RAAO3RT3E/V
iHxxOXwYIPddZmQZ1OpU+K35EYccKmF/QvqIfEaMD+Y9JRDPaMFTdtv+RKDTGebO
SGf2+m4vKq5nvX8PVpx2vrztwU0AiUkYYqsxY6OzSIwkxnlJa7yOx78IbLchhfOo
HxGA+RgHFfxG/Om3gg8MeavdDXave4ZX3IVSvXFcJOv+RiZZ4nDKu/dPXrF0YBp7
7i4TvDgrWLsqpmhNVc6DwnQZ26InImkgCkMMnwFpkUjlJnMoIRP6rKLJ+IFT0eCV
KHr/Ja4z4Lf4kIG2Ysqk9/ji1EN7MDLlPQl/9PM23Irr5MJj4ypsuqmsAsuPYvZi
Se/lYuzTiiRKvhb2+m/gL1fht/p+3JJRLT7EOEsJ2kzCVeqfcDJCCYM2gjpBF2LZ
28PHsMSAys/rcBxbQVmU2/KyGnhgyihdzmJcytEWUebpvxVsGHSF409+vwGkkw5T
lMVmtdJUaf5JVzESGQZMoUqk3bqHLRcQZs3rYqcVZkQzQvYubNgpk/avmeCtWR/2
yqFO+NcYseYNEta6HsDKmof0gkyB31IHGyfHWfGMmPiOopUCTQyJWa4h/Foe0EOi
scqv0KnKjK+Cq5oFnTWjLyAQpw6X1KK9qWeEIGYqAAIqayHHX/pxlVsYCWmEGtro
cASF24QSg89h5+s9Nq+xk8k0Ky2lQW3I67wEotnumXxIXx/qbY9cvsCy0P5/UJg5
uMyKczYOWBcr1lc4YbJjEcM2S9S3KHywwiM/Jj0wY2le4E4lwe5q6HdxHXmRSzhq
BwZr7B429lOiBLIoafWjlUseRjmkTGtuwC+dfvQtQMZJt1T2HM3X+BGcLmSTGsy2
u/fpm3ZC1GRcVExF5MalbdiKajKoRF1+fwEsPQt08b87z8EGjwsriu/lPJYjzcdq
zhh5ALh7RfFCSGcYBdRQy2j25suX8LpHFwKAwfypwQ2aQPL9bT3Gr2Y/KLN2flTB
l3tSY0rkOfeq2qfNnjvMhgPMfFHawEwQ9xNgwKPtm7Zw9rFy/ySRladI8z1VG+6H
fHj+jfq3iWl0XS1n9AL7ZhBw4iFXk2ot5OjxKo73M06uf+OBKJDTwyRbu4UJxA0l
sZhL16zs6ofE7BmjPYr6cpmGfGDH/GNEEiDyIIPc6pWPQEZVqi2hiNKWodyL5zHI
3mmeRw6s6pYXZd1XeAveidGdcSVGGEuxPaNpb73h9iVGWswcl76kcDmUhYt4zLag
COzzj2K+VGmScmUXN/kMxSEvrmrDc3njU8GtN09NKOdVaxWa6ZVC2EZc9GQ5Baa5
gDNzvRZKdWd56RmV7jp5KNjXEkMhTapBQA8WQG2b6qiOfpCDnvqT88bhJDCHTDAz
/CWTxgeXz+m+aq3R88tJQ+TD54qInqWj40WWqp3l8Gl/A0CP+f7tU1MRxk4qa1ed
K0Ij0ElXUE5Bs35JuR20gxnGgMu6HtjMuyKnQH5GzgSLkGGgkNLz4P9OeAgY1Gsy
B5+l1PD9nTg1jWAgITcxmhjmrdQf4Mil5pGPEBcuGMoLmDjG0SGtQHEeWS2qhMG8
AbtjKtcmJ0fJdJgJV8tOuA6CoURUnejxDJpakzmZr9Q13uV2QO13iEYKMsoxCdbF
sEMqzIAockIiZDKkogLP7w0Y8ftvXwELkMuEsGCn/uKTv0e2xOgxA7HgPFd0pZt9
Qjw4jUrgLnA63vN1ZfHUcAMAr8+yoey1jXe9H6fCt5/ANv1Kw8K+mNZmyjQktwoF
fraitEW9cMEu1qMUptY/90tTqWjf1TapkGmZvXTLDIAAPdqxiWSOR6XKW+HkphKb
ofMkyNcOKcePmf2XWc39RScFMIeyelcX0mZ9/NQCIhznj2R/+YNUdBgFjVhWD8uY
Yiafj0r+SZdkNk+yTpnB0B6vPNOByqaba71DozCQCD9im8f3Mx3VFTd29eW0FlEW
M/lTKsPA5YBhpYEfM4TsGDcI2t1qmxLChxEdXe3DFRyNRMFK8fXr3L/EQkfCVwlt
vIkbK0MtFB2xSHYaTu98RrIKyWvUVttSQZG+mHmyIUC9YLJpQv/yMNySneZhRXwk
cPMKdcsRlNnBsd0hLmTma9MdOYlRL3oQ70AItSGerMqZn8nIJRRNzJatwTXc0oa4
jYI+ZlXIHrpC/D3RQiZfyDZIA6OMaGyupqKmzGLMgD20PX4Ia/hZU0FD35AiPMA0
+JLb5EniC0SUcC3mJM9xXPJS947GmJOCs0oH2L+/9BN/f63t7B+R6yMEyITVDuza
NGkIXAAWdVc7s5yfgqAKL6mbldqFPLC+F2V42mIcGiaOMK/kcw5GO95BAshD0cro
yYW2Zs2G0MezNgUEJKMfGWkmeSPwPLpw71t4X1k9B6pVE2gk0Ke9Alhtf1OwklLN
BEXMWcBjz46oL9gAtVj7s2zWiQQb9vgE2sI8gSbmt4b+QHCSuB/VW36OOhNvmbzy
kyN8G+cCg/xl70IAbzfXj3AtBv99vxB0G1FC4LXTJ8dta0qRIWxpbXSzp0BOOdsP
ovw0eXVfRXrAgJLb9HoRHb9tpXsmflnMLaN79JLGbABCbbHKSPDlXttEQXiYcus7
YMZmwoxegV4Xh1TZV81KfjRN0E6ruDIzUrmg4rQ269Vx7+CXBvsV6ZSGZuNSPOaz
4/nAr0o7nwTbZVRGbRhoOUkuXPMpNHXNesN2BES82/+tMgu4nNN3kFQx/omP05P4
0RXgE9a9NWrce0K/vZ95XBBKA7VsFq6dmPCh+dhg2YKvsxSbpt8KOBDblMFXxEvB
NOMk6N4+Gf2T2rlyv9cbOAWSX4Ww/RdWCJDDyJDwxoULU6psTyFT548bsDVHyzAX
gS5sVs66mdy3KkFZi0RUc+94ulAG+mM3ah62/SesQ01qIcs7XOyxcPmAM3C+miEv
lnsm2FhzWNDJ8SU+stHBLP4ta9yhczM9cSSIc6CQt9wJ7eUmV/YBEYZJrdPrwooq
H0IWcbU8QefuZuuWJThZtGAo7gfWKtU6v9ypyYVvPdhI5UgLvTbFGqDK4OUtzXyK
8z5l+8Sw2M4no4BR+nl8kOW4WlABv7CnF6fpa2RnwXOq8cBnIKSGy+/+IvxwnlQ9
v7R/IYAastnnT/F2MUyDahisWm5Dojclu92vRRV28cwj9ntEJzcpxr2h5C9gEUb9
A2jdDJsyPjvcsqwr89x1XsZPHautGlJXLpdeMnEaB0nOs5qyoo7t5Jr++1Dyvq/X
FwNn4jjTso6zcsrdUKPx0AhrOrLsDNT9cbDmF1OrDP6P/QpxdOaDbw1v4TOy8UJ5
nyVmu2AnGZX3GRPBptpBkD2BEbbeicFc6FIl/DxW50VlNPcCJkB02nYo7bVWGobS
+G7NsQ171aoDCHAg4WCj9+xHZkLUzYhzJmZH4/daQdnMXY25suS+miO+UusqNASs
nTbFWSpA3GZAgiRjAH0ZG2S6feywOgEKmhbtaLKmSrLBM7TXCIArpkKMEdM628R+
OMV0MCtrwcfqg3I4sIY/lF02TA1tXiiFD3XP+VpcUraxReNjVryoVeyLWB5Tgo5L
+kfbrzWpYMuCvLlU7/QosssV/fxoJR1X35e6ehv6DoTURgpISjh6xia+ErP9B7wt
oytX2H+gP6xV2LhPefBjyErdt57B+6rFebfTKxZos9pJRo7s2PnhN3BWV98881Hq
OK2s7aF+G5/vdwqYSx6e6Y9D18M5dUHwATdfHtrT0ll6t8SDb1KLBwcICnaK+5+V
E1P8LTyRuDgfDQKnDY5BwfziTSwP1uyN3OF7MGbHjKZGzH/x1OUtRZR5I6P4maW1
KvHHZXRt4xWd2/XjYuKxcA==
`pragma protect end_protected
