`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B67tpRvaO2SvJtp/UKzpFF1Y1F8K+eJYlepAvIt2FoYQY6wplEdhmb8hXKITC/BP
Jp1PpYPtLPOoY1j58EDIsbBqvr5Q14dzgW7pmao54OOo9sSjKws9Xgp14AgmXMi8
Xy0oge7UOtcobNwzGmGqERkhRrRcDCHEmGF2d8m5LaU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6528)
9satM1KelwCdsnYrVi5+TgeNHj4IWGkNTQtwWhg5cPWF4rA6QH+6lBc0W7ZlOf16
gk1d/3nqgOjIJPSvWQC1L87PMZ2VktENlf5lnJT9/kQV6Iiaz/8uHkhLiSv5tHWg
I7IT/rytqe1XJpKb8UVNJ04waskif0o1qpdFnyPKtMwrcBOWLR8jBUqKBplCf1Xt
PAHx3rJuL1zcfoDHdJUqTo3ROihHd0tBx0WWFmteGW0HVsttQ+5sQulmNI3Fwwsl
hRuEbcXfO+cUAvW9RqZEQC7hERfMNtX6YcM4QWZGHrpQJe9Hk23JgQJ0Y1rq89vn
Tkkun/mWflvSkqK5VMRke6k+h6UdkYk4XiabFV9BMHmxB+TUCyJyYDvGbLXBoyuK
Wau/k5pASa3Hu3Uu1YhlP/DxwUzT3RSHYa3CJMftsEkvTV48OYffId/M9n+wIj5j
VrzU0HBjvdJLtcy6LXODkzrXAvmuzciTZK1SV7OrqfIeAEjcUJGOrbG/uK8yVKmx
jiH+rZrz6N0hrAM9Uzzd+Tv1oXHW7oiUpXZNc30o3eyZO0pkuhA0zJAv7L9MT+45
o0uLZctRwQjgTcVF5PygbKaHzfB9ogVUJuuPlHY51zz97WJLm0CU291LaNyW9pmN
X+Q++ZgLSdtjoTqqDfc3lWStHNZ2D5tVIcOlEtxe05hUht9rl1wgolbcIH5EjnEX
8RC2LvGn/TnI/eyHS8CAVWgyl0YweIUXR/Q6W8S14INNM5Wir+gJgSeLl6MzAFen
31GtqEC0sX58IjhmU9+g6Vkxzyskxxs61CpxJfFPs+V+zRL1vrsNiVuA5E4lOhQi
pu/XtWtu4F7yytrbK3ntbqcDHYZGaK4z//2BGMdceUZwq8n9mFbg/iKJUDeoAy0Y
Fc5muwJeeopz8rRpTnLc90jPpbMLSK6Di653mrMuP/SCNfkNEaI1yW4fzM+P/+GB
eJjCcvXAf4RCfwOLEbZFsn0do+KgEFMV1Z12kB7YEusWNotmXhXpJkzg7rHOqwYK
yOjaNtv78FzncEk1wdwOsh7vAtX1wewlJXlOrklZJrBnYesSvOZnN6TDxoRm2k8w
Fnor++PVXvWDc7zf+LCxjrHub1EbvylCUJCCWv4opPnc3+WPliKTMuRnyLmFyfPp
qNQs40eQQMSLbnki/nL91yTCow2cY4fn3eJ7WdJ+8FO/9HVxiqsGptb/V/IWeZv2
OHFX3fFQr3A5M44BX6ffwbb/74DOCEVAJTSOcylsI1AdKjwNu+RMl3EHHLrg8IEh
DrkmbQLhfn1zsHZPT5uxnQw4mk+QywDkZqp3U/hKodUTjFY9dXtCAEywYlghZAji
cREFChJniw+swTVcrlvXFHtmXKCmR1Fbize2X/HTl6HvAe6nPJlE2uSEQ7HVYEza
c+V3OKhXmBe7m8mBzsrF0Qu/5RIQgAhd6d379TfGV8KdluXZgGZz6+mMk1JVZ2DP
EVb9lpACC79poT7he+3Siy3pC/6l0zIzQMOUmHA7sVNTTjYeLgx6b/02JZB4pk5w
ciCeZ3rV4cI5CttiWkqcOxx2+PhtCvDPd07XlpCoX+U5aFkwtUI6ai/2yJJGJteF
HCJWlTDzfZ5iDch7nnAcqNCQrLeOMms1o4+b85B/aIhrD+a6OuS/OCgjLUKFOWLS
/+LmP/CwWUuGwG3TvwG6K90s+5TWPxb0u0zsXH8TyB4q7yHPE4hpUjmIVkzeJUTq
f/txx39/7zPclwERpewqL6dhbYRqV5RIAMda7yaXmvgfDjI8PN6VMYOabDaiy3mO
R3y0vcEL093DRbOaeZrDsU8LQo53I2zTRfE+4LsxGi92VdUJkV6ok1VV4Cw/K/iN
cQ4ezcWDzL57aaKkUvqlg5AAyBcvjQhqx5qINd9TdiK2iKjWIxTz+kzqm7W6rR8G
A8iJn47b03mkDSoVepIKPg40wR69DoierIl/vqCuCAxU7rwI88eUOPAi1oaYWClT
56pCzBwDTknHq9E5PUvvGek3wtrG6RwsNycIiTzutyKwg5ah97QyOKX22lBXYthd
tN3uRFYBi5Wz6wtcUxebRSu1ecs5HNG3r5Huz7LdtiEOfZElYsnIRKLnN3B8UmUr
JfwKJI/IiXTTYbK4XlR7IedIkejXxzbhiBmc2HRezcdAp+v0UjOqGLQJn9Mw2q0A
akak6CvcEFjgez5mBMs6VFRrkspLihnlYjhHG6mYkY59IRvRhhwqIWMOmZmJLhrF
U7TswpS6mcLAwb97Ng3IQrA0shu+3i351qYcH/D2kqvTnj1URBpnNEV3bxhQCJGO
G0VMXwyHvsCDHbxN1upo5GE/RikHxlIUbYG2v+/yHguGRTlKwvDCdJfBwZOpLsaR
NGzdxu3MRb2WoGC7s9LE3nNSrKx30aFcB0znvoTDf/8E56/AUEN4TIgI+l+kTymX
yzchey2/cEd4CxKuw3NWX539jiMI+0OIYtfnDEZzM70JvB2kK3k6wMKPw/E4vCmf
6LFvS9TyF3zvw9usU4PCQgNCKWo9b8Yhlu16OR1fQD8a3oUR90auU+No+t7+EWBF
1fpW66Hp11fvX9ikvYlo9XQRcX0gkT2N5mNK4MbE0BoI8qzEO/lQJRRrWglaS9PO
NEH80wOrQQj6/udqPLrU8FtSV71DGSxV5Djc1vQelUWueiTXUTM1DnJVuN7DNZl2
XwliUcUXwX1xDTW4n/6qoUv5rfF4EXz6NlHG0n/BgGFG6r0t/drPaFL+Bt9q6Wka
98Wq5AomwS0HB5GdWHWPMcuVE4HknwR+lTKERJnJ49z4Viy7lsqFnTM6mnRf448M
rS+4wKX7C7nwXKTjOOdvSv5NJ7mNb5ZoNKgaZA1s7kGnWgDYb/64HwAGSNGaNJvh
zUW7NQSXnwIaTx/4G7tO1gFG3LA5rHfWtv+eCIxknT7wS78KxgGGVgV99ZEKfZsS
zCe0IIFZbpYgFtJIzYLKyfyQA3jmH4Ii2jZfFLTbF9/tOLqoXRuSXyf+544+OXCQ
N/5VTMvY6YP7WQxa5RWEQRHMHYp1P5nl/bkqagZ/QiBCHuWXyfomUHrt5IH2MLXZ
13TmFc6Ir+WQcvp2abG73Cpd3N7QNQXF/JlkF0kQt/fvXqQEUVWLqFYRxvw4xOQW
7UgqdW8Lcj0aiLRTCBbFe00u0DTMqLOKRyBg2l+3Xcbc4BnbX7B0K/xf2Og/hSEd
pWfnogkwWDRl3cbIKo/+kiAjVGbVpAcgz0/q8LyiDz0ZvjOUG+dN4j5PcbAWBCTP
Djy10DI+HN1lYM6mlNAaQO1sG3S4efNAovZ5qTtp+aOzVXvXXO/qoDkdqKHzNQza
dRwPa60v+EACscDSMY9sZ7H+CNgiBHupdnGEX0LnbgkDfVqLN7eUaNMC0cFZ6JF6
oextaHMhG788CCaGglX2H2TQdPi308MEquXjj8WRobwln/VS/lqW+40HRR4+mPWo
hJnS8VZJMaiks0yXJxoJAnjM1QPCYpTVK2B7A58xLoXocX+ccTJCXWxZjlm68vgP
fpcmKLZOnT5oDowFzf5KAqZ/n1RbSd3OKo77P7GX6n8tJbBlprgIZ/XfZlzwk9Th
uwWFCraz1t8hkbJxd5+RZ42GAvm3mvZWb6ruAx4H2DIQVYyxpSaLDj2JnofOQ7Io
BsTHMYfWJumOTj6gZcvkZgoaVnuQZmfJRzljJ/Pk6NIvs5ROovR0mTnSabEUaoWz
ia1pvjU8/UIIj3mv+wuY8zqCYXvGrJ1uYDGgadnCAEQ4Ot3mlixNBHb/4UfpyVRW
8mIph6BGota76v33OSN6N8Fz4YkFRQylGld2gM18fPNW9Swh7JFJxp0p7y/02onM
cBDbNzKDkRiTCQXfoMfStxk087eDRDSyEzGe/G+G9CZUMhD2whsY8650LTK6e2eL
eC8PN5d2fDTHHFvjJzzso6x2apSX48FGKo80GQfkLvy9IaWpZJFUpZU1tmoxmqgU
w65hsrcdLqQ4ihBpCDcOBhAi7ooJZa2A9c0Z5TUtjNX9qX8ibnNCRVJncRbZnA3N
JESLCVUJdb6u+DDx2mxtVhB407zO2JVubIvirb30uaDzozbEJ3/PKqFqlOPOksTm
hsjFo+ePtllO+Aa/fQQsVkDRUc6XBRqfS4gZkwtbd2y079obYqYsVoodahvaZF/q
/8Zb4ddVavpInvdTKVPT4Gh7el36VFIhY6AEJdOY0pGVOfXDr4PQ4hvzQR7d5rUw
mBddcuR/KoNldECnfERjkOo370WxTWBkGnsli2wFiZOi5L1ypjhByQHPO75y/dc3
jxL5fA0Q8K/6z09xeG+6RtQhOimsBbGmD6l+W6gw03E2YonbTiO9QbzLJPwXgfI2
UlJTgxLQrw5GpTg4grD+B1hcrd3ySX+TkD4kkeVlhb1VZ4wG4GydSvmiXWFKAajk
hT7sIXLFEcAS7O53VDUGo7vv0TbNtK0clsarfE3HQznHbojfw0feml1liugynzbF
wItE+gmSkV5QpdQgsLJHwDdBk6yGsRh/Z1URAF81iHo0BlLjHBIl9LuSEGp43kiw
eXjls2vNx07bwQ6Bl4LWeIA2ZZ0bRuRUukJdV3mCANHk+OccuSajrggY9UZhzwhI
79TgnHGXMNgYNhdkzoELpGp98YHVHW0S+XIQJZzLKaI8ou32hwptruunWlnhFY02
nqsN45VhmgfxkykBHHt5VZ+cjOhO30Uhh/PysfvEYQZhBM+XSD1a8q/2ypUWvzVN
8Wf1Nxe16kH12NTsS2m4Gi6nE8o4KX1ppop03pWacOCQZvnqalDpUZMzPRi4lZvg
gdxAkgr3VxroqwxzwLCdiIkN3dxXMGm7F4zh4OZGzlx/nCAL30WFduYsP8JX1yBT
HFebOIKr1KB2Uh7BxpIDNRDxYZXCVFhxvL+44enHFbxtlxfvswK6xm33drSdgpFN
ABb7wklNiAzoRmxca/pNMCaIgk26cps6jmnuARIR8QfMGMVqd3+Wa2j06o+BsjxJ
+CEAXQOYl5VjxJkptTX51TJQJu8Z4abKCTTCik8D9lfVYd3Ej/aNAhx8/yxoHp9S
REtH6WdtjpaZA8dDIOQOfVQBNdWQ3da9lWCFRshrR85TbxG5Xs3krwJ7pHspAYWd
TaiIa6fQtNZasAVogRH4UpOYFKTEw71923Eqg6VpTMfUcGL6eYZe82iSOicl1vyN
R6C9BU0x+AX2Pcn325CugXzLMhLGjp9W/+Sy6im2KS29adL8g25Q04z7ZSSmHycA
KtAoS05hZC/3RQUK77SLaRigesywSTtXnielmQ7uQjHyHPFVBXESFbQVbw6aVPes
Rc1gTJgwyUJNdR59bdPSkoTlYIvYjMryJA5H+YU6LJtH534fa0p7KA0FLMMy3TXQ
qvsOns8vMKpgeQ179x4viI4lUT3h0a8ibPUN1s/Sq9k4K141jqqQvZnAwHMhUvnf
xnetWJcYwAKQbCJhnDWKy9uAmIUThyfrcPrZjbmA5dEx2FR0bgyatdqn+fDPJ/93
GyLIFjIKVgIAFWJMFlbY4ry07BOvJZ3cwBistmtAk0kLz1a4VPe5Bt/lw+EN8iwU
g+t0NKfEQs25N1JcunpxDdAQrRnQRqNhFrP+VYtHddm+yqK3iw1ZVAtKaF8i0aX1
kdF6Gij0pOjQVCJCSawnuSmJ2yvGoqNjpNU+/4bOGLJmgSWZTfBvtU3xGRcriF9m
iqTpa76LtS7dmLdoMa36RTGN1Czyfbo5U8NFRFOKppi+VTCsF7g1HMTFFle0GIL0
RFGGmZkJ8JCT0LHUzcV0MkayhHd66bSyoAsA9ARWfWA9LI7TqDyDfPtKPqLbFMS/
6pdGuAGfrhCDcdpHsz8+qXQi1yZQqEtLHjFDInGnRT5MPjvQ4E2LLq00Z60t6B9D
uNBWACfB0NtKDU9LcIYzCmAXsCpFiXZ5ns/6LV0hTl0XE79AuHzkxB+h+pAvvo7N
sXxO+oJ4lZLlq0CKEHxy4lPcW8sEMlXsnOs+Z87pNJBWA0wu8HKNk5MPx2iBhXBp
TP5+xFW8cvWH5tzmOyfpc+vzQ1v/VtxuihayjS+ALM247n2iPcLB8+ZGyFdOVye3
asugMJlZTn0lUKvnAGX1jEp59W0RMhNX5yUumsz6WMYeRSXg/ztiY5iWbwW6NlG6
NDEX6ElXokSTsIQHbz7f8WOaznpO3T30KHiHFSYpF1WHC6AZhwI2nqCdxP5+HiS2
bkbhij7sth3Z9QvFjVUP9U+ITIadP3CHqG6FyJdOmdfZrHsBlKAS5N1ZSLC9xT+h
+8EUPDPy/rCB7lVdQzKWTvPumtJ7FBiLs8Rq5Sf8zkkXCBe7ykCfS5lOGv8/9g0o
UTKESC9o3/sMWSpMBgyL7pp8ArJIPrPYGg1KdffrtsnfPWPRR/AwgMQ4jeZaFoJG
/h8NUHhIUwbFBVlSdFJyBiTLpysouf4PkTyBU0lq0RcCC2QYBJmKIVbQIAVnrfgs
a/jQoQlF1dYkwa6WaJxP4xWPVb/SvZ6XYlFR/C/TZlZFky4gcpRtjB0EkhMk2d13
wx3EDlrWrKQgKafOHKa6i4/1vsfW8QSvuWkkq1KNvQMJg+8gZ+sXPfp28WNz1ghS
+oEqyig3rJ1RAZge+7Z3Nus0l5HccyftYviGJUqB+uih5NNeD06ghSVWanMF6mGo
/jP8VtRn9W1ucdH50Gf6x4MhKz8EQCc5EXMi+7/MK3oDTspck676xUcfkQV9Rl5h
eFWjsbCq87KnJ7m24JIeBCVCLXa8BiqO2oYdnQxW3YnlERcRL4jfMXHDNdPNI93J
ZNTQvk3UvN32ij2rc72D/qY+tqX1a9gx7QKB3KhhzIKrcb6akkQm9AdcxwQKIcLy
rF3haULooHBDL+M1Z9KOUiCS54a9lPvDrGzduxDAQWhCWY51p24tpGyTNuMtlvHG
kq3D6GZLyiefhYjFTWdLbONhRzbzdgQAxBTvhOI2Z6Cxm8hRZPSxF6fpSiNg+FSx
u6dW5fgjmn8F/+AaxUGc0A1NZ1Q6ve9INf/p6a5Jl7Hrj2GkCCFPfmBwuzRniwzT
IFpgKT4eEwCmm0iY1bs0BQrK+xBoajoCiSgPDE5UL2yLaHlOmwtPfIDuY+BNDMdL
vTf6cEpT/df6tELAbDkGz6sZBc0/b2FKJBpgVS62UMEeyhobC+6jF6prRIHQKrYC
fD/USNWY7R1wmOYkHzRRQnf6NJTdeIH67aVQdgTvefLM9dlhs7KHnqM+aLKfAW5B
QzGPBKT7K6vTQ+vbZnGnYuBRjkNawSJgiam2vh/7mDQEUrXHOnS6TL+K/evZIFI7
/csvZYoQn6CxZWjzc5uTGnLSIr8lBChfe0TwPhqYuMQ3YizWAkiwwpFbmqt0RBLT
7L2rAYHA5hsUlJ5osRCLfrmSLFJxF0eNdlwWgqLIaHp8W9uohvPK2sadxfy37ZZO
gikkIbqT32CuMKrJ8uI/eRAJrZXhPsIR/GPeuZkzFkaBZAAsGoWhgVTg+dExfCuU
QArinCgGNpmHyLvdVHBz06aBzDhjQtoYORbbkeL9gGtC8ZZlUhALarxVvHvk9EcS
drx1vxtgJZTNnEZUbJoaVOrQWkQQjBIqL17kTUbBH/4Ks2KOgRd8UZARG2fUaSyU
7fXWqyOKVR44qCNLZ47Sxg3VnL4LZOkzWf6dcvBnDa3ELFZex44OIdBWC6HooC38
dJ+hS6EOhjwDzuH7leQbxfpyRU1qa6x8zgiWKjtvt+vKxp80IOcuzYO8EIXcuNHI
EfdNKa9qed4kfA7+yVcmF1aKs6xvoPEUst4U0s8XegRvQtHNMTap+WKMLgpAkd3v
Gn/Y34iNe4C8DEHUBlVDZa1AbHJlBKFnDSliZ4G72bU/7E7bEYLZMnFfLtD42SL8
yDe1g3ezpk1EoVuN43ONDeoQtjccij5HpFcMOaIZE/EtSNiowAQPUIWRHponEoot
3UwrcRhbODlG6ypWlU1LDpKqgZsPq0W8TMJuyLncV+7Lv/fuevhNm2NbnVK/9Zln
GVPp17vCr2r+yEHU5H9L9HzH8ln2tnYE9caagZg8yZov5UFqWMm92agZxoU5rzo8
ifBF6J/Ynb6QmZlsRFpqCBIjQrtrHpkLRjdjPIwKMLfieNBtsVnX6Vhf2jDQ9tTk
wP+dLkU1CQ/BYdrD9iCZ+/2Fipu/BAIcyWrl8SJHCfEJOyb8auxQBVskLyir6PHm
56DoZCbDVKCl/67NyBSM98ykkCHCvsDU+3CEgFe2GdGyVs1bhIIGJwdlsMXRKyF5
uwYTNQXmtV+CfqL9PGq3bBZ/iB/rMS94uaqcrTqYLjWDv5YMHeb4u9PIp/C60BUj
8d+giykBVf4ARDXPYaI9muG0VMsC2ZFRievgdiJ5Sq8595PLauS/SVILGnKnG5dy
3h3KmyEwEITs+ODrnrw3RqQAmjjMOPsMO2u/liFntBslanWrFDDxsR9iDhA4Fafo
hO0p02mTmpA11qKPB+BnnmOdqNlWaY8kQduqya5CJq+96C5wN3GFicRyejHbMghJ
goU2Hc0U+G2QGmugVT91Cbz5qhEwHuJBgHIvzUigiIYGuR/L2neqJhqmhOyBZOpa
+Eovs/kiyL+eR5v617HajSVxmMAf5GEhyD0zN2b9aq79hmwS/cRKrk77DcBo13eK
ffD5ljI9FpOF48wHLlnZnnLiBDhQc/afAI7EF9MhVOVa1TaupUyctlv/TyMJLRvR
`pragma protect end_protected
