`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RIPSNwzXPDPxgpCDWevquXPyfUw66W6bl04YNnUw+nGzikx83JLdfoioWlrtjt3b
sm6/2nPbZnrp8baHeQczxqdcz9Tv3jhQBdIIwb3B556jSXba0MmpwJv9opaLMOnI
5Q4nEHwawbL1UBLFllKgRwbTwscuRhuyBF1NBtLAUfw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22448)
a0qrrLcNfJpGYFkzwhVXDpyA5MmWVIx9l23Cc5nYfiyWVyWw9XMQlB3j6H/XeiO9
hDDsS4LNCZJNu+YAyQSLdxfuJaWcfIr8pdWiAr54iXKaA8JDbztH3JM236QX8bbg
P8X2QsmrpWmSUuYTMGLr2mNJoTOmYLBI7x28nkTHC7KGEeyvTMZmpjXbwgYGvI67
t1Lh221bqdtBZTB/JG3ECfJUVH6UnYoLM9OfnzofT1GE1SiRIqSN7sHR9BWxDLPA
z4N59ZlvWAzBwWXh1sExXT4fLrS/6ovDkDWCkHJQh2L3H23HToO77Q5KActB/pjZ
QNXTlF83hCo0h9C6/hi3xL4rwzi14b9BeZgJG+dQbHzzRpd+8z6TArxLUOCfTwLV
6EBl28F+LSeSMAbNsQsacWAxXRq135VdcFELKLwsAak/1MP0urP/r8I1NUo3LGfv
98MUUHRkgVzBG0aPj04pm0wGitmkF2BGHeLUTvu+zYDQaDJ3iK+k5Kg7ascminrL
ye2OXW8rr2n1cvxjb0kvxNzsEk08Q99oyxOjS+sEkl3fBmAhXw2RJ4kYxG1rafTp
FbT4ZHB73UvFj7YLc7807XDGXN/VOtc1ucGzwAide/iBHROAJEwD5lWe4bhxnpDG
pilz4wBZDSQVKyqk/nHblV/B8SS5EKuArGUX0p7ZdddEouWgwitfnqWEFxjIFNnl
0qkTA0v3Pp7Zi9kDkPMfvkx+GX54NwANybhAJTSGFeHf02RMrez7imDsdlSJNF97
UxKZHJmC4r3U1sgGMsNlxB0CgWx6qwDmnH2KgbZ2G4JdWsOfwTlXy9x2nvWWE9ln
R4He48CtlAyfZMJh9Sw3X3LVvk39RTfm91u5nbLnI3PSsI3BBVmvkcemHQ7SFb0r
abK4ef49utobaCvIAFBIxW/UY0eOjZligHud0NA4Qp4FYnQHcM5scShYTTUlGfsd
ciOldVx35SwTyRvFxId6zgYAQbjImTc2LPEOSPHjrEqPmRCFDmHPi2BDhgiuZObw
qEvkLFq6/KIN4qDWZNzowUpOTYTqK3tow6Bwh2PQO/jk662/qU8o9DYH3auvfR+s
fdvRjMEIBR/tQnP8NMkN6rOQaIvUw4dAA2NHmSSwmuvgapuWQFgukV6yCNnKJBB7
XNp2fUXs+vrYsMyT1oFp0F5zaTkAjCNblmc4dGZiDdNLoXztP4kNE7Kji61BeKDe
+meGYtSUmDjU12uEi/nMUk3dVyMCS0XR3RXws8dKYYU76PXmo3y9TDiDzej+ELTd
7K60pmjrpryCAaL9Fcx2ljytLQne0v8z5BI917NY3nNh/hMlQpzt7OKd3FT1OhW9
Iu63ezlc0LcwXNhrgH0pv78c8ADy7Dq5AaaeiOfR/jvHkgWPjP+NbtSN+nkqL7AH
MrLj1zVOW5DOILsrD74vmJPJsXfe8Dm/0YcvQ3iOzw/doJlc2ididvR1mGI/ltgW
IvmiVtnQV5v7d5vKo4LnPfAOtRPJ8r1oxXZwxYayxSYMcUvMfGF9qHrNsV0Ol9Az
IqQnDaaIjwmvaM1CLgLwjXu3lEmhEOPJ+x61Zw2GOfFC728uwABxSO03XmbMfGdm
l4T8RBeY6TAgFKPr+KkU8UmbZls4OYJb6IXCMnHAprSiNawvUe1bwtqfYgGUj7GK
aCOhKIeQklEm3vIgmw7lzCGivABdDXGDMTtEeBrbmj9ZcHNjkvIpGWQh7jrOtlmt
D075LxWIBQj5C6Nz9CHGkcTx3IK2ytLIk810QOUUrJorcKnWVhSasw4BP5kbUp7l
f03aGC0fUM/LgS5zgSf+Ydf3Mt6Zbl/Z8pKnRSZv9BlvLGpYn6Pzj0URFwraxtt9
w2ibSiFL7tD2kl2p7N0mpgQcZ4X3L7QmhcxISh6NgLSYy9Ppi2/yYdknrV5iwBqq
kImBgukS1pvJZeP6VHL2C546IFZ7T4/A37kf/NC6zA4EMp+Xv7s+dSsk57IKb/VN
5CKtzlwY3FGyMBY7qbw0gi60ccxRjR+WpOBEE9+KgfVniJQg3GisZBHYuaHEpTlt
gIzXelvvgGhoDXQbj8xs0SvqHLRuKybZawpBZXRtT8n9g4V0Q74KocTu2YmicS3b
/5/ZrIzmXpRsNahFiHHG23XhenkMiCxlZcbhERhaBBeV/qx3P0GA5zSkOdPa2Kny
FShoieBHQcfp76puwlkNwuV8Qp7LqJ/HtpE1ndOM3aKUAYSTfSG6baYbKytR+Av6
vNLWhj8iYlZh3g8NF76iCd0zlMjpJsqbzp2vHGKZPSJbNlS0Vc4IzdwmtmwSmSaL
0qlskv/Wzg9Z4p5OjV27yJp1Gx2z09WFCQRN2/YPk78LnqSKN2k/9b6J9LyWbkZT
VYiIGI4dVXvhcJ9R9TvBBrS6s7vnEijgvzzgtKsxCukVRcm61WpfTUJHlgZe2iwe
dCUvVq7vQOL0t5BqyHWFO0sgR2gOTzuHCqdA2oMka88TGcPP3a0boj6sMYT8ACAz
7s7C6h/GuFg9ogbmPYmAU56BAUMxSBjrrRynnSW4jV8vdMjpZpzV3kbBgvC8OtSp
t3lTa8s+NxHJL9tXprTKQL8kzgpi/F2FYVm+FRIf7MM1lRhypfkKwFLedoDB8XzU
sxKMXW3WOzpRetTMo4WEnYEOeLrk+EB2JOqACTlAe/hKnaKvLu+OSrdPxF51/eW8
4ELvHJQJVREIdsFYObWA3O1Y8UNYiBVyjG49mit43KPy/Fecs/rNK4Pa8DmuL13i
Xg1DEGAjIfVxSFkcOSH2CWdjfEYznAJhW12EU3/47no6vbASSNmaFffw/3gA1KIj
/xbkSK/FPzNewIoekTRFWFL8qDRVu1KihYJHMWAlrAtA7fr977996SYNWliGnpWf
48SpI8lzIKh9LhS67T88rH0l46llYgxioTSDKDSWWqHLpQR9xcmNUR+GO6wSax+M
nzVy/QuHa8+GNlaN6kwIK4rHsIL6wUXPfMDLy190aD5JZSGmYi9vaM0NpNUG0ofH
7upgzxfShgwIML67rPTJ3oPmhi3KV2OLJQEzq2dO+XdVeQExHmXh5M4x8m6JcM1x
snkqfq5mOrmc5QuRXxJs64Jh6QTjMILfY7TOF84LlPDaKmUU3dWS9PbxLOl8knJx
asz1UJXUkaDXSjzq1vJ+xT8VrtSbCGc7TXHIy7gwlCBptLXGPyvjVuaeS5AS5C6n
gYDKDZscgZ/8wx0nQ5AwqFrT6JYMB2NBgz4CMFKVB53a6/w8Hx9NaXfL1ZAwINuJ
ZTwN4B8B0wb8m2XVJAZZ1SueLN2s5ImueatDFmh86eCoyy7s8z0FJLO29f649CR6
tcpQACVYAIWqqvWC0T0SGFVw7xsvYk5jjogWYelVPweZ9EFmFoPFD11AE/rh+3N2
8f4K5PO1Feur9R+jk/Hpg/eUtBD006fM+uOg7uIAHFtUInwawPDT3V5MevklkxjV
99wuYRHPiDJL4TYDUGiHYyGwjGaTWygXq7C0UQz/IcMfxFaf85gRVV9n/YeHvJX7
4wI6suc6MU9r5xnmsCE84jl228ftdxISlqLdbD6ts6d2AWNeNotcPoGuUv5BtnYu
PSHzeG6ZnvQvSF7tery+4syM+X+fEarZWe8HeZ2R6VYXwn26umqF2aO90lSCZn79
Y/Q/NHP3DrArrLM7UKuX9E77iTFxQ5+HzrLjvjc5b5lIvCTPoLIGKu2989MK+fiQ
B+Dvu0FMyu38mWAtem6R21GUdMcaLpi1XZVqBeEIFrvd8kK8zQCoEhzUFEmCLAG5
mlZZU5E3CoDBLuMEtG1UpmBNyjoGD1t/3Zr1GsjHIrnHBl6Kp4WTulLnQygpGFhA
FJdY6mxHFybseNi88wxLQrc8CFb1PxLY8NSDqWDcVVTBNHYWWE2cw1Am969BGIwW
Dw+Sb6F7jvYA2lKYjXjdmM67mD/4jRBv2QvmjOcGBJ+YLn6dR3d1bTl7ShXI4vrp
fLaAKXNjStmXbTblcy7hY1EEE1rKkpF+uw4w26wXSrLdrq5dsVo5cjFOoDpcLWEk
q/tNrN4dNY4ylH74Gr/O4HaMOgGjvMEvrb6T1xaCt6Ud0qG9GQkUk3YWfaKI1Eh5
PQsj9KfpA7ApDqSJMBjisy3g/XJmC/nz1/5C/TkaXGGkOzXTaS7+At/9IPQZvHI0
mT6Iq52r2uD1MSD9eBjRdzuotTpOiDVYxk63AAf1gAUUYSA8S+eARKlAQHoHDH2P
/FbXv+LOlIucrhYR4vfeVOBtvuGtRrhzdqWpg2WfdLLCo3OiTANgU1TCxWffxseB
HnLCTGnLM04geVPQN7yhkPee35sunvV2qbVm215on2pXQvPW1UVXbgg53aaj+iVU
+Yf+Rrlciqy+KS9eUUCvtdWpUELGOAl9OOa3YUI3zm3rKoTzmkYWV/fCgBNcET20
DhCRndipvJxA8KFHRgGX0C+JcLFySJxKwLz7723pb6QBv1zPOWoJdv3aJFH4TGIX
oX1ea1vHriYzgTn1vokv3mNxtqf035C2583MoRMnD+F20HSB98A0EFlNJHpiLtzk
40ER0eiQ7QYL88uOBY1BXEn2TavK3pyVnmVZXzNjg0bdSbATsXnM52MYRtUeIuWr
WjPVH9MOx/MoGcE830Hy2L/L1YrCeXAuknWGaczlKs6Cskv1Cdg3ESxhLZnT4X9H
Y0AhGWRimwicjCp94UFb6/sUdAvrMlX30hzYqKq97K/fQwItqwFRCG5gdWmElIlh
VURydrDoHf6ra8VoATtpPLikxEIU0o7/XX9ZEad40gY0CCWMAG36TqMXmIHjTRr0
RxJJrgLb4dNH/bqEx/qnpV+Hql1lwWCTlqxnuuori/7VVhEHtZwB7jUkrflg8bOo
1Bv4QcT7HKdz5Dps+UOp60vIifdh2hyarCxO+Aazwii5ovciaWZCjROjprB0qSI5
VnQNgkGxpnFEU5GH9dZxdKX4zAjcGFuNJq+dqgK6vKm7rCHI3ViphH6lpt3f/nMM
fxq0oYAw14BGMeJMQHu8b8TZltnLB1Gq++TyEKpVY8ah22mmTyBbKgciz+p58Pag
ODJP7J76WHyX/dkBWr1XsXPwSVmiR5zUjwWr+0sUgYNfZCuHezhcwtOQXqVihHiR
MQlfhgg3g7YFEaZ2ropEXceFKoyr48umVC1Y06TUAEh6FTcGaV75OK5V+NBGHY6m
Pqc8jbWYjlwz599U7Mbb+P0+I25YU5bCWDnqs6H/QHX9qQXPxrWpjYHgfTEco97Y
NeBPxz4GV8eyAe1PbOFezYAmxU2ACQTZKpwkdN58d+ZHvljepSjJLfwADNCluj2J
8oB2yViaBFIZI0PY0RPuNiCUAXzN/S1omQ4dP5wNwWWH/tpXGlDOKNGx81iXVp+h
c+2s22myo8VIm2ly9YPYlQXff8ymX0ELFaLImoc+BejbSc29P8YvdbhywVlvUeiN
WYx421PH95B/iNe0XJLQsJ5TUUjRQE5DgVQZZQLSsYbDR/0U6Utm0L6MQ7iX6lod
aLm6kZfDoXcBqf4akA5WNLpWBuuB3NYdwWRJ5k/fZ44A4hdspgjOK8MdUpvjqU4+
NCq607L3EtnopJPRLbT+6moDodyXzNlySmfQOrL0PQs0bOpfQKiHiQG3U8jiZFEc
PYLs2DBBin09+9IONl2ncOALugjAwSzb1J/4ET4lTALJPlbiCOGwXCby4B/Nuq+V
ghcnLiozGk3FQGVeINwVXXTk8SzXQ/Y29I7iWuEG740yWJ9pIy+0c6ihcQKtWnwF
+0zSlxYJ8MFBXyVdhYri49c7ueK/ubk2oeK14rhTh5nxB1gQRTYWUezimH8Dvk9H
swFyJvB+LTNZEptvshgO6Hq3hIXz+OfiUyXXDSGSxcyZx927/0br+LzCJZSEI8ga
ug1b3EkKfHINUc2zCQm+ThREgbc0pAi48ArP+QWQbJWVoO7YMhqqtWvIWiCbqnUM
89Wgl8G253aMNE46RmS2spmE7cDa4ov0on7X2ji6hIHlbQwTwcaxUPDbN3tGm8bU
7KxFNyjgfdAhCdhBx5NCZhxr8UUH2zj3ebl5ZT2WG24kake7Vnz8sfKdc0bJ/JX5
cuARA8nd3Gi9tmHRn8iskS4iwKun+SiGKr8tur3MfmDsW8Vvf9sCLDzhbW+6Lpbh
Sx8oxYZkmeHNwLkcyB5Egds6qdO0PzbSspLh6FEaEy36qTpzSPFLyKhl3K2DO67l
UNbTLuHlHSWSD3MajnglUN3h+Y5+hZmLFe7D+qPCeXzYNVzoW886/hwtUBN4t0+B
WeduK8CWYCMiLHBAcGs4jzdz+0khlp3GliTQ/+Xqu5nDDISaaiCfsXN9v38z4XPd
XchIi8eVBOFeQKjgZWLgJckLqew1RLYtXSvLNePBYUkQ3LnZ5nI1fAy4DlmY7DTU
xdRuoVev3XE/GWrz1VMS1+BDpsrRNR59IR3We8oHQLcHNVMrPDbg6G84skYVjzr6
jVL//Zl+HLBEh9Gh+wp0P1O5xmYs4bDJz14tLycdN2wwrY/7wcIDYNpNzq7g7P56
Z9nNZwsc3tVQJxppzmfuajVKxkK3xA2CLs5zfIoDC3aDVW5YNQQAiqC4pa6tzJOc
PP3vqaEHZLizTIN1M2Idm0ObzE39l+OOt51CcpOZPFK1qvT85t+kZAMLixQ4UPVd
xrDayut5fqia0ahdeCK4WZcNnx9S1YFFWEB1xzPnSgLz1ol52N8S9sVt/3IE9MSf
YMXehJDardznI7qQAIeLnt+i8v6GD/nEgXReQMB6+CGyp3pPzTNd/NXB7wIIPfu4
MgkRMPxNNNZEw+vYu0i5yILE+bqeczgp95Xt6ZXGFf0L9ust3hJsJvWcRXmkYzAs
LyU8R3yhAzvyoluT+4Pm5NctDuHxg+JHVqniM85nRtCajWeGczZdbVnx6rrbFIU9
bDMkvzuY/VyF1pK/ANrcEQuYB1ys1bbd2XJmD1RTis9fNqrDgqIg4QOt6up0YodK
z1Cv6ZqpcQXLH2RULIRiS4dpvBbD0jEtJ2tGZUNHfCefwWSesrTNwOdIRBHyN2RR
sYq0JLEoG1CyKtc0PXZMvYoy0EvGz1W5unzJdCblS8DZ7lOElGUFk4T/Ck8+/0jt
cecsq4rKtuPp05bbDBBEzxLbUE5oG7gVN1MFhtjFbOWT/S2cOExnzHzdeAdqBhgr
c3YxUBAcWvEeKWAEw2HLJ7dTMS0zxX2VaiZNMxZ03EF7acoWt2HkqsK41J+Emlql
bTj1+YlUvj9Hr1VP+npaz8aFJGnA48aHTEtMPA4R3v0MJWNpaCKjvxqMQ2SP47nD
j8qMTVVPW/twFmiz4dXDMgC2ojJdPuyszZQ0xz3UuEhZP0YclziPneMlu9vaOtwD
SltQKoWj9LRMIYHuNpch1NgtoUWK0P1rvD4OUPbu9y1UekIueu3FbduXjxraV/4A
fI6kcDxkl7fI8yauLht0EAEMwKUOg+CVaX1plGsAusSxK5ZkmzuQ90z49l5rb4Y5
+4DfoWbaIp26HjWQEnVC2irfcC1Kx4fAhit92KYK0E6bBgkz5HO4rmXCqw/9Sjei
iULiv7lG7W/I+yO6NGD/Q4+TeJzjaZkJnWm8ufRd+ifEppCBf2/XI80Nwm6DeJ0Y
ULmeIwQKBb5rEoYxy/kRZM9J6fx8sTFygHpSsxNkbK7Nr2wUtfKmC6ds9/pVlQ8n
3pui+qPLdI+i1m79SQS6gfGO6L9v1SHy7Jpce+VhiB7j9NKmIJIplEqkZZWc4DK5
vaAv/9dktFQT5zDE8Te5wH3FksFuPOwIUqjl/LPoXI03Uj8e7n2BOV0gLJwn9s7U
yf0m9/0gGZW6zcoNKFTrwPeWyh6RZougoDoVIk83UDV6MEwlsMPUFd6F2jx1hOEL
AU3vLhvQc9n0tFh9e63tofS7+uQ+4LxGPf2CTljwsjtSCuffr4HduRjBvEeZGpBN
pzzN0uxL9FVSvJyix4hbfO8G5iYjBnJcmy/16jHk2x3aZ6apbcmKCqIH1Mp/RD8c
4SKT56t5pDEiFwdX7Wlz2rjW3jna88m6761N9H7anIvSaFztugqWa9lQntWGRA79
XxSh4IYkCJ4wn5drotqHFOYMCVoYh4dWwC6sRxVWLOjvNIcmQEN2jpuR2e0dSJp2
Ua5WS221aUZjWQiPDoqaYoISoAiK+gKZbVY2P/Gfw53VX1woff9Wc3LD3fpCoZ3Z
X2Q4KZ6vOmCIZHcHVXd9CA6GdMrzrtYw0l/8BldAw4OUtirEDKO8r3ACrVe6QUQV
MC5htTQ60zutPUBDj2SJ3wu0TjLXvxV7kngrY5o+oZPcuR1TUtW2Exv9QyiiFaMN
aIb6cUOTB5WgK4tgSX81XtIgYoaIyCnZKI1X3KUn7WHTFOPq3Mx+txj1af0QR+3Q
E2U+5Y3Ax1xXzpY43zqQ361mVZJ61TcECOL5mBOQ67K2qW7z1zpBdc2Q8ulWPMNz
eU/tc+K4xvPWvCs60R/GjJ+WqBJS46Z/Dx13gQ5arF/omc54vE7GKlJ8XuUQJwIO
8UCrm2nRu1brvsX14YRTmhlBayND/IFQhD+W7IKC7GLT1fRjNo7MJ1WmebG4d2y0
INf200he9r+Z/U3oAcg/Or6egAbOQc2qfKr676TjW7Wh/Q38Pl8E0QjkjsDFdFCC
+RIKH0pjki0b57KoA7W/+GiEngNJMPHPkKXmHSM1ynuc8AX49MfIvGDhxmCjqP40
jTfzpl5IZrZe/FWXBXiIWZB9efaaNrzgUBgS/sH/2562hFb+93kmhDkgNlODBNJm
rn3BdBy9tji8pi4TykCOwc3ebz4OOaiLXTmHcmJgCqJ5VI+oYKshQ9fumpKqndgT
tTofIh0uS8C1xKcsIRuDqjw1qwWlB454UWoxlWXFZe2AOw719raVsUSIGHpvBQBf
XD3OvyguopFEuyig32RZzeFb4lkJbrtZaL5/Msa/TwI1h9wAQRDJvlD5TsM8fwp4
f8jxL8hCzQV/zRLQQ8y4E34n9lCJ0mSqL1eOp2N/mw3h+nVO92IMy7MwmeGhC5m/
D4NnOx9ZlP/+1XEcbCzud6kD1O8VvnZhDvbbWQepvcLaROY/MRkQfwsmDloBVRUe
Tzr6JzThsrpDXrNgVL5pIlMcaIwrZVNCm9OV/J+l9Dbgssnx9aOCrvPjfiEiaRZt
e7yL7R+180X/VpgjvhL91D+gVPDVKj8mU0IrHnKcAf9JY2eLjmWeImPzyOFiB/tZ
eqC0EyCKnW55ghwwfJBCys4GExRsmp7LBYSLwsjK8bAfv0LrQ8oib4nUMv7oYVV9
MOWo7ye8rPlTHEQBeRBhbO1OXR5zDSECizipjhFrUYK5BDYISySkR9X4Pdmq2xjR
gElfw/NfsWKfMBgoccoyxnGZJZCnVlaEH/Mzus5aIwI9n5g2huB0Pc8Jq2f8QEzt
qYx4+nAPU0cra3Nw7Sm1JDXNYk+byY3en21xaa+pHQUYX4hDJre6eMgd5Tn1rKhv
E0evSuJTop1vPhVvbbwH5uyocSEOynMlQr97dNh/Nsafv0ErA8i5uZqz7gKGTUqF
wDLb05CEoqbtlYUOb5IZTTckzVem4k/nsfrP4Mov26kM3FZ6Y4QRZYUK53BAS9+/
phpRuzJUeE6WwO4JSOsOlYVbun6nErddpq1qU/O1jdeFaTqIp86CvPNZgmQBagKW
yvHpbmEhjyxo4+gyYyes/BMVqh8FUk9/zVIzG0zogGNvGoSASgfNe5JRcHRaBSws
uTOrSA3qJAfm/yd6DeQ3alETLMeSzs+H/0skG6cmvOmf7QrFIfZ2tsXU99YMsfcZ
4ahhkUFzkF70BG32S2YA5jPQVtDABLbVgpwU4PnCRZ/q5Dfey8lVugAQQPbKWYfG
3COr5ftOGFSySB/MQaqf0AIJQAteXV3HDZBsJPDDYqXZl051tmmXBcNBURYLOuWE
ISzAdW8hMjVlNS+3EDa4TdvdH6HWEPmpzVKMlNrSc2x/GyLBclXRoMGWjy+XAJ80
EonpdIcYY8ZVL9MltjNj9xlldpd6nq9MVQMHbh4QVYCSuk3ryrvl/nVYiU5Lilul
PIzWKAMiQMWx2HjWGOJ1qvAHdTEeqHvCIPrlJqS3Npg+uo1nG5QDCB9fuAj9P6ji
qjU4vAGBb/oa73wq5N4IlChacuf/yHX3t36niN4siXhKzWBSqoKVl4R0nUG/6Cyu
Iz8aAClshbg3qRwRKsSdhUiIW7L9q4VJGC/B8QD/Kwl5MwEXvdY14S9sX5pP1ZPR
cb+os8x8HXgU4GS2Y7jKd67qyUTZoksfUyM3sXsnf2PnNFON2SxAf4rk8QoKz/jn
WnuD6xiRglolQIdZAZhmgx5tNkbDG7SQ2c1asSIXQAVQtjbzQ8w7nfHtFhwoj3Od
F8oOI/6uQRHsSRRjefTDnnoaJYsf7FmPbYC6+IFBbPf9awm5OHFYi13leIEucAPm
gYB5pKseQgzQtyWqHP3NAD2dSwa5BOvvZ9E737lWCuIOGpA2ecdg+jU3N1FcULXg
zUGkLmN0oesuHZIp+0/yvqJDy4+fvmpfTD2VJXYlUmm9I+PnES8SmuvsacjuETTT
DJQAMr2kUaNFEjZF9qgAGwiVfQaK6Me9ZoEE+XQdWNCeYApxD0An7MQwipiiM6lb
re/US3OK5HrshOhQyLt1UjBkaFuxK4K7zh2EtJyHZDNn2WIgA/9eTPQ19cNkyNsR
oL51U9GNcuNWUfy2kp2IR4/q8Ez7xWwLWeXPEMK3JB4HXagevTMP2nBXszzdEzHy
df5eX/f/y1cLTKcnXnSNiF7vGCHy8cU8DodbeCZpL/uHrCoMwlH8lcLZrq7Vm+qo
60bLo7JwTrh501+v5yGZwCbBE5YQRZ/7LB680+iWcG/2lkF8JdDW7McFbX5BBGa9
mzvfRGh5YvCpEf34g+rUrPQtiE1Yf0uTkJ9r/HakNYhU2pCVUOZUPNJhA1t1zZ7k
mmBgK61WGxar/ZfEB/uZggmC6IQYNQh7SpaipwLZLSpPs88QNZjbJf6fLybr0cYF
Y1uMFAM3lopy68ERmqfEwJWQaiksyAQkCECK2tcgNt3lkP7J7ufbMcZAodERw6oS
YDRIBox8VqqmKB8msBEOJO6S2VS5TI2b4+mMh15wFlLzfb0hHoJ+5zPmJIFT0TTs
P457ze7IJos4x2t4uhobX+gYtQz1MikVz0Ha+YCESjAGxYzvMwX764iSvyNvFP8J
Pc3qKY4UkeHb8nwTMm2JG7GCI42SLn3JTcIuVw+mwCw5djOQb/FjgGG7U9BAIXzh
w7HN950VEm6wnRM+dX58huUWZocgziLQqiJ75HCEJJwLEXU4KLwp5BIxLuMLeWxe
cYuiY8koz4Kma9M/ejd2Jo85/7L3bUaCkBRFMsWfG4M/PD/Ja/qxYxh4WPPX72/9
7iif/fhU3nZRdddXjjEepGUcK/mvvbUUq3MO2tb9CHf0zCa5M1+PT1dlK59iLjXT
roKkPm5zYTMNbWU5c/F87qEVq7hKstFZQhak4fNXEfkUaebqWxrsvleuri/H3pna
xY5Ds/jMQJ7Th0gy4/3srge5pMyu2QlIiDzwRpYzdNYIa+xUP+b5TJmxx9ld635Y
OOxszw5Yx5+nsTwbrnPgfuNMndZgBH0qfXb/N2WvazEdy3AH+hb1YPKMo6oBvd2Q
aVScaUhCCawV+KP0K7avtJoDjoxI7RAao82xH6LUmcldm1ioxhIErAjSFvZDehYV
85OceFv+9Mct0UtDGqM8iP3xAR/gbN3JGRYXkNDHOewa7SazmBX17sFzNW4SCm43
ea2ycq4OqsDJutOqu5d5ZuI9AfiEXwtMF2dvC00g/7mM4U4IP68VFWPSbmDxqvMy
xF+vTb8bfsHnVJC41R2ZZ/FZFecdnfrB7X8pCMDWKKJtIi8d60JyQHPAoBIyIa5a
l3uSAJ53vvsvkwOC9DRpkj1qkG+41rug2Hv5tUCg9sG/tvC6SWfk20hvEZYRySN6
kWhd7Up493GNxEJaT5w+ZNw1RpA9QGnToZshfWOak5sMqSrsdg1hHvmzYx8y7Ino
9tKJdjj1k6/ElJAdJFkcSz/zUwDoTGtdSWL7jc6l8KxzvNm4L2ZGSHVHwsrRZ8Bj
l2AwoljA4LX9Yb5Go95A8MOhfPuUbie7+81YqwaNeFdOdZIQhP1MM1Qt2uSirV1s
PEndTlnyGvjcg/ZZAE/3/8Ef2rhFcYUke0eSAwCT6LHme2D/TE5tOhZX/tOqMmnJ
OGEc6nPyW/w2uwGELYkPHdO6FItPqMIo6hnbGmZlP57C0BJ9fIWdrSD4VxtQFye2
JJbueNWdBIscJ/6YcreRMKhI4MVHX9vxp02bGhaptuxN1G5fiFc4Z6z2muclNK9L
5jChS19hbIaXmEpbKhDaL6iKbhIy6QuopKZuSYTkOF61GUoqHD+3QekbuYK2K0Ir
znWXyXxFaBx9MS++GgKZ5BGU5vaHIvdjciQVm55gTnggIO5TDoaehUrsrkWuKt9X
8FNHjfQxSdn9fDkkSaJrdfZRv+18EhFgRQa3LU0m6bMmzjQbB7uU8NKKqdaHR66Q
sKYgM4I43mISjbuMAyoaEElk/JaVb+US4zxwd88bNWplSZDBWJHg9olAdK8l3nxm
/3jm1OYe2/F1EJMNaeb/ioorQ30L3JKyZqByE4zpQnLWB91fyMFsmO8IMzsHTwPW
ha2Hw+OLybeork+R3W6b8gBmvcAhtBF2xQJOvpw0IyDyi96Jl8U/6rvNvH2Dwtpn
JVQQm/Vu5+8Z2roykaJc4JeWdNMBF2sCG3dUK7zUWHzuzGlQ1CW0vZclrM/And3O
zkxy75v5s1anZLQO4B+z1KrIcvVtXr2WqG7cTQT5VWd3d+1B21TIoh0leDyNgI4j
T+XFbQFWgkCog0pAc0MdRcoqpwVNWQ6ja2c1EoVBQigpeJZw3eSSqFHsc3gT2wXL
FEfK9LiuNeIunhFIgndvuQ0P9D9DBf97mU5OT5ugv7VC/RCS37xzHlRx4VR6Ictu
5k15E52q/vINx4DxMsgaa5hXhMIGYkxMiuRoXeqECXRQtuyN2WUmKpNTnBPSajQH
rC0qSn27OMjuHxPESi681nsJ7etHDFReDYI/Pn8T9xaWfhfBdQHdeWSNFqlBQCNy
5qBPtQN2Q2zany63dS7xoAcfq/4VUYqjIzjEQCfPL3izBGcZnVsmfyBV2wNFsAEO
+de6RCKbvrduPGksIhrXFdmQF+wdRZa5b/uACuZq1Vr6hWbhvYXfBCYNMRofH2bu
ji5exG66L1Une+zHAUkcmjykQ8IpB+9m1eftQxLPoyjvL+AhsujTvwcS8wLl0M68
qXzYihkTG3ZOtCOp/Ws3ZLAqfV5VjQBCayevIknIwEPLeTpueKsp7/qxctpku6yU
18qyFhh3hlLwldGKYQPj/ntHkGiRS81NM1PW4NHFxRyMf6ihGUz/cWTfkd5xab2e
w488QjO4qVzqKYbLVuHymbfVc63dfT2BYxCmvtlmwJ4PYlQIeC4lhwwoZUO6h62P
qEOCVjN7BzOaPYf2Faf/sw9Nbr0q9pi11agcdKrsSWUCo0TiJoWCveGTVtcusNqy
9sIXvY8w5+tYAARzNmQ39kkCK5swjll3aazwWB8YgxqBqjTXMZPAF9gi2I6bLQEu
JPqZ6btc57hpF4/437a7lBrjPJU+hSLPciV0+kxu8j4vkmIc5zKaF4yb4dIEh/bO
f1Tmiqqqgn8EfwLMRbJMsnBjkEyCCd7K6my5w0LPz5XDAPHA7JOB1ePHtgDeUOfK
BWMP2TnVlnp12RzkJIUUUDt/g4vSi9doWyTsEYnISOp3q6aPA8M/l7joKw2xYZAU
YWjUstGS7hWgDzKWkNjFjt/AVHWBDCM777pClhYNXwr0fa3rmpOyqH+pfgOVY68w
6xoziecomGaUq1n/VwjRMM/swRH6N+9g0xJOa1Yu5Od9vbKr098zBv/6jv0CEMl4
p8q+nhvWLTLYY7U0f/Iw6C3JP9c8EvYRelI8X8jft0GXD4R0XQX8p6h6GAB1pfC1
ouseSkNhNHe8KzMuP1/IF5WIEK82Fe+BSnmiAo1cJ+3VrIICzNVYx5T3KadjIq/y
CdUMldWfexGUouu6JN3SS8zacQ1sfayrCAbOTCyKFiyPRbxXpZ0JaOLijAYqbWu+
t+1XgP7P737/8xEoQXeBLVBqnJYrDG0IxgTyj3lFN9xAIi46Mh6BPs7og029z1yx
YzWGRj4maMVQFBDFXYz6oe3TbjsQ14k/jWSHp1H1UopQMyvXFKWhixljUC0lN2l3
Ojsqjwu7z4VwmJH2zxoH3D5FGGmZ+vSIgQXX70ELlx9cSrXFuRfpATJPwP6fik03
qwQmBdILIIBrNlUSIc0Jxp0QrJbz8/+mNZ3RBlmByQ8KXvpjlUp6RCYe/D3Ewe7r
qGUDzWMUr8rDTbadgNPCyTpYHDMYjtW5Z7H2HRGUNsG1mvq1tNnvyfipHq5EzlF0
flm/By9+Dk+J1jHCh433T9RzEkdKYlaB621c7zE5dQqBDTAmpsYDoc3EmtDoEruQ
9L809vxfmeNlCPOYmDqxE3jAaAw33e+qX9HVU96t2BeW1WcwYz+Hj1YKBXBlfeaW
DDkuHHJGqLv0rsP7kSnKKPUfZzMSPr7a/z1Im/JI73W4XQkYfenbsUdqiRJU0Wrl
kuipitFZWSsqs2cVhj0XSe2wMrEAW3/1c37CeGMoCMBPN6OkkI8IHHY+vk94v5J/
scpALBfA59cuU2g51rtImQ6dYjYBZbdBTxpwLT3GxmVARumlD0SyP9AvhS0GK+AD
zhhBnh+MQfP0TmvczuFFs7toZm98c86v24js6rJoMXWcLSLHjaj1Ld7pYFL0zGZ1
NeFRd6XjoSgKu2Z4HZsEN/kcLChH44F9RyMFgTRssdSPwdOSjSPyB013OEsJeT30
IarXdjEKW6aycI+KiVHKTDV/3nG+ykkxATqr2cQi1QzJdqxhGSbAOuJ91B5haM5B
hDYT5aM0fUSJQGJzY0Hqp1k/cltPqPfIp0wrzZtlvO2pC0Qqp85IOwcle0WlDa6y
Kxfy0SOryAZHOX7Y3sUyPAcBLYUJ2D0r2qqWhhTb799ugAvNneX5TSBaZ+/POwbs
cH3uqDF7tpZO/kLAlVJa++dJjDmh5A+r6M72DNWfz7ybj9FJHWFJSRzGpfdq2fIh
L3M/O+1f+mhepzB7s6q86f8HJ055GeJ6F5xXmtC4ZAYYl3U/dPNWEQRcT4U7r27+
CuRP23Na3C23cJMZrsofyAFAqp69h8zF47E73PU0REYRHhERMBgOEdWgzwjG+lh6
tl9V5kUmZKBhJu6OZZponKUZQp/ZDpKswQhD0HiUYJ2R9DBYh8aYIZFjMaqel+2Y
70b4LBe9vA+6EyDMmkGsX2qsf2JjoL3wWzLsH1e8xk7O2F7ElCjnUFZqHNZQpeLP
fk2fA1zrgZe+8/o5tK7KyZ++10gnnFTKwVeq2QEEIb3bksxczzUHVb7MkieBH7dC
6je1vBYz8Ik8D1cDrYecNMNJjZ1X1yEeDONJDl5QffzDPSyBXdrCfXjJMi3pV1Zl
1jdYlwRlLRYTEgHzwzeV/lcsSEGfhwWuDXXHxXTfwrdRSuyVEsFSeAkZvu6hIpHZ
kSjw2P+fguFuryju1ZZsnTYjrxEKJJiGg2GOnCvzFMixQjl9NZX6kVQxwvdgZ/5O
hALU5wWySfEZMtmP346nBMn1VR+8+gT+Us1gGKEyKYPZTE9AEeQJsG0PtS3O5MfL
IZmtMKloi7DLYeD+tq6zVth0drE1R6JVcd6vOJmT1z0Q+XhRJs0lSXuyZw06Pc7O
5WIGSSemdb1U+dhFlL+taPvRXIU1WEUhdn2zAKP0g9Fur1ENyikNjpWJoIyJKOKf
LeaBDfYtiYRGyIMxENfmw+fhyQEmu+l3Aj1SUlINKLe23jV7nlsDVBkdSvtNyt/x
xkdYVPZfHhwdN9uQFx9LSdz9xO500c8cdep8U4CoyvplvBwFRzydbo/2Gzfe1+SO
jlhrWWMrOT7hfJK5yfTEXIrIAXlM6f7cnckmYUJBrZA8BiTmzLp4DviHHuDdWNVH
U/V/65e7qgw6GlMH3dSLkxKi6UmwJ9G2PdMclpfGOT7lhfQLEb5czfzwlKx50K7f
BnoU/QCH8y/4Mt9auD8MpAbX+7CLU6G2avHPvb9NPUhIcYSAADidEFD96mTaZpY8
vDtXhzD9EJlO0vLLAlocFumQRcnsS00Bt3pjHGu+nY01wpIwT01RhMeVLGQHvuSr
jyDNcBK3Kz8UHKK1AtTRkbJNXstqwBE3V7ii1IU8nl66/r1PuODV6NToDeZlfiNf
1VseDQ2dk3boWpTpmuFDJQH5tYm0C6DXXhDENauizM/1EHu76Hfr0p9PhcP/aeez
hppE+PZZB1GBXZS06+OdmHqtM1oXIFQ5w1EGhUj6SFEQ3uceGHoPsCBYiaipmWgK
mqlZDI7ECPU02yamHA6kJQcj8p6m9qbtNDfOE8M6NkfZrMNnryOC/561kl3fom2K
LWxl/oKtu5PylQfjhUi1EEfk6MXj8hPxTk2HNNx5V7qr2h7EFg3JMshNa5FgllzZ
DusPTmhXpB/OmIky1iZZDCwg2fgW0sJhlCbf/+YKXQAS+U5bklPdLtlnzHyPA8OM
E1gHZr6l3CODf/XcWNLhfEpnSRVHhM520Ay/XZ6wKV0rRbv302yWex61IF/S0AhJ
Ktd01x+lvTKdvFnYeNBai4eVSLWerv1/m4TrMo0KpJgRS4MGxE6naF7ZOucfh3Jc
to16XzmBgZhtiPnMD+pynyXmDhBElh0TMIsaynJRmVKQ5MiiL10LpL6imYBzPW7V
QQrkS8QJarbvd5tGxt0cOlCjvm7P1DYWjHqSXT0pOCZ5EezuA2DPLEeDPdWiKDWM
nyLDVVgHjulSdoFluF7GlMjA9flHszOPuheacOajh0LCgZYN9ORtCjDFnlHsgIWy
G7BQvEou7vuLg36t2oofodhsCTSaIHnFIr5NHmFHShz5swPAz6UDYq59txSabftO
mZ8Rjpl5QDa962oCld2lal2moKeZPdet4BGoc4AyvwGqaLd91jhlY9M4z2NqVwhI
h15ztuIPuna8+ojIgK9XkWqMM/1E0GRJpui+piiRj3OdTS3a6cikB9Vb8d6Fcztl
NMYjqx9/0QmbPZrIhNeIogHF+Bf3o5FI4Olxn3Z5Ki1iaq16+eSffeBwBzLabOhi
wnhl6gAr3rKQ+J0C9Tjm47MJNw0xJahmV6GOsciKH8HkB6+9N0FDDqNcRQI3WGLN
H05fYEeZpk4+YD2iDqs+CvbTeNrHZG7co9e4ciWqWkmP1EqEeUTw/DZhyixkXsxD
NSjF5Ho0xGXlzoStEdirMe6WDP4KhEgobeWCGW023QsJZCdW+M01ne4qnVpfdhvi
uTNL+zZKbUlWhkDKrn7Sj3DkLuVAWJKIpXXx5AVKDAprJNzkBcqpIonAQeBR/Myo
a+xr7si67mEa9h8YL35GIWl5Jo1L3W9NyvH+pTKODOZD1GTrcgRLG+pIXHbqzPtg
qH1hl9GCoHi5ZkKeJrcEG2S3dVFa6bbafjlDfQdc0mB3WQtRhb8qkz1i/8JHQsDH
lvmlmM0qA0m0GGF0JmuE14p7t0F6PtVATxjzq6LNEBTJ/jK806zaOHQOBz8nMXF9
X39yvSivcpJoEogpFw1st7Xm4vWdqCj81PVpkGzYaRmM1qVElOy3A001aPTYVEvl
Lu0WDvE1jx2qFRTNsBE/dFT+UbVui/qnstdNT3vdTzCR3AmnqoHFXoonEfV98oc1
pNTd2nxwITceYCW1xzaIJLJQtqwqXJ/dyI3RmE3mSn1+mghR6RD/mMj0vnoxylFN
uuI8kE4PMrMRqvJ379pZx7qU+opTYMvQm7aM6+PxdAIN3PNMWylq7fC3hXSyBT1C
74M6KkhhjPTeGE4xz/F14B5dcU9dlNMambD3kIzXKe6dUVsP5BhMWfHlYrY4oFGC
alHGogBgcRSKDcT2OW6pQEjPcboOtcaH9+GTU7KaZR/TBNaKEjB6Mu+AeQBznGfh
p5JwcRdO6yIFmDdU8xVxXTJ+5wrdqH/NR0LN/EDCF7ohWXLm9vq6Due8PpZ/RNAu
CiWDPhRPtlbJWm8x2QloEr2XIpy/V1GP4XuPQr5vObaqwgLnDlFRl7HHphlUGPdd
sXovD6bvKd8gjQQteFiIUQ89CWlC0AD7TxyRDEFvnXAl+dNo0T2R8PHQZfcC/bOZ
eIZbhD3wI2wGymF3NImsTFuin8XiJN4B9wG+RwqIFIOu35Dz96QrPetaZ3AMRGGT
lgsnfHevYiJ805ZoHL/TIJeVePQIL8I5uZqwKWsv7BsjliXi9HjUOEcqrECM3PA5
KCZ2V1bOX6jM8agU+i7Lr31pt/aGiG3JiuJU4wMsbyLfcBwu6BxGPvaqQzZV+nAF
M3UghNqcIaZTpNHP0G06usfZb3WIhUiFZc/jOvUvJVf5DJFS8zYy/8W2wHZVxwgF
1VhsPuCVNMeLsgKEVpE6FpVxd1e0kJqF0+9z880Iez+4WJjTtrujxWX55nndOb65
QXdQHSXxD0shXPLD/T3+Z9axKi3ePAN82G5lPq44N37DwXmj2uk3GI56J1P967Pb
co4SWCNIRfYprJwBrP1hAOKmwnQwD6nKPpe1jrSjiT6jZUxZunslf6g5SYwezkZF
7o5pYUuJgI+ec7ocydifgG62he8loixmegtKVvW/Wp/vvOKzo4DDEaVhHvI0in3n
iYh4REnrCy41g9rlIhLv9De4Z5bDkp/BWb9io5DzFx9Hi9x/0AxasWMz1ca4jd4S
J5TxetNKavM8jWRa2gzgFqljiHh/S7bOwInoxpEnfo+rp8s2lpx504/D8eLVYq0d
Q5XNjFEN7OxWkJd0skKg/thfLBM7l+ePHOQU3pgW6zZaisVtf/jz6JQNX7RghO2o
zsp8b8EN0GoQaJeHIpkjLN9vTid5CuUn5AIbPrkYEo5alG94XMz4mZHOeT32n3JQ
a0NshFzN4vd6AkJhdiWnQiMAPfgXSMY6OzGZTV62kpAhN8uCxs09fOCG9bTC4NoI
zuqja8ukoGOIiXJJuIByI3DM+LmVgXEjnk2ijGSnSSOx/N14fshGuxJroAFgtWH5
ippNBQKZSQgRAzBXfqUA8nIhXWS/6ZQR5gJMck6r+CJeiGvx3vBp/AHlakHhgCJU
Q3E7ezVTUDjLZqO4SymK3pReJ7Q3nuUaYzV1wbkLw/dNoorMpbbUd6+pcKCeaXAt
2oUhPPAEIrk9gVYUfJAUjNmy4uSrHNdDId3KSUx2Hf6wXaG+WAhR9+ZCjSKgtplR
/Nt2HJh9B6JxQ9uFaeCqQR9+eAxN4WidJTcOVvbgYEngeA+ttTNLWMN7Qzi/LKUh
vTnVgrUKySLsGtg2avgovGsGTgv10NFe2YhUeqiAdcpQUcuqofphrY/6eoq9X/BW
bJM9xzLPSJ5+mqKoLkfU51Cyv7tKBHwFo6aVBeaFKCo4OG79MNbhkyJJE+Z1SKjd
AbuzTYF2/5gV8SPBQ+W5wHa8FCRHABBr67crvvNfmMCleT6ZjozPks2HWuZFLQVY
tymZyZXmatpGa2i3m786eRO9e0lf34gOKIDhA1Yo5NuTg4QpgBv+j8XOP8xSvOmn
hrVQMC9OcYWlt4Zc2vnV31u1wPlRJIsysjXpUn93ExMAvkwD0fPQTSmIB87ZcQEm
M2a35opdfjpOZ/RA5L92QAqD7tkhZsQmWy5MXDVN05aBOTS1lfYIG36x7dQhvIEE
e/h3HzbIMlyEwOP0WzQiKxWkMWhARvN2Veo95BsxRWwpT4v+6RDfU3BbujcTn3tg
AKoQvv/rWomwhF9XILSJU2GeG4iIxH00w4v8puPl+VFso0o6/tDg+FwHIfw2qH/x
vaJ3l55R4kkfAIlidgvRSzWy4eLaEZCQbqYVHGlo8/H8s6vZsNqm+VmtK+QgRmKJ
bW4YSp5v3UDXcRBfTdIagMdO6+Iz1e7z0eWrDXR7RzHtLNMl/Y1Lbt3dy85lMcRm
ORDyIhr/70sfuN+SjUIHM5AVjTOYJ4RSQjEQYWBJxNqk4brFBAk8rVs3EiacOODa
45NAzRC6OtCALC5vQ0whN71JxyACXEMnKoaMoM02kiq4GmV1hCGlS/Z3wv6WBo3S
B5cImdezAc0MiL9EDxiUdUg2cck0CfqzBdLg7m8SnvVifeGdkee0gPsVmxnfedtP
3Sp6InA7bInZGG0hvI+ERrG4muUcFvy0sO5SKxLZBB8KzGcM1IAkqTuib9EF3eHe
grXrOpkFuIq2q+va0fyHVOZqnTqvd5anTFRqrGmQcXk39sXUk4EquYX/hXRvZ+V8
xPk07/wBEZwXR+AZpJ2C6e7twmHRAy6T/0EkPAcB1HK+gF/mkLsEyXW4VLOwbw+G
ppLQll4i8vCyn49OQus9hj+KWtJRf7wuiccUBJys3OqT1nQKlSxGDd1EC01+8gwG
UoqEBTl7jNevx71OKWwHChJe4hdlFLyXR/qveAsY9LCYP5eOEBlP3Ni95EwDe7oV
ju2Z5GXqSjp0hcryH6fmBCH0yWlsXW0ZXKuqIkiG9cGSY7vKwKFV1pPSG2kY3iXk
EfjGktSc9YySGeXw9FAIE/PpyWtn0Ehft1LLZ26lpxgy/k/9n53yl2u2hnd5ZVTO
6A5wkbeA1INhpNOyX7myy4jaGpuUl9ozNzkeZZiAQrpioQq/TE1/SmATFKW/3KyZ
mLynx7B/+Zw6tFq20fVdvpCPi4AQtCZ2UZwMxWAYrEbcTjRyZHtrwU9eX7HGZxrG
gG5WEMjZ18LrzxIL8SOGHLsjHa+CT73KavBfh4H/LFGXDB/fUEIWSB10UsManPAS
chACIw28BKMlkZnSPyg9RZPdiTM1P3y8C/v338o6VUHPWSBFfIu1z2tYS0BYoyYt
QrLQHZe7rLTzYwXxi5hLtAMluQxL6TmeJwfi3n22Db8XR+JR2f24RXIj9izs2qkq
kXzWIJPOUcbSn1BTDcdB1bAdj6biy+JcUMBELlZuyxvLCkg7E61cUBYF/xKRd4ii
XA33oRMKuXTLHKw+WkKA4tfforfmHlqyjmK9fzglIng8FqhX1NvOGJ2Zb5aMG3Qw
d/7Xdh7JQvKbJa9TGv75fwMpEqwoTrLfNjQ2rrQnQRDEQDvH6wahglbDo0yJ4+2T
07BpGM09azGiwqiWdJKDnk4qCefm+tyJjmGL04aupFL2B8UIHJiefF4s0+KAu+hx
RPeG8tJzpGWI+VvnY0v+LUevwgcgklKjQpxSGu2xL0/LFPGN9PaAmczS294nPXtE
mmifIBs7vzHTesbYx0Ek3I9vYAmgKtDHWud76zsr5PSYPtzN9P90XVaLOKiyklID
F7+FmGmNiTCCn2vTfGTr5BHusJ0nLz/0Y+zsa/TTnsW3hMT/yhDd3RNnbGqSL4mR
Sb553wJWQVYO9lAzT4aL6vrOeoCMc5Z8y0Gy3UvgpxhVcxXPCC8Ae8THTpIFprtP
iHXEUA0I9GYWSRtk9h0Wnp2YzjjHLQrFQt4nKGPPKbdUsZuGDAUjrj5ZbOe/BBXP
CEwTLly9Z9+yEBL9cBxbhnmSOKLQATVv7Ck3z5ujhd38byttHFGrkEsVksh3akrd
hfZeOgXHdmGPKeszFYVqkSgWxsSC7Qonh3sovxDo3C/TxwpTbDtoAMNkKAZB6ymi
AJnMMaRe8QNng4c01u289DgRvRsH/Ym6IpVhoa1GX+cR1cS0C3uZ6Dez2id5z0C/
KWg7oaLCt20CcPHFzbwh/YMN9rq5w9KKUhFodln3Y/TsiavlxP++byknEJf2GSwz
d8IcyXON2QLbtXGafVh1i9fH5eRtLlCgI6P/zv2k3go4Oi+8TpAiZRmhKxie868A
wHNZuRYDRi+9QXfdFQFdIcXKvZwazO2yQT7nXMmvRllSCNYecKEXzDPjnwoC1LTt
IA8OykgMDiKg4uDc7ZuAMk5N46SrrEgIEEWxbhX9pMgab1rHIqCXuMCKJSXTalX9
2gNl4z2IqgdTlWrPluaHpb2IK9iUzHiHsSfJImXYSgypTl6hfxC8d2qAvYp49Npj
mcxkIEJN7xSE2DBkq8iVo1tpWRL0dt7fqv8Bc0AwkxjJpoMu3DDFeswvTz+NuciK
wkWi0R7k/moR1+/exSpIBcwuDliqOj7iBdzc6ZC6ybgjO875IrovHBMSIONkJCzQ
yK+ZkjR4/bd1Ga96ssNSIRs3a9llk9B52BBPUzl2NnSg5fkgTF9fWnrHnEs3+Y+U
DienVsFKQxxqsrm/szDTfn79Qw/SAf7wFRtNqn9+ZubfDzHE4XXpZ2/3UffaLY/o
xnTseT2jz3yLJfZyU13ptt4nwvmml9AKCznnV8frXHUEQWegXzL/4q/q3zD/dHCY
xnOlsczYupenb0m9en+DzzcFHjZ1Y9aCy013Cr+T14j8oKpHRoaYHBm6Yr+E7R8V
SJyHrZvKSgWk3lREElGzdtHe8SqvQoThd5FiX3lTPKXy6nePo7FAgonLAhpbKC3q
t0YJMDgdVBxBNAUkO78G3Ahfe9j7CNIira1NVNj2Epanmn/wCv9UjDzLTRFVnmtM
yZ6ZbyysiGIMe8NBsrZ1/5uQhXPh8NmToB69e8Etkys2tyctc31AQz8w1JoXzXMM
N29abk/P1eA1xEGAU5arCeJB2k/PbouHdMdpRudMQoV9Uh7jAgTW22v6IL6MF7BT
9bDGldk2FK/EoClfIb2puia1/5UWLFWvHBq4oP/N9cTrMce/FG8lUM6pSS43EXE8
7Txj+vrSs/hL3wIwG+1ITPyKjeH463L7McLiGtQ4rwtHnnSsPzZeL2bYNvp5y/0F
jszvUdJNU8D0FyK722VPpXfYFg7Fj/dFsSZAFVOwYTp8frHZTKyw3W3bVuMTsnZZ
AuXz7a7MqYFP4yKp/b1b0DMN9Ie2C2iUvzLbHc1UWIP/WK34fiDAm9SKa8U+xLLH
cWVjmu+kC7dZmjaiRZXzAZzWaNhPNkSgOc8SkgrUP9uHJx2t2yGtQPG+DSvPabYY
g1tnh1sgNrL25NoVYbsx8p/VBqFltrLxfmBr2zy/DtyFCKPN/T5iwDF6KfT4726+
l6AK+792oFiYqm1zLsjez9d2+4TKavlkX8Jc0fQuKHjs5vaFWmuJ3CuaqdeujBec
Yv2fvbUYgvYyx53zDcTTxlBNczGrliAF+4VNYuZCWJN/1B3H9V+JUbs8FPMEeML5
RB3oiANNGpuKJTN3KvH6PjYLWHesGa51lnb/svUyrTx+L1Df4yIZfaf98wjAPBJL
EZbTdiIdI2AP6U3rCSuuKb20xpSKsjX22iY5+ceLy8JCP0HjPmmJIx8W84FZkBiB
eR7v5BGlCQIvGrO6CFTaRO8vgVgzsDmdosIUjCCi0gZttY68AM3ci8qZ6eCmbQLs
LZBufgbjtXebc1RrbaukkJx62rxTHKII8WJtbRqvlaSrD8OlhQfzU/Mjc7LmJnva
iZd5ew+jKt8dOboBlG+lzwToEkrV5xhIYDbE9sn38g2oGvjbdJtOWl5JDJpI+Vkx
nSVvwuZDQGy8uJbRO1HykYFBioRv0qhCgrFdZxa2HHIgvtX4c1LI9RyPUARdo21X
czq1b6oLsf42C4zFLWjTcnpB9L+9R3wqJYWmxOniN02/eYs1ECcIIAHYwZvZ5A7X
fZKH0u4y8nkuFXCkHJ3b/k8h6Paksis+jtSBDjOx6VTfscNgTiVe2YTV/VgViWiP
FhB0xDz8TuiGiAXosEAe8U5LXZYVTG8xCsuBNRdIsCc+PAeP2Iv+bqxeP/f71g13
sAQ1hH0hPwGOU/DA8gJk7QPKzRmOwAdOMjA70Nq0/q6S4ygYUwckKcqRWSu6F72Z
YrAXxPePxkKV+7AC1PvtmD5cahI4/j0Na4K2IzKEVLQ7VE0XUxJuqIO8W2mDOTyq
gM+iycYXmWB6RN6X9QeMscFjV6eTj70A7KCmSFAYuzpuj7w5WEkshoiI8Z2pJBU9
rJteIE4PPpATud+ddBdJQhNKWzTxnOohrLTuDIMNZN+Oss3eR+AYWRQZQhTKgTcD
PTuuwY/u8g3n7f3zqV1Ep+vtkqsEeTW746KMDEbwpNAmkAAholkif0gGlWmmrQ/1
GOxwQ2De97J5RE5PPKnFSIAnmHIEAfvYER87asAhq/M0NEJqHTvsrsAcsFFqf8I0
M5X3xPCf5lKDgn8C4hqfArRvg+ZZwpSaF9hKw22Dxz3y/94BDHnjIigY4vbEuJLH
u+gCPG++w+QsAUfGoefR2T4Nhjbu0KoSXr3RdnOhkjjEno7Y/6Fcsd9FWwqZDssL
kDU/P1mY/8n785VJk9vQFlDjyq04qolCK8DSqZiluadaufEvmI7SUc8mfUO/Gudf
6powaEYmgbqOVClnLdUgE3IL9ZrS1YTYC9fopB01rxR0DWSKNwglHs4jMIqhequA
LFAgOUSvra59liTAWyY6t+qhwrDtOVF+jG5X1pn8M2Qquhw3Q5SRmWUhlggTgnpJ
1giiWgmaxEMTP3Y4nxNXL09JjVi8xTqx7waJDe4cHqWqB0xzcwZWETE0lYP539n9
eqIiAdNJHEz8Q9NpDRrcVcfID6L6mzaHcW3Jxd4emyt3AhkIl2Vww8m22UJnTJR2
DW4bHqwvMfifDYbrat/PgbaArtcVC7joE0hIODvk+57qbn6AgJYXSNug6LJvlS1Z
qgXNFxJMUtrERse7HFlmgvkpHDOSwRcghPWek3UkjW9By4Y/OUYetMk37LLspWyt
wgEN8QW6mR7iaJ4h8tXGFn076HO5deg0NXgyUVVNDFKZtrI7eEj9kkuGWznz6qvW
7IyRif3pbJSk4kD4zmo6Yy3ih/HVpLkp1wpOBYWEe88rE12y0RXBTaLV1Hv/izuz
+JOBcSfO1yXVrTeEnn6EINV4VM1kAD7hIM/tIRaXPWlwPnGbRBTaKQNk/d7lP+FL
WnPI58Nz+ftDDIkrLnKP+oqM6R5S0zd+2eDwtsh4LXpi9RJRgGNB0sHtQIGtBvWi
2sKFHt3RWYDENrUYu41TT2Mkn+yY/gMmxdcIWl44PZR4hAMuR09N4gElH7erEUn4
+GbhTTMiOafhSgmefaW7xblV9x8M59Fp9wVathBQEk782pUNMSJ0lKfHZcsmCjfQ
PHfVSnuA7nI2oVjqM+ljjllV8HT6DFF/LCQImwmJhfdT6/vNTCaALhPqTtEo1sJ+
Pi4PhF1TMG2QfqD8UaloOh0veolP5n7cWxxA02A6np8zaMqCfMY17bhtJH8Ewoip
3nkgJCgljGSJqzQ5GLviK92P29CJl6U/o9sscXyqoI7AVLhQD2Pk7ZNLJEX/uyP2
NSnGryYVDpadqvZAvkt038IZjmX7sH8Cji7VXuI5GknvXTfrh5HhuTxjN1n4h+SU
3UPYUxUjPuMd90A5wQY6oeiX5MLVRtPOotKAtg9CU1R5IzG3W1ppVWWDQtAhvipB
uUadMlNS9pydJlclJ3aABDYrM4KhFM7rJXpjRAbQPv7tK8flZAalTKjIXU6ODWLS
hutXxvTplR1dKhr78RMPS8/BAQVwku5Oxjo9r1vcGePgbF4woGoS4essU2G6asM9
JfP44KKhRaauklBnt42AvanWbkPmxZuLnngPwA1VBE3inZCeqlsFJlUd1gFNAgd7
ISM1fVcD7icG8eYJfrKPZnHIHcBMu/BH1j4kW+Cf3wpK19fUx6sGCySqZ1Z0Q/dm
xET1GW3gAvYBtqNiqoPgziIwZ0Nh6QOx468A6bEVcyUGtrC+AHpnIe3lvGvwzpKh
nc9Uel+endZlJWbv3KHpLISeqeJmk1UlnTvm3WBH4D6DsFzRMlGI1OahZotHKoLC
87FMrDSTZuaZOKEiYjmyHrSHronhodPW6RorquTo1Ocro2IVBsTyiyARgmzinYuC
psWNoaOaGek0J0I7+/13MaJf6A6nWxi3KXU+GPSL1Btt7axF1XF7zFCmdFKUGRBn
+yTnySctMoYNFLXGu0KjwdCyRY5cKn5cgVP2QURj5jZRWMTjVU1VaJqnxLd32SDV
KePjDA+oBXeeVKw7i0Hr8qOSOZwcCfolWHR5TwHH/N7YML4L/7Yb10f54vofF1DI
1jEXbaFKWHV44bulFL6HgeSKlm/K2dToRrJ/jGmzgXXj+/ZgCXUhgKNitdOQKbhd
a+9rw/Dz3ZdcYOXmyACAfC7VeByYOFAc0egp1+tAK38BlcGBeeSNA9IWAkoBahqs
1+HO7MjVuLQFA/RnIWAVV668YCToD6q/hWlexd5f1q2jbHUN05kgqFWTza63Wa9Z
B/mY4YUOCU4f3SPkixfZwwihiZ2uz/DmsClljHxXWKFBuFcS/bIHmef4ta7qqnnY
wFjFFgfuxOEzlStDXOLj38q9ikcGt+RdtJiqYMGrtm82R80cZYU7Gm4weLvURF4/
1zSclNX1ml+Sm4TxW9tJKyzv/CMaL3d5JM1KcYCXQFQpWOr3ei6z+okgaJY7hqte
CmEAz1SgbcFb6fSKq8YGAZyDmvMY03DekT1bIBzG8f+clTQTmxs5RjFO66wWNCLO
W5Nc60ekAMqkmfd8QZWQIHhKsxZNZQ6T3JHo/UKU7dmyDUxGg3FG+mww5Bar87Jb
jlva2oUDYqPqII0dhu+i5yfa5OH+KAeVsx1KeFjM/2DWpnb5rCS6dTXxzfHmxLwg
PdZlOdXgtRTuTAQl4hVnvuPwESYNrpt2TC+iYp8b+rXiu6KKKxP4st/FI/l6g7jO
AQu28S6EEtI5NRX41NYUIYzwXzPH03y+r1JDbhXBbYuz3aGypynpgpH/9t9vmHF5
icEkDMYIpMxUHsfwJ26eQ66ByC7qTTsHiWFYp3eW3tjCauTs2Pu9unQporlG/ZaT
hr2q3vUyIMxk6t+lm6mfDR/n0OAI2PJusIQG904ue4gSIlbcePeYI7dhRR5SLSIp
rqSzsTekEqX6iPx+yBNNwDqDwSAN3mjkghTTgj/Vy8Aygcn1fY00tQXgefKJWVdQ
QBGuU2hKtd/mTxC7NC4vHJsRlW5DQUlEJR/CjWyDisH7CiSYjUVs+KeLKpIr52l2
x5T9EF8J/X3sEIIClkIZ3Yrs5nwQ1HHhDqUx3plnWmVrfPQ/GlT8Ryk9QjTQBK3d
YlPiAq2Q+iwDKlzGXLsxRCDanwnx5CFfbx8nd6Kwp2YK2HUUu9pJ5ufwb0Qe/tTZ
Yu8/Zrm70SbI06hP0Ym5LgmM6hkJmGGN67m1HD6isB4LUj3EyDUyYS4XuxKRBUnR
4xtgVDZQxO+rRXq78/drkzuPASKKxHGAZg8tXweKNfydZ8jhWMt2JW1ivGt6n9Kg
deC2SBw1hdgKiMTdD7mZTQdQMdmobXE/5YY+RzMyr0dvyPyfyqb3DeM/FtPdqvpL
9gxhqsDI/yGztI38ApSLgaOi/+ob7eOhCCDgWbX3eE/BwTdGJ6lyCUH0jisq4AFy
M7+LnkJ/qZVqGiXlnc6iQJIIN1GywDuBMEtdPLR+76sl3zGFyuUIYV/ZPnBksqT0
M4WRT06UkrJhzAkwj/lcgy19qSKSHlNJbdHchNER0Bk4flqOqzo5OtTmDD/vDgpw
jM5WhGTq3h/TsMIJw3OKCN3GUBgVzMH7zC9+KNOYHRLKu4dnOvNYKFoaYXH7j7RM
2RJDVlpDX6oGY0iaPz7UChdA3vRRHbB30/5C/ajY0/QPsuPrSBQe3nhJ3lWjtXnc
m45hMmIXg+ILYqWpaWSzogi4S49QWiy7h5NfEZLakpqq7YhkClsKPmAq18AvJX6g
7PcO7jDJjne1HNo6UMROufV3p7XVNuQt0au6uMLVaDfVGhVNpWbCghAdwRHZkeme
8ECoB6SpuZLY75glNsBN4klWZr4Kqk8B90h+pue/H5j1WmDsrIg6J4lVa5jqegY1
ib+220UpkEBaOxgMNq0qA99yl40nCjxTqh1khOsogfb29wKJdm2BSA25pA5GVOxB
edz2WXwNfnlu4yQAoHhN9ZUj/QkeeANzLUgceAT5VANVK+9Biwf+yBgL3wFYahm0
0jIRFsJ5bESTaumSxooL13vMDwMsANWJQKdKtQlx8l+LC2uT7pzwZV71Oc9zB1XL
KQEGy7F8GFRpiEhdbSUrLLv32kgo3yI7IRQDxync1fVSGJA1yAu3dYtIc0sDlbxo
el2zrrgwfJMJKLEKWe2a6ymC8vqrBwLJiukCprZryApZiY1zKB3/AmO8jFYF6anC
uaHPQOLBG802NXBVqhggZ3UiOlTzEhPk6dvOhRjV5oErYHyD4nVglR6LZOi8nNY4
ZBHmvr58Y9G+dVs6yRoLoyBIa23n/kCbh/HMSkFPoa/JE45SCRBitRRhbwNKN9nW
dw92wldb/URjgDAepY11US/YTeTNIUgGUlMkCcHYfmnRRxwOR6VxLmGId9XfGukd
qAh/kKvZcrbNUleFVXcuNmNP57J16l+TK3/rYRL/vLB13vz8GRznG3MAfuGSoZXD
ge1lliUe8qJ8rGJHpeiG36mlZ2HV5btdS2cak8tjKNGfmSd2TWh8biV4pDy+/qe3
fkQ1REXD5F4KG+WSkOuDgaLt1KzUonxFhXhC0TpSIb2YR407PGb+WW0F+mH87q1p
59FZMLmnJU2VFaYrTxItEpvRBd0+EeOKKftbxdJoyJxK6SfRojoeYkcvuvVdaAKV
9DuuCx65XIfi1KPbcyXLZPsvijrRnTCVmZiB+4ZDBJJv0ywChniQn917OmnGgLdI
rF6lYZCRDA9BdShDFiQIj88d3jCD03LoCU7v1p0VLLWNci3ubX312AtJxzydp17c
IS2POwuoxA9hurbbarSMd4jk3vWCCaRLY7Bk2oEsMwydQu/HRp0AxHEcrzsEqUCQ
hPSULSOidpWBGVG74x+e6xBO30PkOfbmVjySPVyYSu9PcNc4iLBkHTQdz8bPbHGj
ekeix5kh+Me3I3mDUQoRPRRRJJFu7LmvGGrIXz9tAkesi8ODAzieH1niYhXbMCnD
UwCmoa6fSdAjfLyVVTSed5lHw+4HSVHui/3IT9PajJxIwfa2Hpydj8bzYliCzt6q
RqNv9jeniaAQt2sMhpDzuxKUM86Wb3k7GvZIoB9NDoCLgZZdkcaow7ueaeSQ2wFI
AhsvziFC62mq+RzgYWGdREVzsDrCm3EuiZ7/Q+soEyaC7zFWbzlQnO2clUhq2EP7
n6HwR+G4w2ExvXtgKENV8cE9XL3CqAHWj5F3hjAa+SJr0U+kD/LHHGGaWpnFc3DM
neK3/BKHWJ9V5p0lZFtIEfoYNBP9LGmtkyQrMjmMHHfNUoHgcE46XxeKiezQSuqF
ahaKVtDW+jLT3WOwg6lNaBttE/fa0NQnWlfSL8jmZHnuYFhMkYXsXTA/rcxp7pN9
XnVbVE/EHuVoAxWcCzvHfHzYw1VCBa/PvuYAiIvel7Ty90C/D9Mo8d4Xt4f7wbLs
F4tY75Sq6cVnMIUU1wUZo4IFcTqyCEz1JVxPQDqnx+FjACMFEr387paKoH/dUFTy
uaV7D1kAYzu666fapv3amng+bieDYUAHdQ1q67BwrKXQN3jfC+bmD2tnyjE7b0UK
Zi+HcElTaTE2J37o4hfb8yAlyK440is/hvTR2zHROf6fpBk5HRpsfMN4/MW2YGsU
r9vfuRFCWg75SG1Eqx9i9BGxVDbUoEbBwX4pG070eaERmUVCKqsmOlKStJbu2//u
cpC06oTSb7G5DCNDd07Ev5CA5w5TgXDlEiK1UyGBi/4GtOx5ITCWgO1I0poUrjJJ
bxyj2T5KjZx0b19IT31jFEbRYW3oLSgXSPnIqIjY8LGQdrDPOoaAS5EfJbIXQct0
zYDyebIwPAKYP2Kvjg5DR4lxmD/ri/RGVsZEOsk6c/pIXMSXK+j1e9Xn76RH71oF
IBlKrfnlW7YIqSArJlhsDBJxMieoi7c6yqmZLg+QqRc=
`pragma protect end_protected
