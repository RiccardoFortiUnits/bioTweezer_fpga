`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TiiqsVeW/jdHtXOrMsfG2ECUaqoyqZxemm83u8b5xSsmIoh45gknPxP9ASjgx/oU
x5KVcFckFcwHCdn9K0JxFSyDXIabcrDJwOrkqEmhIAxXIe88MLVnpVt5xTaJ0Uev
YNCsSdS2Zsq6vQQQPu9NW/oecNbOhDkKyMVFflQ8sgw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25648)
SXpk7E8M2P0xXOrab+7eplda3MQhJT2UWN9wbqXHgcnbl0unBXFcM0S4FEkRRI13
pTHaFilKfxtW2S1nHlnDZ3yoELu+0ngCrYuEdUzo5ta59WL/h6lcapkC0Xe9fotE
CP9avcH9FYbRC96yM/vG42XY9x+jY5b9Duhm1yYxQf1NAvvnXq1E/8n6tK11HxIF
Ij4K34VSpEAicRrTisFKCUFEsRRVpovAUbC8R2CLxoDQF9rAxfRvf/qxxm+4rvZq
CughXdiKZHM92Rk4fvFQgxysHs4LKI9mvPdCLPQfbRCeRrXBF3x+C3u3xEDeg+y/
fZun+l3O+840OtQeEZqVNtNas4nIQUwlnsg6sGVie2WvugD6Krma1cI42ZswQuFu
6D5uuLsSQvicByfXUzmjpmIL3OIngmY74njXNMKeP1oHJfJP6jhw3S9WSVpi/PSR
ybLurvNbj53zJbbVaUsTJaQLMcOnow+wgXCpVNi2kZe4af7bfr4H80cgfyF+2i0j
igwzNI8CByL8A78pTLRGyIASqniQUUE44udZO2JKBcK+/sBmcMwslD3yaKZftBQ4
clOqhrFslK7MT6WGUGKapWq4+FZC2lgIZaHt7Tm2PiEEe8loVC208hzIqISgymlY
ZAVafg0c2IEHQ2TiQ2m+iZcLtZjEfjqPuIxlQcndDrjpE4LdXvXy05aCqLu7xiCf
Exs+1CcoC5VSGnpRB6NdXv3D7glpmxrXrVcWmosLisMzfDp+Os0d3LY+IQaUvHZA
vb8+RvO/XezhcQMC0ck5di6luKSp5YVgQxgXc+7mhSVR8KBra/2oEvhxLnXjDLUj
ysgd2fUY3NvLIMwJPuCA0RYeKvQO3QKeVxSqzoHrudJKuukhhaKuAoElScc5f3WI
tMAaNPdDRRx7itrkrugnVoElVMxK3CAGCN14rt4hBqQZOJo1EhmoyzsFhc/1SPwp
kIsqqTjOyvkbiN+fwr1g3WAmI5J3YpD7m47ia3GHWu3afCBfrFKd++7GAUF3i/rM
YA7oxWR/OV0LnEPfqvzbx1YAkKW4V3i+aYAzk2Rert5jGVRT9RAwQj7SMbw9rFMP
cNH9w/yuKiKrujGJgzirpzy45K9OW3CfTy42JDsR1MciwBO971Fpw+GH00S7dDXO
UtghU90RN04WyuVQwXSrbivE2ldALDNEN8ie0DkWdKyd3aGCXo+eK9fR/HwF7R2/
GZglcZ+/Ej5MLeKupJTajY58LZnRQkHJuSyOYG9N1KtWshbq12RdnfkBWYeZfvXf
AI+qOwTrPS52trlIXP26dMFyYEFyrn6RxCLG4WlyAAmT8/X/a8T+ShAICq3SgI6B
WLdpIOPRo34TinGumcYhwObXLpMMlb/7oxtR3SaIFhRuHm943Byfu3ubIVFC9vRJ
HoPL3+ZgUC21il6jGKwOL/bOEV6C8RVbzG+/l0jWFV8ICwYsXPzqnkgtSGHiSSsR
ARLOhr0fB8K56XjMRdcOeNbWD3cKISR7HE56PYZW4UsqaoGvVW/qVKVcvLa3UzbH
Mg3h/ug4SGqK72otT6G+2p/kTsYAPTAkGVaMhRVJZ2c6rr9Hl9XDzJaKeN0FTUsP
MwZ5TJwwe7ffgy6lCycOcREn88AT95PgGcA4vRk/PPhi5AlaZTYSdF2c4/9gDAgF
clfm9nam853DOjnD+0Xnqht4hXHJCnYbtfmMLgmzvdrR1xQkhRConzFmsWFo7dta
ZWe27Uc6chHlm9ATh+HyVN6+fho1i/gLtAMX+8NsF4fgG1zAkDdea3cWcYfltGiV
fqpu5kQOQQMzY9fuN47gJIqpamW/YSAZnBDOZdJaciCFQPRZ0dkFDNZJOY0ScuIc
ka8cDIRUYl7cTxiNOWj/eb7HoS+4RQqJgZKzGTGTV/UX1wqPye8WxJ9pnwtNMClV
U8txT8fBYSjqqTVvjG5C7+tBD36sLGWl9/FqSXk+Pj6Ci+L/zSlL6kjXJDs2TLQW
kNq/xr5VqqAAQka2vMhSr5P5BdsttgIoSWuHBKcsHp8+PUqm9ny4Ot/yRB3Yaur4
kYqYo3C54oDNZyfdRRKX6hxJ/5AeioD+C84xkX2tKzOapIBbvaEPdlYQzOtmTwu7
JnPkgJhhiz1YhDc3Q3nFz2vD/sVazHT4LuAVXBogWicBlev3et2ZYSTIKt/aCx/t
xnKH7hIXDadr7B9oEXlGByLVbKYn3bm7mpO3OtgciRatSQIJyTh8DxzFCImSJujX
Ip+Ng7rFqQCQJHbOlEiFCe2GzAlsln5A8zHMOlqHL2gj6b2Zsb0b8+SLFvCDYZgY
jaykLkD/eqjXhAU/fkZEu6mQERUeKzfxfxLFqw6at/hz5xJL/0+BM7dfkkNMNVPD
sK5lielSE2oQT2wkyFSA0hf9M48WQNLPn4gf/Uptg+5f+bl1R5mTNNaaX2rd+yio
E53TNASfFAyYACppn10qK3BZRqr8rDk9ftHada6nIu+Gsj+F45tI92BTwfY6p7gh
vJQncA2ttVk8xIGl1xzRGMVW8Ot8OJiTE9qw6m05uiB1UWd8yhX7ZVWi7JkNxQA6
g5RwArph+RuwL6/mlgi2d5cGjOQENdOXd+vvS+FyLysiDt8l+BJdf8mYd1qAbbiH
W3f6bkTwtLjc5i3p4RLksWxvAlqCKStJ7vDlGQqW1mnsa31fpJzBF2ZCrLrNa0qk
NEH9cIPpGehk/9l/XTxPFHO0vgTnY/v+bXitYakVlGnae9sVow3hcNU4uQRG7dXI
wHC7erbaWSXDDVu7Bx0ckW2rPZT+Z2qEi5Ggtn2vr4K7/t4BlSbv/eQ0Wl9FuNHA
WmjR4y0CO+bl+hPSO5cZkkOwcdkHsrQPIXGdqlQS07Sz/y/phuUxGsEq0HludJh9
tzJ3xXY8YrXco89fqNxe8f2DiFGd8KxcveInWx40sSknWimOFsIuGkF4Q6wNFvDQ
ix9Ng0nvG01YdCNSljQ0+8xeBuJ4iW9ZQ3s7T/UgX/u+0gsy7fIJ0/aHKUcjPsxw
OlEZdVyRqnevvK1eJPx22xtkE1BB+FpjWv4BuolEN9P+udWz4bIKy0EUeyZ4auar
kd6BOg1dfEVuisO8dDzynTKZi+nZDqxPWhqo3vLQ8ZqaAyODyNeGrTYnwjoQ6oL6
SvpWznXEw/X7XT9BYpvxlmxVp0XslC62K7MsvRouU/7gYIYPTKdRdsxiowyHvhcP
XK6vdjT8mESA/VVK+ta+omuUMq5ZGew21iU7M2H20OMQP30pRsAie6jQuAsJizhz
ohiX7liFyo+86YOYKuTtJWY5SSMf2sG+5QK5+HGwKa4l8KIkRwrieqGmJmq2Mmy0
LASNLuCsGW+wCekLv8Or8ZAD+7jFyDVORCm9sixCmBAy16oqeOOUMUn0NTkak89m
1y8GLe5R4r2tV35JTSz4l8bh/7XFl1hzpUAx7tUMEP7Ae5pfzBIRP9XcdmYUx97B
ULWrLrjWgTI5pa3CquFQK51x3x+r5p2lp8QlcS6ZRXCwQM3UYJiAxm2/sVFGmXVI
ZlIhTZQymPjaZAfB314iIT7AtTbECbyl8cIGpTNwo9+8F2dfgxqlLTNO//SZ2hbL
f6FloYaWHG/jfCPWxCRR0Vvrr1Hw4RizKfQFDpLdlFMbTB9Wag+8RaQXhvg9y0tT
Gu3bP5f9LtCuZC5J0jMfiLEnfe8CmYADqiISZ4Qv74ayhM0H8pTMUYQmXpJf10V1
DG/w1Ymv0TlR9dMuwPGGz4+M+ECwo5eS4m4kM79HO2irAwKy8Vikm5ZLlJWVb2Wv
u5SoLvoW1WhnmE9Zmh7nVzixWuP2K0daIW47ab8XuJwF8sJDpn06bj0u00ASAPdk
8WKmjiGagv4zyXfSJ5SM+BEOWa36D/Nf3K1SiAMzY5+zfUeubfo4DeY4wnyDw3TA
BDNEauGHrKMbVVza2TRC3Jh7i9Pv9q6JQjQWd6+uqmHR3St/nGuF4znr7CUXXkoL
eITDx6lLlDcp6bIlLynMQh+i91hdaD6+gOHg3yKERaUjqJUulPxEqVCD5eoU7gG8
54c/bUt4sJWQhUxrAXuG55JimPZtaibqQh2ii2DU76KUj9TnTWfPuc1jxMBRPQGt
ot9ABioz/+q39njeGq6Nwur7sQUmUWLUNBocx9yn0ckTi/MXIk5ICp98WUoCmmPb
2s3d2WW+PwANrf3D1VkQ+/0U2L8wIw0+9u4xTe/20LgKukgly3A/qp7SNPT6OQmQ
vUEeVM5lE/5wefYuPyi5spULKbWsZ2kQ81POzXYQA+j6vY2nnzXyCc1dfO+qGuwB
bRNuDgR7iLuAuWrWbBgltXFXb7nHqxvENLeNiCQqCbY2Nb7xJz8I2+HHpUx2Am4b
4R+YP+rOhQ/aabebP511eO7hjqTnFYiAfSXhBVXHYEmGcCLuXIm15LAVWvnigmge
jeFb7YCCiF2pLuyecXfEwJ0WKxH8IjcoMWXHGi/LlXmnk2iCh1eRzonAC4K1RqCg
uSAim/eJYt4vNiCC4tBO1Huuuwy0a/de5ja5eqWhzd5SRwoK8xqBThIhnARq+uQG
OiolbJG3oN2EMwCHs5b1bAjPyX+ufqd2mD8PP3LvqLjsKxDCPHHE/ZBiOaX3yYRW
QEPcW/GvN8EOJ7otaeok9I5sJNF5EDhg9akwT47xA2LX1A47Vf5JJ6dWlk0b4uPi
qd8kwsjDGOJQwtQXLQSHpCIxZtYdApt9vDeBKVhIFR64iEo+N0D0utNSWWbTeTbm
y/VsnnCaQpe0MX+zJ/7EgLog8Xk8tfxdlVLPYmfVg4EGeJUHg64RPHaYWMQfx/G+
KIvbUC7p/kU69URkvfQnyWZbPeFpeEK1pY/BZRktnS0puI7yDk23Q9MoItlaPMln
7FeJ7oj+cb9jg4AZBavXshaYslBhbjX49wxibJ9RNz16QditEj6Dl7t+SE+EFXz0
gTueJQNmcP6fpMOF5dAMWu0keHZ9NSE35/TySMMo9uGJw3cgongpcQK9A5Pt6Kmf
YNe3bNW4pz3QdzbXTDFj/+Yp57irrZBSomolIkfT8rwDo9R5xnoUTmfl39b+9VPG
a2RpFSVWoPf/JrBxr8W6AkuMdY08vEjOgRNNaswn9K7ppidWE4xpjF695iyu9Jy5
ocIWE5LtzEQjxn/vhliORVErm4nOT5Et9RLPxEujl2yV0cnIguT1bWSJ328zJUh2
yryB/lpdhgaKBXQjsRDVtrFlJfplxKDlg0AR6F4T7cQ3FNdsk2loQajJC+wK9nOr
xrOiebVG3SoSB96JQ7NfzcyJ5/XoiVBLfbhE2oZLYeCVhzMNLNNmVTMZ7WlF+TZ/
1mKCvqpwpq2Rj0SjlgleLYVbBRKslUWMc+DAiEwAaw1XoAIpwo1SKUBmM2MI/Nqe
/Wt4UOUjXc59LrUITJXichBXi1AbTWxyFZf9U4UOap3zgAX2PRkEApQZ9sOcw7Fs
42ivtUsvQ1qwxM7LywFZDMP7EY0mqM4KvHwd5KSwNfdjMrgO7otXDmlAxYsYuZVW
Qxnh+7j3Y5a4nr4wa4gxsjsNPNSnHrqwEVe85pJFqbeyB6jafmnp+Kja0N91EhMH
RTtuIc+UkxS5MzXV35IQm+XbdmbNXk8NcW7Gq81uzSrjUG2mrGqvQIqfVy9AUgSI
ok5AZFPoDQav8cNYJnuJLF7sCEMxl9a0bzfyR2JWLZ3f9+F5tJPuxtChyp6x1j5C
7PvciKEq0Sj2PlY0aIwV5zqyeFhPbW0ntHhVlDRZmi6vhtu4eKTu7Ehd065UFbjA
i7h0YUkQq1bNde6ZYzkWUiiwh1S6v1B6J45WZwYbPpQqW6x+spr3aaaJpZu7V0B6
UIw6asI4THGpkyj/Btn0CeqfY/EqqX+V1k+mvNGCQ2BhHw71Rqy6uAi0ODHZoS+7
d0sUmGxk7Roj+sbWtDUCoXYFuviBvhwT5qZcdYfT3oEiN0ZZLQIrz2orYTdMp4/V
FASzdHlDciPSDxIjIogUfjBtcKtBJ9hELg6RotOPjvdL3x21+ugbz2vWPP31ecin
dCMByh2OpukYKpV8GVEewRhyebMr7J0sN6IG814vgfYetXOmTNtW5yZF4luPQ5xt
axOp6gIDfMJoyLu496JX80iqefWFeSgQLZkncNMuGQKHhpv7z+G2+/Mn0WBR/OyE
G6Ypa2FTvMhceMIMn8bhgzCcRIUM5li4jSRQ0sRoMQoBl5M2mR+D8weu7xW5qiFe
QNWADGRx/00/wXcDJHxm15fy2BXH/O231043aufGne/OaIoOjY1xrvGGu1HAXIBi
WWJ0qrC/jg7Ic5vGQW1bV73r2QsPFCLZ30MNh1imaD4qFywfWyxD6StSdSakTCnC
+mThQWeFixrXKUzlXslL3w2WF5edIJcsaagUKkRniQHqD95LKWZUPcwCvl0RwzsM
IdWdvxnrtwGLMDrn85wY5sGZOQ63Ps7VvQX5RyWjhPukEdx3ZVP8bPfs7iewFYhZ
JUSFC4A8mrENm+ei4x3ZlZp8tNephRugFpxJEecUR4LcNrwv8fk6ODfCYGhsfm4f
G2LKeW5vRGhG2ztvAkAzojlh4Kjk6UFmdrWLCYbDCX8e7zoJi7Lsjt00Mn8xOB1I
fnNbll85M1V8d1w/wJ41Vh1p60wG5OeLcInIQUVyiX25NjorzKT3UnsBVSQh5PiI
VL3OCJ+hFTxMR16Pxo5znObhDx3DCwrQaYAt+LOfI/PqpuG8y4kUE0kQaGv83a0W
ftspCXY+58b9zHSeb9NdgF7JO1q7m2N1gHe+u485YQexkdM0QlagXJebrFF1c3BK
N1CwlL0EYT08L3Uomgtlpp/SdUoI+yW3ZgDc71b2NiEqgjrbfxrH0DRFwZ1FbQpQ
n0DV94nAJV41mKqDhkI6nb1HZNQbJy6il55y46qXL0G5Y88mAHzuI/vPH4w2/M8b
1rlDALc1qXGYQrh4QyCDAYrmgk20wHjeIpqZ8KJTCMBaI132HJw9vNun67RD26wA
V6MUrsXmM8TcGDiUvwYj2h4NGJgoDE7XyjdLy669WY8gzGlCcpMpVokV4RKw0vI1
oPWrpc5qox+iZReey730ugK1OENo5Hu3PKr3+NvKhZS8zXvsp+dlzGrDL9QNWt/X
CG4CK9xiotsfa2LeXWFemP7v63LU1jYlgU7SWr5j9Sbw5dF0i0cA7Cca1nOSezLX
4kjHMKagt3HLDIFLlzQR5RI2bBEUx2vQKk0t45x4XSgu15tyj2190h4ow7pvAgT1
Iuye6NfmFRhRdxFMfAkJDFNQxrlqQy8lvDelGZ7oTfirN+GQgoL+VVjZ8aDw3mxj
/ciTmf9MBHPrQZSfzt8usqMgEunrfH4MWb3vMoYbVEn2IN0mVr4JZnUlgMeZy21y
KscGY9vhlKfW5iqgbkVcgl1RtLkL+VkQfgkouGDivyTz6xlB2IxqUEMbNVg1o0Ph
jrpvpoImvS8Mn2+4xtCylhV4ABpGB3/yJ2kwMCfXLyOIdVZJYLh62fRnPiXMBXD6
XS5HM6r4kE4yoSRDS0j+RCeQQmWRPiyU8URNE8hlbw0rEhxsY8T4WFkXgvRIqgvm
MOmJydvB1i2vQoGCCiNf1uTTGT446NWm9v3Xt6T5Dk9L7kW6uvrp0o6ms0s8gKQd
4uHRDmKmvBHj+2tnxlNQcn1pT4SFPur1gO4sq+h7i5bHS5V4/RFHZtfe9usLE4rK
jXLBAqdtL/sbe38rhR/g+9Bhbm9SS5WH++YhA+V9lS13ZTIiSEHxCi4/3obx8XfD
n3kLocq0g6oqKn392D3H00BheJfGcfqKy1JKqLHhOnPjCcBHoP10SdbEx/y0q52n
tVjfomQvo/19BnbtDdFH26ikQQ3soG++LtsUKPQfjlxq+wTlTPNk8do85uoiDfVM
MtQI4RzQWqmJI2XqIm7SLMSkq/cEfi3Q8SO3uVGv1MDFgoiaGK22jeb5SLwnqGZT
aKUkpmhuxv2E8ccsUojkVV9SKCxmWWx6qvNzpgsUqDGR73Wfnx8VxG4/i1TIw0kn
9vkuBQ6wIGaaEfAY4HNcc1xZJLfjLyclYce9bDxGy6AaOr9PPeZPLhFuMxQ1I350
Mh9jDQilNvYFptXkha9LcHhnXzI+kmQvkfECEqpM1N1cIOOBIZ06JnczPoUHQKGQ
Cgqg006ZT0qYLTqwT1mERFC3ieRFkY3OxRCuWk0q4LnTxsMXl5AvAUfof6daJYIr
yMB4AD1+NDkZHdmTKTPurmtv3+XdVos0nw6OI7BIEt5rFxj7mPolMkGbobANmDYW
JfUAdttCnRaPzADDpJ6216OuTyZlaik1oVAHnAXqB/OZVABVdb7EkjEf/YJ3BSty
m533P0Xtt4l00gcKkSnpMvT+ZrSFj4tJoSXY7E9b/64A2EU+nR4esJC2XEIxpzf0
OYeC+lZXL5QeWUq02QktCnp3Qq5H5umHY/2hgfmR53KFZewcBSXComqk2L1f4MBY
xe1jUHF1czFN3VPdCz5tFQ1fv99FpQ5OoioeOCtxfodnegSk4HiOR2tCil194Uzd
gt0Qr2Xs1o+u8HZYU92n8GHcXhYPIkOBJHlhuSrVWjrb7R3a7puOfFBtTB6lz40Q
orF8CDWAOAOxGq+RqfBFXpbLFNKwTgIOG32/26uDmdsteUr5J8diN6yYPgnWC/Tq
GqFMCynV5El6G9Gh3+rBlUyCqa4H415RMwAouHqVOdBG5SE4jbkNN14HS65qbC9Y
C9xCpTsQusLInkGfSov28r4LrmYU/ZpuK4jOZDdqbkzz8Zb/mZKSgmHuROCdZv3/
KNLtuMAO2/uFT0jB3BdI0Rj8F1NJgsjHNo9EUi/qsOTysd9SuQaV+9kQio6frH/h
UIN0tn8u6Mni++14R+sd/N034MDOqE/zQp3K6b0YIwsLmaF0uY0omRMAJnjnBBTT
Bb7AAn488urIH1vyAtCW5ntLkdN14W4Mo3FHTAUUzyBuQAYrqrlBHCzzRKhzb0P8
rRy6WK6UQR61C0KdT39Av99N8D71BGFbL4OwEvlwnnyUeKMg+GcGQqw7ZYmXEiX9
YU5KrDskOJz7OpO6DnArhfZ1ioML6f4Ht+La44sk/GYUM7ml99UcYDvBnOvB53w6
PfSFKiyCnN8XID60YAzJlNQq6CqWmlz6jBTjoF1umj7HyTJfb+rxMnY29aS8mwvp
n3vnPqPCpGzI3VR+J6p87U6rTSwc2QV6n1Bqo9N9ZP07aIWT0f30V0swX6wFLTpe
J04oD3A4vlC7mjbMLiTVxD2USaevEUXmkyG2wQrJUlnvaOWTiQylWjPM6QpTcwTK
yeyjdKB70k5RxmBxSmDwkwSfbrh8fK4w90Az177qF128j9uEsoHt4B0ZaHaVQz2h
AQLe61AVMPPdlCF4XFSpbOkAe1725mJe7h97WcIKk+OTbKwMCF1pFXdIdgIeZjV9
PHf0723B1iFIfPgvG/vTCL2MAHdDMRGsXjFXT3xR7OB9F9+mBGqPVWaA6ZGtoCBh
uD5i1XQAo28+vA/pnDsIlEIweXCV+8XRA5ptkd+TO/MD7an9i8XaL3dsZgq9vCBn
kbR0cy6betvbCX1D2zGrYx5a0t5oMJc2A893cpNpRO2CRLmtsOO1HC5t9ps9YZM9
XUqBb76tS/wrWeJlV7D3j9JQB2Mn9/aRrOAARMl8mVtAZCL/1lADugyTGq5VgxNJ
7TKL0o82IhTmpm/e0oHT2QFp9wldGUioRmGCdEAjxW6dxxGPZE2CX3hT6ojKlrjS
FZGQDHIeACVKEumkA7QmfaSpNt39KWL7DmLdGljSxJtGDW6GhdgG0bS8biBDzKFB
m/n5MwLV9WJNH1B08St979WRO5xooxAaX1W8EIUf8Aw/MAitUJmaXhdpP8OJqDew
+Swa687mzfCqN9rxShV6vcFL5bwtEeNc2cLE7ZxIEWsOdiTNHtBwLWHUkho8ytnh
AJE5819sELszib1C4NgT3Ij6NXGhKBFoyCJitb8tw+ARG9wTt0CgXJVK0+/K5tH0
5NWHtAkn+c3LUZriVPOXNEw6v+tIcAzanKHDOft2XF2laYalcZILjKt4xfWSF4ow
Vh1Uzk34Hc8KawiX7tPCuhU78ooBhqVBme0+MQ2U0LdsSItNmxIGW5A8v78HgYcE
ZMm62LHr7RTpeG3ceDPq8C4Wu5pM6cLDGUFkzvj8nECD/brAEW8y1N6yF2mxjQ8a
8UQbLXnYYaHt9WntSQU6wN0/fef7t/ROQXO2+KzbIQ37tPPYdHSArBlvdl8jOpSN
PyXteJH6iZUJjiYQ/hrrR5zbMgW3vuIxr7F5feHD8AfHQZx2kBPsnKvhkCtfJTuH
lk5p1V4D0vlg53Fc8YUmDB4DQ9Q6iMNqdps9DTYLcsHd8kaou1qBdA+G5beGqfQI
TPwYSW8ZkvNpe/iuYLXWSOCfxguTZfUbbq8x/Mc5iVLAQDFg+/a6/pvtkcRq4CbE
cytuzYfCYOof/9mOdRxnwatIDCeWH+DBZ7WeCVWppeAndEXj+k/9IDb/K1YPQEU/
EzcSnb+Z5GgYwgVURs4Xk83A5dpFXSIJ9TkA1eGNML7XCNMwA7KO/Pc2a63FcATC
KjosuvZQovBK3e8WTPbwnxWqbaHuXDgsTu6CGYeEokrBrJ+qyRmK9LjbWS055H1L
jMAQBj+kylez1lUUwFwida6PZ10EOHQex6IFp+z/aksD9Gm5ycty2qiBUF0Cmvp+
Dp/0Y+meBUvU+BSdBnr+3OnN+A/mrxwja39KMVTKdBNLpvRlCd4hgif6oxlvMbiZ
3/kpFdn2JLkoXM8aqNp/qs97aIgOFgCk6XeVLzBpYYAK13WpSGwIJ0W7uAKCEBun
BYd5ratgOaolGBfX/dKCJDbH3/0IYkSD3HM+AB5x8Xr3XB8QIp38Y01zia6XfRD1
nYb88ihJWHQuq4KzyZhGA/78Y802BhaAd1ZeD4cBUZ166HwLZ+wKinIEOYKkZcSk
B7kHhU9Z0UOhFWwQLdAkMawfNU2xFttwNZOBUOdnmFQLdMy+yUSeXTcLgyLPO+bi
/LlJ4Ge5Ik+cWsN9g9nU9Eiiwj+YDIom3IJt/Wcs1HBLpac9mTLiBMJG+DvvUgv9
f86dWqHO4kA7rmqJj2xVclrpsk7WkT5txfrU5yJSaSgZIZHwb9Hvaq2beESYFa5k
Y21hb3ickXdInZu6ZqYiSnjhRdPPCf2bsgPTUG+mpF0EaxofRGndH+PULCWYA5ND
xPDSrL/trfSgayft4LPeeMv6j4bQyxKajgSfaMElWQ6Y8E3eJP/0nzfMSih0v6hE
Ih9laCPOgNtaD2TZJzB8CkYUBOZR42iMQ1ZkA46Bz76fG8HbXmwZfuknbN8JKyY5
31mLjIINbiKEEC07d4sF+6Fc6wZoYoM0JTD/xE1i0uqIdhvksEf5y5mbA0kGnlU9
1h/2iKCkuVUWErHLQniJDt5Lyg7DTSoUJX+cz2VuaG1pUKXegr5gWEbsKbqqLLuo
C/ozLCwk7kbyxnBNyH5lJygqPx1HaOrr8ogqRK54XjYYpA5MiHKLPeMMtbPA/neo
B3w3uddjMOzwvCBtVLjTewz3kKTe3b4ZHQiAT9yqrn+lIAe0hJHkkyXDTMdNRhpV
5hFJOupzqb5ogPTDEkAx6CcA0IMINSOhTcYKuZ2Hpfj7i5uHn4c0bS+3d1tCnCkl
KBovV+v22kOnhdRiwGI+raXCsXOYjTNVlvMSWV+OwE+VHJY9BVVMnyKFLrTrKkTd
4Jlq33do/FTiMrfV4HQRksBQmcDOuXqi5WwoD87211N4IgPE7rjKlk+EEBi6Om4F
BudjukIC4ybHggTczLVCYqEr3HOmXbDAm25U+wp22vdonmObWk7/GXVzIF/3phpG
ddbeec0FC7pvVXiEpwapZB/erD6cpeGB6S06mbnvBjakfdCnpKp6DhhIcRbDVhv8
Dn09JC8lNepwAAwNnLNELoDC9YtU3SgsfaLSLxZYrDU4cBQ4ebRPXTJl652F8yL3
TVhhaz4kidLJ2v4aeAaJBkpKNrezuJyJIEwJSsejPC8tsAgp9jR0oIeSsCKKNlfb
RKOmThFOfcZFAgakLE7Dhg/7XoHpOp7e5YI3T5TfTNvoMI0t4XfpGQBdy6uoa5Q3
LW9rsu9cpVtP2ue02FaWgwA4tGHzi5TIZXXsEU1yUIX3pvmsaXMww3miRVKAmsXp
mZpTNNQQd1bcDvSMAFx9Tf4sxalGaWX1a4RCcbkDBCKbNGfsf/wC7ak6Lf74qiq9
HijRjjx8ZQWVm4Vup1WEl0s4kIFt2c0FQd+YWlogoxKfkeSu7VOKqRmsF8+PjM/+
9CVbv8mq6m1XbL/JuRBSNYAIjJ+9J0ARouJ2e/hv7vV0yi8HSW4sLiBMG9bNc3Eq
X2jIp4+Xcjc++XnXwsV/883+Z2nArh0hU+eNCdI9S5aEZVfHkrvysDBvE2q7j09A
3mK37AVIZ7weNl+mzGCkAiinJBbHvOyLSM7JHQ/ZecMR0GCAUGj8Sb87R2tlOE2c
jhlYm9niZ133+pljfMbtOBjOS2I+njklqhg0HEnw2O9cjROtJtETFTaRsTEhR3mx
HTVfu8aRlxkNfCTHxTzmP2Idoh1rlZ+vCxdRMA6z1PPWHnqwTHTkw/TRY1ggvwt2
V67he1a4iSJEBd8M1hf0z986UjlVktrBMNCGXgz9V/IKjfQ8fhAr1Ja1JQ/aVhbg
imhlC7MdDKH8QbouIO0/4VFFBXpKbJiACT1PtB+tQeFn/qrz57O+oKzK8fBgtxUo
R3UG9/LkqEVIy0u1jYM+GJ13hnb7vkAxWAHyCxZr/DTnKT52wwqazuJr+yRvMW/M
cf8WlECYLE3TOr80f57DpaU6Y7uUpEtcJrvuCLcWBjqwnWowTEYGm72k5k1WYqGQ
r8PDgkOCYXEGXB4o2POmDuEp1FMxWsdpBe4z0tZFoKksI+fDyIjHGN8kbliZJlm1
dGgW/deSx5ftjWMZ656/hFpQzL4QVZ9/7m/jdprL5mKTrnZRd/Eg91OaC4sa0E0Z
eS453uElEzZBPClMcsOGfEG1H4g5yxHc2hg3SPTx4G3UIygpJ9lG85J9xNcapg+L
wCGMLKOIt1wAmRGhaYJFVxEV9klMmJsWxY70MdchDmH51xxyRTI5iGnk5EB/7Xd/
WC9x6lfMb8lLM3vB/V+ku+rU1+LKzheQfrQngbCaWpCIskkLsLUpx66VV3cYClcT
n3g7n1RnnexP7ZaHTp55QFFAdh/Jg11Wioqnq4G8zYPUfwU5cl1E0YK22SwxEjDE
mxhrcl+1jA6BVU5nERnBKRU4WNhSu/XvxoRgBQElwgPRk5mwdnSTTapgJ8uIZh9U
aJ4gZSqXpLG7d6rNePthTvw63YhhSGyhuLndj9qX/8a2yUW8KHEGf+Xlyjmq1b+7
2CM2Yrnnr0pNXx/z4AB185PpJ8yNWylyCQETyTy9+TQksROeo+ALsRTBtsgJ5t+n
VOJz+bCkKs4tmqUu3vjMmoOl87rufiXMu04dyAhPaYhLZqG5gNJcSLJ6rjO5aeYv
5s/oLvHcjisyBNgQ507HSQFhn9/VcaYUB1r/DuN9Ea336rZFdL1OrWhM4ugUmksj
D2W2aethQ+fDxrtgJ+43kMFAX/Poxp6jOJd7I3oGQIwX6c4z4WHAGI04ebVFAO96
qVbhc27I49QQHcU7Fs0cJQzlqNBx9myod9uKuKkkYOCSUaV9mSQHSdg/CNnsyxit
jpVDIp0YQ9U022zyydKgsOj0oqF78oiTNueHw/JLvGOsLuqGC2Hyt8VIAbhYAvML
CzvsX5WulzWbsXDE8AjgH4eYG4P9kHXyDjleUZIFaj2b1vAzM8deUEhOefCA/Ke+
iWCoRZs/h15ILzmUpsQEYmVOYxxqzXT3NUZziFTyjWxEn6aUOIGXVjDbHGH6oWHb
Bv7a2qKkgcehA9NpJWdCe9csCWyfgAfVg19IJrLCb4KqMaFXmMSh1NwGV5O/KPLw
PMAUcY72NzDeqxwBogY+2yWLCdSWqg9vj4JjuyyHIkzzpJWmPZ9SHHEV/aIM3iMq
zkTu+xIEdyE3a65j1MhAWUPxK5idPa5FywDAgEVocEDKgZFLFRcSJjjUqio5hMof
/nLVSCeviEYuQAETuQoCMT8MDU2OULeRWW0rpecK3dObhbhegifI3ul+7lrsm8Hq
bR70jE2Y0Fc+EmSnHwv3oI48uAkqWOAw1D97+UWBbHSDJdU885MgTuDh7ZWmQY62
UDckZLvsWc3oT9q8IPmrN9Q/qtJm6j30jMI5QJ/JCCeFhObivOFarGXcMvzKRx1t
0dlMQHTuXn5lgtsS/9cLjRKA1E1f/ChkzsNO+ubxoDt3VRnaMfBKPmU/x1DPxkwk
DkC3WhYp8kHJmSiLjRpEUwgTzkGhDvYIlvSHLePiNN3S5Re1u2fRUUm8ZyVyhSuh
2U6MghmyB+NrgekyGt+sK/Kp/+E+aG6kQun9/wkAUuv0/XFQ/BU1dNjdWsqo4Zv2
t+l4tl5mcWXjKwZ4OKB2xEYq9sRa3Pra5Cl74TWYGz191S8kTSqmVR/U5Lq/xjbT
I2jkyX119EFbhrCR2bllC9NmKfXWH42PoZPDQnbLQd9ni4sHZlrZ8Ms533YcaDp8
z6pAJ9r8BoNpGbtHGoTr5LjniNO/CZSgS4Zs1HniXUV2V/v5pWP5kIDftlKZTcEU
INxt8y2BGEpzo2HonzbiJW4xXV1vETv0t58EN6ypRHqIy4e5GRINYuvWgL8h+v13
ML3OKi0PKHg9gCt0NZinMdTIdNBE0VkW0whTOnE8oxwD9tzURvXqM6huOwbc34g1
+DceTuns/Ztlc8i69zAY+XlYyql+pKvGzjPMMKY1E/KGemZjEPH9+iISS7d6ONt/
XnUO83+kbfMCiAxC0tU88aR+KGVLl+IA6dZrwsvpRujgEgjLp3CdIlW39xNCTA+4
e2MXNDmfthhEAijzegse3T8r8xe01Q1i6DY3wPMmI7q8CFXX28V9X2zEv0HLYwYF
03mmJoicPN7/q2TgSHc+kqg3Ny5es6r7Py7PenO46GMAOEIvMAZnxNoLBuSREJla
pbboR3TZXJDWT6QiBvv4RQ7nK6Rs3awgZrIcZCchLP3NY4vCJ/ExIrvBghBwjCgq
4QOctAxHxoTVvFaO5popaddU67uiNGCJXtRkasUvR66ob7scQr1M8ZyUqEpi9r9H
m8DJTK8NKgUPA/YRPH+5YTLUMSPMphgx/WtuOJ+L70vn2/9Tq4uU7GZ5WU/g0L6/
1oI5PNCWzxcXyyLukeHqwWoCmo/9Cp7dU7U+U7M/6DAwjvjZNdKQwhY7sJDX3JX4
W/rRY63RaftlBeabEaTz/lRkyx2UKLc3iTl7xWCvFrmQkRj9c8szMphztvb27sGV
CxZoMDdCIV8GBdiAoTIHA1/XM7BuqsOCYFbRbuoMGTgkc8OzyPfpkj01kCei7wx0
2aG3eYPEtc89v+w9u9LsAwIPTcKNBoTpGbX3xVnfij4enLHTg2njAmgguHFQNpQx
FqlUVvxjCtyOAwnbCZMOGKKzcSKmUrdjnaLZ0F0m36nOXQ0S9gbzXMIZJJsWcl91
QZQQP2jBFYJ4eAvIALLR36WZPMmGoYRvCY5c0+cmDOCls2uYPwhuyMtHNMdau22P
lt43lWJ0fZJ1CObeRekxukV8zQDaJYEM1jMuL6zmDC1/8Q9cL+IFq5/F1Vv91al0
wFKdySX+L8cS857cG2Hy6YJfjlxfmzMcXEOG5BbOWud8jnrQlPD2xQXWcY4rFg3E
G8xTERg7mJ8nyd04nXdB/afkkC2hDPlEZf6mmbyyDL6J8yqapIwyLtd93cxPr5J2
faTljwIJRqtAAcQ2VkqlhW4YsWAlXoRcLzebn+qUEVFqXgAlFCl7+Hr3kYFn4mzd
XcpxfQN1QFgYAHs2V2GtmU0MOcUKvz7vp+/FZYraPNCVl+iQX/PLkIf59akPta0L
wMMs4LJ8yxCaOxd22Az9t3nhOuc3fpMqPF3EUKZbPrhuWHxRPNR+HK9ZSuJmTYs3
D3e7LsUPxCl2fXKQTfhEOUnvvBEFEqVL5SCjOs3pd430HmAGic/xk5Uql8X9sFyB
FJT5IRvOWE/2Nei85iRoTFSqYmcF7Kp+ZwVtDA2OdJUK8KkznCxk2rXzqF6y0tV5
HWLIIgEJR/a+O/+zRN4VXSOEFY9uRQZFl3Qd+ahXHNwRx/Jr6XyMI9NdWOw8b18e
j0SKix91VIKINoB5qe68+7oz5TV1hThDuIOVlQWkHPAKX4gd4aIUGFP6JMb2JIm1
fyqa8raAx8bpOKBvozcOlL5JbY5T7Up7ZanN1s7hSdmHT0ktdJkyGYNNzejD3QjW
MyfDxRVAmnclktlyYfD/Fo7R8PuXagRFtQlkE7fveNTYRcIsC5rBZrFjkmJ/LxMD
V/VAub/5/S/oGFNsAvoxk+DZYpIUylOwufSExalq+q4nPrtyULtGtOcheYKnKqc+
iInCDYjmrXClB1ReJ0lMfFngta3ZiMeAkuDmVC3ohdcqHAgkQWqyjUNUn7MIRNQE
dRXvoxAdwoyEbLW7vZAL1NZ22VhzshAUAMvO+i6VcS9lxegt7Hb0k8dK3CEY73be
bSoOch3iwCX+glwe1IeqOIym+3hvfhNyS+nQyyb37Yrba7ClAw7Y1KJqXSJ2PUe8
bd871l/hZ96/X60aXANplxmrfWu9KLEFqV94gP7gvFumxd4bPkdx03MaTn4/O7kU
5Pc8H+eXQUJs4AkRFt9UwJw1CLUCUENG7bwZdEpMCqc5+aL+0XokbldniiGS/IQE
KxqjdzxAxVOTJcHDZK+Cfhu3Iux/cBWgkedascS42wOcLFtfeT/piwtylXxDCn/G
OCrt3mChwiKm6sOrcYZm6F85AO88GbrxrEEt3ungSmTeRXD5JSgB9ZWfnjYNcRzk
MBHuAINOmhBDUCKo1RVYNYh0h6SEVWGl/keU7Ovi60NJBqWU4ytCL5B3qoc+KilA
QU5D5+b3wa/kJP5QJbk/AmJ+n14Oi7wWy/p/UA5WbGwdDxjHPpLdKSdAP4bKlZf+
rKV7d2ajOQpHUdyf7nB5dVnxaBMdJSDFeTnI3ikMYOTYvA3lX3yW2acYMjLEMQ6r
wTxz7yCHdTWt1kx6wl4QQ/Aeor5GGQ5PH4InRIcVHejNrxNWKGewqdqiTPvgxP3P
3YarP6cHCMqIVnYyGc+iIrkP+Zehbcoqy5tyNEXM6UGEBqbz4SQ8oTrOYHzvvyhm
dBLd7tn5OS2Ri38r0Hh4oxeMnXG+4cd8pSmJa6kXo+p1KmnZUSqc4hGmWd9M5n6H
hhv7MTPc5Pm5ePJmMTOpOgO8w79xMFAmOa95mr1aBQB6diQgYWV7jAYbMakgT1bS
YP6+V28G/Iibwm0TeT6f0o/59IMXMDwZFQOEt37DGw1nPigPN1BPF1xgOt+rp459
LHFxPMUoasc8R/fxOy146gm3OU9T7jCMH4haAZQudwKfyFg41/u8KTul5f/A/RaK
SUYZ1qn7SZCjrdUe2F5HDF3UtpCJkvJp6RysFoWZ9myihVKS3XVsE8vSRzhwRnGg
GXVbzEAOi9XHJzTWY499STI4NdW/9DlzOW1WoXPV/aNxdwQSYvhUCTEVb9AVqS0b
/uaCa1cU301ccx2GO4K68ftOR5NXfbT2tivOApCAFkMqc8HPtKQVqg2VnbLQzFAU
eQ7ownJk9Nn8q0e4bjSuGC66M6nknrTJC4qm9ML9OLTSQClJNp/Fj2OlVRyh2CHz
IaG+Y5lt8lnj6Z9NPvFbv90m7x20C7Az59oKfxcJrzYzAoVs4shnxn2hw5jtao+U
bP8X68GJZ+0CoAhNxOpfyyKfHT/NR8jxM/dXfsh/89D9Gv99wCmoMCFfNCBVUxYc
e6hlS8OoTlS2JvjxFZ7T0W+jBPvGP6rXJlUGWY1HvkaBcIohNWIafD+noyoR2bGV
K0YohurTU77LqhsyU3JfB1nW1iVR5iXs78fCYTcAOAwpc/s+Et7ULCHMdyjxMsWy
/MME8INWM0Z82XVpjpoZEPMmbuE1gh6YP5XeZOdfhAzqkfdLoO6Fo4OtDXsOqaxS
KB5miBP/ruTsFKJqE/zp9SYR2gJkZ1GGyvfTFdhADmb7XqQ1Qle9tQcLUSWX14FL
IvuAnB3MylQ0C5H+otMsl3mREFtk/Q7Ia2BXoz0d+887GyPAY3BjOU2fb59WFbVN
CCIIIPdiZi2wdeLdBJhNaQp7n8LiB1+X01jsCAwo2vtzNfH2MFb2LxG9pohH0gdm
44k/1pYVomvtLAG+RD3/YXaP35QUHmkcDJZggZDt4v2R2mh6oB78v7eBDMGdkgwi
MV4N5ls9LbAbXnxRK3lJMX+//yZT7qVfV8uYxzHWveKojAa4zMqZQAha06snnMhl
blwn/5tO5PmNBWMtm9fLDPY0XXd1THjHtV5UIsShufAqJyusU5ubkCG+BBd0VheA
ZC0IwKw/It3P522oqHiy1LhF56WPJTBDzd4pOHb3G+YYTpInzwGrh/Ncx5F30UhZ
HP2189kfDo7nVcTS7s6hlM99rUy9gxaN/azIRRMvHhdtvatVl+LOgcFHXgK+Pei1
YLmqt/fDX30M2x57bKp4TycEdkoq3xmdK3VhiIfDras0jQPn8Lf4mC39/rTCtM8K
nB4I22gYydCsE1AZQQ43t4wEurry8ODdn7/n/i48+kEaJmN8KzzToVviGZBs6aCE
KLeIgSEAPoRLIivFxBsUL0eAtTqVTTT/o9JXmlaxmfgJmiXpDMsPZWVTOBdhu0aV
Q/pd7gKoZLEoYW0awQ0TJloz/yXopljdPpyUKZN62txtbwkhNnTSkYxPlJMdTMMf
VD4MJ84ayPTb/h6cHEYIf/aKRKroz+WCON67dTDHdxJ71O4l9tMbAjrkmUm3vgem
8LKuFGAVithk7o1dMhkm23AprlsMgQ/+0HikUNLD28w2LcW2HWK6Pni+toHzNWF+
6evAatV/o3BXZqHQ5a/zZvcYCowgDhgvrK6XDpyP2HJ4+MpgtObdNK44ZsksyRQE
zNNkkpEZVVbh59cUNeMPOc5AzPZCS61xzsRItyr34hi/2oB+PbdFBEfYSHcHYTal
cBxO9AN+xXctdgcKXSOISDVrbUnykL+OeD0iG37WJahQhOCA5Ev14PSTRykufh9D
FJCdQlRPbCWC1ba+eJeSBfGx3tf2UI0DdA2FNfGsAVadqzCyBFQqfySUdJA4dlTk
s1Mc8dBJxR6fZCjhBdDiX85uqgbiofoRTfI6Yp08mtmh5k5DKRmIIIh0c9K7Sdz+
qUjkZsFEvG7gtnAxWJ+O9Q3BbfxdPB+tY1V18dP2wYbIisfDUPR7Djvn7rTeDux9
D1kW2DqA9a76nAUK+NU49YjwD2knwo4cvmW7AvCI4PJzNrpOshcZXpgLd6Hdco0m
NUtmqygymxmt5Fn1le6z1YM4WidknOzrMuhGJ6zLrcmcsgzfXFt+SFSd6GJOGggM
PD6Qx27Y7C8+Xw0PBPiW4EIOYBplYhZibiGX9pzP8Zdf5ynYm86HDifrwfa2eNkO
hjRBAmwvlDipGQF22yM0TdDZFCFQ36jT05MtpHk4/JtV+H95uik7Zg3OTRFLkjK1
n1h4G23w5Ssch6VNvqQFeKaIy26ZsDS5VDSfv0B/3qZBW9MFx3WNykfTUAF0Oa1W
gOZUAUrT46B5bV3vGRSSWkFuJFCtpPywXeqIUvtrPiuM7vSvlfsbC6rIyPPi4bwz
axFUvS0zn0R7I7aCyao9pCxoeM20f1FoXygGm8fZQwj3pOzQ6Ey10F8VzkVeXb6r
jnpmu9SPl3BzGrt9O+poNMzLXW1r1G8lLp2ZAEjTPwUvqF16YXvjxTAMUQTwCqlC
bQNUYLtS6rrv/W7FipUM6WKLxksPFflct71c9tLgtbzqgFQupqVW8pMtjqHFjmF5
i9juo6sBTbcb32jW1R3rnVt+W43bneHgdkLap3zBIpPAuSUGlH28dVCtRGpZzyYN
8MhVf2FVnEI8AYMgkTpuradw4XrGwuVQca2OsvsQQC+okLsl5iT3xgR8/NiRkseN
6y7TXGkVQDa/MW/tjJrILIBG9Nfv3BcP1FO4CK5HTGTyC9Qe41c+Xi4rKJ2Z8doG
/zYfOipxtM0DQJb2Of4T7x6HCNYMYXbzWGfCnBgH4xVnYKruAdsMGzCdXXmfhhNm
coVzNZ34RE42/lGDLmKqK8SufstX78SHljdgtusr6lXImBdkxAlw8IfRPSJolzAF
fr2HhIV2on1+EkZ8kq13AG+fwYoSyGh+hrX+MvC07FfQzIFFG/ecym+1QzIPTrC6
dj7abIFhHfzc6pZOY7gh3tobQjPh/QFWbG2M8MV9oH7GkwIcEevxjQFoTHsqqYVV
o4hL1o8rS8xsxKftLjIqPEJzu5X/bl1ANEDAezMgrRInM3JxnGDcnS8vfM5VHqsl
q48Poab7qBL3Z6TuRxVBOlOlePKwTyCbMtobpqJ2/cTHY368RIUT53zM+esp6zY6
tSIF+TyvTxowflVK+bXkSl5IsX8mCjm68BPUjIMBNjvjJ/HP1dCHEjqe9XS+P/FN
2K5BcKz6mpvvAf7DsNwThnVyW5w75THxFfk0FJ4hvyacqsv/ao8ZeuAwdYCohult
Ac+eVWrPmfLWkMrWwxBJQtyoKaoNun5vKNE6TTVeNGb7VOEgHZXpI2FrUIvVTbWW
Eo5vcMBPnrOptrLX6b6PlNsD3+76F4PtywEKDSuTy9gdP7n1VbJe5MDR4GdDPZsc
Zpy+loPtabbc/DI3J1O1KJMIJoUi8yGDCrPA2I5s/xfWH3RWR3/tYcTRRdGDIh64
LtH9CFXZeAUMCsFuut0nyQz3fw3FDWBVlB/jWHT5/FBRfJtRyaBi1iUvJF7iV0lQ
MOLJ4k89v7rvDxRI4opdmJTuGXBxFjm8JIA74j/Vskz9TapN6x9GPwP4kZLhjyZl
DRLAv84obZR0tGa5VecZydjiLo95FEOumMBJX70+MJCPI4SKARFqFrnm7Pr321eF
c/jxCzyTXzerwJIJqR5bw/OuZrFP94MTYxiHoZ8iyKcjB6LxarHGpZol6QklWnky
OtJ+rVvoNNbOydw9QK61FtFhUP7F+TDNjJmQNAnYpZboiRhoSCG6ltiFsW6CYVJh
bi2AQpfd3IBUFPBqxuDH1SKdv1VsPY8BLCNRgsWJYZXCWTnCB43R0TS1ZodxU+LG
sRbQFxTbuy9/sgpx2L5r73GtYShJB9whm4LsvVifR6C5YWukEuNAwkQ/EY193Av6
T+Nc7FRD8nYBZBgWLqsK4JR/JhpT/OaJjQRAkXcsaQXsnGko46Ju57ApVCTcvYze
0KXKaBJSLn3I7pBWCMgo8Ugqhlh5OlQKhW2+UvB4z1tekgx0vfFX/MxwJttkWcVq
D3QJFFH0PGixeOhEDgAdGReNNnirM4YQk85GgtkffmfNcxKMBREbWu4ztMafaGXB
JsqMVjJI2Hw/Hw+caEnN0oJq0MW3a0gI+k4bhVdLwohC1TnMG1eNk+khNIlyMzHX
mfX6neY9VxCOwqa6kMaea4VreXJ8ERx2K7FlwQpKtc4lze0TJ2iodo80Mz5unuba
w0ZWO1Arz0WxwJjh6ClgKRJEUHgi99N0XxNICoDm+y6V/q8+/51tnnug33lQMmWJ
WdTO5f4F9DrVMMkdByoMy4ZwszvJzgNUHCYLgtkl3LSmHHkHI4GfYqeMgx/VIs5r
905b+tpNVA1/1E43mnVJAn+uhSUw883OvlgMLrPGSMVgUHBXw1MPyarpG6DwfoBb
RYQFNGFvR2As7zaWTUWBp+dkvm7h01/BF3HkzddIzdHz1wkgC8f+sWLGqKIdhFUu
Qx3wjUVq+IzQAUjCBelFlMyZoOypZSuC12NgxR1fAYFjAt8WqBfOPbnLpzsWET1H
3TXWzmcEKKIDZLkasMG64uR/Y9TiPxX1N5XLnnwOXM/PLDPToSgmJaBqsWmkjiyu
sjApKIZPBkGnxS/oENHZSVE0cfNdpU1NllV5D+s82dF8rWVRiYi6nvN/AXgFl6Ak
0+sHg+H9iTW++D7PiRI4eaqRJL/WegO62YNtpFrnc9Xxji6NO5gc31dQHmpxkchx
MG8DU0VCvPY7H38h3KN64EI9Hc35lZURjns18E92AL7o0RoJ1sGXjvw1g4ewK71l
/jeEgWjLg8dFzAfiqZRJIk/qTDNWFazpMhP288Win/m7ni70sPdpi7e4gTgcBppx
5A2qdHzIEB3b99e6lyjLdpagn7rlod7fiFfWUNzmicweauKsyPkGOYTn0Y6h/I+H
qVmMaxHMqvVLZ6IYb1Nzoj0oEUukwjggeJ0zDEayyuYYpFJ3LcPXweqacp+XKlrT
GbzbGH6FexJvbsMsUlDw1kwXAldb5qPcJazgThk+H6yNSzHmcuAf4mPWvGDx7hxF
LsqSlb86EwODGOjVxaVNepCHBbhSRvWv5HAqfUGsvoLoOi1sFTv24enAsmC3WQom
CZkZfl7qcZ7haUkaLor9LiahIo49xmpxyTsfFGBIMvpm3qrf9wzFXoW1nmTVhhEh
5Xe3T/5VuVYQzPPh9cyhwNG0WE+krjO7ACEBepyuToYjwkouV/Mdmfru5ak1cvlD
V0M3xe6qrRzgAu7SeF0iaXwX0sYJjxruQMJNmwYLyNF7/KgdqbooYnmcQA3WbWp/
SHrKxcz/NACmU6WDmlBcUQbhydNpS8uCaVqVjmCx/RHMucLboPMHS1mEb8fRefpZ
8sycDmN/wclKnhVY7Mwq+UOQrZKA8e9SJ5XYwAlX1gGh1ww2Z3AZnmlzDKxEhw1k
B1dptRssF+qJvHVGpDwlYx7GROwb3KIlHfzD4Zn8zsCxhAiGF3FdY8El2UwFZb3I
vsSeofhCuvOazYon9NkTZH48/eXhKS4buiQLVP2VZAuSOa6i7nT60UpTSyJDlk3c
cKZSL13yfSGHnMJDVKHnVMa5TNF11CnJ5TNOtfDR0AdgHhHmdpE3bYo4JB1eS4ZG
2USQwed6iwXmizNLdeMlv8R/gAGY6X3zIL+l6w7WE2+DTBIk2C8pJM2kIoaSTg0O
1ZR/PPfGafbtbBM3lk/ds7pOnf80ptbh9eGLeYi/PbNTGe8h9rs45EeHTNC4EOqz
SxyZAaWzTkseFF004M0C8TO8s13Y1mqY2vYpu/5hlH0GzFyhGAx8UByxFB8qAkKS
8HOzLfu2NbfCNw5jrghLmHpgTTVyTD5Ca8RgZbQepx0+O9kWZKdk9BYzKZvVcrQf
ekYg5lEy/NA+m3nQ8UmqCvK9YvToplroKrXmyyXOGaZpHoNoN+wRC3iQo3v2Yg7h
0VP6Ziel6rrc+rOfHqwLK5WMxtjONzflVdgEwNgG3QH/6CHh+lkrAqUJ3nhNACEs
hRBGDwPCn5M0RPMRl8s+V4IJmqLU1or6e26+IVOYb2xxoejnnRQX9Z80m84K+Azx
rMcDmUS/tSwEhS6F5eOogzwv3bxLkKnBsUUWxmefkmQMLR17o5tliEZ0vCMul4/1
RfamICWR6TbQyBIB69lHI8s6gvMrjYwiotJyuILwki0mqxYd+EMSGu4KoQ15n6L3
Mmu8PaPTXLcaIEDodAzpMtB65p2zdQiol0pT8Me2sDo6FR1LKHZMEWflNzkOhK17
XeNhloJmdh1+kwSTA3I2ioiew8IGavLvv+T6VtAsa6raDz69dDK49fGlCdtDlvqb
VzUeFH5Suf4KHNMF/6y82FTlPlPxPpwRVyOHEGegmtmSJpVHgKyIPIZH7OzGOmrc
YSlVmoc3UgQLDdmIaDYdbdkaNoPVxcaqXvpGPErWvA1sSSSRTBTySo2gTzv83paK
onQQcM8v+2eMUWOXRhqsi/MvP8cnp4RQMrOgBXzFEKfxwcrfBniNAg+WcPs+ahdD
eqqyI6uySLoKvGBBVfNlnS40kDD13M3kGlmHuXya8Pw9mn76N0GoY1Vasmr5w8pP
vBGGcI0+knzL6xb0IPlt/n7sPeEZMXpiK6fk/e4WBzAa/cSvcHzRKZaR+vclwA3/
iiC+EOUj16jdraazvRBNnZEOSJKrbdQ1NrmyKS9z1Rl2NQpWTKFltJV+Da03ALcM
e4WOYd3KT1gNgPS3a2tPIfi4ABKJd2zPzTP+xmzZz4/rBnb5VleiMF8WeFDojvjI
xPhp3Z9ZX7rgJLhg2CDTnHnhtv0S9ihqXO/WruwResObS7GEbXDNHBtVplBQfuaO
e44VVvJtDz8D54EoI3Wdjlyx5KWDCGKgeX6xgM1S+bwwKnpID5X1kafXkvin+qMT
cJ4nth2VZCE0IMHn8SCvjOh47V2nY6RVCXgYbuESuAaBvi//5sz5DStM2tD6feh9
cgu8JQYQ19Jz4pO84KtfCqv61Mbi/xIpspZHxK4dBQPhO3AJhkDdNotgIO2RyYGK
dhztGpgBL9qj1l1P7tYHqcaZNfeZejKxa6ay3nD4O28qoMKlfRco5GO4QA/LC+7W
po1gZalT+Hb8vAiovq3A5vCthkKdp8oBxP/kYZlz7E+g177wk429Mc98dTiC8qdV
hOwdIqTTUFlITxRUWvsVLQU2u6R/TTfQqeTW5dL3GXFCWzXVhjOi6G4kQb5eyT9z
LVdJPmK0ROQxOWDACDTF1TOSdq8mqxaf+kQXVk9d7xTmXA2DTgsd4faYgsIoA6oB
Ch/a8TIdF7j6AcnW4dotpp2MLUTLoX62jwyX2U7sirhf/tt2JrFdvdg1HHfcSX2h
ui8Vpfgd8JFEzsECk305jJburNbXIzWYLcTyJga5fr3gS0KcNR+0F0D7DHGCiKOx
cKP1Mw/b6xRgsyzOQW/HKqjkFxvHTnppkqMX6a9QM4R5sJSnJwG47+ufTh2bjVwt
69FEs2G/FCucVqBVU97DXNQz5PUnZN9eNAvLfO/FIopvSFBW4L+xTB2JcUHx23qe
hlUnMcnAeq185H4wqfR+YgcqrvSdXl0uFzBj4K6yYHamJO+L8kISeBHI0Lv/nXzW
JUrSr5MJQ04VETLyice3QlMjsROfVXUE9maEhKoZQLvWhoPiWYLCn/CvbD3Rpx5H
cLvswynxMeIx74e5KGmW306WalTWhRFjHQrDr/DyuLV4YQcatyOQVjqyvhBhxv+F
AX+tMXGIZn5wPA7CL5EnDjORk5Ael7A/HWTbi+vH2cDYEpJEkQw+oKp4T/DXD/kB
ZFNLFrER8Rd2gbF15uSsNQ8RCqBufZt7aIIj//e0QVNIY18cyog3BxvhrUiG9TqG
LEaxpnMWb9JIH2PYDJsh8/nyN4AXkiI3PovfBo1JKjrTHKSMgCqbse6NMgxqyBWo
anGz6/WCMJK6HpMxOwh2xHCmKLEn7U9LjuK0nc97JDnMs3jW1Y3cTHHXooRFJaRU
h7/Jg8UqlTju94q/CwTQzF+MJ6CyDEi26/QT9nJJc5W63N7YBed5Dfy0Tb0Koan5
p+ClDKy49gSO9mMvqEthPZ3kx3CfKctoiCD7HN5VO9kh91S3a9zDjHTS36LRVfTw
bY61x4vcWet6sGTKHGTBEFTNmAsWDBDBy31n6eleh8Mt9gETaCD6VJFT/QoVm4az
d+U1dd9TfIOJ07EHXJUWcaMbgeN3Ny2W0Hegne7X7aRAZDFaukLoFQW1ilpnLDYb
UlfsczbdHtzk/k2hyZEbqnh/rJF/H/qWM4lRYsTPTZzx2rs0PfpYXqPMr47l+Ccq
8WYGZMdlgwHLDPCUhc6GmH+gQ82yPEK7PrNqDtVhcJ75VqsDL0phpiqVB6Hqc4mS
DrVY7zQSHamgkSnOvh9vbl5WJcT5z6flR7z5rBUSCOwT3gpflF5JL6uPl+85xq6O
i8YFw/aQBWXjnLc55IuKeP4yeda/JGMCPcjV54/tIaOLFFOBhblAKm+JxYX34f+r
8Og/qbJXeZKRjXTiEEnk0FqtGV710nbFkUTAUQ7LCkXP3wH3/eMFwywq8J6mrVr+
l3CbRDwKH0HYR6NfYm3j3Ap+Slt6JDjOjhJxqa1NcYpnNl/LiIW93OIesIN6LMb4
o1ri5szAF4kPZy9uu2AMdGcEDkqoEpsyKPBAO6q9mqh71Mdy+rJDRCHDpSNffGD3
FZgTyOiHqjA2+HjcqEmp/sDqCI/+Z2OO14Vk7Tx8lYOhHzcfAt6UU8D2Zc+7WgRc
I19V17tXHRTqhIX2JpXOK1pyIPQ4wnfAywVqW+rsm+9HaJJObWDMQs/uaZuVI7iP
kVAj+2DL3VwF+QGrSXECvnVz9ua3UFMxnXjbTud4DgME3pbf6HVY3vmVSYolQX8z
MhlG1hH8xpEKp1+hqKbS/gYAQ8l5rPkpOivrNDDP8S2wVqMMJtilIuzyxkYaLn9g
OWlOK4WNc3RShBvSolTu26cppD3H9WAAVym/lf0VPxwBPyxHqrw5idojjNYds2Zy
TWJuAxYrBvKUSYWfoSQu3o3NVMkMH5qpXQ+Hm7BQ06NGOJmYmQonqGUAhwUM6NXO
hrQiUX700ENEb0AW7UHeWfJB/kWoPELWv0/xep14X9mFqfqYNz3ibLsH89rwsGvm
DPqP599z4xP9vADTor4US5J/vjRR4QV+vMUV9dqXnjxslo2zQZCWbAMX+rxqdMC5
+VyIhgMWILcq94Qy2wSkyFrUAqXhATWUPABHkfwgfEX0Ktmxj194+jhxNr4RbFug
hNCnIQuickMhka4zKpdypdnr31X0n60KzGZ11slQrNvdx/dYG5+UpItTtZj+RNKi
aqA6YDV/9s46HkCBzZ5FIoVMTDZqmSUTgmUwY0nOteeY7H2/qEvgOiRjtQv7pjp6
avIjZ9DsgtVVQr7HL4MPUxq2uBEHEbYAxvwsmq9NVKpkbjzvSWKPXbA4TfMOHzvJ
ohPFPHJTOOnMwqgsMb3TrpirmaMUYiPnh2S0ZoxUeXMaXArXoQ/Om5KjtENx7Xlq
6/WCfH50guwuYESUa5S9U1FM4w1JzfutGGhbZKsRQos3VPzDnqHL/fm5MSox8mBq
8k+Ed5lTEzw9xMiuEA32BpO5WuIrkPAMazyGuq39vuM0xI1zub6rgZwDCDn7jsMR
JzeYsC4V6QA+B89SBNyvRwRcGFuGKfqtfuNUVVypYL6QC4aVdZQqxaVEmLj02Mr5
EyATG0zCNtIRIB6lpVOcABHTxYwU2Cy6zVar0SolQgR4cVI7i3s6QiomO5iZCAOA
rQUwgBQVDmiTRt6dyB2VZb4BYatK/kUAagFsvrDjiMHkFcOpNM7/EJ9VID4HtiTF
jBqNKnXUeoRlca6f7DYTHI+PL3WtQORBCuwapmy6nfPsF8UkTGVWbKoRWa4/0HSA
SCunjpFhBRqJ7OKfcYJYjQOa1Xpx9RXhxUBi5wIlnpujd6QGTUw6DkvzSRe5D4TN
d9hyBXsULWXfYByWRR7WDGSVFLtuKjZ4OFcd6cM3Kn6rD1+qHJQZiggThb8b3JAP
midGSwwLa94XI7PPEkln84WWoQeD163lVC0uPNn1Im4bO3l6YEXBjwjTGgWRUHNC
qij5REY+yMRWJCQcz+v3+rjrZ+SxCpAWi01cGvNvJGDSOQbFUI4x3eSrnuXdrv2f
nb1wt7Fephu87pGrJ/bayhhoKfT4EjXytkbFGazvn+hsepQNFOyJl82c3sL/uNaY
uRTODb1ILO7s2Txd+FnGwVr9WkYKiTQbsQB1HEn8M0yaXZLho9crNdQP+ACNtZak
aqGO0SzycMjUgHzhalqLeoJ3ylvyB0PkEzXW+Y1hwBzCRDICsKMbfQf5TN/cgC92
FkQdpBLKjf6RFi9uLuk74rHqO99P6G+CpicdJrqALrd9M4I5gO6owpACP7Hh4ZRY
1ihroPhdHooTNVZWFEpnwo+6k6jiOBzftIb9JHlLSxeEbH37IqfcW6s0vvC3DJjq
5OIvdO0tAevjgvyzFrEulnZoPZ88v2FvwStw72JF/oNcFdP8n8R+s6IhpAAnDz4Q
C9asRnFNnjN1CceLnyiQiTjdv0FBaZw2d/9LAiVUzdDougGQZABzMfOafOGVuXLV
y/5bMzPag1D8jc6TsVL8NUau5WA3DcEenURVR01Bh0MvRJF5v6AX89a5sYnmMABA
Sgm/cp+BBDtVsGVsbBo40G3O8iyxrWYR+5AfILA+zddndVjPBgFS0V6q9EFAX0FN
F7YuVDIrehBPtvVmvsi0gaUAulYJIDhUL24MSfgBWVVWrOtPTxRk6I6w9IP3MfY0
Zh/6y8bBx393icPpSaHtwcUdyWfoxZieyRLnTTXojg5tQtHvsM878NjNV1tZysf0
0FITBM0ZhsmZpbbviq9bz4hMfpPpyllv/bJl+agg7/t1FBpR9ZTpZ7izZ6u88wpW
Hj1skm84fkJkVfB9NowjqHXC8NY7E5BptOHUvNu6jyAThMGU2DhbOe+sEiO/g8ib
sV7zrUuv3BS1XSojdy9HibB0gIw7X2ESViV0g6W4OOAF/RzNgpVItbcsbPpKT7vO
9sIAWXqga7lKb+QQAXOp08wN747IgKweNvCE1STqiC6pr988L3RCQVAJ1FGJKlbp
Gx7q6fSyB8k8FTvCk/PazlEUriy18EDB3cRwyt4AaK/U1wM3L55tgEzdbOlPQwds
GwdTUpsvp+eyxeqo2dHhneQXCOAHg6vbSoOnuCFh+EYBzCdPHhmcvV+cBrcnFEmA
Uqpw1y38S4w1qNQPBEXtu7ZByMmHp3gQYQZIaa0wPbjZhIH0Wpm09mPzOwGWF6r3
nTe7yRKsDYsniL5lf87XTqZq+W5Nd+fFPBaZkaOSZ4sOM7xXUZ1vwoPg+pZ2f42y
tOj7kjgpFbNQjE8L9o7q5WqJGhTBwA3rSMz70F6VCyXNNuMPQtZrC7FefLrMT35Y
lBCd9aCoNw6oYe0x/SXghIkLdwO1sUKlNwwJWwslkj1NzTatTkDsVOpBT4kIP1Lc
gAwM/gyYsRH4kidKLTizcyR/cSTDmymM4sy5pdAY+9K6aez9RzkMC2PbjPRS7v4x
D9v1+OxwwAP11gQ5cNCnwlpzh6w6YHvfr5uI/0DVStl7XQMjZM8CtbL3uoOIJdzU
sqedSlBfWH5StWoEqoPagpc3z9ac+uJi+7Cf6zns6plzEfC2dOFNUtNV1gmaNWhg
4XiccxFcxfefneRhINWvV/IwJNhElnbW3B6rBgqUXS8X7RYUrtmJw251ffo6+D+N
Yu6fEAE7hZiI9b42HKY0S7wokpxPkjR2wz3RJSgLCjvGLsmDl8sDoLMl06Ghyvqe
3mM/pNK1H54Tl1jt+CmingBhP5BZU4lWAw/srkUatbV1qDvt8oURTelmyErJO20s
zQBBNmBWsT6rASuVRAmyqQLCEUNdjWYAmSh8A0Ld02EckqJjLhutC2Qh8FF+2XWY
jNlqizajwSgPOHEER7y5tOPm0La+HdOHJbzZvLaDXJO6bTFGUGTha6hSNeBX/mqZ
UwpJgUTJDE1JDH4Q9mznlbdShOnP/OMnXMMRcICzOfl0P8rFhDWpum4Zbckpx/u9
5IWTZ50SlPax4X1hAfTN+nLRTIm9P7FfElZHjoEb4/kHs8a1zHrpQqZzDACLQVoR
PlP+SZ1bjRjPlI5tPX8qJzR/u13xeP7Vr9QlUki7Jcebhyrj4L/dAogznesZa9tJ
G8i15IsKPsuij4noBxupczJYiwVgLZsLLGMgJkbEllwjgzEwBYvRTY2naZ3Kt8IP
YvdRNcInn2/vdMjtARBE95YrB1E0cHhdqdGA8bgamzXX11KG/NeWogYir4yM0IRN
eb54yx/+UfiR6DHnEX7gz30r/YjgJHH4IhU3HAIZPFBcQCTvIc9Nnp0MkPejVIYh
MD351yNxbuQzRokQkchWvPA9ldN3HSrWOeibp+X34w/kh8Zrj3EjGT/g8e25Gj/C
aQxiXeGKM7+xnzcWTGsTkBoazDls1YV6PYRC5tUc7BfY6ddVoKLdJnLfF1Yi4BJb
tys+UrdWxvTtziTzTevK4Nyv4saP5lCyptaGBv4MtWgVVRQG6Ww3oSPrAprjjmxF
gn5X5tro5jWzJEaznG0P3duCJdUA/vyAdxfN1mYMFh2uFqMZQEGGJVniiC3r3a/W
Ul1jc52noutSt9fpHyZsCpypi8OQfA6vWgmRZpQ0yOQalCH/4TzedQVPdrcaCrwV
VdglWWWshQL2tBYZImJabbbWAhkOcK2QE09DpiFCuV+z1dDc/ufH+ezEGX+IQ++f
7yFrkdySmW2Bi6y4/vk/2xR/tsftw+tWJ7b0u6IpDn00Dqux5GuEoZBuluTjKm2X
G4c9ctomHwx7+lUTxp2EApKmsOpthy/21WjHW7KIm+1kVPPdBSCnSbxXtB3EmACf
1WeE9kIlYF6qiDcfqhxsFxKGfnK7RcaShG5W72ShnDhOYrtdrvM2bRe4jjvzQzoU
A2xnzbMN7Uug8T/4R4UydTG3dngu4tmysb7wcOjZFkJLwd8u1stTGCf7mlLTnnom
Po3rhbotz//Dq8Q8hoU5ugllwLf4sFXNSbguwTE3f6yzR7QwVzx6vPXNo5Rjsr16
q0P8dtV1WB8ppN4i/gnd+GiS3EysaA9zdSRflSnTwRXii/+6RAA3nSPycYc554AR
3+G3eqozM1WbA7fu2HEkYEgEjZ9mZqrsgrWVgUj/+qJDjPMEB/tsV+XXofraAYSd
lDS61+AFteX+4YE+PVCRhT0uieFAklaLE87TourI/w/ObFVj0muiWyzrDhm95xED
iz2iisn6ItRxOuGRi7IHxbHXwSOyg8pYOcBJeQMRly+qv/n8dRG6MS3MiH7RiZGz
XE8cEIusRFFcAcJywUEV196itqQH57C7NUh4ZaEBj+vN43z3sjudzV3SjU7JHP4B
inYKBNNEPVoStpjt/qzTyQLttvalmxe6DJV8w6J6MxXeF4ESZN1/oS+IoCiITyL4
LdZygroYVb/eK6SeW/8QyXMhk5P6zZwzpN2YR5RUedsaytVjm5QhepxhCB4n+Qla
35GZf0MdnRIVkP6ObdCEz7VjFrfew+b3GAs0RyFeNQqUYQAki56a6SROSwoz0d/+
bBoejHbeFPd71cxqjYFPrMeQc0XTiZMwDvXbkdqw0SSrqZIbl9SIAczoSsclroiE
BjSbGG9rk5BvdGsL3WAb2VsxbcFXpwwJK/+A+5sbsrxoKpEuTAfEgOFCl+R6+YMk
a/1ANZqbnAP65lDneb6aZokEQu/ImC5FT6ifp7qsWNPi2xusqw+cU3zUW2dS4vjd
5FaeZV/+TLCRUxpqpDoKMbQhlwkcpvrahcmDhdT/YTC2sjADdjs8kZVBSXcCJs6b
MS0qrywQQHtMMauwsj8TvXrfjsrYxnSYNaHpFuBHmQkt4uXKqrnCLdDb6OO31GtC
ulMnaIi7H5fV+P43ORrv+qz8Ink3S/0tAPcuf+TByg6Tg1IqORv/hm/mCQhLwbVS
dnk6BCRm0lzgMkoXTIl3pPNM4ndFxIqhuLw3faPtF0r3hRopN2fFctDcN7fu5X+6
XLGkjIrEpMp7NEObKA79hDM+kGIMx3iLodNksbzzUJCyFlKwGLTxp4yLYGWSGBA2
pTaJobBPCaMrZlhErtGBK5Gj+fL6L5T4wwpAev4Yj5PXk3rqkYKRDmI9wizGjrDN
f3EQmYLCLElAXr4klxIolX5EGzHZtJojGjtxkDG5S5E8x2DERR75E9GFCBV9bay9
GUa4dDWwTtDWahsGN2N9JMZ7tjTfW1LVkEzMgJn4wkXEWg/27wim6udE1p9aol5I
VaTVB5R+fMhcK8aFg/RzbStK6mU8lGnPTQ5X+CX5r8CNL4rT0GSKF1mdB826Lq65
yWlwaMsBQsoMlOTIuaibLVcsGpAon5fPKF4CThgrKeW1hN85vTef3NGYtVQqNCbo
EUcGBfDKWEn/GEDCre72URklCKcze+WtjXDEoz8lBo6O+VqzZiccOGRQiCpaVi6r
lqKzcYMQ1R+nIgoY5a9ZnSngidElqIRqaS7KaO0sg1e/RAzbfFqJPVrT2InBwYdy
cVjxBEUSG/zT3yBUx4CaSjHuC8jpGWB93ojoLpSZKu8MfuCaEKlkH8SSibeG8WkV
bz/iY8e85LfcB+X4UtQ81YkxNxjBVPRl3avjM4lZyPMFR3PvKSuHBqgN4nCqhSym
BeN6bJB8feW4NypI8boLUHVN8bqUyVhUhpQIEcd4a4hcA5QrqRJAs+w1hzS/npPp
h2mJy7TRRulNItHEIwDBzVLfyJ8DXXdWEEGQUqKFVHY1i9tnhyyqIZSPLqJqQIFH
fhh6Vqwjy6lUnQGYFsbSKuV1b26C7IA7p4SmXZ84MmOV92yHeerEgBpL4s04+cgB
40+TwvsTRRKWD+XZEkdk1oYsSNN4AUnvhAtvaNfd7i9kK869f81LlsBzKd2sDOWb
YxjC7YobixWJxMOzNM/dxDlsIER5c2Ti3tqn+0bIWxXdwWd72Z6/24Cwli68nHKr
SqrTSBcTDwCyfnE7qmfMIMH3DOme2b0vOKEpa8TPXl5vwsnfgPkofFFUXllIOjlc
V4ZAWDo5od1JcQLM0PamXxoI4rKdRADhhYc1rL0/s7CUF5+qvlYD+AEZ5uDkTGCP
NbWadEdun4sOAw64G8J8betJX38eQJ5bdumdGgJFMYMoUXMxokV6EBhjcdRKQrbQ
qm0Pad+AlJb47z69dRig5h5H10Vd+sN/W1J6eEZlWVby2/6oIj9xVgSHyzcK7ES7
t0Sa4vlYkegs67Cvh9Gu7P8TMqXS7pv4o/hYiSYCuXX1g9s9LCepl6a353mBUwuG
xF8Old9eUqusJXFi/ayed6Zu6xYPD9jzpd9KfIaQ479LiOeR1DmtuXOVXnlzV/9t
C9NNB2kUvhI9dQ+oh9Lr8Tt+P7DLXj6l1187v06fkDnEEBCuBE0K6IZUQfTMvTv7
78LCdpxdbpKsZ3w+cBh15vRhscOT+b6ArRFvFMgMstYCi7uUqWHh/8hSSed33fW4
ybmSvUF9Z8BEgnS5OLBJcUWnIpCDC6PAOH2TAfjwcpqAN6pZuNaItHXMjp526Q/R
sG47nTb8C65L2yhuOZx85Nrx3nX/tcmNhw1uO+MAxasnsMI9K/dBjLwoYJG0exIc
f3aTqJeCuSIZ3wDIqV3NlqM5wYfnOQbm1dhU/vEDzTY3AYADtDWH34LuhJTj/shI
OS9dGpDEtwxuZmz7r0wRbZwNTUIfdhrrdn5E1mBQkpHl/NpbKZTR8WWHHhI86k/Y
iPUiJi+IHwJBQiGltqna+sCiAMtvY02Xx3RoG6o/TQd15bxJqyfOSOaQBhhkwPrn
LP960yGxC9NvgJRg3F50DgBbEkuFnH5qh9RHve5CizY6K4UN/eYivq4JMIPG+jdW
TTq1RJCq6ixblv0ZOShvHgFh5gaSsjew1iGMDDpdmXgB8GhbWNGVg1zkG9yc21X+
1wLH6LYvJ0vXvMU9Kq9p3vs7qaZBg6s3AE25Fs3UjYFJZ6Wb3f7lpDx4+m1eNejO
ws257BoviB7H0Z/u7RGuigaHbIE1olHowKt5osPEIKIjeWoytV3s9iO9OdYhyOed
pc8hjUQQIieDo4gH5Dk/fhgrdJbQqyBIwhckmk31l7GPszNejthYWdXiZ8xokyuX
buFcXwZ4ViRLmrIHAiv3pLlSMm6mGu3/xbnScHMryWHx+dKXtbEVmgsEAePF7yJD
UbVMalLUO1rxHxGbHtUmuLOx7XImZ8aTNflxISdR75bt4jnZpr9bmGPSnmTMFrqB
7oMVKS/nxSBJu1aOHRoMTbji44qRJ8iEJAzNrVmaHaMIxqMmCt5ye/JTIsUkBJdR
WzlYVGPWWyQr4u9zRjeOzrbDageyH5mZnEFhMaunribVvJkOPOOVFhRLttP6q211
d9+ygzaW1bt3DKrRq5T9KTBlnnwbgtuM+wPgYSdEs/vt8QXIXGwQna+tTNQEuRlM
HTPGLAHYDKOk4pkhsmfT+spl7QNMlDcQYXU8CnfzaMvyZ3TH+B0XEqfytJk3t7hM
kJtVK3A1qiEJvdWEzHsW6KPXV267rf/GTcQPnpyzVyb9bjDZf1d+9dyevRBd6eyJ
tE9HyADo5uqan55w5UhKqSw7MbNeMdposHXoJeQKpFOdBQDw/4Wh8pFBph4yvauh
tdlz1nMMBXvB+LQWHpVeKuSFGm9hOmCati1lGW5y7hagblCpsgXmBdorSxWr2W1g
yU3Sv6ekG6GRFw+T7TDlibOhmpITUxyJjdSfzA/b9BrjZiH2iqCTvlQ8xfniwI7F
qV/UspYA1H2X3HB4a9k/ZQ==
`pragma protect end_protected
