`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g+kNeEZfBN8tG8uS7jW3XiLDgExZqaK9wHxgageQS1nI/9q7+vfi/d0qKRkuDWF/
t9IriU+yGzYxoAQLrRtWdewIXwutJFeyxbLqNmbAv4dTnkDE0vqDAceg5LGlk7YJ
oEEwq29RP6ai+0QERwXsZSvuQC4QAI/6Q4ScOvIUin4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4784)
G35Mogc27IoTliSb43LPUfOZNCcby8LIsUcwI+pNM3DtTrBsESGghJTtmKemMA67
1MH3xPnhvOEa95cQgsc+90JN8W0AMtKGaqGngrWuWGiWnQVihERKPf5ySAX6qAQx
0xdQaYC6ISPLI2JRL3iRMVBTOzD4MB5PvFFBN67PzuuFrtSftvEVZs5bwQfMsSjb
PBBfKblPbxAnCxJxViMjFekCsOfwR3z8mdw+OQrDsUxj7gkp4uGpdOcKvzCQuVsb
dJXMPOVpTKWP0OaZhsX1SDHbRZ/ByYsROm0K/Fpn8KPmHoLMBmql41dzxEq6xIXP
K4H+X8O4xWMZ9dd+cY7IEBhcEyI34vsyjmwGFNrrC+Q2Fl+l5G3xuuELV0AgRtLX
JRAfZ6NQkyYov/28WLxNKuWTifcuoO3QIaMVGwUVMVhrxBXoLvWu3xCyQekiphmj
se9z8UhGlgNBnm+BoZ/lh+u6R96oLSR/dQdkxpJJBkri+cuX1X4GfyYwEK4PKmsn
tsESYq//qEK9AHFhiniudY7q4bQwJ8NNM0YYg/xUHywOjk87Ay+3O7kR7BrEMe6v
HHXtc0GAvFgn4JfXiHBBGJiLvRiE1nv1LS0KPCTvHaFHNoH7zfBY9zMOTftXWJs8
XiSa3gRUnXw96OBF4ast4Dkr0HEj3+ph61FHZBhTw2z2IiKJHowWu3Wl335p6fVe
LppqlyGJAnbKKQsrsXubHqfkdK7DZcVOS9a4or+sEKJl2fMzkybZkv+PZ2NgA/xO
8rVISpvDgjMLp6VSPdI2xoXZUHP4bNO2Q4B+OEqtfIpMU6xoCXvkZOzJb1fl31i6
6pJNC5Wns4m7hQiUtX0yXahmLHz9hQi1xb73vayegg54+n0g+31OD3LdZoIlKY2x
Vhj3QvuAvpH0L2umdsi7uWXizE6OLJHsoFTrBfIhNuAt7RUO1mLUYrjJFwxOoD/3
bDWk8SE8s0/cRdyUQqJJTu4ugF0wa/j/M9eqtLIW5O0ww3ijUvOsDC/uY3apfMMJ
nlE9RwpuCSR61i0uUXgunw5pm7qiTKaT6T7jzU3mJd1u5fJzVqRzXFpOk6PdZS9O
8BbOajJ9uSi99c9RnRhRLs5YD4T8/JeMgBfhFdwcidZoNihLJiOtJcjpCnGYbuRk
zr+adPWRPOztaNav+1BfHWZeBTvbFIRnwx1t0Ep6beGEYhoxREsYlxRa52ePgbs3
7UbQ724Q6AZ5Cl2d4bb5BR3UAkCCqK4PE2B4hs2RPwNylwlug3PIXYNbn/NTOuGM
jEweLSpi5up8pY7HNXbSLavV0m+INwDS7ezXFKxk9hGC5CudoGjZ10HTYHQvg25c
m5SwOZpmRrLdtkw6UkvGo3Th6EB/1V3VU1DzHd1C5PWZQKmVtN+Ujt9CsGZbC72W
PR2OYawM9uShapu306h+A4+QFeTfIm2/DpmkC/8QUxd3WblZtYOAOeFOCdl6ruO3
/f45ng8fyjRLqsAIv11371nqiIYAYrp2Rg92a9Wj1jpJvMdGUMCTlyGMPhSdWVRu
9WfdWFcABvgh9UVF4PgUzLUAy5f2xUlAYmU2op4hWEdZCDpisOjzdkRVRZLgAPgx
EBt35PN0ByTr5TtqWtXPif9caitmGrpsVmXtr2yno2adrXEHTmMcHnWTyT+UwszS
JiblV/bTIBupyFwOoQSo80weZDg84dN4mzEuq8aKTghKd5QdTJWIb5H/5H8iz48r
VFfp+j2zHsodoSmqnjG1MIbb5umUDpzEM91cREprz52VgZzSsLe0god+fTVtvaLd
N8Oj6iSNrtNwglC9dAnEo/vhyQHUvsGH6yc2Ivx8H4jTC//WJt+F+4JM2TKELkUn
vZyoLm4IEgyF0ZoYY9KJA50mTtFtPTM/oLO6QbLGeJJ5H1bfniLtspRDWX1nXiDy
DVJHHAYh3EfqfiLNTJowM2mkpUudPWG6/42p9b8t8BWxx3JZVpnOXagBHhZsYmuY
V+QZPDPGVofsx6Uwtu/dNaaQbvgBA8U58MC0agSBfjHf5f5Bq9sqEqHHnaI49lHT
A6JQoutkV/nZB9mJsCgl2o4OkLYdSYcFlVULOgUaEEYt9jIyHN4G33W0CxnoDLiL
AVru0/GBCtwfCdRl9oppZ1TMheGPs5tWOSyZohcR+5UqtR52AGYWJI1p/kwO85LL
WX/gVHVi8F64MTCUL6f3Ofso9RT5Pt22++GD+ZrCRJp7gAOfwIbRMGK3nTow9C0D
EFKP4/1E8eY/MkdwKc/WyG3ydT4LVpavOQiN9WRHN+cSOvwnYLG98p/KjphrU8Aw
dyrAMgTonIw2lasrLzeo3Fc4yAZcRecWn9WstN6m3a/NnTRpOUCdDdlT+z6k8FwW
0Wka78osVBebwRUo1ky+xorbWhBKjbexHTlWb5E+frRtJ8HjNkDs2EQynBgd4Y5l
vdKeWh+YPY5ehtORFPx6tLfCwpyi06SBcehfaSa3g7GFSv04SGy3i8ug29ildRtj
W5wdpj8un6UobCrQEA6YaIIiP2zWcDkQJMH591iSDD2xt4/aOfmlITLtK+HCe5Cr
OOlTpNgsHhT6ypSFZiPRA4ERAGZlNJeXTDSyltXcY1EBfSVM2ga/ascXwennBUJe
UoHs2X9voGV30ZVrd7lTHcbq0xv122tuqJs34gctZi2sV3EeInWpYvkzMPQvyk0a
+ysmPC39isI4zp5Y6KrqcHshtsJkB0zK/2Lu3lseaG/1E97i+rZmRyeMQednffH1
bd8OGxh7nmUPxrt8hvdR6xLDvck5KO23bQnwLJa3B1ttbdIFGN+YXvB7Hlmuhj1o
6LpdqbIazQ6tEc3jdWjaSu9r570nSoVK50aSltG1tYOCjsNoCUP/t4ZNmDr/mIaI
EtNAiGXsahcABiPPhFiSk1YpU+bx9rjPCia8WP5jW2KIRTvutELA5pXd/etFKywy
z2UV4lYiTqcuG3+LhMOy8OciTAPY++B2TbEUTDmPClLeuomXu7P8WGgk6+sZWYFj
am7gi629UoZC1nrgPBFoARkSZz/asl5wwT/jLG6kUQu88fapLaLvzOVpeM8yYihu
/ZaumbtN/oVmcjQU2Zl0cnVnJ/R5fGjPWV23FnnKC2YTITUecjCsUOp6RIl+CiI6
bBmDU85V1Rml14874d171XaRo/1Ft/aUkwFOjGX6juMQfoedT2twtioLSTKGjYmy
k9VhTJ92EcY9HovKJA0XvxlArFgi3SB4amZa0jVwbezHSMZn3UE/X79mIWvVB7oD
9tmrHMNKZUup2RIvLrwl783NN3peqZnpODaUy5iGwZZd+54hw7prz+rfEbQSWKXO
+riyyA478RD/oFv9C35SeLzKWSHCfS4LDjV008lk+GKNKzJHmkS+1BECAD+xkRSd
UKbV209nSkb84LxOa7L59IBHX9aTycIEyrHXnaHoIjhYmxf0LGBitwB3qd6PCmfm
y6qNGrHyKx6yQflqupXhSL41Gg1rvctOoHZV4MrKMhxrdSBru5mOBshhj2qnfgvh
CNqvRL8AVYvZXuJYiDQYJUAGv+nAq7haj9QhKz2KDApK+6JGXHlkwJ+ICfOlZxzC
xBHJzJwV3T3wnkLxkAw2qImMnCZjkjbuTUvaxWS7TcRI+ggN70VieeOquXSa+NVz
t/0fEgXtcnoCQaXgHhsrrqF/gMsISMxd8iIbEfE8Q5J72DsdZuIGN1J9IhM76rav
lBhUF+CRGeyDCy7SO/GyUN2A5tqNrIiZXC6/5tGe9gEz7qquj3WTjyoKRYVtlFr1
8aC/dbl81z4YSGvWJ3KDqLLiN5OAMmHo42GNRLvED6LtaM6d7sbHvT6kEb2o6tbp
qbsTKxbNsddUH9mzkk1ZbAkN0sLniu6fLfVpBvfoA90951uiWpRISZBNTQmDUpE2
lFj1qvnVoJyD2/5zzxZ2/gQi0NG5rggTU4FP1KvpLyM89jTcxEK8/SJidd2bv1vr
muR4z6QmVM52rVA1T77WQOoBqOkd/6dTzhSuJsogLe55//1WvRrpCNBBri0kOFxb
KRWbTeV+2aDydgoFBxnfnZfoSFp/vqpaU+n20ukyLT1OFb2WBe8A7cHJtwBcD53+
wZ7etXVh6YbfgqMurOhT9zIuIaxIhSY6P8h4AE2Vc/s+qSDxF+oPdgv9desfusUS
37j2GOFk9yoWefdvsVtCpkbYwe9LJgih3+m9ztkwK+cgxQuUnvjlBtH/wgZx6LHf
BVqZMohB6r7F9Uyq1aglUrSux2XCGnfqKUL5AMuoWh1fQzuJStcdxktji0xSEk3y
uW6odhynXtzHJHvbK1G00MdFezlab4mlUdbbsDiBlV7C7K7TNdkTiUlA/PXcnK/h
Qunt90jI4/dqbftv1WPCKnK12mv0frN3cHC6cr9fZbGyWteChzFFvHJI8BMlbiSZ
b7JBhOlXQJsLtk3CRrgcrlVaDntbWC2uNCuw//ntKxmG4aAMLAqWq06vCRgjRUzs
4edwS/7bjzcvNLaukOhIk2p1c9dIM8GUq6kqXELrk5/XBjjkalgHJdsQrThB1Wlc
R/dMrWg8TiZnCKRG8yHPv6kg2DOTYTD+TT42Wjzplx4X2JJr2mqig9PyPctgnqL8
xitRWseQna2uSkJKdjEiGmarziMrYDUeE3ldZ8B7io2yZWgA2Z0KNi/3hkLHGR6Z
jeBGl1y0L74lCqqff8CYIPpiIeg/eRxFbZk6Loxsq/pMkdgZoep61nW6qfIQtxki
6pW1aS7fIhMObrvc5KaoeNrfZ68YAGVM6/5zCZ+BY010+O8tz161wUMHUBxW2e4g
fF2q88ya9vRBkFh1uoL2RNgAmr2syvXb6oy+jFs1/ufe5lFLhOjWfF5lxueNylKV
tgwSPWyaS0bibBuHoeZcY/G6XRAa0UvdPYQi/3hHBGh6ec6cG8bzx9m0Qeua3abO
0k2cPbjeRxOYMlFCAmPGhOjFtqXR1Vydqwd0v8Rb+YkEO8i5QCtLBqZlAJN8URsS
OfCeBbDnCaa2VVt8g92GTCCXHkMQf8g09T1uWSifg876bFRx+tN2KstSssiZKfUl
r26YBDpj/niMeDgAZvjhAr8k7jXEVv5QOk3XIDLtqypJVMkjYwtbwL3WUgCmgu/j
pROmUlNcTTLXRuuHvNl3eNT6v75wTxTvW8a0Ypa50B3psskTviV6sW57i0PQmzWU
knpFEaTA+EdQ2ledPZyp7ZTTCAj0Hadild2mjMFln4uoglzxxVSn/P/iWD/jnZg1
F5SNaqmb9Om8McmdcQ5u+R7913XaQvZ+Zg/8P7T2Yuj4UrEkqDDbsLry89yRILGm
A09cz7woaWv+hDPUbDSaHDJjJi1MZJmHF8DAbriZ82DFRJtHP+WJNM+N7+T6MgD2
jP1h3laODg15uR/UHJ7oAC5N27cbrt1UOORJ+0HKcyC9boYihpxx/G/2uYwypCGh
IzBBZS4SZ63pwPlMJXAC6li8Dot+6A3C90yo3/rwOBImOj6+29M3gNiwZd2ELMyP
oTK/CFkPFdIyikwEiw5HZZ1k17yurLi/OACQROEG6m2b/pPilIn8IggfxEAK+qbq
uvBkMcfjmKjYyjSBNV0wr6DTGR7Q21R5CiXCkFRmukfH1J1w+yi/kCQegbRKJD9D
Y0PPmN02qv0orXXQMTjGE4wpw9+6dmlC4uyq3YkM0zLxeYkJq7X2SDd6Hs/iZuz9
PfDY5nkP8T2Q4WEDgcW1LQ5YAfMkiif6ZhLbUfis0QRPmERjYevueRfUwdRpEFC2
S36iuvlFdqoAwfWYiCe7KG/jm4ybllzOfoWtucRnpjgUk8lbwzMS5gimBWvoQ1VQ
G0FKo1yHFa1boQLAY0uKWzVs+EtWcXJdWts3WyH4AEQVVF4TiZbO4v/+XGdA7vxS
noFEim24GBKT49v9NR7/C0GhYTfNE/N4WOnLkshI0Te3iMEBK22HTxYwzmCJnbhC
G4S/6L+0r3i1TyxfHyZtYSVI32Awd0vhYiCJMY3JqBuLfhdm0isZ8UT5255B+MBF
vq8HLy92GS6hukz+3H96fls7e/rplsPFpiNjceF5zMWcQ+QfTpdmItFUAAuysXWl
m9dX5/jQh2MvgJT3jdEBf35UDujcs7NEZ2dY03ErA33LmcufAdtdBI5shZfKQ2tN
6cziLXndeKHv5E1Fx0JZKGDjOqAPcRh9jWHiUHBxT75XjCfwkigH0SnmLgheBJff
ZIQkDS9s4NcOu2+YUjPu3pWZMm7Jv91zqogA19uXpAGAw6vERUdZqwTCQocktKTP
W6LMCXzh1blobsaWYPfDgtI6uOiY9eQRCegWtw8eToRZ12FsCjBUidzJq0jLtm0F
8La+4c1hQQASeX1f/csPKzqe646wrK2pTZDhkzudSsQ=
`pragma protect end_protected
