`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZSIoMke9l0obTCC4tRBUpS3FGhZvzFynEd84sohYclbNMMyzWtDRuamWKAGf4tpL
nXh1oPYnlc2Lt5Kag+FfEy+60X9GsHy6tSEGkNO2017OX9djAmVoVXWGCGM6RW6U
P37iNqiUhU4mCCq/a4msWlY4iG0mQWtw6eM8y/N5fSk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48656)
hlNg6ansaFD95DGx0lrlf96qaqU8Y86qlAgnmXdno7pXk8pHVvuaLtZm9t/2MXpQ
3UMsv3xqECZvk8pyrHBUfa6LW0QYKVs8TuHnMaZnyShkwbQhRFIxCb21bTQrg4b2
kBx3vpvpBsExIwb2UUCod813SNDA5IAFh5MFNEQ5wA+o4gfWEwcgzF6QWXozCe7t
4+1xpTkwxthM9McUM4h1JHXovE/W28VlREUxbKo0eUlfAMpsMDwU4nFH3MEBtZ61
FlLL9j7HyPhfK4FXl/f9jLzYEIOtw77DMFh3Hu2RHwoEvNTF232o2jOOuOIGTi+6
AT5rWMZWZ597Hvgkcrn52aaIwRawp0a7wqEHmJckeZYwtsg2idsLEkPAAZAyCoUs
2jI1+gP8n/k09Qo3mHHdgx4J8+T9JqFrJnTQHkMDE8Srg1mKafEqUIB7c357OJum
zHtTm8d+iAUdFQmTJeYkGZnvAYySYxTO0EwrV82AUibVkN75Z4xzde1wjTfKQaEk
Ps/TfHuBfb51z679MH+4luvwTdK1RB4qZdNkjXA41bHBJlZCKbK2KJdkxhUC+aCu
TkOP/jmtlgNBFqwyQye7gvqwaA/Y7qf92wFEEe519Rm1Z4vX1HVdiKZtlodzawGG
NngYnKeEhkT13l5DMAGkvcmLVsiouYnC9U0mf50U7dj8Zpe7L4Ptut6NVldFSKkI
fJidmdd3Jn5qe2TKKh818Z0DNdy3EWpyev9ZUFsVrxb2YEStqW7k43PbQHRc0YnJ
NinEbV5oTzb8r1quK+XT+CtN6aNa/6CkGWxRBIBG3UyWC+1FbWnlpRAs7sGIHFQv
/15RPodgamRMkGdOosyWF+AIQs4X3UAyV2FH2UFGb0fDA7Q9krh3GHKZ+vPGmugO
wl4wy7nr3PoC+vu70u4LOFca3DzbuUX/3aOUYZNHGJU214T9ytKybZim7e/EsIN8
8QB26bs27BLbbncjBjFQ5gv+1tMps09DmJU3Zei9CJCg7DuaFKVv7fCUqSv5P5Xe
fXHLjrnQ7VhLP0QG5eTOQAmzMXaoe+BKR9y6IjtPfXfs1x0vYFoT4JxKmtqNIWYf
c5kbS4fNVdyal/z/UAc2EAWTQR7Ai/yOCVpPGToCeAmaQ0Ep44Q/IdDrCp/60pdx
/oM0/1QYRTvf+PjB5zIgda/31p449vrycf9UiYvRftOVfi3eT1kGokLfZUZFVo+K
pC94w5HKIloR2JXqt4h8mPd/Vhh8ISeg0dJc0IByFsH9+catd9r7I1wa3RoiFCoL
dVLmW/6aTl/Eb/QvneTzbofcIpXNrJuzghf0Lk64w84zhEc//4SX3799P1coZrFh
9jPRZ3/1liXdUKUSDjMD5t2oxEOk+fVv9TsfdJO3e7GroyWiA1btIoHMc1vuLIvM
PlZoF28jM7vdAcyTqOcAw1Q8u9pnhOUw6qSgsazrNgmEgzooVNBia0hU0K+uKojf
x85PKAPE3rx4GcwgFb6lByTBOVBLeG66tMjwHhA0so8B9XH1E5nhMyDw2Oz/p0D8
nwfiI7XF3SOARiv3X+1smVYt5X/oWu+BHDmay0ArY58FyNWEkF1x5r4niCWdJKvD
fQZRy0f47a47ZmtpOucC9DPZ/tPaNmjE8vbJmwEGEgOY1fkLp6ZBF8gK5i1foq/Q
xZdRyhkuQ13RbcWM5tyUXJr2J8p3mA0VAoQ91uoC2ZtEj55wRDwG3Ezeq99GuqM1
kr/WIGWKfzQxpEIF9Vn5kpIY0i1FC/g6FD99MszhkiFOrIFLFyMrmPoAYp1bYoeA
2o2nX0Xo0KiOupObN3k2206tWXfxFKo7470b4MS5m+ZBDT+mHxfIB68LEfenMMLK
lZz3jfjleg+/WU/it7UVChzYBDphLkKouuSO9JQVubrTLO8atAZFQyO1UYZnmitj
AE9HMctVNnGUwYr3dXJDLQUg4lKpo2MwzUTK2rSbQtQa1zNgR8/Ch343Fk3m6DiQ
E1CiKu2Z8CU0Uo69vsFoia6DqESkO5cs3WzA/BE6b2gKol6u6dAoaLqrCeceswAV
yPMpHKaCgnvaVXtAg2FV0lUz2VszFNXhop9qERJFDHVxPBbgnzJ/T1nUFtKX3W6Y
76PkxSkykgI2RLzTe4VtlVgybL1zAmgDR1jqio/56DeKAbfn4h0E6/RpVbyfc9Ij
2eMI90zhLI/e8FqZ6vXgskQGyz3wBEf3E09YxAxsdkGA9EdYfnrj6MSTeNiIFs7X
bSenmIkOR8oTFWG5uqcUyiMJHl/r8ghmbhanQ0vkINVyoxe/ufNbwyw9NFSpdqPY
rv8ZDOP3AXdNB9eFhvLsdjQiUxWGtJ8kgKAVP2pWggHffCsRzZtKhlQIIWBIyh+0
+HEq6PQzBvVIZcC8qQfpMqk0UAq62Y2yEDNMJp6a+3w8jCRcben2ubO/oO5rNBN4
/v9TyTevGTidxLdGhPgN1qbtAeKula7itPbw2S7ym2xzhY5Lm7wRjEj/OrD2DFer
/zjxwMJZuZY9co00v9PZU8+9obeL+XUHH2ZyohXEd8FCeVJd0mpsvd5SHRzofWzg
qXntL6IeHzglvJI9yZpr33AWjPb6mpaQcDCBCVALbZVk3OrzCrqL0gkLeQY76vJO
x436LgpY0kNiIprIlp4nwUFjV0+ZH0OYwHHqnL5IOxSLi2FPfxZtd0OkKlFDiyTU
AZrX43ER1CbXSnfNFaJjHHnrKZ3ezAiQfVs8pUOpSSSEMY9/4i6gRxJIiVdQRLIz
wbi9RB1sDextRcqdW4izUwF23/HVUKKsUc6BGk4IZJpVRqiGPWYp73lRLEgRIPGS
OLpVw7gfk2FjoHt9EJXXEjvtA15m73FGsqtl4sP9JNfKyHN3cMHvBicFiK3qfpf2
ceEnfi2YzEcm0MPKjcyGIg7NQuzUITDp3DWNzvqKP0xy7l0WqW0rqT6gUhHyvHvk
JWCVJhthDIOCpZeZNJWOtkPL+3ocNhC2s+n0n/rg3XnOzTkwDkhvW0zO0vTiaQey
aN+gFbhGFup37y7iqgmJ8YRHWw+pTSpRQ6wXfilqjWQBAAIsqJVcuwC3ZlC3PsL8
JjxX6hyvWNOvu9vQeaVe9A8UzfiCp6u360cVU+SYVH2GYKN5n6S6ckFG7IZ70uqZ
eLznrJXX7JqEUpUw8sT8O7ZnK3MdgfcJ6JlVmwzT5CQgkOx63op3L2alu7hdWnmn
vLYkN2I5vH05YuYcYGamStnvVofJsGrdb7ZBvdr1SpiktlGFVt7yWf3LCfCo6ReW
3IkatNuiCZTjypGegc8qx4WLBy3MGPYiwF4bOkVRZh3oDOV5ApdLf7wgAaZXLKH5
+Wr0JPT1EbF4L0GQxSyXcyjf5Enfl+DcyWC13BoOrHNW81uPIdYEYLxuju1zsh3O
bxV783O7Spxx/sD5CzKETska1pJVjtCnVuBw/e7Az0Kak9nT3kWo92dUyQlUhtXX
CgK5sWLiYART/RC9UT81pdVL85fXwJmLUDBbi3grTtK2U95iEAQ6KyXUmXcQSATf
43FLW35FXywFLwviMQHnEGzNyZ93WeHeKtdOf1Rb42ejbHDKJbnXc3pRlaXejmm3
78JnT9CFnV6jcSxpZB8sc7qKbnCGbWlOsqpflH7YLAe/3M11keUGZ2i7zyQ1H2Nl
hr+NhcPBD3KvdCkis93gT6vTHzPAiqmxUGEz2gU3OXGBi+hdPxb95T0kD7ekyfqx
Sb7qkbapihNxbTkBGrt5fjVhQ+czRCILtqIL/KL16/0+DPQcXa8XhPBeJQdofAB7
YCmxUDjNPbGHM/2zW1gtaPMMJudWZybImSgXCSIX56l5tb6o00r4gTMUNZ0yOD0D
dgs4gOlfsCy/YqI7gJ3kKwyHvhmuwc/1WZKShReeJutDDnZm/Ao/rkn7pTEaW1JE
r+FcVgXBjLoNza3SVZElp8r2sdo2loecXJsjk4nD40MXmh6d0ORty/C4zc+XPQ6q
nDifG6lUx0nsq0auR7Ku0lpSaz2FsOcEtjxxfbLxM3aA9xFsq4LuuS3C7oyw+S/C
MXXx0NNQKi6BGS60slgRgK36b67LXqkaHwbE1wL9MyT0c1VK/glGiXeZjrkEQIjw
vHg3hKQ4BgmyorGlaM3KO/QNw6YORl6oohdF830j3fjGJKkJMN3bE95/yEMo63ND
d807jeFBYp9JaMLgCsHRbrZa++gGAG16XwqidfRkjvciqS6ho1W+PNg+a3gsZXS9
9XFvqj5Gja14GqD78kQLZ7xQ3kZEUzaifIf1ik3t06XMQCPvzVKCPI9lUHILQPa7
Y30n6A7XD9FJVng8bZai82sWLQgD6LufT2wmp90XVBtjzzIljrNnRjCVXvGMQtuN
RSJ9a1EmzeoTzyB/0R4b+X96qJzTtefuzIYbYVe5xyaIM54sIjj+224G5otlBcYh
xCWy/dPg1ms/m4grlBbHVcYL5xzqOLNSz3Vt1kGtu7fKgTcum5u2FMfCNwkc3tJc
78NvKY8756ZUI6ceT4Pr+z6fdYAEhgVG132E5t81qSTy1opoy+DjK3MEaEC50ZsH
JTzTtJGda7bMVzZCdTwNvw2iHIcqt6wkdnu3op0bgfhRMRe8fjLLksMrx4uiIyAR
veNh/q1052cgWGvLZbCM1vJZFjqFmpnADDl19El+qLoCBRKGyhwBoTxWY92vez7F
dqXZ5uZYPDLSINy1+o6STYZVuOmXTqPms6IFmAkMxcGK7x9eOoUQNS0r1HZYpH2C
gUBzfGS+3RFt1yjBHSGZ7U1nOqmZ9sFiqeKYMg77Mxhk1/wbyY7yPxw8fqB/O/CT
zNbrqW3TdxlEyKckcqMdD2E5K5Vz3Er0KGKqdJaU1CCgav5MJJl0FhAL3uZUrqT5
Fo54Ebqvt8nSESBmBu3dvfnNvhWlkHaVAXomYyL7TjFK4NLF3K+NKmV5Gz00zOR1
Y+kP/ucXE+sXKarnWNqq0QYpS+FBx4hxWB1YZshqVAaoXeJVu4Kch8l6RGKvfIBZ
Gxlehg2tP5pPyKkgci7IDgJ9UpVKGbBLCWbnuP6ZqGNvavHd7Y91Zv35Gor5LJmE
fijCmDGADA9Ql1qmC3bzXDhT+r1GS0h0MMjryOU9+6jv/1mG0etNofKV1/ajT1j2
cYHxeVs6OmEXJ1Ay3oOYfpwLkjzkLSKwYLvKhdkyV3iLAQu2tE7VgaBbDhtC3BB3
zElGkH/RCIYONmTvGO9L17/oj5dXQk/fmD+abKtt39rmbDiFMuBKQAxYrKqcFFPV
7RTaDM1jcNx+cX/CfgRA4d4ySaZUTAdOnFPBHxGr4eqqr04jGW0awzT7a5t3Hy12
4gvCtgoYreLazj6RiAOcGRh2hdtsC3Qf10FQJsqbEbrn0O0xTCQpgtYG83V5uWWP
6G2jw93W05JTOS++0gdWY31WWuW6yyRhsFngttwWpKVZJKqMGa6O4q+Bdjd3wbP7
qXRN3udhvceRhQ860UH0CMD0xJfxpQpEs25Met1b85gs47XRimgziqkNDvtyZMSE
ynTwS+tRfPCQQ7fa/TCrIMVVVcNO8h+E/X0Af9+eoWXEzLft4/hKTxKFvRGfM+Wb
T5zo9boLMcX9PTE0y5HewptDOxf9M/a1dD7L6KOQoszevwqihAZmfpQGUBCpDAmG
nvgMOWWh/ESNPVamTVRu8FSnHEIHQvT6/zq2g0vtGHutp/tQpUCyGnt4XF7Xp39B
HA9H6RrcWSvpNKOuZ7evt9DeDXborCwzXfFBAa4q9w/7i3IHcKyM2EbefiBuwjj8
6+ZQ1GjcFgBycDtbN6UAL+Y+sxTHW7SMjZvawdPn5+Flu8Evy8LUqS8e4bNvYNMA
mc6eB5OV57010OY1h3p2fPPMO0m/4gO00yDbzXDF81MEBBCybry7ixB9v6Nl+t4T
2PUpLIA30eIGD0r4ZzGYWSYZaxWo7DRCDL97avOeJrzIeDA7vWU5H2EuuUP50UqL
yZrKhD+NezT/8ixRVfndXn3k/cmXHL1kwS/hFKOYJA/yxXFvi3dRtrfFKD26n3ye
FP9g1eSy2PXyrEH9jDKdpJWGzclS9d4iwgBI4og/NfGRweicnC0uLl5JbW8Y6VMo
MNaT4s54nATC/BMOyfI99TaneoWPCQbQmGg0USW3Nk0KulihpXW7SZ7SYD3qND1p
C1BQ4T+zrx9XS8EmXXz4471Rc5Nw5EpJOoTA9GIY0aC6arK08o75y7xyGW0EpQpi
j2PkgCJtoXXgce/JXN97xZIA6Pya5FLiMN7y/4frkM4MrDvwdo2j4+330Vq4QfjD
9GfOkpZOANf7zT/HEUb5ImRv2bwy0Izhfa/3B14CgVBjjSj1WlmpoEOUw5maGzIC
JNlHFMjD0DDBEkiRHOPVYgPVApG2PpgdCvmIxU0aI0p1ipNR+rJ3txFVrdcBVoVO
uPNUXUH5q8ntxo7K1p1g1TW+UD3bRxjDPKPan9OT5EmSmbqhbTLnsN9ySuqrBr/T
bs2MjDpU6CQ0Fx66zLgQwyDPYRF/LVjwo7cASrAvdYvxAJ6HT+hdD6TX/aNZCNGm
27pqqVTS2SiUk4/hUbyuhAukHRQZtO8YpgAY1k4GZKXfGDU3uBulzG0nvT7+sbmJ
BsS+NuhEvMVlLMv9W1OdqnDXiRD8G5r59xlDlEQAKfoXpAHDowmo9iyQ5N0fL4Et
PUwqb8uFQbSeaB7g2T4XPr10lwQZHD0a3kYrZSHOGJPvKLAQfsdEjBctO79zPKj8
F/2ncOysRYTljrjKIA7ei8sZOLWDCBmXQqo1CD/uJNuVz/4M/AYAN/1KiIAyufa5
6ldmshdZgBp1/KP9Rl3uv+HLg7gk/gamvfyZVNXfsyToIDGvbIu+IhcVfMiuJcT5
QSg3B1700HLkJ+TlBd+ih2y0BIjUzMgQ0uMNWZTyTrbRQx0g7bdYQhfsfyhoQ+Cp
GXsiZT2XLCXAOx6CGSMroxbxPYK+vm4eAOM1LLwYfCDax7NoYAL4W+XNkUDqdeii
Tl7BvLLSM/2wRfibmvHGVtjrTL+Dep7e7ar4XPIe6QtTf/I4cpTpvXj3B/K8BCct
TWj1xdqqAVfZAFjMFT34J5DZt1KUvuqSM5Gr6EBHNDBAkj5Va6ux01Z0NP5xXqt/
lppAYvh8ebjmOR7TP4geJ5HXGD2ghhGdQyRX/SwnvhKamy5fCFmfCwdm2DLGxBmx
3J+C9dSF2ismhj/MCZNNthuQ/tBEXZDN1PcDt3ecjxX7j0NdPEiS6oFXjG/5pvHK
EAv3Vtd74J6FRdgiM6I+KFgajNeoyRQUM09phJEOGFi/FOQqy/eWsSLyCqle62SV
gCCXjOnIRtqA6SQ/0SdRhA8n298tSybk1+AYTJcqzUED10ZWRElAK1pg+Im/uHwS
se9hcCWqhJNW8PaBSJqsEfoUJbpv9G9cXQv4wFFt9ueEl6sqLXiQPh/WwUafLEza
bqv+x7WM6Dy00txPZ4Ci2i5E1FQH3GfHB6v+Sl3EYaIxLGh2zy5TSeYN1jz3CGdG
zIpAuBf31yEzDZY/sMduVNoR8l1tOtQJund9P79UheuA+H69ikS5Pyv9N5gtzaeS
9mD/HBvu5AJdzWd277MNE7ytX+Ruhx9OOqj9CizdX28ZZPvkGaeOWIBwaVy788oK
BtwdquDRSqMx6AZ7h/eRcgqeFds6n+PYY0yTMmOCna7o6Kli4YgN+bLGsfsf5c9q
kY4pLcLmt/Fdq3AuAClQOCiKPZ1qV7+hnaGDOy0n6T9hcJC/xbFbJa2ecqoeUCKr
ZfGgwG+lRyNrO2JrRzDKkIb4p1aKEf/2gAnt6yi8cl0tGrLsNoWAcuxco7ksB3GZ
YAEUoNyjhWEUIPsln9cswtnjwvh1MgAqsrdCUyPZNtq1ucIEdLm3B/Gj2t0SljiP
q9rj1CU8rJuLVElbHkP8ChLnIZ1xSjTkEvYk1WOBbaWLSFUlPXQd6sGMMXpmwEMh
sWEmWY8yKRMrQdO3/2D+5YczfP5WZQCqr9/sIBZRNRaJW+hqgLrWTuvuoI6FjekD
A88Yub8ouymTtRpbxiCx4uyqsQpNhFlDpZDTjTxPlpohkWq6xPJJsIcnPGjRIS7U
Ovy/VKKUWC3Z3AaQy4FlxIpITvN1GIjGF2yurgZCtL3D7qnovitVoM9Fk9moIwZf
c8k5UxaaWsYyuvbZl6qeoiJD3NXZPeWPAaV3gP33P1X5m5SQfpWnhj2uHDzt4D4K
K+cK3ZU0Nwxw5GoeVPe5FmfEmHKnZ4yQTO8Hi2vMZmh+n0a6GoFY5Nm6YcNu9bzF
TKj6K3LTgHVYZ2WTqeK6To1wt/TstTOiovYKZRZac3/j4At0I/hJXTqbGR9Byvcd
qtD9A3B/L25nnSuwzKb3gvwkKReY4Hg7hVmryYRfezvWwafV6UfozezQ2kLKQN+A
IQSsU1os31UK7MQ3bzasT/HIXqf2g+qR7QP1CefATzQ/yortD+IyS07ufT63PF0k
tGjuFNWiOkTSs5munHJUGY6exYJ9AKqT6CvK3xfEyXV3BZk8w/ipNfOocXtA4zhS
9mgMdGu51b3cJyG0AsPtOWCY9LRzl+riKIf/0E912UrjfQ0RtXCzgUA0Eazh/NKS
nIuFHEmQuKZ2SaZzMy4V2zMgMtzJAn5fxYy5ZN8eIe15Z3YpeTzcv5/w2wDWj+Zl
gg7uGX5zu9d7Hot5vmMo9YMi7vKNVEUPpv6Q61OPYrSelluYzsSyMc1uw5Leh8sO
JqXt1/SDXS3Wma4YR0pTe1G//+ZLx3ARBYEE/4jmU/BazZQfBBYITkYirN3HY1Sm
5iIV+ORong9A5ogeGn+CSVyueQuZh3aUe0Hm7eCsrt+hjmdgU0+2jXGfMP+hbRxL
tgOM3lvKRBX8wRhcq5aPAhS5BoOiXe0DDkAl4UY4HhG5FD9Hh39dYkOba2E7AeNY
t/rGCd72UebRlQEGmGO/k8ZbWGtp75Xhye+IA9iHl+jC2m7YSZi5W9B8gS6/rir8
VFdLsoISdrNaaHApUBozssI9mL6erlwonhchVjPL841oVXHM7eXuASv5nepiM3Ft
/jpVZkoQNLB7qgdppfxkketiRf7C2aaAXRttf5iFV0OGeFWQPm5MADHbWu9ehWv/
TLBAhZXwOd6cwLxXE0nEx6FuhyALTszDjSRrHUvbpESUksJYSCtpn4EPL0i4QS1q
6avljdma6ySSl4LqZs2aXSfydZX3ZrEbsJau0Y/5zoTOEqwPRwuMSEA19Y273nzZ
TRR4jWjsgQQ0vfsKdLi4eB46pI57R5qSCi6evFJW08lpa82Exdus3+IG+bXRoJmS
nBHc6y33pDFjImYHorWnrMtKnxZzfJjE7qP/16VMdaLfSYpgG7hQc4jn/rMk/F2b
WAfn14gU5XWrUQF5pLARi976u805+sdPTFCfBIlbLfYosug3KmYJM4Hq0wuCRj+G
zT4zHTN27hVMDe5GeeW/buGucMARfMRjieXvp+m1yU7SedccYypimeaDapnkidUw
zOMXKZhQw2cYXqgy4cmfmKe3sjk2pIqFeIzzghc2n8sDMiTKszW8OMo9zNI0kMnm
Y4PMnxIBYcUlQrW2P2FNo7rxkB8Ad/nVY9zAJxZJe+cW2X72W5X4KVHsNqT05NXi
NOrxMnuwjfZ/UIe7pbbmeAjquKLZNPxMgj8LwFPFZ/Z5tD3kv6n5xHxsCERt9h2f
wTTPZhvQ0Q1G9WTYB9E/xcjAx1PzPMt6BpvQUi1+Er2zOgvnisWJkOobWSex3KDj
tqgfWitAqAeb1z4fRvWlz0CrEXJT9Fp01mzRs7PctUBs766A0I59DgO6yXL4YxUV
FMLZKnl82kITEIZQkfHqZ6RvrSQ93W382wCXaErU2/Yk7pmM/WLy5528S3rZkx52
KJGpzOO8127QL7iGhX3+cagkikRTcpfu72JM63vMLR+RoBc6dxKnso4/shcKOU1a
rPvmkv8nwM4Vrq/rP2c8rEs3sXsCTRFnIHHGnCBKp/KsDMTkt8U8Y3ZxuOWEIVw2
PIaVBtp0UKrypbnBl34HqB+UwST26zbWu1UdrSAEqjpKU31R/Ef2P2AhcK5GMI9u
HeAEHF8ALcwiokdBXK++MkglSu5EzQfnOglKs0iHUsp0G2QRFFhW7JUwdKti+41+
uQAQE9lbXwjV+faOmunNTOF8dpSPr3JGYUAP7EoiYWB5njkgIOFZLbTWzq7NsEDr
XC2DZOQEpTUsp8S5g1J4k+OJIw3qX9M0e1W+ZRhJVuSGV9fChZ+fbZ95VWlDIA+x
aeWAUSoXCjqt2y1fcqqVZxY8pHcAGnNmY+2CZlKUarM4kCG2G2NdwEAvIy4GHycc
NUpxzWoSJFRYvkTXn5r5gh9nt5CvcRj+VA4DqSbe5uewNufmH2AhiDSg3+cfGO9x
OFf1DyrGAtGRpO2mu/tL9PhcbSu/wmZL8R6Q2wvLdWo6awT8oRwDlrv2FuW/siHc
/OKHDIO4XnjgGmkCoOCufTqYZFBBcNqz4NwrgnQxU8oEbgoHHa627FXqjFaIhaNp
Vz3WZTaOuguYSw3hIVcoJE+Ftk2ibWlkc8VjYTf8PqSzzsYnTL5HJbMObIpnawQg
1138GV/tZO8WkbloQOlTI0vcIrsBVgXvPb06KMiufv66m7mAxNmzq7rZVlq27eKw
PDq+rKzAYjOdgJ60npovt8DF9CvmnZ8y7xNpg5LjYvygs2gyVRynbS804ZTcYzE0
jMdgyNm5oAJzzbR9rbZgdcVQ5+PCIyi7cy3pC44UPsZinAWtoPoJ24CTLZLVNPPt
Ee+D3bThXSe9jfRw9FWd7mPg4G60VYbzdFuVddmnT6N2rnhCzfzDKc86DouO50bA
5aJn+eLM77FAUdTBNwWogE2PwE7glI7MDi8hIQLQOJ+EmKoVj12KRD5u2ZohGxj6
4JOFE+QbrcDn/1R3VheJSQr18ixPByQn2No3ww/DhBajlB6wG4zNM/oE11H8Xnxr
BClNF720RihzDRav1YFWiD6cVYjTChlg7zrolYDV/7TzsjFf4gBr7AGAGtBLafuW
DFSZAaldoq6Y5/xnmhEs+C3Nii1TwqJrWcJmEfNk5fFz+5v8/a0HSlyj7rN4iNqw
0D8pYsnoQBInXxGyIjiGmKMyUeHLf6d/NDWjCRPMqVO11OUxGLqbia8iOk1LxCGr
juHFQzr+P7fXMhZD4LB1KISchUKK4kcZPimg5RCTScXBH5aEKUWZCPvQi+tTLaLg
BRWspfzz6WXWDnB2BpZdLSaUN6dQZzVsM/OzRDegyUZUp0sxGUUJGVuPAN7/x+TV
3nLH5vri9DhAHt9/AvMqBK9nixqu0cQmpn1S6OWCQZw/RYQOIu55KtdsSoniNde/
vNVoXn7n5+R0IAEnttndKqVviN2aU3/xSsHoZ60CcCJHYv57VOyhDluDkRwb8Fon
wj9CibRqn4gQdwG3eiU/l2AHDcXFZgMY02jtb/e4xiB8mXFdCui0+dWgFcimzJs9
ppdJ1pEwd7vsvjXa95cxiiZz/uTNSqm166rICb6zU6mAqtoFMs4kA9UFlW18XIjM
cNuTa65zK2mdHHrpX+ocQ//cw2yAmOu11tSDD/TDVi14LCPuBMN7LfC2D+tM6yif
GT5i+7YbNK5OBEsa8p5HviOI1yyGpliwigea1gMEH9Mkwbh0oO3xRfU6MaiOHxK+
6w9/M/Z7zbOUCUvDQCzPCWstX2FyW6vidq5HIaHjwtCyr06bLdzKO/5+GFZRk9lk
XPRJhjDRoQtrCGuwyt6ZvBQ37YLMAU/SOQAN0u5GQ3d6/aKF1RBWaW5guoapnea/
sQrbuoTpoxtL3jgrsu5svxEmvanAkiVDjZvNbInXeEpGaZQFh5+v9D1mf44mT6TV
9nFgwqRqW5yr+yxZ3MmSJAM4v1HaFvqAOPB4zvgl79cwr9oXu5dgLZieIhGZEzkh
YdL2DrgSobcjLtGllJu0uxpH3E4hFtewFdwWXwMAZLpSkhnX8AL4vJpUuSITfgB+
WjOqtbpUgM6457m2s9v5rqGt6NLFzt1oQfVkG8yiuqhqreaJ1u8SUY/G7Mf7UTsR
YSWWJzYJ2QPQsidFVt1EkQXazkGnaC4/3fnREi69OxxFv8uT+TeLY+MkFQyWQitC
p6ms6lw/P+4l2t5Wji59+YCihS0OV0IZdZFwddVJitAHgE6iupQHzxgbKpXFh1RK
6KK63e7qG9dMhvj1zWYtIft1tgWHOAdOP7jdrVsbAbU49zGOS7z14hkC/tXOdge4
K1aVBtO9+BpUjMC4v97blUYMMex+GJv61TkAIjiuXG9d3D1wqEhh+5cb68rGUVVU
65vg29SCBc5xNKUBYtxQ2Gplm5E3jeTh1UkzCKJimX0z1VWra8vDE6RYjnEoxYSr
5df0ntsMndjSnfq9QrGYkWuZRS4U8Jr8zWrU2AOoRTy3kwBvE/8tBI5kpoMj8joT
L0ljq3eTa6ldDk4FDWKRX/369V4OthMDWGDOsI884952peRo1TB11Jt+zQasL3vn
CDbPjQKB8MT1E36cVaYQf04aNmQaYKWGr3LaGVJHr32hekEZojZKMPVMHt47oKTO
tvR83EJGcdO/xCqxtueSnxrJCBFKmthPWjQLHdd4Y5IfcRDqo29Su4szf1dGIL9N
L+WodBogD8Zj2rMmXezrC2GYoDRKhcMGLpEENmtlJ/+OSdJKP3fYcFbQfMmdYb3r
dLn96aQ9PRBu+whYj5npC5IqFVP7GERjNtLISTgDWBh0Aj8xt2yM9FFlmxLPMeBf
CklTwo8X4MYP7ccpKbYbUnIFwMfoTIM33qWOEzL7EnqCKWtI/kTrb7sAUQIPwx6m
vdFmut3iV7Dr/bVUsQ5j9bYFPWeXMvvElghMZAutPwzic+eX1xhs0BzOJ5xkFMua
ErLM8D8UuVx1dqnjp0b1CK8ACIUeIt7bCGcYQvVYDPQqwIpqdDBXmLci0KkeLs/X
yzcv3j7NWhLYO5gZ5P5SFjtMdLR6IDoueWarT0GGkf0ZqWOVKdzw/NucaKjEZyH9
g98qplnBSWRsGmhnA0TYgHFupIM5vQUkFiDy4FwjbFIVThMCGLjKUEqtYQDZhmn3
/za04Cw3UJLvxMhStFb9Vn+v9Xy/7llqQ5g/x0S+bOO5t0uUEzJhDWspZ6BVOKU/
u5x3oBjVu7k5jrMQ3G79YaBMf8k++FqT6LiqutYWzCOsRVIJiN9Wv3WBaH5xJht+
mXir9A1UOSsrg6ljADcFGaDxRMbh0/+C8PY/ajAOnVP3qYUY/rt7dnafjrAQiDb0
KVbRUpCP44jlPb35gc52XchhgArKxEL3mEjoPmJUQsb6cfjie8y6Vh9IQxM8jTY3
SRo4CeK2TCdrp3+20pcGuTpCv9y/u1A3MXpkeOYAKc4dz3gaHDaXSyguwqk1Arb3
60sq6X9XVkH9OemOW9mj3eFVp7ZU8tok11eSLfE6N1zft1gTEXNZ0iQjO8GPasOs
ihogjkmE6kQlUlshy6t++aC013x4t0km20keTrxS6QLgNhSkmVVxAg0lZi32RmWZ
gHwIbzfWKbDNZPS7fmRW7uAp/+M60jUhbVCXkeRn6VQaIIbsJc0fsKGeIPZ/cQLE
Z8FdaeJERcYGmNtNFE8aVmwuicO+Z1WZda+q5nwHlGiVpgwadRdNL/tRk1uOHXYx
RwGBfflArinbHIgZyl5y0yi7JH0i8HcZjTnc1HOqdti2NQcqJOeKCoH0ZtCKxqqM
OopFBdIUHTdDPhaSBJMplJsCIpKX7Hcq8OWNwcgZcVH2qa06j9gWl3c3iTqa+Xlv
9CYN2bgRqirJ5caG0wv5daT69jaocketzjIwggKaIYVI/+uJmrqJYRMCjanaIkBC
Gtpi5Ef8oqh8adpKgPH5PS67m+aWw3s2iyQ0F84BG9YJGY2+8GbMu6Rc4yhtJFq9
Hv3/41sMTITb6WF+30KFOsfHCsA3R3iN+orLmTVca2cNEW/735YldWHupL7pgGjn
fa9jevJ+YkoJQZX+A1PVOu7Dlvb4tv4dUofqYnXSRwtVyJlUnyFihl9j+eVo+OZB
LjdsD1pSwodvMrvwwC969mNo+VJeZ1ATF1bPsH9bwwjhXP9ZbQpnjCKez7kZ9+5I
4MfmFe8uqw1niTUmXd6k5PvCajnovsXp42aHmCQqJH+GC4WqqmcpcMxy1pL4KS4n
CZCmdOj7AjSm5d8rU5JN/f0CkPpMsBHgOK2krtha/z4PPkkeeKXr6AKln/6mg/6k
TxlnNHnRKSRfKyt5d//PrUIJBmnuZMBOd7Xr5wv5nj5SG0m1oG2N5lhL0QQq+5Ts
G6GjHwco7z1Oxs8qjweiXK9nvpnxsKVD1wRjAidkOnH7loz7O6SyCadeyel4amlu
+wbp93tsro6Rl9/sAdUKf8FWn+nhE+SSDiytBaEKj15QW+lX7nz88K57GJsHnchk
23t0nembf7rIsLd9zET8uSN1yALENubErLxSOTNOMpf62nMMJ4b1IqDxtk8v970n
ICC1B88HaKwg1azrNb9BGcSe2TGI5j/V1d4u5mV3E3M86DHvkMDuJs6utHPfWwIJ
ButUkBPod6hUAaLHuPrhpKoLMZ2X/WhOEd6SMs9teEiUhTsWLqfYTl993WRSDtof
l8WI/NmILM8eSIlI7OBgMEK4ejqtfY6//Xc80XrnD0xbgSukYcgxwhRA8FNxQHHa
9M6v68VHGKMkQi01fWq5ypxj9Db1lrQidiyrwNGRLljsePvnNU7otcs8+8J0qrvr
pg5vB2rmgOkqKhwo4wmdAnKmeK6Fkik5pBfqtWITdYoJOKdl4pdtw/I8h0IZWGr+
Ddf9+r2gEhcaJifl+oVzPfVmebWW2ySpj1h6I+6UO1tNbn302T8HVfgwzZWZPWHW
j2hQBzVwvVufyTiofruSc/iRQZsM0AkM591iFiRIKeVqTjL/D7NXRUCE2AbCqXIg
oBJgaIR4QQIavOPj15IxnPEw7e345QDvAJUm3x1DAJZgA4JscbQc/tkGElaW150g
Z3veH2xrI6JedQmzjQE1O3xK/2cw5xlkY1GzgF6kBSpyZEF7j8kiugk9Tcao1Tot
TjjP6qQWWfJq6Bi6BFpJFD85YUmbD1lYeGqhBS2Ic6HCucWsNYdM94Ic9EKlrQA8
gaBac8lYPgy4i1zoT/x2d6gpdiuF7IwAy0nrRZETaszINBgObmaBEykwVEvMCBFL
z5vAG+noEU8hYpeP1uPr+zx+7NIr6m7pit1pMXlEhwgctSVBbJIC7U2JQ6vFU8b+
bzU2/dtvPzKCqOS9hyxP5bMwnYdKiK3kMeq7epqWerxu+YR9OsrsT6kw/NWZRjPz
NnJ0ptFUItUqnU/1UeD+euL752B2LY9Q3QbIJo/O8rlOK3wn/hR3Gao3Yxhk629d
wYKa/qHEMommJjmTMm+dEfKfWdCKzAxRbvf1saAhSiudqDmbU/WikCz52QV16D0O
RgBCn2qycdBlE/vfSQqN2l4pb9cYMUemoRltBzEx/QXvLmX5DiNXAw9hIgf+jTRL
OA0vI8uWM4e6pxx9dXGCuO4pjCFXAWNNmc5PfnDrJW4xdgoDIgQl4fdpjemU76Fs
fy/oRFd1i/3AqEr9mMkmHtEpBDCzYDPk53Kp2RZPDWqhhsZzzSkH4HLwMQQy5i3X
2YFabYfnGklWP3qQjLfB0og4jKXKEODAuSDvOpJiBRwF6oVIOQqDngb30wh2Vc14
hjpB6XKo8vg8WqZlOuQXAKYgF/KjU8mt1ij2dDPFMFUovkBo6aroOpSADLypLGyV
wT/OAKiX0ebH7ckvh8Uhue8FkK11Q6Ol0bA85sj3e8dSIZOcZPPqK7q5fDyyibg/
LuSmb8s3Pmo9TosH6Sq7Y/M81Mp4Ryl3L65Z3FHBkV14u7SgFm4RVwxBArkIa5fD
TDy/FZ6NexJ4fKKNOHBDNLorUjd8g//LV49fFkdNVRm7m0AJDkfb+sHcNlfd2q8F
sMFxcj87GAGEhGIrtY3A4lWIxOdgZuO4FQbTtA6zMkhUtmBorEK0SDkmWZS6JF93
fZMagaV0wazHdQXiEUP5XaDajeNnGU+DXkTdpw7w4pttHpvb/LQFcGIDt/bPtOF/
vffom9ZvYRfkWBiri9m9kwv1WRyJHgpl59FNjmF8ZPu1J8ybMjPV/BBWdNL42IQ/
OE0Lj/szbI7L6WGTY83CQQUJW1tvUBvnrs/gU2cP0OpljosfixLtg/xM1hLQb2q9
RaRFPPNWjbaFijukphfuEAqDI03lozKue4XfzSGRFpH0DZV7JiqZ5AJ1y6HjyiGC
iCDFllk04jxEeVoiD0CRSrAz9oHcqDDndhd7FAldSfruyQROZQG/WQV/F75A+ZON
KKIS+bJx7Bu2SUmxE2CXp8CPTJ/DrmJ2mvnOUZR5W04dPN5m1Z2PLPDmOStvjcSF
Cr2Aj4sRZ5dv+Bq0RjRWHLqWKWOYrvfpwd+VHvKHTHfE/lTrfpJNbuae/5jNt5St
sljIKIli+QJ1+IY6Xcc+p2A7rRbPLht58VB7Bp9JoQRl52CpE3RvHMRQ4fxoQc+h
pqYVtqYk9drrjUjMBh1sMOyRz0dDHDYpJeftE1n6onHRKvC+qY6SsNFpoMYFBujT
Y23tDne3UvGUBDyvk5r8fW/bH0db94pPjxmK9A7q/hs/w9yVH4a343XJvMc/J0co
X/Ca9XwHTk0IVNlTJQ4Z+s0jyvXUXMyK1RJEGmPx5RO3s0etphHQMQ3NdQX77ahB
P4A979Zy8KAAgrf9A9QV1oWagJgXHVvcaFuub3M2gDpGpZ4Hz4lbXo5I04t7+xeV
TdMUNzfjBwy3/YdfNIP2hivWMu7JEVeUatuA4LvOhJuLyJpbHCtACJbWJXo8f5JD
dorCcgO9tx2VyfnDzvbA+mlHdvAoZxATiqNapk/hi63dW9tScP44XgrTNzKp3ZGv
+rZODbnNGqUA9utjTWY7+HuANds+p6MTQ88sHUoBPKRVZwYqhnaPF2jNxC9h7091
WMu68OgnG3qgpJdBhxdZ+GEzsbSKtGoZy8btA6GH0R/m1SqUccsdFjKksDFHr8Dz
Rlotc/Ab8fU4E/E+ABhctCiBMFuYZGsTe38cxde6ptpjgIy6fV7rChfeowz5PQbb
5jF3R/wdMdEH5arHrrvWjkF1u72TtUUpSjz1QNruJEKkZLJLsRqFZu7p9ZHW346s
fwigb2mGHuIUWqqTAcHGjSdTZAC60kYaS9ry/czRwGG8gIztEWDGkZoIUZ/Dah7l
4eFXQ85fJwL1Dc7iFrLU6TQ4LHd+iX8qhVVVW0C7DbNYgj0EcM228Qe6cpqXKGVo
HHYywzl7giBe1lUaaMAjI+2S34z2k7MGUCjglPDW1UCyZEdpKQUh1/bkE9KBlnge
cyX9RmF4S5i6elopqjU2I/hzV0nCQwEF/zMadccVVz6vkoI5+Opyn1v3gcCxkPqq
Et9q0IjB0inGpHWEL5qrDRBPN9714gLqsJpw1ZccQmn+9eFR6MxniRL8haS/TKUX
anDuNBF0RrXMhr6rMDY1hW3VMGgl1eXB6/82Xatq57tvHt/bFY5pg39F+ZL2dgx4
h7jBRJU8fNhiK4XXZzoCyHp1O8qap1vk3bs1LcirX0fACpkaxvcKpgwHDlH/Rp/G
t8+TuoL5L6lkUkUIFevYlP+idBTZauGzifPmhe9k/Df6lKpt1wKRyP2gfK5jovLL
YKk0F+hfmVFKZQwxftQxUuCnGlXmDCJLFl5cQ1z4Pmybf37WokjRQezRJJJ4h/LV
eiLSpCzhqtPTZWOgpu0vN/d4k3SQGn/Fqz2EzjkLhrm+RbZLBksnpMhrE2HvU3cg
qZ1d3GFcFedfmdQJ02Hi5L0mQEFsEYKDNz8XnJIywCOr3k3CmA6uS9O7t8XUddBj
5Sl9dB+0Vl0NVq4cgiVqpHjUBcektBX3HACkZgGJuYClQsFj0oXeDLU5C0NnDSTt
nMmKnd7UZHsg9WDWwaD17Ka+girbkae5+FgHIWQYqH2FjwThHeDP5oYA00iJ97aL
0JPtPuRv8oHcnhiGR+27wOc7SC/oXro6TITRBtXYnCEJb6Ucq8Iehd0bkzG2RcTZ
kmvxq1YstowORPG/Sb9qL5TbzVbRN8VV6MNG+nXBgiZfvXCazmg6RxruI3oYk/Em
3odJgihnK7ttaXD8jM+nDZNwWs1loqfd8s5q26dEdWAYmTJUO4sTnrRcHN+I1UMw
wVlMqMu2BLBDcQZ6piX06dYEVukmO5nMa7v1si2OUo9aos05QdiEXmkutyVaRaeL
+QkY6L6q3jfSfFIxvxl0XqaqA3rnMVQlwJFNJbybQCeopddsMkV71CtKKDpm5MZt
V7yVqwYzBsbXyNhg3EBKBKArV3Cj+Aq+sbu/84Ctbt4cH/RCN3s31kwVGCdVZMKa
Txf8JDtaLl+uYCBPRZHD+dh1mUnHDKmDJveTAeY/o5nCI/TZuRU9MDJaVu7Qr4Ww
mqkoFHNVN5fLlmph2DbisdOLqk/F0n1bUpTNcd0VUp6QQofYas75OiJ+35Tvaulo
puk5JmPcEtrlWULV/bPkNQPngJ5XtvzQaeW51cCaIuzPccsEoWcIt5Qo4Xima43F
9wTUStsiA66Co3/Nk8EawuO0faqV4uY55G0myOXRenbdPcnYpO3+xSgwfy+i/nXi
80ocmZ4DH+F6gXQi1KGfvOGUR19/nNszvN42rLumd5U05AscrP0vUn2F+k3omHXX
+/+uhgHXKLkU+0N06zAZ/w78Efsrq0Guue8gHI+VN7s2ljlrDItrvDVvmTzNqwx9
22moYQORJB6imXHKuEpjIx0ihsOFoqeYQ5QI+iFLt7g/53v45/4ZuwlMBTEmNaOB
yYzdqUU8gM3DkgaJerFCQpe+P/DzNohoiR8rCOsHCRIFM53XDN+/nVQjp78RHSNk
R/PYZQSQ/ld/VaYh4mMo2HdgdQ/+4eFqMpxAUtyTWvSl3bxQSU/IfSsjwL8RUqDB
v2UUwMgt2kmjzOnKpT5zpKZkne9CanizYNMs3Oecdinp6TqWRIlU51sACSlvXbFq
0GzAHV0LINd8eNs9ReS41pZhWqmT+/D7RAVgVf9UTfAewlR601pxY0a7GzIlsF/D
HGgwIHyf8vocd4lowSL6n9pCOfg0U8QlsCBgMzUL2qJPTNyhBNcNXvXTgjkkpRLJ
zH7eW73MwC8m/1SfuXErQ+8uburCsKocv51WkHLb5X8qCJieivKBY01ygIqhEDTC
kpBrrOax+sUzqtQ0xnvVPhemYbNhSTE6EnuF4BhCBDwEK2dpGkxzLs3jxG2Nfh4+
cTtxnlkmReNAZlnaBejTYZYEBQ3cMtglmTt9/k3org6AcNlqkaCJz2ITu0SZrZgv
gbsuEBr0GtLQ61PBTpSarOqPDXFd30p36yKEU+OABxOmjfh42KUJyx48u7bPu1SK
NaA15jcW/327vG0vSUkuLSkTJoaVpr6vf2jQ1tZbKTha3xmZ/wFDjIAasWoTT/HI
VgpXLkre92QdLmk1z9+gozfS7g6JUZ+3V5brnEmx+dr2da234z7GDHrJVsW+Otgp
FcTi46B85XfeP7iJxfFVvhrA4ZiV4NkMC0th0JqzHbh7NGKnDdSDDocPzGvQFMCa
QZ53VPCaC6lgcbFVr9mEsUHK/mBt9seNuTrlabziUwpnRgCQQ3/tRCRzraDForhl
mt6NRdM2sxMScPUbhsuxk3uQc9V7iHFAZuY57BexL9DT/8YvENRaMbThOJPeMvDh
VYiOCrL1FZQqI3mOVzBE5f9sJJY6DeTsG9JgXKEpaEmbRwcuWYnYInuIPGz13fup
nv5Wgu1tVv0uBbGpNp6NIB6fvDS7k/AFEeUDzekXxJSeLb96tcgDT7CYdZdeVXg4
Ac/VTd3mBe6UJzrgVSloKCijndSxAL3940A+sw4qWIQ5kSAeTMOeKp43zOHIOdoW
KLrPv3lCelKGk/v2Bzt32ZOQomlhe37esatMTknraw6ANbYSNRMco522LCtUdo0U
CDvEY5YGffwQIMhtGQaUOrdvWDoHO+aKrBFNpfBvgMxOl7FZbkhJZ2OjoePNw0Dm
ffT5PEvcSeVVUJ5JH6hjsKJVsYTWetMOSpFQzYrKJ0pi39OPXpDZ2Yo2pYVEIFCw
pgLydBI78POvc5ZgyBdLDJmg4FBsdH6fOjubXhgL9oEu79LEqBLRJU6zZnxbbN4a
tF0raM7ngolTlJ7cQm7xpxJFHPPQebkbQwyMQKIOwtMnTlHC2RLjvoZVRD3TZZpd
1xMBTu5wf1N12MKEZYng+ziOw/6XS6e3/0xsnK63V3/T64Rb+6g0IHTuoQO4BUS+
ViRYMVBgExXuDFePRcQCgoJxw/E+Sn1tmD6wKuS+Bq9hW96yX8M+0L8s7pKT/qe9
96XpYcLruzwpzaF7TDmwpY/YwtMafFfycNpiLFIuLFm8s55s6ikQodx16JW46rM5
NYZ+r9ljEUlnyMHKBWW/W+RaPscvjril8tgLcTQwcfOBz7YMfjvNypRKQdHl6z1A
OeRkGWHlD4EyNfrwhQ+ajqU8vrVRzF1NGVYV/NJlm8W/9APgSEKLHXe60++Gydft
a8KMSWpwzMUoiTmkoxccAcXZJmAPSPVAU5dPzfcD7Ov5PVdrbD3zDnSqAonUR2er
KpPXlCcocEo8N5sd6syqZtmjc2pv1G8j/Nqgjs6xB59guji6taOwPmhPZauZvvWT
jWMy6MHWb3/SVMdAe8AfAimWjImwKwL/g+dMM8Jxizc0H8kVwSYzQUUfV0eA4Kod
dS0EO47B16RgziSYzOaSCBjo6L4SB3yWyMN7Qq+XcsilZTj92qdEMp2YiLm1vI4P
bwUfuCrxS3mi9FS63YtNohMNS35EjkLw4uJ+Eua4LXRI77H/nKEcILgFu4hYkctD
EpsngBaFFxrRTa06QYuO0Vq2zhyNJjFiOtP8yCLy6XF4+o8g5E/OYv4d3IhtyA9n
axVi8pUkshq0tr64gYh9+mAa+fKcxL8oRVdbdCPwYEU7ffESer+QIs/TRBB09kBA
odZIyiZNglaw7NxwUlPAP0Hke8lGHG9NhYQisAPtYTMK1b68zs78ONt9WLu+Zlao
AFFE9MGpZiy42S9vPNRtOUDUnUkid29p1nmVKEKCyUuOwqo+q+8jOKSdD1UAGCLs
MmYrWl4ECSSfVpBFBBfapArDASRkTd0yarbIJ5idYq0A8z0vU0n5oCnzSz/yQ39k
GQgLN4nsuVSdY79uIdXyGfUl7afyxefaoIr46yT7/ia/s0JNFm2MmCDPSQmC7x9y
SnWpAODLI+amy/shRV62ropxE1mkDTAaC4drf0YgX+PUr3EcdEQu6GzTns5RAi4w
c+Hu4PI17ZOd/XR/RROpsmMsPYfi3KfSMuFpOaxjFTLoJb8Rt1lqAJegn3B7smRY
l5xecibein2+lNb7CovPgu2vuBq8qpe4ugKEjNv+Z1LMmTTobLlf+TzHjvw1kxdM
AqmI7MGA0RC1EcGltJDfzLMH1a+xiNAdLJrN76GaUfgXcazgWALjbhRX42yFa3B3
8sVSWIoeoSOBPgcWpkYvQQDvJOMbK+Eqql1Kj5karUxwuB0uoGaiixkT/5a/ClL7
7d1JbdrMCybBiWaK9ZvD5FfMWaBleGSRixlbN1HekYwLL1mx4rc1Ie8dQ7EtY4Ja
NiMsHeCN3+B0N//AA2sv8QFVo0VwyvUDJruGFxV8XyTttS0GUp50ETWunhyef4Ag
/ngokGABeOmY9iv+h6IMi1ZXhr/P8rga9FKs6jwAdazXCW1HMJCcw5Pdcng/YQzX
G4z3vQogqpGX5muL3TtFTfiAcdkWdLcrMcfpDe+Ocql8bk763scI1y1y6O/3aqQ+
ez3VyMHYpDhqjYq2Ol00O/JSunkSMHSp9z7rrimgRM9ChryGVKC5LjBWsnulqX24
ZjfmHdY9wt4wH5y8Vj+eNrCm5zBj2Bupc0bwCRXCRXdfH9nS+5+7SR1nacd1sDMF
er4NeR9AvujhPV6j19xYdgUiaMas9k/pb/gPRwsebSg4YRglv1VxJWGl/ZV142W3
gI5xTE0Bp5tCpPNUJCE0069i4XrcYTtkZ23jfsRRbCpjujYjM3ED0eyj+LTEXA6a
MZtaYIoxi3fZP+OFVS7+jBMaNer6zR8NRY7LzjWKt9Z/Wf2NpISDij1q2sJqNa/4
tOPEVruxaKDDerYbqI1MolZMzc8rEmZY73b+Nt6q3scFRKXbDtZXrtxf1L5ZaADG
TNsRwDvIw4T6JNomyMDAk+PUdZ4yBivQO2PAT95+gerX1D8dJn31eIQ5Ur+xxIyc
4mzA3OJA0CUyeeroMEEAyUP0ivXO5rSHTaMUUWdl66ICFo+87DxcxnPWn45Pk2qX
8VpCRW+7zpWlm96A0aErCgGpIQeW5MvlhrhcKk6v7cc7KtgwQxyjL0t8AQZJdZg7
1gKZUcRLjG1LY1EKFAl1tm7flc82gqa//mciwn4eAqur9G4XR1uCBFbFknjNw3dv
KmB4WKa4NsV45C/cQ30MhUfkOkhJqq/X3D/NCYB0OPsrzvq/evsF048+vwPYseIZ
UX262CXI20HGlQTdI7c5r79ZMtToDLAzTQjQjSeXGYMrO+W0oeBpR63d9Uxv4rAQ
oiobkpAitA16uNRJzwjoEbqATdKbVx0AnJlb7DoEbT3y2ybCPiKhZcsqqg1u0RlR
NlFUtp0EF8zqR6Wrn2+VMpBoCG9o3OyqBa6msRwH7Cb9drkMyC1wIFRija1jf9jx
OEbYXOq2YZS80DdJ/n36bYbiU15FAEdtXkeeyHpMVvGfgRStI2mNkjddRZFuPIo5
0O0Wwsrq9Udma9EZGF8DajeqC0aZ1m7FOieflL4V48sHqH/YRUpuhVs1lAi2RZp9
LMZk4zNUZYlXW9n3tieSkwdjeC8U4GdXYZVgUd3F5VZJrO7fm1H0uY4ppeGYepGz
bkmJOgU5YwegchXgPfeyeq1vqsPB3zrzuIls1k1X+RofL5AhB3AxjqYnDQgTMRTk
TjGQQTPwwy/8UfHkR4lWwmWvBg2LF3vSg0pG1MJPHanxmWAuxVIUr3Bnj1pdTOBj
lI/8BrivXpXv7dSy5+/4OHRnxWM9gVzedQUR/hjjtB1qbUomMwsBul87KbxxD6i+
uuYjfihIcPBLn48BCDWNfiujb8HHYiJTAtsBFt+njqYQ/5UNbnMKyEdlEXD44/mM
Dyhhe4Vre+1p/1Vpu3FkeSPUckxmj02SRT/mEPkutxA60gEL7XKom3CxaMONf4R6
wG8PYelpdsLPrqLaYjBl2tlTd0oSYp6FywcS5elyYTwzOzLVLxL0cPWZSWZ4Q5X0
GVRxPnQHRHD64cgVe2k+PJn71olDhPJYYed4nD/Cr7LDidfVjbg5HMhIqPKef+r0
x8UKeQ/4nODFstDs6vmIg5omsxq+WYHWGVg8FVmpgAkFxse0uEa0fK3SaxJpeUpp
ecaFyYe7AB+6oNwoACDwFWUE/8zoiNb2PrHCfvu9DazluNdhzVLPZQiJXR5meKYd
UOtgS/9ux3XkEdGUnGnKLug5CvKLBX7XRrcgoJdM4KFRQ80NotnvOH3aPI6Cz0sw
ZEfali/YgBFpZrv7aJlV87nWD7gVWVQoLLOR9VPboP6VqFH1eHZRCzpXNpYgv9SS
aATvkpCYNHnR1twQMZ/3rXj1klOFyffvNkuxN/KUQaBJtr4YLO0C7k9HGJBAhuax
c20FyK0GCoU9uI9uQBnwUxp2ETTiBmOvrpN1oqhx6TJZisfIWxKybGo+MSVRINjf
iISat4i4LM9Jdd1WCA2PbD0PKrflKU0gKY5JlhlC44xB/j6XGcOBBscpKN9+lrQw
78zoDnywf0l3sQ25j2PlBxgzYBeFPN0Z0e0JbkjWO7+cp3cXU0ucZcjC2cvpgieO
G1PaQuzvwlr8AaWCLHmr25lLk8IZooonVb0Ht+QfFLuPZAf2yXvFFVHYI+mm9LSk
ck78uS3JcHnAevPOlN9JtfQ22a1YPmU7jDlz1KuDSHumR47GJvU3anLh/P9qTnSg
B8TJmEI7uZDgDbamJPruezMzbIefdXVrSDGIRIh8uYC9yZTxGu7tbCEl9gOrgo1V
MuTRTCiNsMhmbX7bPT9PSUTlPTT+8QO2ZhnYT9whO4D5iGKcg+/c/pf8o4yqp1aa
9XJn0ohB6mRQ4jbXfLblkFvejCUfD6QMXpdoEcpA2n+6VrphtKitK5uZzXtEjw5F
p/Cw/paUS4e85gUDEYXsXI+baXJ2AEk7bd2g9CFiABujetawvwh3CMZAsg4u4uNQ
fnfVLC3WgXan5hsIrS1v8KckdJTvipKUzgOCYHoDarR04DNARFY5iXf1VDaxdFxE
pweR8pUkpNhVs5CqODV6hNlONJDFQmyeZg+kxu3eISMrvhAGwBli1bPsmkB4YMS8
ObOKKBThasfeWfgv8hC5GBcvWvmCah4IlUamrk0+LcNZuXZwEDEWPL5CxHEMJXF/
3jNOMRNahPfzMAmrqtJ9bjQvTE9x6YOHPKTB7TxZm+t8+pDVn2PmWLAksu4+R4Oq
esQTLQThK4io9EU8G+myJ/3EAjKgK7xDvhaASiDMkVmRz8Dv9t4ZmoBn6m+9EVfJ
p7d5auyGaXOFKQBvELKLsfz3Iuz7zS7MXm0jyn+UeIgpgLtZ4w/pZbPXFQ4LbUb4
6ORvZXsgTkl8CcQ0T3kcsgYwPuY+ws7IttbqnX15TM4pJn4a7+JmmaqErhTI67VH
CDVaawpPuK6nSFbUr6fbr63r9yT5ObJUsjnl5oUq5GXaV+YvAuK6OwP9PjjRn2SY
qxUsMNJLnr/LHiw+7V91P1iFglh/LbOp6DLBwnqUQh+pPQ7st9kDY3srLb4ROTKx
vs2lYQzY+quii53UnmGbUNY4GH0VMnmVIis8785fIweVr09TF8kGM0mZxuDa2Ed9
lAg1RJoDrl45Xbh9/sdNeFROnjgGQncTossihW7nEbsXDn2OnGZdDNQesoja/ynw
wHepN38Bofcpvga1gUY2D4UNFv3j/gMA5PgFMNvPN9D6eJnjnikS9ikSFAfbiuNh
b2x6d42yBcGmxn+IQl2S7y0chMeP6tIFdyki39nlNEr39xXuOSFneJmvZTeTiks3
mDLvGJp1ZXk42mllgY1yGAUtD8PrVrZAWqa5OG6GJ6i+IL3hvp3t0snP66Jt9jfy
43tTRB1iPWWWMHOhYHYMdWz6E9Kh/EunZ1Er+m3dEvoGTsZ91FzYVq+OznsiRcBt
lNkhoNaXSwd9ec/AqBBPmQ7RcEP6yrpPtOieAbrIeQIDlVQ+qi9ESDn2U7xRBfyl
Vo0GbAULM3baUugQFI/rIJBMMLSJQtxRsH1yeb/D7ldLXLUjSUoyqi23ABBddxRE
vX6fAzkIuUKdybYu+p7mGrEN1XNoObXb9gmexExrAxAyXVssC9kScuRRBzEUylUv
AWu7j2bwnwqI4T6/5h/fz6EsnEUd8hZUGVAYBZObdHkG3XwvdCl0VeA5DxpAZfd3
VJfjOnwNPTJplfbqoPQA5MobY+SeRz4rROsStZHR5RK93mvXAqQJeU2/OiQwDgsr
QzyiyWw4aOiFEzdPPXDFyLbnEb1wEcNCHivRbAMrqPyJSoRP0bLI/NdnAWBXwdL5
cj9p6bYJzeuc+b86UVwPsb/k1IE49Gnk1RN9Gop4Nlz0Zk8ded9UlvGFDw5Lj9z9
8BZROxjrykmN6O2ptTJLrtMqFcfmXNogdEudTWV19y8WLvsuEIFNmxVqzHlyZu1m
/bAxhccULiBQaDrwxTbBeI4haaZKsy8v3y0QnIT8/B3zGxVP8KIkuOOlbQZxplhv
PE8Ht1CKrw/jMGVu+GBtJUPEB3HQEhy04YF2D+Dd/drCWEyVgYzhWXRy4ALJEnwT
JvoFOPF0Xvft4/nSYSTabzTyBJkiC0c7bJeURT/04hs5MMdskwAzRCpuQkCRXadO
xunhgCeaXDskip7sp2f6AMC1ITUpvv6GeYDbf9SiLJ0X0PY1ONlLfZEfMIwNb5XK
jwYYAKuNCc/IJdLe+pVAM3RYkN5uPRSwb8TYT+bOW3sDULxOI4BCAlHLIvZtnsd8
9TTcLPdBStm0SObuUUVnA3UyS5CZNkJ57YX+cdPhaxJA67zTd14TZbmm53KHUx8L
s3FvJWo/bP6bwZ6f8mlJp03Bu0RlJVRdpJlLWnHbKLCJfffbGno4bJmouePvr2Qd
WVyfCIMzqZ8KS+bFm31ivgT0r/8K9v4hI4Pdyk+7+fKV3v+jTI/l8dbgMlAG55SL
7w4waMMUbabPnClrgNgFqqUhVXUitD6ZOkYxHCTWTFvjAWhUzeKncAe18eFOrocc
JSfM/Yma9nTF8PBtoaTlnxDmJDGnA56c+kYsmifMSWbVQIQuWKCT6x0cBIOopiEr
tfIyvq+pXS61OPvWdQWHZ4pRZPTs1iBhAloCoOtN0WF/mUI+AI50dncxmFzW4Gve
hqye2x/tTCv1vBIJYwpGdiaK+fVYnOr2Wb3TaN/xHIpWLs3NBsLeRYjefD327+nI
vzcsBYnTS02OGODtTWlmflhZe8Ot/aN3JPLX4CoLI3uIImXQaRRtJWotmw0pG9iA
/WdnN+ppLxW3tg7O1vVrm5xkNbTrj7ntkJN6Gyw+n+ggDcFDE9HDt49RP6qtflO5
n/OtvH275NPNMk+Ph10fQUL6AYq0cwrUmWBt8NAc6xliPbCFDU4gXFTgTR+cLqFC
n6peaw2Rw/+QnvzjzUuhM+M9bAbDApA3HEbcuLa0rL8pxvl0vwAAEU65b4l86z+s
41qMCIDjgjSEN3ypwMcMDbIdtkNyuaxRMPcvvHPA+cznFJUb6t9ryycQSRVD6mSp
PwLAoJicJXkeGDJsPAHVyqwjmnmcoAY46rJ7NmbOKHRpQ2Xynj+H5sDJqJMkSANq
9XrZR4eQs+Y8juSAJbw94N8qpoHP4+yJM1Saxml9wBKsC3CyeES6I+JbmWuych6u
d9yyhc3BKfIKWCAUPkAfiutzVd3Hqmu8PJLmutokGqb6mwtgCAd8z4Du7C1cz571
+sR8aXotW7w3GI9FVTpDVcrvLrhj7I0YbEVa+5u4oVK8oOGJzQcH5T5TYseAvWC/
48Eb2kZph4HpJ17KY7j+1D7+ntW3puXzj8dKFA12rKQ0Vu2MjzWQkqJVHokqvrX/
794h88RszhhHH78sMd7I8FOAcTo6bwKhiLsILsUR5HrneyU982Wckp439jHkT64B
ALHlRzgIuQhYgG9IFj9/9BK/8AfIYMOtIBVPc68VgSnCbOkKovOIwwjV0JBBUtxV
w4qYjRq1EvJQRlmix1j1W39s9G8TbEJRGPpZX5Fku5g1WDe9xTSphzNFJ/keyPmq
wU7u5oasRh4ykrqrFgBdGsTwNObkapwxooD1Kxb1d0IrEKqY/4vGvqD9Km9WXgeD
k5v23iT0mW+d87/Q/WIY0kkAbxVfWMF1p4T9+ASOvtZtfYyKB2ijI6qSSaG8ALGA
DcJcPGqqD4RQ3u87Etv9jsPztUiZbqREzq37yXQ8WxpPOjGY4/PZBBFvgo9981a2
+E2M3mM94t/9xIw00tbw9Halu2vrLnTxSL0s2cLgF/FPKKs36PCiAou43sfvPoct
lG3Qd/dxw9BQKHRPxqT2Un8pv6cbqRRaeE6adYXM65BcuGNN/ij6g8Y85WakuvZN
ugarM8xFeyUQsEkjbUfU7R3d2l5uZJxxygU7Z6w0wdOGgTYXbBX2jqp47cR/dFQz
miAb+suNr1a3xtIeZmGAgOyxrwTkH7W2OZKNDInwoy3HlVkped4cvn2baBcfppMV
VP6ymbAKBpWvZyEJmmVpvFKq6a2Cqt+A/TOA8OFrqS00j5Dep/PMy8UsrI6a7pgw
uEA2yjX7hQQ5nfyYHlP+HsZEWFaaFGN5siJx12Fs21P4fh1hAPE+OmBy+7q0vb/M
Yq8naI4CeCNkloe7HO7wMoyHTrE+8nzcCyQdx+ax6yPTvwPbMYZrWTIntPCoiSFv
8emZORo6L5tRoJaqDRiCNjYM/FGt5wpIPrcG5LTMpbybVaS2nvI8owWnIUBVlIb7
gkNJ0Xro8eVYT12tbC3KDxc8JVMQ8oKa1H3rhjuWE/3+P0n1EjGRXvbK7iTtw/YL
CkhiNQuUb8jFStNw3uYnG6QxCS2q9nWDbt6+yJ975YjiyEkKBqplUZF5E71XXkRg
j+RQbAxb66caFcPsh44Q0QxFqQzZE7OA64AK5oG5tDFsYLTWMUOQCYesomLkQbrz
3JURSIoK8gYLmiEvcZw8S//XGTfqNxTXEVVLFtqtOmAxcE8MZABQahv1h3CnkvmM
qtY4K+mdUeHEKKzpQqiGYzA5jwDs6zFvzgE6nYez8CYBtPvR/GpinIZ9NOaaj+uO
Ija1mHIjM5OS7gvkTdREex7nPRLlaORTStZiWcFzXRk8TVtCw52OXhgxxdSWZ/ZP
QWrSiB0I5raVQY9dy9Ia1lLK58++oFAmRV8VtynnWWqoa2oFWoRsJa5CcjLq0f3l
vdw2y31N1q+0kv4pwPP8K96bnN3JTChcGkS16Pj81N+GtdunnBRfXIRzRCwZz53q
vqrKvRDXy26wCnJ/WAMZ1lan0DjIGmwzkPFWCYF8YpDZxia3U9yP+wJp49aRr/jT
lRlUfhnKBFm2z+ZDSWoF/BU0rVmA67os8nDNIsRTEA4CIYpBVIS3748QMbsJ63zU
2iUV+DskwofO3apKJVRT+SQEqaqg+I2ii6LbPzZJoGHYZ8B/7lVy73U5TBgHuPPY
LV6sU6SQs6ZbGchcWqfFaRyARNDuwP2OzKIRk4EF3H9Wf8znQPKQ9ti48ZVQ+EvX
KPzRzQSUsmw0JuMCSNTPUmmuZsO1CEfibpo8JE51tOrIIVRap9OSIl9JAtwR4w/c
q3phIRWexoXIVRZmOT3sFXCRufrH5yPDeBRGTp1pT86B4eTpze/3WZ35nHuIb1Zn
drSlPlbKmOqWzb4oTMAsqn7S/rtLQ9ywUnf98gM7YoVYkBxNzSMA9S6ybKYAFwqy
n8VZhE4cpwen1XL8nO9vDakw4LNvb1AdBkwxmaaAv8J6ABpwnS8UCfbIOOyU6Mgi
Wp8JLSeI+Eg4ko1DIweb85xsiSnpHuqMgFEt/NuDnEGFiHyZ1AtScK/nUc51DCRH
mUq74eXnlmFZrtxwQ2zM8MDn5wDqPNfaKwa1dHmuCRQYCM4Chysuwb5ea27lpdx9
1LKQFFTo3pgLrquk1vBeMl82ggKPZqs5eAyJxSrloMDh5fMrI2HbZVwwttVZBWWx
BxqxMybTiJMDlE/U5reRT8UfKWDCF9YD38JLf2+atORxcxMKchBYY3BoRZBfY/ay
JRXSK3CCYyiRu+ExPQTs2iHspOy2nQHX2mrBGY+26arFUrNUHZfJVud4Swsab3yQ
ZzxfFh5WvNoivkQ/E/6wdjoxmejZFpg+EMdGEu4X8Sg3F5N5HCBHPPtJkNZBbX1C
4677YhqMiZYCeSvig88OqEb11Y7S7VQPw8c1qp1W73cdMPQGveexkSTKDjLDQjYO
SlpUn8yU+iCpqdKUpsLTJSTQ1fDJDjZzw0zZCnDFmDDMNmV9cXrpOXTovFVcQj4W
IROs4Hvd+bzTS79fYfY2ZIExskZqt9GAnA7v9XZzVRg2ZPYiMp/7UZrfy50ji3E3
9w96Ku4CIdwXsd86POwlnBOFfpIgC6rqMyIbg+Q1hmh/ODQiyZio8GpTf1XEjzfa
GAGOVfqnGwWlLuYwVQzfefDRczcWFrRa1/IPBmT1rr3QGwGallyLugFKhm8rBSAq
k67ZkldHvGffK3AyuU5yp5dfYnHEgNCilkcAv1bh309JKIPcO7qswunpUW+9a3es
jppH3rohQSurUjLHOmh3lScKtpT6b3vpZpFeveYXeChswQw+77SZQ0g+Zq+5Ca4h
FtKCTdNT8Zl9HkgWQfvSUar13BencLlHX9WPX8j6s4CKaYMdX7Mg92P/4ml2r1mp
h/qi/M4jz2qh+DAA9hhjnu5cXjFJgAQxqhhLmiSlQlrpoXs4wEtIVVm8ypSuHdyS
GfUhwVn4PtRMW7jkqQMExQpcAX3ov9iY87Zek8My/HqSt6Q33n9rQijiX17en4+I
qFwv2shvFQvkQTsIuKX4PXIwPnQ8WSwbkJ/F/WQD2NAVjQNa6zpQ67GxHUldGLJt
NFGEQYyr5cjSn6iTSu5ZsCIia1ypEu3tMBI4JODM1ftTKHeY9IDlzlw374gtUEL7
MJ2H8TVMIP71MPw90PSbeE6od1hibGO6VHCD54kh8C/ly7cBXhyXzzopFapGJooJ
I/sr4sdwNZ/WbhKX1z5VyX4QZrtRlPZ0JMT6Z6ViisuCc+SfEErHJpjZ45upBybX
3dkPTkxcSdNxk/Qx6bGASQ7Y/0UCxyZVrZZE5jlspxvPg01emOcwttI16HcYCrrL
lO37mlgTFQ0PE7orBbk3CtpaAO0xt7w5kn9styyw56hCbjU/yCIpcWHIUVr1ImAc
PuL1RRjc/JDApmSKi09uvboNZNlpvUGIipk3dJZjKDQjtbOKz3K7JvxfGhJAv2s9
WfCMfkZcFOKave11um8j5TpxX0AMeko7m8D5i3LwQrHd/P0v7+hakwZsN9BmWjXl
A5XwF5EB2M4A5lXX9LHWxjGOQ1Pao76Lu6Tqvp7Vi0U1wkqT6SqAOr712okHvPNE
9U4TzNg+gpI0DAfYOdQIOvKDMMyur6Lt1xHv16LEoxKX3UCB7+N9OJTomC/D/Ts5
TD3S2J0MTpBPN9PznYa9NC0LNh4r5ZGbThMODYzDVuFP9hhl+uN1MiUrMv76lLGL
jjeX+cHwZBQtIK3mDuGc0s6CVIfBrqZCNGxkouOilKNDg9NK/W0nvfAnfgARZ0LX
sfuUppffVBEAEqBs1BOW4tglHKFN5D5dtYzJMAKLiwU8/mopR8VSJuAmL+vwZOfA
Lo6iDbLs5+obDYffScAo9/x171iWmMyYykjdIrryzsaaYz12k1qXY9tbr7pS5Kmb
NTmmt3lLnwuZeKQawBOTgAAmxMqCJ4tiitymoRToWiSp7HFDjJJKt1c5aP/bnc8t
acSnLoduYDsWobgqgSRix9e/REsfytIH5wMPUCbQSMtE7QUgiHO/vYWMwCR7XWGp
Z30juUNF5czG4LQoj4B0zeLMzhQTG/AWRoZnNqX4ez8biYPefbJxExnpFj6M2SRH
LmeKga6YepgzVImtRNMQHIb/nCFdb/qo80ssxTcvMyy/hdaVKoZIX5JzjIcKiyIJ
uTn2LvkntOWqpKczV7LdcgXbrZgsRwrHF41iGqihEq8YKUfSLjMRUuyKW5uTS1+x
75vueYXAhl5xHTGRz2WDH7hMoS4zKlAWtzNVK2+T7etzptLmM+Be8OhKob9h40I4
M0DV/WB8LeVbgMBxYLsX5go3F/P3rq6zWT8F3UxlYTHeAZvogez6eI5rj7jcRvTm
B8CO8tGUPqMy01OhMUpwNI2qTZly5ubYOGQAk3F6MImmhwFK88wYK7+qTGwBwx4U
X9k9i0AAhTdlHCG+fQNoAb+9JOI1EqG+Aft7F3UGay3qrhVElhYzldkPmcVZBSfX
o0QJ7IYTviyipkWFbq9Yy5bkEmLVfCRBpjbzAVBz0RWVMVUQBkfOiyKiB+RHv2cA
cG9d0OV/wq2OzdQyalRAqZZoOWKmP4cmc+JhlN218+sfJFNYFR3Y0gd2YKk6hdYo
H7F5xkdHdFpjo/59XNlbAKfzox8ieeXvU2sDd8vvFHwBwvdP6ofmzbtlDL2b/NrS
3RfK4g5kScactL6ozbZ8veHegjeN/lRAfm8EnMZDWAGftf+awwizeiz8ImMa8cLX
X6YSkbU20qCSGW+EKB22OUm3+maCgHzYT9WvS/9pSZPCjdvZoT15e+F3Fk13hftl
fJK+gyfN+FEpzj0N27NBZ9wEACe8ApuGMAcBzmaJN4ObwhyoYruepPvlePa4fbC3
mm6bDod8lcqRAHVJ65YenSsRA1IELseOROFSBn4eWoYK6fDYwPIqo69w3/3l8Zod
NuAIV4wnK3lySFfjR4Msw4m4UF2tDx/wbsqj3iiW8reQbPW88xy+8LAoR89zYiTY
lCezkHqoA9fe2VmTNuOMBnRLyEYDH8ZalJ1FVenxJgH5vXY3uBaFMsajNcc2sprl
OGbVQmktTRAn61Lm4O6HpdGpvnWqOVIEd7tarP2w83ZgF231KUdlwxJg2GPXAg7l
Y+acUno09+sdH1ikUHMC1brjrcFA72DQk8qQhX0oMPUWqzIrsZ6vXKkvZynCNop6
f2JGIomP07m/odYIv06vfAyQJo3a9Ds/yoAMjDhyGINFdpL+mjfTTgPrJSOs9ERN
20XOxBoyuJl9CLuaizskIs89XpduOLoMOXIwmi/Oi5OPkLsTivPqrKE9ogcdIUHd
Ei8ASFURTCoEDaYukCKOl4HBS23kM5ei98RAqI5dGlviA0bs16I5BqxtNlrG6TSG
/JoVQDcatot8KuwKSsbdlpU9Fp2OanpzzoDRPbgztLcRy/2Op8IvPyz6ERQuD8Qk
9p5z3NpReO+6UuZrQrhUCfhkuuGZhP+J8MvO1SC/jp9AR+WA1x0GLX9SmkXXkIAA
Wk+2ELI/9nBwrdh/uLUG9XSpTyT6KPWsL48/PclUWGjlcoPe4Tvu+84xhrGvNLMG
PzDl30cxuEL/alcu8k3WECsMZ+muUtGQ6/DwYP/+KIDhSNA9P7G7ZMAiskRpB21V
DHw5Nye0JQpyEt3lCeBkDulZh/SEiL2zLZTrftqDIkkPP5tfwPq6mulbIXf+bIQO
DaXpPJY0UWi41PUDS813RFJ557O1p88Ix30xxbJiOExl9Et+6nMQ+Ez1WmZiX32/
8WWxfRhPWzUJc2oof0s3u3LP+uTcGvBYzE+Bmy5aAtUZ9mLaYrdnJAHQmzDn+Bf5
KoX0IvhIUL/YtX0mhMtp6q7dK4einkaI79Vh5Lok6iZ4p8dEyOGj818FRjYOpeHJ
R4y5HabZxtTO+kzEzwbg336lZxd5V+PhszJx03UuH7ctJ61Hvj7eNEpIX9w5JnGq
YIHKYgKi+8PyBCoLdz/PTvmSoLmT/z9aM6BL/gaS+SQj1tkfznXheoo/ut4alPa9
cXisAvWGXCzltnENv77e/JG05VKB1RD4JSJy+pLZ3SL41mKjgGCLLebbeQOhzd4N
FWkn3oUa7UfvLQRGBccSmUc3keaM4BgJRDB+m1K2ZU4NWEEIs8rjRCpIOLM1gGzR
X3RSbPNurr79QMcJUcK74KUyGea0Q4MqgXAohBSxbJ84W6tIk/PfaDl975Zt+UTq
DWnbAGuTygw6CuSO5hyDceGsiLas2jo/SLujGYPaBOlNIM/C7Z5C+yNt1LWrs7Pg
7UDsgbvZYOZv+CfUcbE3knX7h1Ua9Q38e0/rikdNJ91gIAymJc9TGyt/5w1Ej5RR
Isd1B7MoMXROEQ+kedE2yjBLBbVZZtcFLv2gxK+QKGPyluII9dNeCMUgQvZJ7nib
BJ7jTrmRaFkQs3t5UId3mjp/f+X0dZ6KM/ljQgGrYf0TXMWEvoGnAiWu/Iy8WAG4
cWLWhu18tFHYeX8vjU0WZd4UOdEMpLlIEQ5J5W6KeYvTKZiGqmdkJs7y/m9A+7m3
kYq5jvll4fBoBYasuN0POzeTxTlrm3sXPfXqiE+zULRtGPvtkSKgE/5kAvKMCkDG
ew2eSLL9XfUMQ0NHpHKlIY9nnk7ARMcrQ0JrfoIYGKvtvLfAs3xUKqn9wZ21xUeu
If/wBBRRb+hV4uLIJypB/qWk72CjTtZG90z/WHZljmDrjyPNOVv50+lUSBCQuM4i
Pw7ObKnQl1xz37HnGdaAdCVdpxhe4stgeSN6CAImOzpYLth5ZykWzeDnFFmznryl
Hxa3o217l7enOlLxR6QI0qNV2wtYoSX15O55OF3iyFm9PG/UfWE7sHC3B0xsWNqi
OWTGw1ug4HcbTUktna87qVrSmbqpelX5dE7VLE1O09TR7HmW43PI34IpxxcKQOxt
OTLGdTqOnG5B0zCG4QeZhWPQZ0YhQhXv8kJGxkjj++AXyv/7+uAc8yfynhnHrxpm
z6e0H56MUYfaeRwqD6txIyOewXyUDfxQG6Kbrxhh/4NCAEF6CDbl5e9H2q2Po5cw
Y/EiSaIVRQUYzdtLHSpeVSZ2eIQz24byzSSGp/Sbvp5zs4MKKVD4uqKVB/X+qFtf
5C+4FBKq8WNEN259QJOynCh/igDtu3E5UBVQkadvV5NT1VzbXwFRlyW45S6ob0TB
+S2NGprUsvZQhyT5zvrN4ztYA0cYpvmi2fOp6QXM5XjBjHBAQMmdZIO61tbZObfs
Ns5SKSBSENQZSMiopsstFPYp/LDWBENCGzXCSo6qU2ISre2q++9CCC+ryXby21C6
8IEeE2GBxc0CJAQFOLnh97fx9rBqQzLO0sojsyG1oadrHX2Ri/tF+RhItjfXRBqd
eplOnnHS1JPALAC++QkmI+B5YuSSAMvxXOnXJJi1HyJea2oqI8JZWvbpNYYqH+r0
WO7iRYBSRqo6qwF/hrwsC1q9+uwMWrx5Cw6yiqTewxgu8lfjMEpADUjJ+PrA2PiR
7HO5GdMgqPSg7aMVGgXDnIlJHmr3sMoNrRXKkxkDb/A1KT1hWloLo0xlPM1pm6XF
ozpkBlfA0nmbfqS0nBTu2Orl/lbl2/Kk+1FNpxG9HcirH8lBuCtRn0DEQzcr/CNR
47AMwJ0KnabmmKqflLaQl2waxyqeEbtUp0ktii4mslTdpwDUCQxgGa54zIEjFTJn
ecYdTCkLjwru2Rq9VxLClTPSjWURqOiSwnS4Cb6rMkJN2OrT7VP9Y59jbz2IkTe7
AXzHb4CzzYc6D/DvtV6M4n0F9YzytEKGOlwXCGMLj9J4O40dH8btXMefZsWDfOSM
BPJoTwroggzGAXL8Io/+eHbzVqv81bgOz5e9XVLuTvk6kBWZ3qm1G58ykQoNXVcK
20bVlMhd4RD24Wzj30RTwvoFMYKph+eskRTF91AdwSH+aCij9OOF4511T3jAc5dL
/yu99C5Ft7PQTHS0CQCf/7R6W9zdZ0CDGAtONOaRLWQ7GFd3ZKgwphhFRh8yDtYl
N+iOyXKGDIEDDvpY06Lf69psEsP8loD72OQRTSbGHZtNzUdhdJzULkAywQlBNlSO
NPGrRE/rv2MwGduJ8Exnyu0Y6w0Vh35V5h2jcCG4C76ZX60r1SGAakHYJUUj9wJG
2pfZ1meFExzGkPiasXRgWJpG4ApoCfZ0/6kSa6baVdllgxc+IB0pYTxjadzcsf5e
gNyT3m9kCN6KFah4+xr/b6VYMNnnlUCGO+7sc1xToEMx1wnkGoevzmD9cWxpFcCo
1pX1/iMlzXBM7Fqc5p1ddZ5Cn4yuSODWw+Drm2qsBs/FvbtS+vaJx9Pd0t1cCGai
0z74NlsCHY5kna1bS+vMPIql2JI+kg8AxcQLpFwe21AATc8XIxSWtNOpQlEObrwM
qrX47GaYtwYyvOd7/KI/fp6SxSf29loucvK15uCWdjWt7r2huQN243Dp8/RT0/n7
TGQwvAA2rJgopcE1utPY12ZQAt5/XKBdOdHSkHwCCDRyAbbJ29btYr4s3Qumya7U
LmQa/HFsncrCYL+EsoegfBR5cqC4UCNd0J4R4eomTp6SBCebzMBZuODDofM7PmqH
hAfXJzOYRfif5+FexaHwhe/WvNXiEkvvHFyiZy3ElkYm0E4a1xM9fhWRbxaa8y0U
6HD+Ph3vpJy8UIS22/d58Xl3KAcEg/kj5Z56uQhitdLEohqQdQO5sgO1WqFfCvg+
YX+3psTtdkQcyAcxxaCyYSxjgr6w6/i8cCinFiOmykqo3/Gcyy+Ao2kRFxTtyDEz
+dLFMqFubfXn8eMPGJGrz5l/Ma3cD0W61SgB4X3we0w2oW5vtrpgKjjJX3V/XgE+
VxNZrYZ8sOKDaW0A8dy8kHn3/4eUmEGNX0xP/AX5UJixh8Mr645uiSMgXK60xSgE
tEbaXeLjStx1amvszt4bjasGXWVJY/TkX/SJ8Kbz8gbtPIOiu6HG+Ba6zBCk2LHw
I3kp8Q+eJZcuwrroW+dqUghbScFVYpahJ2LPnNrB9DY2SLbeYQ8dcDHcCaCiNKXe
dhE+CE4lV+m6VH4Wto+sBXldOZsjf/iwemVbvGzFFzoHHr4txgWWSdfUDX/i+h2e
o0ZG0cn16Wr2C/NozambtK8Q3KMwcrTBzh94+3uQRogT7Iy4hl3H8NttcJsP3Vwm
eBjPnoTHZhTWMiXo51bx5+sINE8uXG6FGU1PWRDiljcGiyPZ7ZhXDhNxKpXFq6BL
WpnyQsnny6HTIra/e5ruKlnK2tbFSe+ajdhKupzPq2dnetZ2avCBM+4zqyEXf92n
blpnm3J3gsYsATPPahl2PVCp8HdPLbxI0ZT03LX+djsgleKgJQ4x8H1tflRI9/d+
lckI6SaetXP+j//QcJ4VxafX9RggkTvMHnk+DkW1efyqrr/UICzvV4EBlbGV7Jsk
UymCj6euIr71Gj2r+FiqNzvDzxegH8g7GNTqSuSE2s1EHvV9m3uqKFAjEipTGSz8
9cs8fjlYtfoLd9yF+tSSdyLylzUzRqRyey5HxW8V+1rHzsoc7qfIhllz7ZiMVGdY
ozb7R4q1bcm1wtBWqqDn4akgm4IzncHNy5HxNcdNThre/eiPhL9vBeriJYNpfiWB
e1KdvuU3Mtnv8FLtmmgvFbSWa+a0Jlopt5f9JAY9nIjTppJvhnQ/97K1Dv8nd1aN
ROf7QX7KnSnuTKTyTvyZTmBf2kDhHqVcEnJXFmxDHp/ipM7rAIS3KYy1I2WjY09R
U74dCau+Hbiy0JIaKpGXZe1BOB2MwFO8z9IvkFJ+iEqakh2VHWM3GmqrKE47d8E5
G75Gj804TM7sze5N4Wf0N02+ybZtnyZXX7z48thuTTk/f/9DIC6pu2++g6VWq9xM
KLo+ZtXfhY6R2n0Wybp5rccgPSZmgNolgiWSsodgvLBGHA68jGQMxtXwxAyeQMp2
MIfjCaJcP/iczMcnOj5JW0rX1g7Z/10UzbH8043GNIDiaGTP02vKcW9/fTNvty6W
MXFmVQiAsn9WcFLqoEGhq4EChfaDldLks+Z3YuSuhVb6MYnmgInzbw4o3o56cfvm
NKRX29wSjhjp5lauXNhOFztV/1yssQXZ+83slQTAEKMDVAIOQm079V/fdopMmpki
X5jMC89phXVgDW+dMapOpgywgzoYqpUShBQQgrmd6UNF7UM0YwqDkLEWAGMvXZD5
1KnrF6uRfnfJAtmbKbkXCr1VH9MEP2WVRXODv01VZQxyxECBkudBG2aaPF5sgItY
MUanz7MTyBa+xAkIN4QvjAY/Bki1zSoF4jW53iC52NX73TQX4X2Rcs6D3v+pHCZ8
ZSQ/W5/tH4UbKV4AirA322wJAXhpAEaXz4a+8kU6qhydepNhkBrLb5SC88lc7RzO
yl1/gHeCxdf6AXehbYZ5Kgw11o82ElrOFhe5Dn/xZkaBMFt3CBdeeUAP066NH/Ke
sZFTpIhzElqXuIVJtJABZCTwn2nZn387D4zlfgLLZWO9oZ1s5Avrgqi8inKN7Zu8
yhaLUUDceKtV246ekWlY4KOungDIjkNIdbMkcXCh7TSRzkZR025noSZNc0jvFTKs
vYK7tIuwr2KFSfQX6hyDz+ZK2ZHGRs7ep6CbuMq9W++I/hoTHZp3Pv3Q9p4QtIFJ
PoFMM1tU07l2Yf57+jB3ss0VI44KvDYEq6pps7ekLqGBQjzyrVAf6MWCkcAwBn4j
7SrK9d/sPv9+9MumkFSMtGsA73Ucl+DDokYm1fgGRgZmB6iqWY5sHLUozI5YKJJ2
zxSwgNpiNw/c5ws728ut/ZhKgrr/UBgRbfVa9Vb8n/7mxqjvl2WZqwTv32w74FwT
I6/fCZljXBidHpoHKRSiLSu6FZGtckxZSM+I3c3kG6VArS0wNdKZj7vh40JU3mQl
q2hS7jpTMVloEGfDByHtclQBUVf+8u7LkvK3uvV1owzAO8kyQDpTj+n4pYMroqdW
EUQlcDoZar67xY6jozF2RFX0rLA32jFz91MSsp1l7Mq1zHbtEWtewXuOdTjKoIaD
+EuGk0ZTgBAZ4lZOs2/5vSZVMudDgo06nX+IfG5rvRmHsQJHwXY5/z7CxNCwNfhF
mgWUZ7MwzybVW1I1zXO82jeDTvxvyEdoz4zmVovDnCGE0EKsJCyLsUJB3dcrfeJ9
ibHqscsW5hg6cvOjpMRQGK0jOYBZODfkoN/wGlv0sPcLhtseqfsTfWNGgA1RYz+D
Jr32N3i5C+NbLxuxB30Kc/Br148894hMdFXQnANmkeU+1DBhxCBesGn+So9/izY9
uHxZVDHOBcI+Kysh06Mu46l5sdptyS2XSNuhNM1KGYhMmePDj+Qa3bXX2m472+Dn
fTBZU+mN/a9AbRpM95zpS1WyiGy7rtp7qds7q1MrLGhDBmdKQMS2iaRqoJs3Tpzp
VyCyPktLTiI068INRMX2YBAMuCbDAOvYe7mmzSWPPJjiUcSnIjaijMFNgoYAxZeH
SwA3PQ+IxmJDvzOU5Jjvm+JwjIuFq/W9+CXE/gj2O/KWsrsidBBtjDLKvbnicHI3
CrPhh0hZXt/d/ssSlb6ffGrUgnVAQDJKj4OLLDQSoOGsNbv6cFEvJESwGItlQy40
5wfJWZ01fyAS+XLwi0a5aYp+DQPllrpzuOXDn02aFEKzqaYK/NF9bCI0xxVDMt1M
oop+wBQOwjR51BDBSJOUrzWaIhutvSNN6R1hr1xioaOZURAZvZW4WMcL65ZrjwYs
qPvT8wbn7vzj8NKsMu+lLW95AvsUIOnsZE9pis3FsUPJmyHzi5BAN8Z8hRo1eg5N
Xj4PBZW5vOzs9PAR5GmQwCvvvHeHG2bP+Ats+z5F8S396TFXBhcGAQBdbCGzyPpA
f96v01SGVm418eDKFBW0lYE8XI8+qKSEqppDKV4HfSOolRtCCi+Q5Sa5YKwUIV9e
CG/0wa5vdlgFpe4zt2Ed/h46XkvXIQnCrYTlSCll6os8DK3gmkdVBQ7gCJhrIyIS
pakQrO5zQQz8rNLYf0Grcc5wgVCIio1FBjS9bdJHtrrwljrk7DPsfhjGPIzLLk7/
UAt/A4MkWWyXHfYUFAqqUizLHB0RK54BtpnKaunmKSAMFiCUxgI5HA/EXRA6VXEa
j3PrQFrbVEiDjICkiIlXfkCCEWXwcXxhTLCqtvuVEd2I4AdthFjPb9rxmhKUQOWH
IfuGul9laOqDSZQ+S4xzuy0XZTWh44ZJjfPbL/Gju8Qlf7w3n1hLLtDn14yn2g2O
mWaAUq7G963dKvivr+/V9S2ffUWB48n6tGfR2Dj8y+n12Lshy78UjX90Phxcvoym
JexFzCzw3X/4Gh5cs3Ju0/fD0DFYXyVhuvhl6uMhnRfvctByXHB6fg/at7lOpMHK
iwQCDyYNcUnksmLz+LhCXNCW6DPDLAl3nvtvWBDB3xL4Ei3bv8Xw1YMHW6Pc6CPR
14WdHzMFgdkUsoMkQ90rd4El6eMm1gimqpJ+9UKcT4+OO418HI/kdv6OYmOBjFva
0YqGKliaWcf+HDQRnxb8yTZtHTph3U0aONeihgKxIBwubqIeC+q5mql/RwjAzB/a
2/Ot5poP7u1lhn7z5vVwzlb+IqhUF3ohlnChKHXVWrCPw7SSRY+9cnQ/JG4MxOdh
BctVsOxuCQPLkgVDo8kRTVlOkeAC4UxFYaOal5ctGWgZac482I+RZtiBzK15hxwX
m15s/HYfAASrC6o/tS5m9XM9qc/QpxTQJQ5Vso52R+8EeSff6LJliImkM9Cct2Ie
s9BqV3n5gSG9LYh9egTDnz9qXRHqacw7wcW1lOIoNXWY6U7hsLgTd6RwoIfZeWTb
Vf9YFeqDkZdPPvgxB/RVQ1n/gA7QmxA/TJq5l0+hPMZxOA1g9LFu4ViNozgBLkkr
HBykX1yVsfPuaPeajv10oPjau7CvZqiPsnr+zXG/lA8iwfH4XzqDnRLrNC/RrOEa
+CxadlPWpTZ3QwDzRRadMq/OxZ10S1chesYyc/QJaiJA33uA2VotRcVLdDIzrh4P
P57Yj0yz4NhqpGtXjaz8or9Vw/eWKynOKeT++GtygG5tjAafHNRodzfVUf1KCfmJ
ma7JReFHWcqenakUhlXNLkdyguzEAK6FYYtwq1/dUQusw6SrfepGEob/8miEShZc
pSKdKJDCK2NU9zqwTveVYtriIWyJ7bjDCuoJtmZHN0X/nxkXjSBFiiOS3NS6DYcr
eeJ6qnU4weeO+UGcGIteGNsanWkqz0PydMWGvFr8NNDAlIId/sO2sdYA8X98VQ3R
F2D555pW/HgJKuY0b7DMQnc/BMpPNVuSjiKxldXPIhZ6b3YVmDPrLQ43fap8tcpa
UgyjyaEwknjaAT6tM1FWXQZDkw4Udcep7KDuLyjSOyTgV7tO5Oc2cPFzl+mBOrWr
2m8l59aWBiKLkJkkdIdPufgHXd9ckCnQ3RlSphxGoyDM431n9+P89JpFOpJCxO65
zGyEjJkoz9Vq+HdgbWYtdhzhS2rZPBe+rYu3RinDijqFS2CI3fCsUYwKsoO2vhu1
jvdBMIo+l1CSXsH1FyNY17jUT6AhLzQxpd7mFMJ548oYkyqucBY6SIigCJAYxPZt
kYbJ+arKThtyJSV6bGr/AAnUKDsczdiqceJ2uf1reZb1rfi7wHsGQ87Ga8p/vPod
E4F0+9fnPWqEeBJ+fTdcwpIITg0jcI4G1W9kRc/FuSsHuJ8fgfRtGCGzuqzNUxho
p0e0Auwa4Y9r3vSo/PdYos5Gzeq4sO+/t/PX3o428rl2p9yJz3QZULph60WchhJo
6tMIlYUtayO1u1xBgXwmw6wOAne3JeE6c8jnQCsIoKHSBY7WPwPFmfUMAhneieCA
lM51Elhz31EgFl+jFLBi2MZDrPHnkSJ1anNeZLQh+/hs+7vT6bxkFwDl4NdLrM1I
QhnqqltuSgnDTuMBMXwFi4GqxKFGO8YiFKO3f8xK5ToEDlK1uKORDvTLJ+dP3BH3
CyPeDxvziqu2GeQBLWxT4O0sFhB8RO9+KXUdzbceaRnmSVLrgxSeyC3WsSD7nfcA
TFd1by4Zx8mkbohF2GJS8DX/EdHK2F7zD5Euj2CkkNF/rN7ewxwTHkULBQ2yG9Jl
/fyiWXySOFreMbqUmYCVXnBYncLSpIYlzq2ZiYuwm+Kck+2jiE3+9Qi6b+s2uVoJ
CsXKHXBrcFvZ/nC+cJGcE67lU022W5tq3PpSpXyK0wfOPmPnl3pXa6JTlOGZcQ7a
vTEKvirAJomOvx5FB2g0iRrsou7e9zkS+/KH4Z3LKuF2N3Tno+9xMfmy/olkuenA
hJsIKuB3ocAK43mbkA8pDsZm65yrwyBzQxlmr7TBIgl9E4qRwwuqoIGTCje+OpFQ
3z7bpj462vAZTBczqrp1xX/C+pk2slNgKYAr+RZ2+uExGOqVe69D2sp5MPnHqysi
40YaYqqu7MIrcckW9HxlLdDV6MbRcjnm7r1GE+/AeKr/cpPj1LM0yLTEo1B+2izY
Y8zLBjIk3vb+kgMePvYrN/NsfwW5uQYTvwiMQSojRSlHAHMMDiFbqGmCjw0mQImL
GgiGluUmvCoI7lC3E9pv0j4xQd2D/W3sNoaR6EAi+cHzVz5CV9I1UCOfN711mcQd
mCZBIkLVCqhvQeiZFxPr/2V7fKEmSVwYLUhRjz/4HmwGGHh2slSpTosMg4Xq6eD6
GBmPBctzL3/29hDDEQ31beyKvs4NiHgByP9gXtujDzjDP+R4rpj0x2f3e6Zdvo78
8Ky4KKQDD8TG74l9lsJklVEBEefOmFgZ4OmMVh+TEQyarjTXLmNuMK6PtyghKIpK
S2cr66pmU0ohPOhJhweLJXmzy+AC+BQOxDABQV7ZCC7G7n83ceooCEQy/7KkGGcX
VoBEk8TXvmlxXxZBUg5HTLpuSovv2VzX9KTG90RscLH9ymV45mEQsv+Fs/UT+I4m
5uCbhZ3LSbp3/iHbFFI67pSRhHoZdWjfbsFidlt1y0SrLJtSlwkWiOBqIl5v8kRx
ZbBLl+Fe81SI6iQYeZw8Yaf9Xb9WJ0Zoiq2hmI5fUCczCfj8isUM/RkoSjkj1NPT
TpOk4xTD8cFedvZK/eUwQUq/TMweC4Zkyd9zYWoWgo18S4f4mWKVAO8mfeZXHYgO
IKtNsxqHTwkLOEvMfNp5ldeHiqjGFhAC6ajBDGsj5QzxD7UqRVXl/PmU7sG/lkZN
CY4mPA1nyJEb9JcQkItPzxejUyaJ2ZDD/kJinXcHbTDO1Z5N6sRrIWW52s26LrFt
U9tdSwnZdivZFcOcy/iQwjGeld0t+iEQdjV5DadtTNb6GJCWvDaEspCT8OaA94wa
J86SKR0Szvekoi/uk4W8rqp/0U5E/JmtXxhqYAT0qDnY3K70uA2DGalV7l+AkMWG
voveIsaoJeP6hxNAFJBf4cLQHKl2H9anFs+pFStmG+ygDQDudv5DDfdQVACFhz6o
MQnUTzI8KHhSj4FgH8bGA5TeiQ764zERGVYIAGg65CVhXf0iSuMbaMHFPi6SnUxk
XOJGIFSOaX10F4EVnpazFXhKv3ZQLBYCRPIxAfhwnS2JcAomzFSt2ie3XKqe/6D3
hi2M7ELc5u3TYauhwHdh4Ya9kyRdMUd4zMtlOpmvwncym4lwMKxJ2rrSkgk9AdZh
X2vltVXe5oqFncMC30FKUJkOfqNy23C1wI0X3Z2zUMR29G8GZByaKHWwJ3tFEDno
IaeGaRKz6WrFZvURGjHUFYEsTt4LjGoD1pU+oecxXUtsWvC8alViMPcMnI6TWwK9
gSV/Tt853juxW+kftCNGaNxnlJvaHtxSFa5PVVVp+9am/E4FhZVazVRaTRPu4nXr
LAJsi6RIrBlCBFJNuEo5qAZR3EE/6E3WDnIT7r63gpVDGLIOeO/xjNlJnBVtFfs6
PUf2Tbv51VEI+F82pCKxaKDO1Td/YgnrxByZ3KOzRPINDikOA/wt/ks0pZODbGHI
OwSY5Bu5Nou8/5vzBv3SfLs3BhoCiTQBMl606zmQ9P/3OZtMgTUBNQsIAYsvXjE6
cHDS1ySYAlQnG3WVEPNoQc6owlpB7LM15cMWZz4s3rwP9oQU8TAE60JZFIUB+btb
WjNqugqdJmaB4aU3AHomlvVwKar5GeGkLmfCFAHw+3trH+ELDucpVfD92gXWwRd4
0QMW3ZDPW3dZiXhAbTuUgOLWn+YHHkbiPV6lY7Q1/soDO9takq3YE8LQWPgCW5cQ
AEBz1CiTxU/vRaFX/iHHIOe0G/3oz/ubOLZPe1LbjxNO2C1+2lhxK8xms4v/gU5X
+FBE/iTrJD2K8qjy0zLE8xeSHrgLR9MQeraldCYHhNSlvSkCOYpvr99d7ED1a4c+
XYr1vv04IygHsA/Z8kehzZt3ZWoQeg5qFcEV5dz7BF/QQSQYV9NC6jhW9+PwRMF5
00W6iolxk6bKurMPG9WbbQE2qyP/v2yPUJjsopx07CGv+xO6EVqtLjBdUdxoXRLl
QABTFUGUDrfl52S9r9G4+2aNiXEtYKOrxp5mOT8bsbXsAd+OsOSE2z2p0kzKMaEM
PpMgnECTZx6cNbwISwrz8e/Q46KSxHytFqlYLYRMsvZedtDfNHk03siX7j2UJ1IV
QEsFJkzOPOs/xDoJXbvUvdCE/ExOnG8O2HiJBTZxxlvRe3nV80TtT4zLj1l8DMh8
N8X6Ki22ZSHpVLjLRjpmRBeD7Kwd1HsecXawyWQ7pI8Gp0hkoxeT5v43cLpQZiFD
6z7GdcHQKeIsdzNBiEXmzqUZnFRHaDBm9sWLa5bVWySlN+kqkag7C73LR+txIEdi
L/He6QjLw1I7WxiXfG6tHElKGf6JZnG11BoHLzUa8tkpRwWpxa7fNNxT6PCaJO+2
PNP1E7nWzj8hRxkQTkJrsuEQ6Lr4mM0HqVtcd/WVqDaKM0ir4ngpSyu+6v5YeVwS
EGr8Odhzm0TgLZtnNYZQAcZ1HWhd4iITyIdtU54ZCLlbghH8Sn3QejXGE6vaPz6h
8yPTy+9YDoq278fgOfYKSRzS9RFLxYy76W5FkmyjNfRr4VjNUoFuDqvC9PPnUqrU
YzuMTCgWsLS+YNBxamnk2X5JnlMsOHna8aZhEsIN0JjgwHIDKkvvR3sP9wrWdwoi
weOOgaEIG1iFqq1H/Hg1EIqrwQmJxVfNogy2VEAvDhp7RtHnm1lOD9HXUfhSu3s+
lhofCk+ScHXFDO03c7Fa1KeyavISC2J8yDUFFRIZARPFkZ6k14a7XVqNTyFlLrg5
C/HLu33OFaVmwZav44yJALXytV2O7MW2X1aY7wy27/sIi2dab/wurxzrrQ3qELPl
ePaCWIIsir94i4dKFA0ZDrEfm+Moo9wkNLC0WVTU9uYAELe2Or7t84eWNoAya/nq
AvkeRiWIEWUUnqkPVVIOuMs6KF2AW2v0oMBwj31qfOO47SmhA3V31UvZCEh1K1U2
SJR/7YJAhETENT06QWWY0gxQVhj9H0UnsrwoSDtLFOLPkwTvQXQ5A1YSexg6mdCH
36CpOTWqZU7pG+rjWGuBVmulFMgv6fY+KEMVQFRfRnOfqRr0TBBrlumJICCKIZi7
J5m4VbItqqgH6lfJ6xoTnnEfnn7CJGFh1TG8GiQ0c/NerY5JVzopfoz9qrQ6C3vf
pLTjzmVYBn8BlSJEP4VufxMrz3C9krFypkxIlBWxdcA4EjXIic7amIgYOb2p4o+J
hTMkeGHCvrrczh72eK/C5ii7jMp+iHfclG9MTZ2SfiwR73ox3cQcsKKAQoS8RZ0A
3kSBoRDpjgK/lSkso5l7eeMX20iousCKpWsPCbZ6QzpcLcuhftolQnkhGAGEIunJ
ns+QVLAbJptxyV5rb+lxJnsfhG1RCNpAX9dtxKFSehznMA0dD+ueYBL2tg6rBsH7
oqbf32ara1zpI1WffwoIbdZfk8mGykUA6z2NTY973C5t23LRl4DaWL935cwkIXhH
M60Rc/S3dWaRH1uH+DxG3SODbjjSDFBcYTdZuVjo0SUmmoFIl1xOduxKElu7I9zY
VvE33uQj1j1itvQJJFIiDU/Dn4iv50XXoEw9enR0G90HZka90gmCLnQ+SetU8UHX
dFI5Nswl90Ne+CbsTOG6AHOYSQ+yrYt++nU7MLuKzFKQ7OXUj3PnOHoJfFh/8CE3
xS+AZwrm72iyRiCoDdsQYDBD+LRemhf6J39//RsIap+NKhwpjJ4lm8MLAItLn9gp
W8LBHrCp6bsoRHAkPrKgLqLZR988WRsW64LBF1byxvReCsA57VUHeFVylOn+l9Wo
ToWFgNBpHqgwRJDnWKMJnwKPLX8BIef5xBqAyQHpKwq+g2UCgbHm15mgjYc0ESY9
qYiyorPI2wNSSrlrXo01m5IDwqEpTGlTMgPmnnbdZHrC48CLMwNprJ1HZKzV/QSn
AfAa/7RyLRS53aZvChY8UkGo1gOWQgPpxiu2OwGxz45ISyByMqD58def5rA0wLOi
3xuJRSBxikoOwcY49PnVgxlmcbOODR3QG8YdHPMrvU2+TyjZgUj5CJE8WlMrkc1u
L8vwKKjT+vIBC2GO/PzXlsHYjZ2UzS70fa/tcPWUSDSi+FPRgb4kVNcG82fwn1r1
LW3vVvKE7vDD1K7ZJvYDqGiHoNLoVQDuZpkte3Gpx7Y2cLgJdn4LGs4jecq/+0R4
eRS5UCp3cP8fr14u9/TqL450txbSRqEZscOcrpb7mp0AsnuuFJjEilMzus0Fz0Vm
JAgGJwxja/eVuQxzYYnUNwNz5aaxy5mZVS4kTHOCOwoaCxJZ4cYqjScnOisP8+jd
ztjzxx/qukmLhLqd6wR5sMtXrF8W5CgliUW0BhcJ5+fIMgTM6tUthVhALH7urhnY
ePmX2nliiqjVG3o7RigscTSBMY9lcvqYUPOytfJAHUoCvm7kuFax/1ja+OYiw+/w
92e3TIm6DcXeejiMSK0qBuTIZ4l9GUDbQwJSaUnHGmxnqMDxMGVzVplFJHAJfKTB
MbNukEOZ1JFXbKlMKds01xy0g81hDctzew8+EcutcRtz8KhmVgICizWYdG2WfskQ
vGwFx62QjlF2u+M2RXqRejxFve54S5UlB3XK3hPdX4i9d4q0mUpJ8ak5pLGjiCyK
081UCJ1otk/+pkEsF1SdgFKbYSHgI8O/IeOPAT/DHBp95zv1E+WI+ogqJ+YHSCxw
S4kUtc5R720NeCocJnw4zJfWXaBTcnt/S92c4dX2S4RZg4Zbb+YexeiuE6TkSTkj
//F2T+DI43xRYCQtf5eyQAgX3WLad3XPvecp3H/BTuoKfY3ESIbGXXls5Zon/3Vi
N1i9jOFDnSBpOEFC9X+F5GEfg7S/k6UwGB/gfYfr/DggDY3MVbCQo2WtOlaZDX3U
3L9grb/+0Q+bJW+OwNQzdyaE2vl9axaB403HTWuSEfiJaFkLZaIuK9eVmcLU/QPd
AqJ/mU1Aw8Odclh7RqxfoWvxTF1EsAwft/E40MkCrmtCi9VTnUQv4gZkrBhaANtA
JVgi1COuspc5Pl2jn2ewquAYHGI2MLanNLi9Adv4BdwXe0pghnzI1olf/jBFI74T
yIoSMU1At7dWs8WCkEiDTNlSa/NSWrcr/FqRBJLZJ+asOUTpMSjBSbdx4htHN9ng
BdBzkzBVO8W0kKtR27zHJOgFxec4DMlospc7uTdZzZzWcR0V5q3v9fHPjg5oy5us
bH34dOtXH7/mhlU81qTXMtURV9H31aDMQ684518L2YTXjEafaAVv02PlM0H1J24q
mMSCfsfEqyNBhi+205jztXqJ0cxv3d6M5pWR8l8k4Xf8Grfb3U5Q7JoMJTCJRghM
R0tICtHaRO24tBaVkBjfy+hDrkwl7pHzbZ5feQN6h++U1CjF24wYf+g26SMKW0u+
+H+c8Sh14cMPkUjQUtgu4ca4daw7MD71YtUA/u77+yTZSsyZTmy7TCobjF13sJ0K
M6jXiHsnPvBn6bsDFCR/5Ht81Y36E/bRCDK6zVpJnYAd8sC6Ed2kfvSq9oSdIr+e
TNfR6/lW/5ysgy7WP7y4KALE/dAGHgYUAPX3drCJ8YtyvBnuwXlOyiqGYJs4bb5i
odRdCM502doYVExdBSFi+MqUponxMQe5zhG66J8yu1M0iMc71eWgnRfqnWSo2TmS
2GOWRx1HO0rPvILOZ6GNAjxmbyIrMtUr0jDP4xXeOcLvZb1ZNrkIYWNQs3E65AgK
rxzii9Jme61JmjlAitRsoM7LfE9cdxiGj24urNS3/G4Zs40M1y15GSccZ5O7gjGz
yE+yvZYNT0YObctB4fWX5xmKGjaoYntqtHnNsgImrJoA3dtODER+LTu576zKBc4T
jshiyiLWGJ871ZATLskWqcAjVjmw0k1ZSk5ySwoe94S+e7HymQsPcpmiLIP1wOfV
8trvRG0HlQ8GPTVNnEGog9G8QHYDZbrs10VaCI08aPgYrhS3n4b5aIfcU23Mu7LI
p5CpBOwPb+Vt5yE4W8flSu4DdtKtNeHrSsODyMTwAfMWkr8NXGiSjqfj2D1YOuBM
2fsRUYeIPWyQmGX1zexKfCX/p0aht6fAENZbEnQJsprH79aMfKKtAdoRri4grfD4
V+o2p/lBD3Wa/ahpuYQ/7cAqEH5nj4GWMHNjSVoAA6XzDOAwesUExHtVP0/hP3pa
KNJJ4g1YkHOgWW0eR4kX8LTbYZdqucyTcw57Mu9KRqelWPUux48slO8QZ0XA27n2
QIAlNk/57Db6sqVNkT48Orwit/PwAeq4RoLdqvqzT8qgrZT5pKsMEKkeutyNg/p4
2L0kmjB74by8CFvC0qhgLZAoqv4s5GnO4ZGSFvM/80ZwZU3RgpCED03bzID1VzZ/
fLSA8mypQ9vN+7STXPz6yftDwYNc/WFh66iGKNHMwN6CXcycPr09/0hwAByYXFhx
esaiiIWzp2SPy/roLiS2JaegZTTylnz0cRM8wmYMXfGMboPyrD+Y2THXuXxawkGq
xE8hX/s4E2EfJQzLmg+NJImBiUvWa9WuLu/k4hKFOvjjj1P85jUQ62UrYZmBFgGA
dHxQKdveullnriPETa8uI8oIVwEsKGaHdnz3R+3GTXcw+7ppTisBo4D0Oa8cT8sW
Y3g74RB2/d7iWKyaOQgPCJGDbcZqAHA13YmgInJcYf0IAWPui+OSdxs6TKIM8F5L
XJOwweAtuECaulxKgZWMV+yk5ul9YWcvkjmEdAE7cjFOFlidmqyvZUt9GbTrfRWG
6Ty9wlWXTIAyhhvif4L7229n53ADtuRi2fTBg7Ggj76NPL0VBZ3zy+0dRCixyVF7
ayYiQtJWNojc1urVuhp51ltSxlYJNYsZrWFibzu/qiS/dLBQW9o5agZ8dOitkTXk
rWSThvw5MGKNiIO5hzjOOF3csTVfxaOZlX7l4Z6D5ru0qJdU9hsUptMMOIEzwDFp
m3cC0ssuV97qxNihKeP4rfwB0FToPK1NVB839ei8F8AMcIiCnU1Sj9Rez92CEFPG
xKvIkqBdqEF83m1AgFwFfvbc0usG+aiBl4kI7DCj89vyQCW1oANbRIs2RmZUzRov
rAxVSI0oX7IkuHS8QJc4kdvMikWd1Oh2IJB9hUe/Qdw9g8QG2gNmzREBnjpoUjDy
M2Fx3axzasQKtk42hlgn2iWFcJzfnzKUK5xVbHk1q97PeWK6v9YVHUfRbvt38qh9
p6d2jYFNRFFp5s/+9RyV0AntG/OliZpiC/RGIp89++rEt11mUpsoeDv30jVee9p2
YDMvrSukvHDiAHjPe9N32gvNdpJCLvyq2IN82ZeIm/13XR9pJsn5/eg4ScLM8xFC
XfTce6R2kikXTJv/ng8WFFJuhusaATflM0vJPn+iWYdo2c0ISQmLK9H1XSLqG97K
JZBCFp3GM3n1JBv0qkOCi0UF0GBqQswJqDZldbSpDucJGZDtdc38NhQl34zjp6Pq
TTBAsJxeiaWTT3CQzwVyXuitmxlopocaawnHetWXB1tAXtdZKE/TrSUH0Z2zO0UU
k/SonDUkrgj9TvmFP2L2MSn+Iqifae+ko389+9FpnXHWa6onXO/fkYpsigWcAG7w
sxBTozCvAhGkmFu/hBX5rDHv3clKglTP5JzWv98dsCNEUg8wyN/4z/HtehkW5rlU
lPVUHvccgEPXVnfSlm84ycXALouqe5J4PXexkCQqV+n6XOy9aRqaJUsrsrwG7LYE
xJW8A/zuVUbQH8ZqNfmba8GkR1jPg+7ia/CAYm0rBVK0n4yKG7r+BfYfbD5ISqF6
AOR8uRwUKFWcbkJfXFTN+NR+qsUWQojAtdQCWswFhl4Tf85Z7396cheBMcuTBkER
3bN9os1Nq6uwvixXwUPNSLUzPi+Jce38XiMYjTzY8vLRPve6JpW7sxzkQsiWZcpj
bEWvRgpdqRN4NP1LQS9Cea+Mz5bTkBEOaU/zTIy06CxYardhaiY+PTcj0wbLswkX
APIq972RWC6oYejC6S7lX3Lx4++14mkZFkC+XVEbUDQ24+wwoXk10AR9DitI9pPI
EOX9KLucjpa0CHJIgkVezJuJ2bxy8qCYfc7lvOfWaTttbGxmLUwFYhMad4mQKgC3
5pzxIJ+FzJIv3fvSTbnr8L1K7iEsiGKKA3Dm/uR54xcyoxrfSzfruOGWuu3w2VQP
QmPw6dyJym0g/SbowRplJpGBXAaR1OIbsNfwD/fbizXSZY0sz26vziQ6lJbE1i4/
bkjQIpicyIy3wdXjwj9SrlXlSotgKmjOReQiEiQGCPCMnxc/FCrJatIUlBveaKaD
iQ/ex5Zlx7l2gSE/aPHuOq+FtBrTaR7a58NK9ewvAkIFfDqeo83XtD/Zi9+LuE3W
7mmLK93Q+QhL+Hi7ORi9kQlV7N+3nGE529Cp96WpLuVNpbAmjSJWnSWJ1YzHsQQq
G6TW8qOCr82m4bgNFUwAHaLImQfYuOXFBnhk76cit6Itkf20611O+NlR62gdpF9T
wGJLelM+WW2BpTfKJEkH5WJzkaPLRDJxjDu9SDCSodUEi7yEqWd/Us26X4Qmkd7W
ET1lfNx1se0lxqtiDEtwMB4dYeI9Bpgf78CuXsFdQRBAeI/vFjuvKK0QjmIGhWH1
pudUgnrM8OdRiPsgJ2PFJIJzchuTh6NvB05GIZxrsBT/yE+WaCS1ImOSptHSm0TG
I4ovyZfiRmmgeEHxgef0kquOzIgZAbO3LF7oyOT0GWTXAyfQF920/SEi0bw0xSnn
ixWFemguNwa4oFnJaBlPmXKX9n+MzEbjNqoHOTX5d4S+bb0SMu2g/3xCFuqsGsZd
yV8diYx4skWRcFxii5ZaYVdORyqkq858zTXDR1gp/yzdVrvtaldWF89dFx2nCmDb
JepgewFR9ihiwjhufJ2fANJ6lRrM1fPw1i4Vhy0OtI91k7CJou8WNhBknUluknts
3ZZGnJNKiXyohjgu2m7jX0EolHKrvTZ2wcIPH4+Zcjrjdc8jTotv8W1rfJM9uLCs
d4B/jBxQjQB0GgPKcwWMwCgG9LprPCcDe5evPVg+As+EpnocS/XVcO0pvduWfCFN
avq8oPu8AT6DooOIJXmPIHmxNDujznakWCwG1ObseJ7pyER3yhU3hfw1J7V7GkpA
njf1gxirbu+yneoMZFyQlabC5BIS9wSg38lnk1WZvwYBidHDushn/7p0tESvPaue
mTC8yH0AFMnGEfxFmtkr3uhb3+NBCSf05TYzvrk1eApyWv/PbiMKSDlRF3mLctLl
oSiLk1URKto5gX00u/aIYAzcAjprHBLYcEfBUPMRTQ3LqC9AJwl8JQd9hP9MUPxR
pjRUbfaD0r5MDQH6863xkzCpfei/0qygxeCPSSrU3nRmbcDug1ebGqey4EB//+F7
EUpwSOxbaLFYirAi4pcoWUogGKwPWvyKSQo1JmOs63XIdu8qZGx039uTrXTFmEgf
Xn3GxhspDuOxjKOHNp+rQd7aD1T1fK8IiNXJdhKC9K1+EEYWlFeisWCJAykwOwII
0Qr5tuJWZIjdsdsITuL1KSX0cHnhdpExfcmLxO76VGjjRFJXIt09n+X7hA1Td6QY
iR1EazyZGR7XgzI9VLtF5hhlznPV/FIYs++Y87QIgqsEtrjRbQllxrn+hXzcmzZq
F8M/KuSZ4OeukvxNvZAv8rdBfkyhsGPqOUrdmqspFlhL5nzSS51KkENxn6J/wl8E
5ilLY/COau+7dY+/5vHPZ3YVSNFaLh/w32+DTAZt5jTChJCgRt5rOSfGqXwYNtBc
hwf6tQpjdTIxtARfmKKCK0AXHt2oWjcJFQAFFzWLy9D3ZO7k+WFfn916pWitJHOC
Wcs76pI93i3X4iTGTpA8e0I8JF1rBhw5nF1Nmk6UlWdGrf8X2ZZ3uf68VyfKGWpg
TsBRo+MUsGqXcjbt7Kr2c4hqOBPrMLJVlmLzoKr15wOSZDF9ZJYuDl8GFLyq2oc9
YjMWBkDfYmIfELD34ZwJKSoDoNBYWAS8EVFKVfkvDRfwCTv/1LswzL21aAd7kxB4
x5hSo2IWhKWF/M6Ov+QIPbqDhDXfI5PE2FDHoLCLy7XOcjAHe/6F1OblACVrBVSS
alPn8zuAqa/wrbf8ONeqz2djHZ6O6bfQBTf1wnHl4OR4Ym1j/luSvlykdRoU8k/f
BJ/3h0oe1HXq8oxsUxM0svn2BtffwRXX4kpfCpfvYElMSjGrPXcj+QgDxye2sjK2
3tsdvIvW2vswhETH8TAxNH859SYnMUvtRSbDcAvdlxlMR+DutkYYnATMgoZ1PhSO
u00Jdv3s+bZdXyt7v0BRXtf+1SYRcgw3O6/CF7WRl0uL+yhofpFA99LGKqqgfYI2
HDCuKNzAM5k5VHLnulJdzHsbaz0UKiVhU7PSzqpgkHadtCNwC4k5415h04flrlaw
+fN2FVNHGXNxKgNlJKuhKwndaG4KXOJLcYb8unFUQ6VM0W48EeC4mdwxpgiDGdFJ
DCNTyD43c6DZKv9nl/+fH59E1Vk3LLqAe4Pft2t+RqNpzJwD1SXzpUF5cfcC/9I2
+k55pGUTjJKTUnf7gpdq4kj72j8MGxIQxRKD8ROR6Y39B8wb8hWy/OROw+a9knHN
qkebbDNBTwfsBUNS6vHND/JX/kKU7UEABZlVyGSmSAJKoS+iUIeQFs6VGB1TNIt+
JcVF0PhAT/FijaodaQF/PgVBMxeoDICx8QKNHU6RhJ8Nf00i26QjwRCfmyrMEDoA
4rpTyIrQwOkD1NU8YhEfmIr7UTcubQB8qTSfdnIduqpgGyXYYT0gBBEOp+wwNxea
BnMftY1MDT83Gybxs0xiDzMBZot41b2YOLr3awQM3D/pK4AVeSKDA8vvxq0yw3jt
Itj9cS5Ob1WWrM2EYvgRxTs27GGh5KZyPNv4dTwZe6q3v5wWL2CHTSXSQ4xmKs1x
3mXB8XPAcvq2HAI8JTBCiwnQUTqw7vErWvnXTh/lVMAyz6czI/4nJcDy+tv96iIb
zBX+MRES8I22LdEE1bpVE0iulza8Pu+CmFndNsxV736ucde0KgrHNYLuHlhAOHvI
qyUcGmvfqk3tOER4lcj43heQVg/2/RWNF/kPmpv9ZYkvimN+iapHYUIsBMZQyErd
uHtuFaWtfhg81DOUkQsZTC69T0Bbrc5ssdxE/Pb0qgB5LVGScIsQhEAzjErvHOzm
KcHI/E7wBP8sHR99lWgRT25pS0I+RZqmxjUcjN0zK30OUr3xvcKDe6FIXTqV8Wgr
hlmYV0ezUbtjWAsD8m8S/5eVJT7ssHq/Ttmr19p5WPKO2HQ/dZSvotPFRhVWb/do
e0B5sUTSvxUhSEGvF5WmzC1kt8eVLVS7JdFXmBRWM+oQpvlfs4CpBd5J4rqPAxUL
fAJLAZCiGNIF7Jc6q4Oea/UUBzgVDlR0++/nglORCmYsjAQWoG3aUtHXIA3a73ok
P1DCyVPTKIun1pC62JQj5BNb8FCmbOOwUo001jcvlRsHkEpyE+KPYJyfen+xNGt9
jWvqvvS/aAs4gklusRInJEByH+8d3CuIWqUPLiFIFmE/xxY16aTakoi4lkBsGBlD
HzTfnQKrFfnU7u+sZShj+7iH1+LHNoWhdTWsU7r7hC6cL+bvBWp4j4jMT98Js53A
NHiflD4OHjMtMGYKhB9mcN+BXWnBR85XU3ymdC1OD5Po8c5yUFjyt+QtATlU5BwX
nR7gnDOeuCLiN92aP1rXh5+iIUnXx3p61b2qPASVX70d1Clt6MWnMmYsYdAqr40N
clalh58er1LJqt8nDf/kD6vXZv9/ephBT8W8KMzLWt9FetOktPE5IopLqz+lGPvZ
t80OZQekWSDEQHjnTlU7YcYRXYM33O56V/Xq21KuPREfXSP35iRv26Xc4QsTRZQW
emcZtaRrcBLMnq1cpF0pYgPRCevlfFOEdJPefTXDaZpxAlxYPAkP9WsiU36xEwKb
65OW+1x0y3fsI3wqSLAWT3/4VXtQRyAdnuPANnMDgSQ8g+/HTvw4OEx+sXuIqRxi
8r5IUeAy+9GpRV6UX5kLodXyis5YoqJklpF6wmfA8ToxDHEJTN64jFUlZoKtUWXt
ZGySA2QPJP6lu0WFt0+mvRdEXDSR+K4oOa8lYThcAX8xhTWj6dHjjsuL1DtFger1
x5mII8SO+kWQH1/DvV3DBn92V3lJyWjKYltTIRaB80JvL/wHHijcyVsfqyDC3lre
ELu0rI5G5XOIdNrMFcptHDI7GUr2Gx/QMU9C5yFsHQ9x0tOkmLw46zk5FsUlObZL
5HFci7pJARDCaGn18AWZA2KYxybZJpXdpD+xBp8payOl03Cu7HpcH4r3quQLGTYs
Vi2uAfbQRwGXbf6TKwaHdCgTYpVVuMh/BzghZKiKW7Y7sPpmUezdTV31oY+XxkH5
PcysJ8c9+0x3A1RIfjLMRulXoyx3X13YoEaJzPa6A0PU4sJvmwg2Vi4b+CkKO02C
j7cqNUUBNL0tz/RsMe+WNCZ01AJPHdc3uy++3egBNPs5/ymlgTZ5BXgIYmB9MbHQ
8YrLKalXCuv/LgeU+OfpwjQ7kPhqLixPPkGwGMbampT/AY+HehXR5UZEvy2nhjBf
KF6yA+8VBsD+oFKUmPdDGG1ZrGn70eVRtQLXv1UYhMmoQym5dG1vTJPVOPqOQktD
+AL++okp7sdLY1GRW6aycMFjaVsje/5kZEGyoe/KtDQsZjRtDgweujMRRSunnDz9
QdlUJSVqPm4HJHC9u/+AKXn/esrbshTwxE/yC1scylNVQ0lcGAe6ETvpkr1kzGSE
OJbqBNSq3xdFX8l7FzfE71Mjub+Qj5aBbBRV0Zk63jmIFyenOJ3NkM3uRplOFLfz
x6C/XYrHlhsZxsj1fvuPx8ScQCTq6jhku0l+PWkcRdTH0dip7qqzTtPyukPRd5Zh
PyZpndTgxjtOKw4Uy9YtRiVT9AOawVPxMRhh2aSF3d0XhEAzmI0Trl2tZXkU0/cE
WV8OkyPov8Jfg/C+yJe9sblJ2cF07CunOffif6pca+/CoPBj0Kp4JisIHOELzKpa
YDb/f6NC/MdgtFnFBBADSgsoKAmesWLHFQU5tLv1F7gffdkgfQKE9OAoiMnGUGn4
6A4c8UI99FZfocPktQL83hAx4eJVqMeqviBBFTKMAW6u5cAkUOepIS4i8/xmMLmy
qN91S0ljt40JJS+9On9HP2aDheKSbfGVvvxmk0n0ySMV6BH9RZAt/J51Pue4xHXv
xdzQo0bbnWfd+RdKODhCKdLgEUkATDXdZ+5hLpK5+ZujRftQpklgLJ5irCf4OA0T
VqgTasPtw8aFZ+O7RBOIBneZcANruhMqNNOaTnHIoMHTBiu1UfnHPQ3SUfth9fEa
mHUiCc7LskMF7eIZskfqwu6gcm2RqFDC8dzvGWbY7c6tQebQzul9IQtthUgY6HNg
t3jTX4o86Aj/iUkDhClNPDI4jNqW2Nz0PtQhe8Hu70Yym4rLiPWPl9wSFAtWI0b8
0RjjZlezjqY0vFHF2nldhpochOJr6/y7LPNem7vgvd+zmrd3bQ58leBVYXMWd3BQ
VlithMTfPdq6cdQK8yS16YXjfpIEkngIg6qi9gUIcu5wpz8hA3wTw+DMPpHIja95
vFxZ1OSkoicI1THaOrRusPQ8FnHjquqUSac9M+/ZC/YnW2tPTCkpJYatziQ1xWcq
T7qy9Uy83FMyrDfy1l7kL8bmEEri7+gH6l80fzUOHvGWt+IUJVUB6TSv+if+xCPA
xBTUGdT983VGK78yRhUDa4Css8e92seVVCbtAyHjVXqtDlyYAI3YisB6eQpCO8Cm
oCVnfvsvI1VZYqa+ArjPwEgdzoAhAakmz23t6xijvNUh6Bwjdo443n21dkR9Ngix
xQI1gOIs3H5TpJTNkoauX2jKpher6cpnm4MRy51VhpWcCFOD0vswi6qXQJpdehcY
v6ld09+o2/O24/f7ZOlankMdO++1VSNRYc3s5DPFdvyW3T69bIS7du3xtMBRzbe8
vwyjaLoEAfnd+tm7jWWvVcTAUG8HmudXPVW2GaQkbZ7o9vHr+j2+XEBC+6SnUDDf
9sWQqGu+pW5xbhXyX9Ofl702mDBC2JfWqVwAzVAhjCfj0TLKPl9V1NXsVPfPJMCJ
YGPiqrwaAnTsAicJbsRWRT+7NrCd4KFibyeLdNeGHkLTI2V1r2RGdSm+wxIrBobr
6NOWEuCI59lekzC288bB6Rt1h87GxJIWaMnjFUEcyaVtVXzKuf392xUAk0Mv2c2y
++vR/uceCQwTAUnNZ2EKzGCBZXbrmrFhfKH/qG1gAwx1pTcxHAsp66QU0gnRYujo
jFF6Nu7I9giVTNHUJivbfoIjGX5GC9ueocD4Vd80cSp927ukZZZx5Ks/3MWLyjdb
SfobSg1bNBCwbc/ALup5KxyuVw2K0OYMSkbb06SxK0xWam1xz7GqeKqlRhiNU/s9
axLvskzJzYSdf4r8Sefcw1Wumqg3aOloAN5vqYol2r7kE9u73nISW2HLbe0KY1Ky
Rcc9D9xDTWcFjKlnxvpYtOVWJ8Kbavj922KoLXRFpydiQfapVu8Ge0i4eWAKmLOh
XcydOZ/3oHpqI2BOERZCLCBLqj+EjjtueamVuqqGd19fzB6Jc2WWen8VqJ6cOF0Q
O9PM1gXPlMXiWGFMZjT+pXrEK88MvFBTqaVOhjIKpR63LYVJypkBY5tkfa8hOFlp
7ySaa+qjIsxcaadSqhHRAV+Yp5vMRAcWKDBqVNhLJL+T54nDmbHJ3t1f29tHTFI1
2+/XVIjbTraecLi78pFpoaN4+2odJ451HxdpeMVy95JYk1TQI5soBQ6jfawuBj74
vCk2JAJWG4Dpj9jUVArsT4ctwJvzdzlWte6t8EwIwwhUEG5Gf90pE8GTva3eA+4a
x/m9lMKxYrJqgh7ek5GJrS9sVB71Aj202s0hiMOkPyT46qq31YjQGqgSv18MqyZf
j3hxiuRM58/+zKNHCF9q9JcliaWknahBxxwRD3h6oapaZvoAD0c4mYsJS28xmU3d
ze3A7UtfNg2krjJH3ouIkg4nrwh9E3IJZm/R8sCiDIhrLyFN4OuxEobrFhPsOfn5
zmW643ICnCh9tVFqUJJsUThLzU5OHasrCNLn/aPBqA4D/QO6u/vUDZOB2ZFxt0qu
a6SULHq42u4wMLr0zEClg7TPduX6iDtNR/KuizasnFCUOcHiilUP+TJs+CIwjZ8o
lPs8LvcSeTEUFMBieZVpbK20sDfsd+KR78rsqRvk22zErJezvTTIG+NR4/AlNZ4i
51GTv/Okeh9W2USrJqEPVL3gytiDgZnAiioD+ODdDMG+leLGenlTyYVsar9AGVPK
29bGO4eCCyEQqnhPy2q8DOrZjP3onFn0hz7tV5Uia0CmWwQVKCh7nK2d7xNy2vYY
KtzqqR85sQIyHqbFyTYsIDY+Eh7ksWEQ+9e5KgVk0s+SUvpxPv396HKCIbzbtIee
IlGSiCeryvFVCiC5dZq3c8b/C0eOkmppXhXjFz84xgvwz3OCUQAIvX42wiHXaZ8n
hkg9xc1/mE09INT7bwDKQdppzJieyB7mdmnruy687qXVMlGYZDc+I7yQH+FZtTb+
5vmegEf5FT1gAKD3qz1irLhRsu714Yvkvcq2jl3SVfQzUdf0Td8bhuFWOmAeaiuT
3/jw8zW0gj5o/BOPscAD3M6IF9dRjC6RIzJoGf742fGJWho95pHLfJhoiVYBP4st
ifLQPmVKEmJN0xUWSsgMxFBAZC4U21gtsm6z7SIYBx1MSh9MwOcO6eA7PsjIfJHX
wu7ORMRjiKnviPmGYuUYNNXFflPkPD0jmYgFhuFEQ4dbV5zxMwbrDU4EhN/K6lJ4
XGq+/6VvqPiKccoJb6GQVX9DMJXniNMRNa/dgDUeu4vjICEDCgi2eaEW9BlcBTYT
JdzgFNLZgxeMGghhZfooZv8nKz4p48kg+gSpg7Sti/4sZVW7jPclQPbiFsMKOI5c
PLGbyAeCOqCYQFvJR4Eog2/M/voVa8nL4oHjL/EOhnP99xGusY1efrbbLTv0dT1G
AXbPshA7pV2zdpXt739FoL6UdeeZNd4Dl/gCR5IYK7u+yALSN3SS0ZyWIfvMndY6
le67WQeF8ChgsDnrKa59SGe+2cOtKk4Vvgw0G2uKxSib0aH/UGQx9yrZPFQhkvwx
F9iksbxraMAbmriQjZBAmJ2lveKx3Lf63mwhs8l25AqqbMLYov7I4hTjD07Dj+JR
ykA15TrgzbKRxmMn56qmVhmEUNW3/4KOPaPiCZovS7nNam+3/7WDroSOlLZd7wPl
UAI9h8jUym4p2sc2lRFbEJOarxC9u5iL3JQBp3UpRrHGvcmCiuqlMDnNNT2Fqz7h
QgGFKaICtiTp8RqW27UQfPgQ6imNyhIbfP8GlyYg3FLdbhpXN2ApJW8sKSI0ewOx
vomAqsjig+0leyPDJWC5lcnfzz6biV0hN6xmPCkPwV2TqWpvE5gaBqQr+NdYawc5
xWZ+mwNL4CkRExRBiZGhRtPuG/fEYr39wOhgXImyRAKBV9afPzqRWp6K3vB/1hci
WF61N5QUbum73rQvcqUMF9Ln0Bgib9dUeCbRgGXOKeOvyKAQbjLSF43uEbYSrQET
MIQ+Le1871N9V8VBoXXfJR3nJyUHyHLyz1mWlulrCUkeTPmBl3b4uG3MJ2YjQAeG
g9FSyFJshN/PRfo9yThvviSv/xztvEJ0RrVWzJR9kl4i7o+EKFp7A113g/NPoLpp
0o6Ac4Wo0DvWLXSzFIWaRvE3bRBuuYXKKpdJAQu1DcUVf+8PL+zGT6/u62GUJ9C+
9YfhfA3cvzIHGFKpXbQZMJl8mqSyFqretkW/uWW4IQbbGT2uf1AX3gEL9fdZk6gn
6Qe2hQ22O+qeG16TJLLT68f1oPithdRzPgGE86XK4WwE8VtNRDfSA2IMKTe7rPxl
8ff9XMexnpEkGLsp77MPMl3as++HOWQWn2V7Er1sKnVVlWdvxQQGbSdYERPtCwRc
pU5DsFz6vtGv6jSeMG6KWqalqwBKOk9XSQUSmPDeipLBJQdIuaqCiCkJdoUBmg8J
7g4FaMv7JdTCJgkxSPMUXHDA5viQB4iyn+MieFYEE87uw3ew+BpMgoVv9JOhf5oW
qp1OCQl+x8hD7oIovg05fqJu5YD5X+ZkUPy1RLlqBla9PgdMGuTs/nkjwBs1srii
kwsV30lenQ3JTXFy4BFiTe6++ffXEOlCO/N6+3sU2zQ7fwIDooehN03Sb4AMVVJT
H4RfSJxchbcckda4y5vGOuLyE5rcAeYvbR3X+DotuxKs3Qg8Equ7ahTUmHZ1Tri+
++ulzoxowwEGTIQhgv1CZiVFZcIbxz72JOlKDQgHsCWhtJPmNh5Qsh0E74uechYt
3r0+yksjU1ZA+qi6fnv2XyeQ9L1ZPnAlIfpyqQQwNfi7D2+VCkljNxq5Gztj1XW0
yuv8BwljUAHdeK6b9GU97s/T/oHuC3jHBv8NG4jmoeQvEg+olT35yXrYmJlCF1zk
1cj4m9m/shz5/srgnOkEzWsPVvYqTorAJNf1r5meSckm2szIeUqkzqlV9WcRjfcq
A+tc1pvH77hLwy2MurEw2mIyShCrQiIXUOeu++eWZzgyzryEscxe1QJl7JYhQpX8
gHyNo287ogOR60Cz5Yx/2ycfTZ4rCR1P/D33QS5IlM5sWz3du/y+AvSAOY3RjzGe
tESP1TQMS0UgpAgt+X//Q8r+xTqM7yP1ItnBZsHNCrWADaIiQiHpOKIVw+a2QO6h
LxT2vYI95jRXZ5H4l1rQODpON2U8oixT1A/5WwjjCPucliw61iIuSVfaywPw6ToF
gckOpMF7jWjFDPBLlkEOzHeSffqja+IC0JOjKR6+OF5wBIoyUvyv+ILL+ftw7vg4
6HNtbNPL9RDxyqyrrLzpZM7gtl7hx+xg8pqw8tkOK3k9iDSplMo/xDeI19BCyKRg
TuspglACwuCh+Ch1DKoEQfVJpf+FOCeamArOIPv7EhlmpHQIrmAUqVCQszc3rUgS
YJFsU7EJuDxEY9cCnF0GvqIWVHC+CNUkDWxBNus9ny5ZLjle29JgvhE8s+VcLhQY
QDzvML1fZdUq3jw4F3WBayDiaHdq7XNQvqgeqbSeb33RgWQ5mhFu5VtEqAp1rytE
WAlUI37tKo/TDvVT95vyztPEJv7EsNp/hkJGz4PzUcLANUD7Emf5iF4z6o+yRrNT
jp/ff8QLLiAQ0Ll8e0pkjiF5G+IctRct3HlXHuFbecMfbPRDZ6/LTBNwcLqfb+Ys
Gi3boATeIme7ACBIi7VRtu1tAWgZad04M/yV7Bb41d6Au2JtrKwogY+eN5maAt61
n3o9ffBeQ8kPF1QrMjCqe4Oa/wAQgp1lsLNbJrOQUpxUPA1uEpLqQ+Wl36ZyzlTz
wNxWFzyu1NuRa/fN7MLjXE6VbD+nq6XcUp1921qpGBkZ6zj+edx6mbqMXkxVXY7e
TKLwWAt+/VEg+/+1nw0vekkzUkz0cnyXWgN1sTYh1ndNSY3XOscbY7zuvWehsI89
jq1K1BJFbKl9qVXsgPPWRB6SPeKpTiHwgDL9S/ItwY2cEMouPWK2qvnWHrw2Tgzd
SPsMlKeh2Lod9dpvrNz1ikJil6MGY2lCiDyqhvsiMTNXN8dJjN7xAa4iITLvrf6v
nkf3GqKpTHI23AiYiF5JIHHwwZBXN1mfvBmksVqCFLDRRNz4w99gBmB0xWpfU/p+
plpUn769ixGIBpT7IlCi55KVvhsC1YEuENNz8w3lFZ/FZoyIdGgjLVOXYlQZR7MR
gho3sTPKGp3LVu3qWFZKd3Yhd6WjneFjYF+3uyYklmijKYMKrLxTZpA4NR3BObeM
mtu5hAkEteTVChZ/ZAYoTHLSD33xcCw8Z2HmnD5GtSO9mmw4kOjELZSITCQX2hb2
4OjfuJJWuI5NQiuXAzTrM6Jn9hLRQnVirX6bjnmqbtdekguBBsZLy8Spp0Zm3xVn
n5CoE+jP/6qx3bXG8f2nhwdwhB5pvmWrsq33B1BRgPCNHdeVHY5wgMcsB2/1nTRF
5ChkNbhNPTfSgQU8c7ibY8AFhph1ufyiO1Nr0O918Xt9rb5RsiASN9FEvSW0zC2K
rCULdZq5OUnwElHjXiN5oR1ukY25XOOcDn9cDANWXDVMbYWWP3Y9S8BBXe0hy87h
fJhNvW97gIqPMcrKJxwAPY0LRBU/V5WjFqU52tce3kdCXcKUcxQZ77BoMh5xUat4
qxCN4hWaFbIQi8TcSifA/Z9BfZH9TaJVP1SSVamd4IG03+3ggUj7NIRug0bAbdLJ
YcJH+wXYZDBaNMOXvnhJ37UxAhWzkRGZJ5UCJzl3xtq3bssW2B/KmPqZM8sXlVBm
QMFEtGwWzgpas7TVSDdDsHH5zsqxuFylh7SVbXDdT0Dy/ZBxH0fNPisiXLNQp7/n
EqwVWf8vIev41zDyn5TfWJcQtr89iT5X9nhORbFoXV3JlMOReKsg68mYyY8FEpJw
N0B0ewfKqmWhhLnY9iNe7mWi/DMGTCJSdKHYzZOQQ9DS87oR63FCNMMGZeJFuttF
cmOEfOTktmcVse+IqdWZHCJcsdGTT2ZyxYt4V2FlbcgAMacjtwpK/5xc2yaeaRfS
GMzuQ6aKKcfH427FAQLNr2KgFnUWanoTJ/mFSz3Z7DMYyarF4vAHeoNIzguxpul7
5OtADN35pUY/0FaaT/26JPbUU2CRWrRkvTwUPrtFbNUpcTOYI01Bwo9ZhZPRR28T
eOKwm3o9be+pX8k08tmBMVXzQxr6Dl2RApBvuzT2gDkop9/HWJpbcBm1P+qOY5yG
GZ7XXD3UHFRucNyhorcmmqAJIbYfc4bgiNRdG3H3cdzvl+j3sh9NPszCYzsben6I
RJJ8fKZElgGfV71m9JAErW+pcdFtJzlbYzD/ZbBX/hZdgXz90LKM3UvRSpT1M8Qm
fQ3uO/dpptqUdr2Fnro7nHG9b689pDyJ1mVMhxM71o1uQ/sku9Au+yZW6DuOaYri
qqBJ+ABuaEB/ChIVNtFuJXYzvbr+tg2EOZBMqdELluqPPUx+l6x6zpdIqec2K5tL
3dRIC1IQOFJEZVVj9rbDgunmhV2Vg2Zc7nwdzECq781GV3m1xpB674jMpx068P7i
44Cz8Hq8KARNOKFcAyoBuwqQQjxRMobllaQTpQqi15NPUe7p9lNNnf4YBdm/chiB
iEvllZIpTrEaxGtSGXwKNwDVlkjEDe9/IH4GzjNSRHW65e6naNOdZ+1Nd8LcTfxP
FmnePyLOOKHI2ILU4Xwtq5VQromDDGxNfjFoat2ndpDwOi6Z4e5Dr//ZN/AQzsur
4UneJZjjjS52IAb4KTZ1rgvU5RDd05vfbCKpNTNzz3+12RFVigC0S5n7v/b+6XY7
k9nS+wQamWOPWkZc1itYtMNvSeeBmSATmF8t/g8K6/M+WMcNmEXiSIlOBB0ZDlmo
TrLOegF99XN+AxA0we/5b2Qu6no/VPbLa1wzSScaVySMsNAkxpGNbZddlbKWmiPg
/TgBe3i5m1ZfcEl60HCOPeo9H5X8YVlPVgEufjq45po/3yacX6vMmxD1q6JXNz0u
R/FzNFZIuDj+4xOClWWo/Bzwr6++p9x1vxdX0kflOuTph4dbukkD8U8W7Jbxj0wS
jfcZvd9VsyF66Mo7A2sIcgmaM3E9kIil/YYWo3gtUwLCJvNV7YJWvbxfw3OH6pMb
bM+7IpUT1gzjKm/6yoac2VCxcw2qXnutXB+W8jbQoqBJRZJSm34z0fOuialGPa7R
rAiStHlItkJW9NRV+MtzKfuIyRFcBg9S4oO6mhCPu2vn7KvIEZpnDkEo2r1v1sAm
QeYCgs7ATGYphSKjDBAuKWx21k2p/Dj2hf/y80FlLbnd2vTUeMnK6CrDirXMWCo/
5LSNKS51+f8H0cFo5r6hglR9PS59mOjtk2neB8oVhFXzHD3ewF/IIGL7ZM3ZniD0
BkYSNSX2HeWPT2+nI8ItDgcjZutkFDzNL0YnSN6zPra7tN3QBh16A7HYxJicUJ0O
w2v1hR9mg1MBrmGw3invN9+ej8eCqWs6QLpZ4p4cetEr/9CwSg+mGOsgZlMdEYND
mo4liYJpC5t6pK9p1Ylf6FVokr8PgoYeZZ/0jLT9Mo6hWufuTylM4leuU+eX9/04
au8jTbhs4Kh3Gl2g4VVXDBFhq8AGcvclOkD4SFKLaYoPJ5oXK92ew0tE7qduSSdi
aYBHHrwdGZA7V24Ut5/bxOHXRFvVs7W5sxB8slMlsw6aBvCbAPCEOys0qo82e2+P
fWDsib1zzIEzVAYFh4cgTL2G1mYAI1wPVrf2lp0bP2zBe142STVRxougArgaIM9p
zPyVaGgTQ72cv7Aq533ZZpzAXSvoh0jYM/K385Cg+4ZBkbVk57S1dxxjZqab53nT
ap88m7Brc0OK3VRnrhRBMVujGCUEFCUn23ek/yTA14Zjnfs/Tq2kxEca1DQhH1BO
+FIIQG+lCMh2lGmsGESuKhLSTbWKCH7mHGyhzNxKm2lMhCwitYCP/eYOUQtILgDs
qNz6LoDeLnz8w6080TGPpk+QJE0pkqmx4MWv4Fm1RD9YoeoxGDMOElchAi3+83Tu
a3Pov9y7YWdGI8g2gTWA3V+9QMA3Fiv4MWZ/pXPGl8lCcdR69cHMuyiciBu684UP
uZ7l+8vzhkbIBrR9gdeHI49FsDUKNW5GaCqBFLW7Shoyy0bVyulMTkuUHso7i628
H9IrBlnVViYMyw6gmUZWH9W6D+xbonxhhPKjzR67U/2E6IN7XjG1PeON/KMTZPcG
eyYvzVhu3CZvqTlQsq03n6u5S2sSsIpMgLhg+at9LSf4MwGrGVW+0vpff056Lrzu
DXISDYTQMeo3e0SigSSwMh6X8fM9uV36Gb5kEdy5LlkkKfCJ34AGbfMKx6OrPj9e
AluNJDiUQo+1KC9AGKm10wS5zPOCRe+ol+lHuCqcXRFiPAqfaw+5HntXN6/6i1gC
dUhoDeg/Y4Mhto1Bpkk3Na8uOuCfoyRhYnhe1IqH3fMHM4e8DwJAcFtoqxSMk4IJ
m6WdpnWlCfrequZKPfrFGMimGRCv998Qq736cT5RkEfumFhMLeEgw9UNqu8N/6gZ
gfnTU1QBi1jiqy+N3DVuf+BmvebhMj7ZF43YR0jsXm/qBm48WJMX2bxPbqJdpstg
K+aD6ll6AbP6O1/uHJOGtZepU49Us5Se/588jECv9bSvuIHTK7KmAMk28OzUBOKu
3mJfhurHkCbrebVYvMdpgwaPnAAO1mDlV+N9VYWMpUtSVSFG50sbK8ullRW5ETnk
w1Q/Qbs7xKogiFPL+RslNS635KELOwJ9mVgAMdSa4uwUT8oNtki1hLzY01sbKdAf
CBpr59t9NH8rI1H6XVssEA0phOeTzSIABg7BVoRmqhAUaHtnNNhhudTgappyJE9F
v6L53OBKRvhP9SjukHBsPi78y5/lDkWJLULrARQ7h02HX5emz8BKC1AwSFeWMiwG
p+xgieM2sEq+BDXsJJKhBdTVtLTdXNBucnAQSzbkHT/RfRL+mDlc5aaG8spTtccz
tyffc34CzZ9S3If323hRoJMUO6PgZTNpSiBNDjakJo5XxcwYb/jeatdqnQxMEbuU
Y8LxW/O04IR3OssGRMan14Lc1Tsd6bvW3UbQZEReV24efky15AtRi+TPxoMbSqo8
cU2DC0MoSyAr+UuYH2Q226OmeUJvH1fsX7Ln9MV3l0gUA/YoialtX3cfPBBFENZB
fODUTHbG4Hmj69nT65gvdtTOmNZcU2ntk1ehaQ8h+7+gEJS00wlnRLFKHpOsXMiM
qqiccPlKZPYln4KjEhfHuiRJ1hV9YXiBBtihQJsM9GoAjEd8n+7Kdy5+9g+KTxZn
74EpKWRbJGYlk7zwNGd5dfn/hdtFMtWrE10Wubsdov/4WozFgmMO7+OQa5gujtjx
uTgOSCU+5DHbGESlfKovV42QzU0S5wP4gvEbSe1HC7GRxY2oynCiaGqAIC1fbgAE
r6BwW7dVBpKaJSX7Z71m2VUjuKp5NTHn8szXThmB5SqGg8juQNJS9SRIVsQtB3cy
NvyHdQZUJlOqxY1ofNcB6tHkMk/KfAXjEDWVw+OmErZobdFrx5RRBXrhum1+2khN
4OsUiVOmXXsCjtkqBY86i1qtAIAnFKuMj1XRO9i07fzWZ16hjtg5AgR4NDW2HAHw
9IvJ/xwbBMoR08pOts39H2OQgUUekY+sYF5iD9nsudaEJM/vrXckrTbrHcNu5VSa
TiwRjKBgnUjNUwaJMYTBv9a1xBn8LUR4ISxaIyDraPhAFzE4UI+10hiXa56b6Lrk
+owoz71lJX6eEQQHlf/UsTrW1iZcsSX+FAuAYcQ6hUY=
`pragma protect end_protected
