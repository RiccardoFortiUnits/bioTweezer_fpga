`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ei/a87MqUUlxXvg9r+xbucbQ6OYRm7xMHlAS0w8Z9Tt05cfC671SGfRsrjyXzMPe
YzL/7tPmeaSTCGNvwI4M9nJajXMpHZkDpJsXpIORdah1YlbTHWM191aV8VOlUXoR
okM0Q0mrwWRYMbjGvq8uLWaQG8B5yaCpgeFMcKu4LkY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7216)
i32AEWYIGEdvqyBwv5wgapMuqI6AIvCznmloKxWAAcmUmK+F9x5fV+OS8yrck7nt
uJOQ/rZZsP2XoczpzuaI0PmkQlQVbN6L3D9QLrhsPuKtFVFYj4BZzaxvlpq8Flrk
E48wc+gK4ZuVfMQR5IHo/daQ9k/HXvxmkKPQQ23bi3SQwDDo1q0vsya2jnyCZmiq
aTiyYGFV4ShzM9tckNAl3nrjRNejYFgsVHod174i0uyYTIrkJJgRHOAfS3Gyq8cl
FfE0LCWxNLQsL5AMaSsLISHyCxmVQFel2Q/+BPiCHMo2xeqsIgFs8WqoetjMQ8et
W5TwvCyXDS2aOJ2YoHthlTbxvJM7g65S7n9/oKYJttp8EMVXI1GJLLEk5tTW0wiM
tFdifUo+u5l4nyUY9bYFAoMaugHYcbna15Vaoswt8tCCAdiOIamEtwV8dT6z0lOs
+2C0/0Uwn3iignGw6L47kT3P0nsvHVPNzy9pu1Q6xykinenMCJAe3Ql7JIKuqopP
0hioEPmL/Jg0eDV21K8Wob14sujYOFBAnW8F09Xe13V1k/dC+VBUG3NhZah2bRPt
v8HjIP0go1WPfU/cJypKoG3qmnPOP33kWeA5xTJUaqUA+VsMtas0OISi0ohsjirS
7geJw60tPYLRT9WDeUKc2yRKTwVsqE+HxPA5zMsGWbk6R9eerFPhLu8leuAHkVVP
HAT199NiMxfftLvWpjjOVbKTQufjaDV7npqpnY3YyTjdRmameP6ImMyra0epFhhz
EQoMpa3/KBMiOD3qKEQcAgjJVSrbh8ZHLeehkhwkS7L/1YFYuPCIyVs3rCp1gql8
gO7ULKwO4hsWLTowmugzERzolC94mG1wcMw8pIFTbC6Xomqsd9FQbbDA7MsXTfyh
g+OmttYnP4R0lmuW5E/M1yK7zgmCsrQUVQ8eOELxqg+U5jCmiZJRiC3MBdCjxPQF
CKnBu3wZVWNws3RMnCaujNb+pqPdJO5VZ2IQaifwsKQS89Cp9R0YAtiscFurwDSl
8Ya6+9R/TXE53+J4BsOXNuYUK9D52zgQ3lILN4JF5mLWnp630Xc7SFbGgtOEBcQk
gn2TtwKHJWSUlsZF9cXdDXETnDggFHTeAC+5R6WE7M72a5nMFHcRgPEzLu76M9c3
qRPz7k/uZ86DzHLgPTVbOKX838bU2A9SPqzNJ5DGGI+8S8Q+Wl/mXJUTZR41GhdL
/Z2NGx7/Ew92K4D1bAb4ZAvfBIa1ySL2rnV2dCFVc+lJ3H28/Iucl7lHOqdWm0fL
+b2ONTBLDmoc7XSU7nT5Eu5qBBjEn24qU9jY6rxUClG90kk4sKMzHH4L4Jl24SKe
GrI5E5SJ8fKqwU8RymWugnQ9oqIuFUcdcBqRwUitYEPOYXoy/fJIr9uTIHOzm64C
mtIgvdHcsZSoXerbDcVGdB5VGaIvn8gbQE6Z24w8vv+Y+AhAxAwjmpn920X9ra2M
zXPV0ZBlwuZCLZYssLFDfXRQqGQq+vUzGP49CJvyhee2A5WM3/ITRyt0tNmUbE7d
bOtSGKfcmkK842Sp1X2niJpcGpRBnfMsf/qhVXS9ZHHEyX6nEWVv+wZtBLYCVhrG
6Nke7hwi/6Iz8u72sDCuryqRZ4YT2BwVa0KUyChpq8cWsp3dtzPC7EVDn4PhAzpT
ugC5uuMqn6oiX3zhN0NknccZEtXml5Z8XUR4mMFGMIzLzAS+yaYlpPXBor3WCXeH
Wvrvppj7RxMwWiPv1K/2/fcj/k8r9l694sGvgjOmIl6l3eeTFK/7WqkOFmid5jVE
32sbo8czGKDKKeMgP2suNI2/pCsND8rJ3Lk0x90vk9NsPEB+jyVAOwIVSR1Y289R
FI/6fw1QBwEDbnGPTyJbBeSQXNEBJ3s6W4G21uFFygn4vjss4+9A13WEX1EWCZMO
GxzmxPWN83gWo8hcvYh719tfsVy7cNTFes6/NIdPQnfXRzI4Qe4oyf8LoSGQbgiw
C9NvNb7gqEWGgCEu4mjqrF5rcTujdnaCLzNN4pcE/ZAi4ph/G3lnFceN5S2TYELn
O3H8ZJxUuklgn3jdiKwtXj1BjaZXbWNt2t6VFtAZM5jSCmLzA+8xscjkPlrgINHH
miNk2i15+BKtraSw05AA+AVPU5DDYcW77LUBhtWhf9XpqMEeWyFsuG+ik//1BO93
97CCIcnqtnl+SKzdvaSD//dSVoB9mymLfK3FEHHVjJ0zffHAZ5O0DoUrCM5xdWmq
MKYrH5tYZ322AYVQdpfkZLRY2w4iuNAWyG5/NrkJrbtnOjeXmoX0ZS2KVAU+HPZZ
ox3RNyi1OdbDzubVg2m+t/IjWKU6+kzVHjf4pNbm55C45YD4Vc+reKEZjHWY7oWM
r2VnKcpJwd+lpENMqizs3XQzppqgkGmdWBCyM2Qq7v0jb01DA0fb8Sjg9eyQDVR5
1mBHEhN6K4IPyWBRUUorcPMFnbc2hjQwQ9xU8Pgt9iEof+XCxtkQdXQfep3HuCcS
Up3pkaWoD+bMUFFVS3BoYy055NMog59xl/xMX6TVGaW2hklRSdveGe1Nl/8xAbe4
2/ceBl+SeqJlDlCXUzNA8nj6d/BgZ3xcznNt7ZQBQ3S/aKgNqwT26Hm750qHcgu9
WkKItgvxikXHxww6l5gCgpfxK9tZTcludwamo0clCUWwU6uYG+A3N9mRR7cU5Hj7
WtQt+/DteOYVqmSLWrvYwUhCWNkc9tpXAYfwwyqIzi0OIkCx/TaPR7twLQ2Bn1ct
xbZ/lDJt/dmO638ZELQqilQg6/9y2/zOyqRm8s3UPDKLyW0LCajMbp6QdlOGSh/R
g2Om8fI0Q1OuPU35SaOEwkSz6VrTFBUlypJs3qIIjf2N0VVbKSUBxHAbzaexAZAI
8Z1c4UiiZSNnqxaxQ3jLMr+b785feEj5McvGYBe7VDToKyff3dP3rVDvujrGeqAj
0bn59IGctJbpw9GICY/Fq6/bx1BKpacYp4xjJn3nd6jOEJ7T8gyPSBB4ZxF2fsf9
D4gvhn/9ZqM/fC2pgI7omTXWwI4mx1aS3nANqsXrv/HxWS8Yn+cUo8UhmmBQWfAN
fie76JkbivDWAWmNa6nBoh9BajF2qdzyyW0suFh9VZqzqtmbVXCe0n8GgbKHCSQS
yJNhdH6r0AjkedKfdVPuOJubA1Culsyg8Q/Did48a9kwUm5ue1gcK+gDATnSWT46
VWgTQMMEdnd1BgQ65bCBaVZKvxVuMOLf1GhaehxdMaBjESmzUnfVw/iE5LlTWHMm
l1MxiXGSOVZal1EbuvGbL0Kvum6/VmvuXacSlj0nH5lPLjANL5dqg9nmGK4lgEdN
82iKNDRvrEZrp/uY8YJ+m6wWA7Cv3bkSvdnGYyTxND1CGq97JnqPzk0or2cmRp3D
IwiCHiv9yzqByC0DBxJUYq41nu/8mWj25EKyugst+mKZ0KIkNsqEftSBMT3oe2Hk
0ujiRb/RrB7q7jCVyKtiqwPqUoXzepJ80TQ2wvXngjKr8rvUytDOSYr0KGeHgaLj
sW2N/5PrkO2UmevJZNbDho+7G/B1nekkxktJsBKaWRZpwqHNRpJHR/zC2psQuS2t
wBoefGgko7BF3M/yH4znO0rp+Y02bnsdCE4hGEx5Ai0/NY1u+2ZXlY9e1OHLvGeo
u4odUBBpzK0LCxoprUy1LH/57c9NUc0CvMrS5jYwUIDGNUgzzrpUsbZDZFzbVt0l
p/1Q+T4BUMFrn3sA1s4rGa6j6JaKjPUFvSTeN1KqWB5tjbNAw655M73nqmRHp89B
NBrEJ5nQPfh0JuHVdOnA5nzqERO7T+37kF0pTjqDjSsFwp1LVkBrh+0j/gQ6YtKJ
6y5LOAR89Rx8JNh5VzTAuzNd9gR2yXV762pXNx8r5zCGTAKityC2kVQl210xSWef
BIRshVHQXtmC9AihBGZRX8tzQ9ZoB1N46Hak6gatNLQobqtCOUvCyBultB0kGqij
eKcUbCxPt/Y3zHh+nDMeEcDj+IaEgfZJak9+8IpmgoLLLj009/5us1NEmMStOVcB
b5PW95K1vfaV4sV6RnDqomvUI3/+8oT6qKMaqDMK2ZdVmaDLj4eqLpUX8IUPbQwu
V5ie6tEpPO0wYUvRFr9ELjMV95+VEgke59oEgwexYbI1hMQOGdAgY6d3A4XdFizB
kHBeelDDTtRbn+SeOAoCwk8Z5egg3ODt3uwxkRwNgNlezn8ViVeXwTUgqxQ9H9xl
HVcqhcO6+tlpyKEEVIYh4dxX3L9B2ynJySq6rPq1CqsNFgZGzsE9bMEGRrxcYbhu
ICr4qmdszLRepa0MllRgF0arMevEcTCAkpY32gPS3Geql8bhqPvjNLL1WAi33iji
RmGEcjAXzmdUzlvSwAQt+JVkUCmueKI7R7Gxor/eUu143Zr4HqGHuqRs2DlEA4Mp
Z2Pg6wTamBDXIAyL44pE9IRrFTGxFkj6blZ3m3+klsUG46fhXSQePHlK6zEOYyZS
WQdnLsgBepDP+EIjrudi51K0FwLENzYHbUYYCD8gC4CBlVMba1dnmcEWdxZM4XkI
G3kr3caCE3XdClSgCDldIWaMdO724PATRXPiJw0olc/ClOv0Ldo6RLBl6/MjbHNz
WK+avSUTMhYxg+lZpabCFiHnCEbPkLjeNkDn9QoRBHQWTX0hqO5Q+ddGzbXDAgtJ
o45KFf/kRDLxieUP4TmBjHb+EU7pO9r5lrIZkaIpYE5bjT1ffgtrKp42I+NXNWpP
FSMHGHn0NS0oNFcxZ7aR7FmiI3Z9BGqT5sORCm6W59HmdmGeMM//wNSWu8VM+MAP
jrRJWFRgCbnnVgQPUXTfovy90ZeFnOTTiuzcHJhHJHMlHzgivR2obPo3Nod+/sow
mbhoU/LxeeK+R/hSCeyxtR7k+KYLHdA3tSgmSjJciUYgGPzdw7xBhhvmgpY0ASSp
c63F8TL1MNtNDe6ksNThJnapgyZxG/rSNZFV45nvhwJy2p3Az6wA/NpwNzeqcUiG
Lf3wHRQFmbS8BzesCMWolGOWXv20tzJA85Obp9NTkt3f7uivczILoKQiUrUYMJvx
spWd/KnAXwt2EVMHwR/xk8kj/ZWS3uGVBYXSg36V71vPOMeaKQI3ZNsADkA/UOO8
kkGxqKbiz18GVj9aOZzwyDg3THRU0yI4JhTw0JOpPdr3D1wqetG2wNEV1KDSQ9DQ
W8llDXl2T3fkPO5bMW6b3nZtTQNb8CShf9oEEP4yZzRdRXf0QN4GrHFD3/tPEfoE
Ro91281D8p0zcBU8aMSd4v0iTYGt1suVqTHXSKz+NHP4TEEU6u1hO0vB3zvIl8dl
C1GPHXZ2jYL2QI2aAGChCCN2TeGA/rpeK0r2KzPYBbU9DxcRI1hntJdGI5LbQRm3
cmIcRX99JWuqFVd5BRBGoost++xkMGTrgg3tVAwV6MxQRcnJElSpbIIeSPtg8aQP
BP7lb869lRr8/v1dqMvzJjL7BW7+jHeoIidtT6RW/L9Pu1TF9Ez5dSLgwZYJm0ch
lN1KnfOl0kby+RtpjFbD9DeyD/Fn/xQbTe8DLQBDX5NhEAyGAzpysS/nhlfChAL7
C9SkybVh5+SkQf5wF8hxmNb4rktdqZPIh1FiJFZ+PMIBdT7oDTbRZRop41CxdrSh
K6Xz6ac+TflsM9CKNqR2SrelGlz3Y9L+zEqDzRkMYdDkr9HVy5gzF3otL2K5QW/n
czhjfVsU5lZYXVRh3a2/YEGR+CIaKFsGlTwUz0EH1jv4DUVx83IHDo/jeai6g9tK
trTyWkSlQvdauzlsR5ej+hAHv0UxrhcPupTfOBtUhtRESuP+2FfWWXMiUS5DeY4y
T7daoWPDGKIA6exuwIVX61usuAbM/Def6tAkF1lx9WujCMCIpwf9eZGiN/5HhrOx
PJabDwC/u6V6Bdqfrb9UTMWIqBWn+OslY3qVFOI9s3QUNwdHaWyHzjz3I0WExXDK
47v7sbDwvbP7mko+BLeiqoKIvft7QFICUnAz/23T5RlDZR0T4NbQ/7tN3k7Hy1FZ
rvtSqe99gxxhGGpYDkxg80F9nq99xOPuYsz7fVq7wg71l6xKdV+OciBx7veUksV8
CjIX3HMcHE4abNEOiGSWwnZiZOYGEnk0hzV/oEm+Ycj+Zz8dEjNOFYkgRdk7DbLj
RrfU/hgAqUn+rtmbgbnVdL1HgiuwWGW49HWmwewRsjK3e4Goc4oWVbiWyJ17Oi1a
6XOhLgdDkdXjNsHT1fp+eMrWztmuE1wGhwnW+550/t0Kw2NEgy2jDHAonOvnqQzZ
OdS+5mqJqYyZAEkJq6NaboRMRttpbKqA7LBFwbVjZ0uqplOv9i4vDDLnlOdtAlcO
EJzsb6dVz0vbwDP2J8Glz3BCeBxUUfv9SokwG86eHwDm6oKDJlKyi1UOtGCp6ZXi
uwiZbx+et3xbUC29R0gSkyz8zpe6s0kzaSf+/DzdG0ad8BbOscD49SzxB+ycBKla
1DKbgEHuhS/1mfboElbu+jNbvJsD9aFYtme5VOAVfWTmkKLwKNwYZKzJwOACYx0P
a+NLBuVd/4IfwyKUSNYuHQPC6TWrIVFapn7L0LZ49bkj+UjhkOiRfcqCGYnO+So4
guZsXWPwl5ptQNVJNsEswpvpWsTvMEOOtqt3gXqXWAXP3AEx9Tssw1/JG0wJGKxW
kLIhU+nsJWE09oTDUort/QaDe7p3s1NDaowfk5Mwe8aySexKwRh3GnfuNIfBdwkh
M2rI3s45SmotcEcoGQzaVbI5Bv2kfQSy4YCbvRndA1Oe59AtGBOSs6BXML28lSrB
QmgjvpKgGAi3pvas0ASIgOMqDG/NIXgA2Mcz4oBzeJgVcL2Avx8Oq+tDi2lLHh/6
Ko8ae2Ghd6rturNb+UMG15k8hG8ceJQbYo0+ZYt5eVo56VQegEaNDr0UZWwmzDap
kacHPJsGHER5QjOzbSGgEkcuTspGinIl0pQygBUDeyHajd1+zdWy/nmGIjdKf7J4
5cEMdHNsO+iyd6PGHcrjv6iNg94YBVesYG3+Wiq/SakHWrTa94VxZe9xGWFUMmUm
vaDB2fMOScLPvg36bH6AIFfW3p6PDA3Si15/BRBX3+5FOm9USyDClY46uJbMlfV0
SqSF4SQl1xUQ8n9zdBXnRK0S/LhhvfMWUlkEGO1dQcocq7qIWamgKG4aymwETZOw
Q6vjkqTtE18esziZvd9h1xQNZOCFrpldKu0sQSE/PtC6/EoKJwbI4V5iYY4raKgF
arb7oR2E9+T13vs16EQyzCATu1h3v2Fv22j3zGcdm7sB3GP3ioLu7UFwZUbD1Blx
CL3wP6L0d0FRzrz7eKBIk0+3G8aeMLOxX26camphCEXAoqNrDtg4N0JIH/qbqF0o
zdHdayOYjS5I1rhTPREsXYWwoeiLwC8joeIke5amc0aLVZGfQePG/S/c7KDz1iL0
owoZYeuEXrtcgSiPnzlWcR0aq1GGzxgvXRq3rQet6eWR2Z+4buwbAmWZ/wSox7bV
J1NrGKkpNkgbdtjhIWyC/Ztq3lrpLATRCU2gu98Jo3bNtq+x38IBpY5x82XLMyzz
gAyl8hbcY9gaCYSG2EkKtwPACoFDC1UwySlH2Jq+gBJvFJ9Ak6vYRLB49k3L9IvN
9ds0kc+9heIUVU2a8mC4JAlNzzvki6zF8uhp13JARe6sFvyGWSch/dhxzWteazTy
w5vPtMp8IWmQLg2zGKCS71q+nVdiQXwAqSmbYQnqlfND26xj0aAFmz/ogl+7FW2J
7jxPJ0+j9e4Z/lAO4RmVsqFhkoeDpNAwaOlDVqLXkp4Yk+Ub5NaLLyQHWePeYVhf
ce1bIYsZBVJe+/dpqJxX8+/CM7Huc/uq25Sl5rA/om0qCldKf8TTE40y9qSa0Pci
bNUwdjH4IT77+GtFgbh0SApSj2XSCzBh/scoFJ7GvexYV2qf/1b8sZihWs4Iek0n
vZBaVlFnwTUcwNPi9oK0I6OjM9rUEWQh4qYbtsnJPyvZVjXFJ1krl7/18ILV6qEM
/Z5wTAYma6H7JNAMW+o7I+SZ+bpRfdf8eeQEtiwffUd1QxdGvk3cxoO6rgXdRbEe
Gp7ncObVDFM92+PMwtzb0SPDJgiOm/dGWEEncFxHMW7DSsUuD9Hkx0QBDjA89PO6
o6opzZbH9X9AVYDbJF9GM6PBBbcZI5CBJ9nkdwQsfXvGZboI9CjQp7DK3zNaSZ+T
6VVL3Xs8Sy1vgDjs6yx+w0lzzezCrMfGMjadMEJ3vS2dfqM/9tg76rtjn7qSQ5CQ
a33xr8gcUxs8pifS/9/du/AD1F2ytHTxYBG0HA45i+VI+v04fIjjqGtXPp1mgLsQ
tR/z1qUmD7zFON7zBZkIq9kIpUZcmLQGM/qW8cDH7O7pgtNlO9jDgrDWuTZvfTXm
QasUk0BsxAK7+Xn49fu/9JR6JqiP/dVuYnJYQMWtYX21pDV1oe/zNVYJInUhbxtz
9ze6Ky2bzjUugraTcgzaSiwXakLXInf4Je3rnCFyBQZc/Om3tV871IL/FbeS1gD7
6DUQ0kb+XLs/464/7MvR30uugWA8eM0r10O5oucqfNpebG1MSkPi7HYYqzv9euH9
XRiXjz5n+7EstAi6ndrdx/UPJH1wVwY7x1p4O1gYjU81hUSK11Z1wZSGldQKstXT
c7qmVeIHNJdbLAMmIhQwYcj0u24z+w0aUXlmaZB7t13aDcQ0/V9wdJ7Dyy+l0NHC
HTjjuZ7AU7zV79qRSJODFk3LvhK6kvj519TEGEDCH1LqSzh1m+5z7wSMM/ee0BIU
iQry2ahPIl6w4WLpxA+RAVLo4+A3MkRq8Tz1fqB9tnxK8NXdJ6HOjYvTnmw7YpK4
OHwWVm4owCkVyjtSkGHtyIba3BGkyG4cDFeDudGF2FuYoSfLh8V4K8+maowXYQX+
8IaCQLtXI0pMw79VZAEe37ly0nus5cMI96pjJdcXZjgPw8p9LCYyMqq0gmzhTznN
7tG/83tjQtKUpLEh4+J5Ck0B0N6CJzfnW4lpNAghI6M9mK3LiBVjntncG+jbwoxc
Eb+AC3q4CJ2irw5lJujpUK5JskgZR2SLpoYQxSQ+gllg2sceKlsGQy+KZopQp9uc
2r3AFKSRFT6p6hQxgR8Mn4GrPFhzYBf2kH4QnduFGGS52hEALDVenMKWJnv4kqzd
+kxb4NrhTrlky2Hb/4YH9SXTxHhXCCYtGPQ8s3xcqKy8oL6L6oFwp1tduuxGTMv4
OHf2VjnohRbpLpmKBF8OT8ijBrZUcYZVQC0Trw9Ei3z0bi5LtJvEDS1vMxwGIint
QrJkdQdV6yvM3avo/T3PCGlUKT0PY+uguRHF+25Nhv207fFFfwewBPHmu3n9jyeC
BFNwQ9i08hCfbHHFjVfcRRs1kHU0s30p/8YiVw7bMBWgeOwRgs8QUpKq/Xn9q3bJ
PDvcoj7J/VrMOce7dhB76hE46SQ8eXv1JqnNtVSLgSFiKLu8snMfekESKTulJiAt
vEnG4nY3EDK7ihXJbTgEcHVBCDQCgZQMBOzX4HR0Y8JtG3esMW/ub/iRClTFpUyC
eEySi0Pa3oA60Ucb5zxC2njK6cmKNMr7Xvk4wyyBmdJnu0JpqDpeueGVFjxXhC7+
9RbcZF+2CgGEPVgfaYJb6Q==
`pragma protect end_protected
