// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ZmSBtB8dlsL7Z1W8ULE/5yY38WEGiCdAxflRClOEN4gtVAun+0XqrXHxN/H+iNmhZEO7zoyDpjgw
gHrURfpjRUppA4v+8KJmoU4mAy23P9MZh59DY3bbY1MCxwhJnoH/xv4PWzGD8wpSm4tKNC46HpoZ
XuP5GgvilxCgzkaSPzoOLPxe3sR8o9PH3mZTvNdn3A61Ax6v8oiWKNnVaOqgPYxjooC4sY59b9vo
P/66T9QvtIE5jJID0CFnHstUsfBL5dEGOXFsohsnZ1PNBSYF9p3eV+2RFd0YRG//DwiTEwpc+/dx
dCo8xUp2yj2pEJ+XiHFy1+e1qDIXuQ27qKlRRg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10944)
EB/AsE6NyRC3dekJptW//g+eJGAaxD0TV5quf84wt0j3htis+kxWGdtQoqNxTO60+56xLol1O2uW
RuqbS9or/1UsRkBgYtgRzHhf6D1mHrmwBA1AXHUbNNwdikWlJIPzwd/u/PR46uUkalUpKvCcY5GQ
3aI+jLPtF0yG7ttKjDRjIZHg9pEX1Nxclo2F9tI9ePoeaGvBj+ANFgquV+omfsoeBfl0PMUznvMe
rGqbWRbg/mG4NIxrO57GOQAJorkVaE1/OHPfmm8RAvk98PbDjwV77YBLlByXwIcdVrLp2G2ZcWmK
wXuQ3GzHdM0EuxUwoN1S3EKB4SXXaCz5yyHX6Tw9LF8i04nPZ9MiiJQOCRKNTFH6POHwVhMyiIxI
NmxT3G0WEkezgJVa/A7qzRsfaI0rowgbCmE1bt/aELWcXWFo0bX4NiLdiPoFmLj4ET1OJe1H/HYr
odFkFp2eiaxz7sNND1kB90BgD0g9aFNe0IE5J3Cte2o9aeHwhcRhstYlfxM7oms6VwzGiorRCYB8
JRQlLMqsYTpVqROXPK/f4hgDkIg/gzl6PSk9JJtS1JKb2IkpN3ZonvWunwNqZ7SFap48Qgbf8+Uo
duNEGIoOSDqxzL14UOIXcJ+Cwd0vp+KvNm2OdAokb0ZvKExtr9mVZZ+D4XJU6qXt+toKdr5KOjEd
nDFqEyBc+Jru5xI68rfQXYa9XeTpwPyhybuqQLzdOi86b9HZmTj6/6/bfMSih/z8FRnyAmBM9s/E
ON5bLqbMkXtweyl4B3dAnAPSzwKofikoBlkOWCMAPIWkYLPAACn+xvGbJInVJNl7IIoUg0BzKbhZ
Mz+YbHmm5g0jXvPQ4bNC8BLpOtJufqADWiQujIcZiQXcTa9wmsgm77hi1Fp5pSCx+0WAXDPyjcal
beWJrcctACHcuIR9rDRi7sdTrUNzjuzJA6fcDrnixeDgIp8ZiPNOWIunN2bnFt9jYtTNQbqmrnCi
rGooQEeK4o+UiEyXLBfYIrn59Xz0OSoVT0cFj/ZIVqFiJjHNJdNelQ22iswmXMhxyisooQay3ZIL
UorXTEqqS4P4lU8hFMiGg1BkR7mUrS83evlm+1/WHfJ8Y+5vedFWBxH9GF1wVfH6LIsnid5/Q4C7
ody6I+vKi1wfMwtEKX1ij5lgM2DTxAh89fpc3SDswPYocdqW5fSb3KYWKgHzcxLteWEcjNyYG9zN
moP/RGUd0RlSwJ8YVnRN3Lg+AqVfPJ2NS2rHaNcGTPgXu7nTGRLS9MTtNY1ORJVDInMGKMDmkmEs
q5NtViBKrY0D2c1N3qg6w/Gd8NufzAPquIPpo1zgyDbN5pUeZhL780zqQruAS5AWWgcSvC/bvnhs
6THqXBcNMJNfu1JaOPerkL7JWjauDtqmNfc9aORYlFg4YSaoZ3wZGSv6c3h7dTdlkjy7ZuNxjs7I
/MEHZI5K0pzed7a053SPkp7o+TD/mAUwQIShvkjmW8/8QNIJGSjKV8VDA4rElEsosA8iDz8rX2S1
8Iwe0Y3JG4GWJjko3fQLe8dMMxtAY8VfxbiGF5LpHu9bfYvmRmzuXlCmZCGf0UEehuni/WY5fBsj
xA7UFB1R36N9lvQWPIeSuCf9FhP56bJ8B3WwYXY59u/5AiWtu6A7BWr/M/Awdpn0xZGBEknjA4n+
n8ZOFr1yE+X/yGAdZynMA7WoxYckXVZCzmzWMPdPAC0ypgbAw78OD3YMOzA9mrMKPXZ6GtFd9Jkc
wNhS2TqOIUNBYFiEElF3K+ftrUpm8Uf0x9OmKpmc+IujvSC63uxUKklnyHB2HFWKiqhX3TuRQUjR
pHBuTSG0WpClzKankE/316bArzzLCcUIB4H9XwWnAJbbZjmDjTkZg8FUlLZ0Jph1qT+39pcrSPOZ
P9xRt09cIssTPrxrq6GKmOmF4AFKGZIAmaDspvQIbiLAZeAftSX/WMasVo8gBFc4DErV1zRahmM2
ll+ywgBF2bPNdOzOzKhLpvbd6DYK5ruXjSsumP93nxB/ARESuVqYcyPtlWR7nhuMQa67quiEgJda
CifHJBk2CRLdlmq0Bx0GrdR+juSmEpJtgbEVyKQrw+6rI4uJKEp/6mC0jaBM+779Y1njT4xEIqMk
WjyoLt1TtFObBOgB1yTV0WfHPi5CCQdngRiB27EYjPPPtkRUIjsqP3/f8na0DP+rbo3BGtKDTG8Q
LU0kYlX9UEIjsXgtQZ2KsgHq3Wix7q3I4AVZWRs1DDpq+FIVqqlzvYBBRc5IU3hF2/4MQYMcY2B4
QVwD1Ie9eqNO72yAG8xR+WbWJQbEdUIMqU1JlUW9Ia4i8ORHbx7wMklBFGPBWk9IH3+PUzABOvuk
UkleADNB3DcdrZHvqqtM21L9fuuQZemW15A3VAOI1p0MBojnZ99SpGLfaEsItRhyKyWQxkHy89KR
mg9uxbF+iyZgY5i4BQKdEklKTMWcmEdf8dimAUn4ovqnzan7rA5vRoJFixOkra6NL/Nzgpeva7t+
BExL5S0Wm5IEDRikYOyit58aC/dc4FdaI8qLHBch6XVNYHAlvLTwzhO1x/ANLAgE3pSD3rlGSo3b
tEdRdiL4kuupYrZSkdsm9W/viS6xk2VKkJQ9nX/EiDuMMGNHg5NnptoKa/zoq1TxwlNPK88U5AU8
h3Nf1DW97Qwz+zt4aimCX1+aRgova/CBlqHrqJ7q6wDzlItwiejjqkYt7p1+q0UWLRhm1jZEWwdn
eyrHZgdtReoO4U1No+ehCesQ4DOp/fRT0+kK57XcdQxsEDEndFOWZ6/W1f/O0D2GpQpzeKl/hAeY
eF7eotgPASc2q2bvS2C9ZHB6LAZdLtaaXsxNGPBlbTG7wWEWMzMHOx0scwvp3MSdGVdaxh2YzQNs
odHhLfQ3WBKzRn7y3/P8/Fs7eCG+Fcgfpk7ag+6rYVbTC9l1qqZP6eW0P4icfbM+LoRsxdVYRPoN
hXZ0q2I2tU02sZ92YF9zCOxU9Tqg2IMBMIeSGwKBihS2L7x6l3mi5f5LLhso4vLmXBanCursAepO
Gaaa53r7p9VwSXa36x/BWydiD6lHlMYtSQj828kr46jRGjWg7B3efAZ5Td2W/8nbO7kXc7yIAoAt
0TrJutGT+s52XA++tP0SVbFVjIjOMq7YLqQmRfhPzlPQeogtw/zdh3vPZeGoy7SKyDZJKoG9vtPg
4FzBGwBTAvkPWxLWyRbDXy5xoW9llLpzCHuwRld+zO50w2Xo57p17R8tBX44m/tXC/JdGuRnpxwA
48wFQpD8bcXGKk7M8bvgICxCwGLjmewCr+1SooF6W0FXetHMZ387Oa0Dx6t//rva1nNNDhidgP9k
fWUIxG6JhoIpJFEFwlrN2BGocWW5r3/5xYG5QpHY9/XWmYjxq4XugfRSnrBfS3i9aTZv4ernSfWD
pIcLEPI1fH17yLp8KYI3NuzMJUgpNPCN/h9yTM64uHe/mZwYdfTtOIJLbRrLXK2I1m7w9cFhr4o4
QdOONr120l8svdqmSmRZbyEoeDqkDbZWiSVyzg/WxPvA9v8q8iVFl9yoV3pOhscUS/FODRKOKJ1m
kigQrvOdq0dnXze7BlEe3EQo/ikWM/nvqdwsPlgqzNGpDc5pNI94OQYMmGm03MQ0EvutnhkAVZD9
wTfN0s+SCqGcILawKxkajN0pT95Z1gutUR0NNZDE0v9+hzGoZs0p0Rs3gb4XfOKGl7vccEtZV0Ij
gpy+jKh0Nb9WOfb2Ta2Aziavoj343uyCK79gM+KRkvh5ltDc79UOYYHF+03s+t9q8jkj0k3JMfU3
91AiEiAy8HgcXAW25ezGYvnBnRmCevkttnSoyQHEfhWN1ctnA7WOmE8BOGgEroeupSNETt0ikOsB
tmMTncYJy7z7t86l4nfFDtCIK8CO45vXASyXNsMF78y2q+dsSSz3tmYfF9d2I5knQao1zIbKiLYC
jkxIiFBcGrL4m3PSquGV+UmFEse8hHkhUTTs/oIzpMAu1NJFQRTg6/YN9GdxlIIHyxcAVxdkIXbI
FyKG746kXdiBkgl0MlcAWY/1I6x3f7s4QcM/ccfkyc/SLFPclJGU8m0Wm+eGJFYRQ0w2Wz51YbHC
Ecj/NqPFY301R0ss14J5/qHmzG1pBPU6M77/9nTODfY6fO6e6hIryeB/VbLvsAaXg6RAJ2WY44Od
jHnf0WURQ0yAGac5xufgOqqlHrTmr5lXhpxhlpHk4ranG6GLYHeHnge+nxo1IWGm5DaRg6wz0SVo
Cb7bTd/7JN3Lm4VRRmJgGzhaPFWkux3oBAXaygMe2iWY7ZjORAc7drChFa26Wzp/EWUIEmF0FJ6X
SGh0UMSz7KnA+a8yCCDCHrM+V++MM+1dV/LMkUl7NPPdDNiaPwS9to4/v+nqgcwWWxx24RtH2IaO
UE62PvCiJ7ObiBsw6L3IZ6/hOX0+jEB0X3pEY8VKkqMvbbkmSc/sKN8QMdfNGXOLqv/Qt2Qx/bEj
YdHB1vVtJDi3HU9Kn0+GYJiiCT/9DkCcjnDs9jAJVKDESkk2dnWhOuxKy44XqNxr2B7K6+P2xWaD
C25Z12mxK/4TaUmuS5fqC30dymXY4QK1Nuni7ZVZRclsDz1c7JHWvvzVvhhddlU2l2s0XDKJRBle
+giJFQ6PstgbCgi9kSoxy8Znrc3VECeO4S2NoPwmSN59C5Al0x8+iEIT6Xw0oBSsb4f0fN7G39AD
/BI8tcdUyegtrDB41WpqiF/SseiT+DqEItgekKNe7llRfHEy4v9OZ0I8eyN1BKjScAe79bEYX0bN
bpOnTvg4baCz+wc64Qd5M0D+2t6PO6YtZDEf9y4xBS1t3rFKcocs5scPJk4wmWnkR9sRMRSYn6A1
sELBymR0CuxTN5ZPZufCuCwmFwh6FmdxrL+TdRtFHG/2aJYSiR97oZy5lCYV9RPdhm/siO32XIr+
Ns4+k1XT70kBlym9Hp7OrnGicmOeRKl7voLvOGXwY8ZvOq7qUJfQxdOQjrNj0UijtQSesEBfqfQ3
1CTshayEBRXWlxPvEiF4jJq/D8DPmuhmkoBCzw95xPFwnxBqmXqyVHoY9sHfRDp8wIFCYqBTt9L3
A7WGl0ZSpk2LyLVfNzK9xIDovpSbBTRYC3wB54e9fR1mgNZqA6Vp0sJGsdf0o8OAttXlel6ropG4
KJXvUXaCnJMShHrJ7d8e9fI9uIelF+XMztsjHY1G0tu0Lk4YAJrxk4nIjNsWCGXgZktM0Bp+p8z6
Sd8ONSoZ/FNLKH050DHGNHNVetKSqAvjd1MClTsm9BYoF6bSDNNryChXonWac09trsCxITL69BQc
g0YSDT7W+DffKmfW8PyRlowhtIWj+SZK8GsB9AgulykzFbAXmdqFx0ZHujjjxIE0fipk/peUFIdO
nkuihM2Q7P18wuFKzMxsysTX7glgJr+EolAg6vyvTBNg8d0gmySEV9pFYckJWA3Gz0OlyUlw0fex
izjewtxlIkavoI44ftLwQT5Vkr9j+DBUIA48jU4Eaf7s9iQFU+0UwXrLfhEZF/UF++ISGuRypNYV
lj53/HqF7peOFm5nlRIJZ4/xb09ebpUtWTr8lvCmztifeD32Xy+YFH7rx23pHuYlzFnukf/JJaft
ymYMjxH5N2YOfSqubDF0Ld12C9JivHZiWXYSiGkhlpxA1gkArIvml7NF5nGM3NyxZ7dZYn/gqcAN
4x3bh6qkUwsEoWo5cEQ9uQEP+Q6p0AKibQj+DEnz9yAX21TE1nDr1wm7PLZGuqQiHF385eZcHshH
lPdEYEbwtRYxkTgf3yy1IPgGwLSNGOdFpykts4cFw2EDyS0QSZCuWHpdfiiuBgt52lfVRLEcNgJk
i2i0z6FL1/ksSTlzxzaf0t6DGMQqSKWaGqN41E+DQw2RYF8VfPIUTOJG6VBMMdt4cw0lmmOgfuAJ
QqFhcoZvklaXOl+i1DU/YawNTZNaZe2dcrxuWwihbyg8hQd3Bsc1gdVRDaYU3HEea0DRq0bK7HQ9
edqBTvEr+MbmzGYPLqXe3ZtOEl4NvYNydHfSgmQQo5YedH+MfsddKlk6EffO4TTwtklcacMe6pj+
joc2OoZbumZK12ntNzvBAwogCQNAje9JevwL9EtSrZcsVp3os4nl8+2hZBCd4D/bzLTelOTIqXmd
292PbEOt2lPzBLAeB7ph0gaza+6r+jfn1JXZsLreBvG+eSIkx1qLdeD8uA/JPN/JuGBOrdwz5r3q
JwucGmhZkewVctIo0i9RlP8PU1YixAzHach6HX/vjWHudZCCPXjBQZ/cq9b05CVYZ6vUvZ05I+8o
RIr5+vmakKxRLx9hV70G2C16RQLBVkKPoQAYxNG4EbudU8mPHexCAYKwtI75yoSzx7m/8LNynLph
CdHVDWkTi9GunXN+gqZQ445I+iPUGCsuWux4bBvcbDiRS/qQIb92PsSqdHd1M8Th+hbbzfT6HR+A
PntsHnnSdkFPEf9isS6Ak8ooF36e54WvvR27xLJ0ql1Xam2NlAB1V39zyikdN7+leDuvljw8McO7
/TpfP6OzrjW29V8cgk3km9LL254JoV/YKj0VQmXLuEasXoQG7KfGWr16K9dBvjXGOtECSC/xDTsL
Q8FR+l341Qn3OXyiAqdVz4hSYrKjlH0+IA+q8dvCi10+B5MrrBukmnI4/Py968sLRB3K/Y2+m9F5
3UWxOvI63+qNJbWKaQXzFAobrmKpt9PxzLNuZUcNRZ5ICVI3ZK+TDK8p2zZmP3R7lOe693x2tD87
57iWnAPUBcO44PtLz3UEAyputgOGL17NgA3UQ/0X+fxqXAm4hM46jELHq/T9Ap473M+scZeR759z
9u2cI6++apG8CzhAl+WmnmAXyKq0e8sVo4p1G/P5FTUVqUHeYQEpGGvizihZnCCHTXdN6He51ZV+
pZxbj0E49I3pWW6PvSOQfbQupLQMH+9ttrb89o5Mnkzt9Vy8GqT4c0o5k2xAqsiFI462XHvrWVi2
Hpi/39VAQs6fU71pyNEktXSHG+PrTcXvhsKDTzyzdqN9P64nvjdz6i1KrIaJV4fkt4xRWnJO+dHN
kEBS9XtRg8NoF1igBMkPSDXW/UbDCy7J2Fr5IAoiv55Eil6/8b6rszKU799bYlUZZWTvLdxhnAu+
0qCIjw517RuCul00KJ/ZKXg3Q7LWzhuUJX3Kj7WNknUqT1lahgJN8v1OJe7Nd0xkjp5eiBYQd3ux
hZFNbfmwib9kat2gigHt7s/USaFW5HLlSPjNj3nPHzGQvtM37LRY/XvN5KjSeKLioxjG00l+U0oA
Cf05nauVKmuhF2QoflQ8gwekEH3bIif/74Epa9gJZiCJcInHV1MnEDMr3Ith/wcmrmV3/829Aa0n
BfCqzDwXWSbUsGZQfUif7sch0bxKGNSGsrcfiFGdmiRmg8xSW5AJNFFqYIey/KaaDPHYBSV0xKJt
TnrC1fl8GOL7vDNe3aFYsbzsHDPo3BShWcsl49k04uh4W0C+Jaiq6G/f94/B/+GHNAFZD52nBLYt
LqZ0F7y+om0RorJQiUsz4eYMmUEg9s/bNHNoW0AfoDyzUPCICmNiJzUXli3vdQPht4Ye8r6RZ0pk
4JMoIT8AcYItJimrLlic9pvW7oUkMGIwdrckZnaiGUEDv9FZ+YLvQvkDDEBXmBkjCUCD8AIc3YvN
mwG7MpxF+ku25gai144kGUrxdR0oiax/DdcwfaXgcvcCMaaWNigkf3OFcS0T9yIBPbORxv2Da2R2
U8xMe/gObzPLVNCOsEl+6MAgm11PuUkZtUOQsmKqPxntAr9l7tcNr0LgsOSptCkt+ouPNZIx/ri8
eGVmZTnil39ntSGKPOJLEBqTJlTavdvdqZ6MHFFffa7db3clyh+eWH5Mj5LEG7kDlzsrqsn7Utr7
U9be2mB5/hOsBDLTltTo+bOfMA8kZd+Hc2JCPNRJ3LtK3D3FI+EUbQGH/t4JSPcODcAF+MBpqr0/
qa24JV5hwSWbYQdmJLkM+qm9UzTLWp4nEpRjUPxhS53vVKM/Xz+yu+0ZIhDw7qOzFXmozoFigpTv
xaganrkW+i7OsJ1ynMaH1hmINxt5at65Ccws4KhAjLLiCkMMm0eHTkr4qfJbdin9lR4DpjzwBH7h
whN3wzYp+giQITGAYG4chF1aS6AVLFAAG+8RWkwu6rbf1MTUO+RhrqbLs39YI2JGgpU9yAZglsuc
M2hLTwFa7/DRv6X+3H1UjzmNkt7HNOVQMSJV8I1VBvaEpYaUsIQ1iicQ5AHfyIdN99weJ027q95c
rvv5nekLqB/olCUsi36KO1TjjqWU04ooc3tqS0CZcGwpRFWb7Ut2wdcUcUGhMrMtYDeFZSoPROBP
6BXEmSuPa9NjVPrfaRhTLrp4WfeXlDMd/Yis85eRWXAuqXuua+GL8uyaSOlhHNGCbhX1wix0MVE7
VJPj9jIyHkuvFjuf8UcDYnNgO4lUyfLXJCtjo3e1CyUyjkOYQTPlWyI/F0YVAI1I+C46+lWu1NMD
Ufavo7/8kLFyNrP+uf052zwrnuPEBcv5+CsLQ/JlDeqRRfKwwOxYhIaKvtRXNyN7JC9iswCNNrnw
vkV2QJdsmnWSR8n8jrx/44npzBb9VCC7BRbu/HtzHYd1TOPDQVDiCDRyfx6B+RcgyK0cUbX/WUtR
pwZD2b94vyHmPhwI1BDmgGqm1xJFfFGbGlJViqaT2BDITkKYU2WFS1FNZCVtZYORNpuUgB7PNNAT
oNldOgA9Plh9+92MdRxZr1xY6XRh6EMkeTlSre3jdyreeOsVSdBDSjD6QV4eB6ycHjcK6MuAhtCi
fcSD/P8BYx+lO0qTg4Ggk4CD4EOadryMPLw0RZayCl+UWKcFX+YKVPYWKaMovNC9xIapEANebHPk
DySxEA2n5NUubbaFOcu0go80Gc/iyWHF830m8ZTydfSjxIsdy2lNdggPdLP7523s+wsH2VMtt2j+
FXky4l7q1rKwQV5L7GRPiEsh5EoMN1LsxGBM5IDHN8dylzyV0kHHkCzeSLvsqrX7vrppkUn6DuRK
PS893gbownmdAA1+OAye6JOQecqCORO1Dvgnzx83YdJuxnysGIUmNRXXnBPEJV+qLTpB1r4Pezqw
cr1yuAATrJYcDlFuXtTnBLhzpISmscfLVl93a54daDuZye7FZB3HcOy3OztSRAcwKDlS2X+Cqnqo
sX8p5+gMlUZgs3Ii50MxO17aUZsqb/xc0ezAHc5mtIqDvsMoO6RaNeQYI87jlg7E6VuXylAz1EpC
uHIdTIgNxQLRqNnKuqWPYWOBfG3HzTXwoSLdeL6A6DBKXsrbCMd4kOtskpXsRqqUFzXFPzlZ9PgP
qNtdZk1mX1bSSdvowq4FFLbCkFZGW1KPQoUt+LnSAcN+nZ1Gjz4uT+28Puof6m3JqE+Rowcc90U7
Yx+bOM/IL0TaSDW2DdmXrRuzmb7IuAMPG4hZRMDNY4qAof6EtNbNbwi06e56hnfnRuO/rzGlFE5n
uJffUwuGmSqUEfvFwbYoNWogNdwjvG6KRU5GldRP3FCTz1/xSlVPthMGinIFQkRpYjFOI1ZgpS38
6cOWwWTGfjmxuW5A81mp6O0m/jiKxipS4Pr+zFmngzEK+IBraBucMC70fEUu+8hM21NggnW0W7pX
3iQweMcZN8lUs6/OyIkZFWX4yt/Ui1Nz7e+TOgCPV5dMIkKL9mos8AQwvXLAwq+wMOH39t8rpTLr
nDoKFUo4FujB8DfPAHqnGcyjnSxxSTSnDb3Kuko8MElQ+NM7ynko8/p5Q75mlrhB84N/r/MwFVcF
JmMU9R8UDuWvo644MzibnF+DQFS5+wVxSDbxsthBDbc1t0/r/AZ/EsQJTVIhSZ8nHVAEerlwsYb1
uf4tWOzrx+9z6GTE8NuQo0UHf5Psxm/wPqxu3VAeNMVJcyFB5SEbpkzwsRivE5VnbZL7QPvNje+B
yF0/Gz5Q+TmEDo02uwdjHGRHs4g6X9fOeFicR/P0XLaOSJUYLge3FllCDiZQPgmq1g+xCFIR1F5E
PHPKfMpdBHjRnBUhDYq1/YS832pA4EouYctVmQEz54F416YG0ovku0Ro26SaRjQ8MrIevem9prjd
5HYFZcmEaKMZG4GtFNju5la5yCpTl6i2KAtJ+lVxSqQVNvGwP+efKhWD44eDnioaAq1rrupVVVJN
qFBPXeolwNKoOB2TeoOJDVX47nnD3sONXzlVx9cOuklEhb4l/m0iHGngxWXmOIla+JoP+HSZmv0y
7insHnzXhuiVDTF2Ko/UTK8v6weRHLgj0Im8vppphR81czc760e44BAN0r3FhguXWe0AtsiKnwA4
mdfZbOT8Bbx96sxoTw/fgGRmBUZeRXEPrKobRHU/HtcrujZPcFM1swSnxm2Crc2GjpjMD01oao9g
Z541dlMdwENxR+SppXqAFPzcTIdz8XDjYxL5ovXi5OFjGRCrFUuoCrMJm+gYvUSuqcJ9fqv2CpVS
3eZP/YhAZmHhqE7Q4YtN2D94qMrmJ1DBAfyV2HLNvBKoAxYsa05GveljF81bZjhXBfgJMWJdOVOJ
EF6LNQV13DAp2HTiFBXGogaGQ36YziqMfLReI7WcaD9RMpT/c0OqPsE0HSVuAgG0Pl50lAqxPR8c
xJnKDIxPhbrfJ2eDoo0wH33sp12lMsoaVJobuKg0ocdt3mQgiIdQA7Q8qIXB8mvU3TuneNAmBSna
NuXrl5SC1E35cFCIdAtcCT2xH6DH9WJ5x+miBFKiPnwuppxPTC22XJ8ZUuqqBITeHFYurqTKAfYP
VmSY8jQMCbUWYMKjY8n2dKN1hk30ivDaae0xwH4yT6Ywoa1ZAj1WuEGou66GH9ZiWytvwGDM+2E0
ZoJJLQTTmG0VS7e0sbA0WvXd4aD/o6Hf1P400DzlWbdijC3Keu3BJLLMBhPdOLS6gJqWX0PBB3Ie
j9K+EIXDBqRx6p0/jkcyKJ7XfHnWP+BfzFnjg/z92N7JM+8R74JJ576uYdRmrx8b/fPwprkYstco
k1EUHDoSe0tm8V6WS59Fj2uVZ7di/CJ5j2nnRFbTOXzQHdzDQlXMAwP30FZyhL4Pn5frA9tnH2+k
M3KJxqNqei1LmFvF19sokmHBaxrcol513pTfXwVszUWCNcKtKrclixi/ccQo75WYw9VIjDHVeC92
LyOtWR0KdtNAu/36epiNGPAi0eodPkU71e5Hl6YH5gaP8H5XmUWEXffRcJ3A8PWDoTclTma+yxkN
VRplZ1sM2zYhiU8Jn9hK3DpgGOio+2Qg4hDVHe4wO2rxi8Xjr+tHnXPTaLhAEbTDy52lTxNasey5
igb2+mHL6HpcyarwcmBoRw4Sftqbi+9x2JsujvLneGv1dz2e/8YcPBJNJjDjj/hp78bBCSJ9i7iW
K+sALluPVK79XbqwSh6FcZyXO0u9kgWF5rLu+PAKCWwnu+l8d6KTwda3DiKmb8fqdXbeeUQ+cFW5
9ybYQlfKXBGaXL7/fqWLMCWNBTy0rBDqd0n7cCIYKWNbgyR5A11l3or2VoNZcWC9AjtmCAStYhwU
fksk0nM+7rt1lJn/wWpEFxyrU5E/rO02N272MbTrk+fVx1B4RBHZ+JQiqH8Xa53sLoaFcQGonqml
KCmbew2EvarlmQrYm9g9rlO1cjhC97sG6J/t0kgZhJFMDLFDQvtA0wXWr7d2Y4wN+HHeceildjLz
cPzNsWeVak/G+u9y2zWQN3gXIUEJjPEPoFArLPXKJv6offeRYj672068th7oRmBUo1K/1Yo45Vjw
GdNrRSfq1WiN5sPHohahAjzAWBnsLcurqL4Ysgej9FBJRE4EeMiRFhf0rTuVY1ab0H/7OzG2c5X8
9h7xlsjMVCrT+BkyMbadLNH+YfDzOIg8/RgtW6gX6eMwWPKO7383MssUGXsv42tgeulHe+OB4G0X
laJSe7sUQctnFpnR2ukjETeQk0rSREj4H5jkQjuNL98QVDNyMTIxOjU458zzIRfQz7a1ofcP1hq+
BwxsYUW1dIvgRFobYzBoUG5sWzPodm5CRbl+Fi5IPEs+Y6dxB3D1PhR/+ZOvRRLXRVhg4H7l62lZ
X5lR5f1k9bIa6aL+BkG20XqMHOJM+GuJeO8HYzIeXKypDacqTQAgpIF80n4NpeThBvz3JybYhc5Z
XvQ8Egzk18fNLhmNE3qgT3+53zCiu9acjFcrkMchpUXgEdHtPnhNTBp7AB+G4jecJUEePhCNiouA
tZ/GEWoVKL3rosP7y1EZeE54Hp8cDPxh3qQ3ngSUj35vrkc5OhtKy+D7WruyiJnD0wCY1ObTlUTG
X8aLaPIIAcS7G+SxzYTzbpbCu/MNiny0ri64R4e66v6Gx3SzcJbRtRsjE6kpe4jLXoHn5RjLcghs
OdtzVVILzZDvARwlef4PsxT31eRpO/WF5MEH+rG7d4a6sGW74hjwOKW+r/n5jZDE4O6kcvrYhldU
dnTp4WwVJM5WCizHNXmSbXeG5ABOtgVZ2N2Dshlf3xcwCDRLaMDfJRRF0YWxS0HY3BMTcNfKND/q
0YU3bneAawkMGJUvtg6uJi564NKmLFUvhkXwQhKijROUXF4WI9L8nLOxZDyiFQHEOyLemjszjphl
eZIqQsJ+NAfvfpYO3lGSBxOkUn+Jj3jRrcC3o37bBXtiBZsGLQF43Xi6jXHa7MbzpFb1Q85lMC/h
tjB+Xf4/3x3tuzfqPTqP3JSZ14QFqw5uQSZCtBVZfYUuqr17Oq9tdpiCeMnHG4/gBj4QFesuA0ik
0hNNVIMqTfEgUlPsQHaTN7KWa8BOCnODJ1vCnAnv+CSyjVbmTbR+7lwBJcvjPlt4J6vCbcVZVoQl
6o5kGP6AibEQH6OLl2oNoCElkLDe38QVW6Z+or1+Pt38V2jn6cq13OcOMrUi4dHY1wKyANf96Fz9
ItiE3OD874RqguYtEbKx8Q7ySY22UYSM3f8lV0GiYknxg4cQy0MysmQxuS+1BTvLnjnoNgnU3GI8
oRbsppO0bhy6p5s3L01/pxPZgUwCrKK0mEbsHBHUKEcpApdBIFlWmpmIH0HviP3p+zdwCgWWA7M1
2M5Gy8FYDcLCb0iNcE0aXBh7e+zXchRhmkWcdzyOBvwdsuGKB/7kjjPe/D+GTWa8kL76DPh5qymS
lo/eueDdgtQc8AGXZrkplKDcU7kgWDhJ3AiwG8ulhYjvvt6Od/3Mz+K/W15IaFqCPB7lwfqEQA5+
H42BTjJxkazqm/8bcZ8IyAZL2uegPJ33ITUo68s8Wucpz//hrzEmzbCYLRRAvNuFPal9ciZtjBUM
afXbYeszwBPpQ1a9uQZhjJi52MPsc5zN93Qjwb4KHRLneXzYXkandT4A2KHr7YduI39rL5R5g6Is
iV8NHvJjzjAsScHHiIXPY8b+FfKZNa4mLytx0gSvJLISY+uZJtvo/+seHPvvRpnyRCXv55OK6TaA
ln8mXkAWRSNmCGsh+AKHccQGH0vhyW+jRmLrGN4t+7Yx4R55qwh/aU3Alz5mrcp0nxzPNtwmCDqQ
avpaNp+tgc1Ylo8qlukrg14R2CAWnPcvWcdKleflyllycSafYQMLeGG6YBEWE1ypOXqTMoG7MKMW
y3xReQ2LBmzqIR7sO/DtNKgqdo7H1Zvf09BQK18hdZrmGpCC8LmKsoJTAHRFaOdQ9u9JQXl8ic8b
dwAWcdbYNQ/bETLiGTxHiG/Ib5q9t4y4o3en7SlX45hUh1HQogMjXMNSvxJKAIHaKR1o8BLQZyen
en/jZKWTyvR6Kf0dyYyaqxCIEHFr6hW2DCzd5/yz+2JD/3pda1l7Q6+niH3BiD9U1j6yTC4aRIpW
rm4753Gpr3IXVDedAbMbyRcKp/eIFrL6y6WZ6H/3BAJhAqHSXm1gkljFhCexb23PEc3RXlOXiCpK
gEDhNGcoilTYmRjWh5Ser7Hh5dWJ0VP1xCXkWnINmCJic0vFtG5JrIt/IClSkJ8aFU34pFpVinIt
kVX8dVeuAb+SGax5sgNXH5Fz7L6qRR49fZu8ULX4EW4P6tVhf0pqI7VQi7xf0z3igwHVXHhDwvH8
TUsohxfFNa7sSLH9EdMzBkQo+hJD5YCRoDl4xjypqEwiT7pHBR3nVnkrxPg9scOIY+I29igEax0b
0ppqC/8b74+FpbLtsil6+bYlKqPzGs+Ae/TkI/FuAkfJXAjbbEvN7YQ92mTB0r6sZHON3WT0jEPW
zJyHgB80MBOI4S0OfGhIRqovswCr0RHsVJ/Juc0pG8QeTke1zyImYMRobUpLcD805zj5pq06/9Y2
Qv4VbRi4WErPEqkuTyF3QeAYHJjbVzezfaMRqyvINj6eP0ARJqnup6o0Yw5D62tkJGMNkoIdx3hZ
Xo+6VsRruiQvx71uJauKngWTE/MGbwBOf5iZh0b+Jryq3QFH/7Mqsh1LS2INraxuxfdr1HjEbtLW
vHwOmel7aLvP+UvF6XHuzG3FEsghrSrCizFGzxOVky3H2FKZJsyN/Ngdb17u/1+q3ue05Dxt7ceO
evd2hBF89ndTV1wvJqhQsEgeN24eAG+H4SMRelPmpdKGOyfdznNkr2RnGZ675qjviiiB2UuXKlXZ
`pragma protect end_protected
