`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sZ6l+zgQ4TApqqMCVB73nXgFO21ZQDRGi+0fJRkZqsTwqX7hDof/yW400a7Onew/
2xGs7YnJwm5gt9ucel5evW2A4cV+j2JZE1MxcPmWEivAwUtbTDoUtMgEvKrObEP0
58sKq0qlyCAeXbpkhyo4SlI1teNEz+WryAObOuF0ivc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5200)
jXhA7l6gq2/mZXINL1EAAcHvIPTePQFqyOokY0DUdmsqy8BNqIdNHlDQxmQ7ZkSS
C8MigKLw5WsJ7T8hhS+j3UlcgQ+hK/UtPLnZorhG8Dxw3XawopzA1Uyw9k3Rhitr
aOtN7e5gIp28b8aPZlMp1fmgJjnkClEpD2tJ3UeqpflVeffcnrdYayxxRhx8c7NX
+THa860XXTPcIwbFK4ZT3GEOPSacInXq1B/uht0luc4/qn48FltssMlSC19ME3m0
iw3GWyravFyVPUZrlOvA4C5q/ZHutNe5wQR64PSKzLzcq6D0+U02qYfYNSSTpCH5
Po2poEyVe8FzfChjMXTpw0QR2Vy1Nq5fcbjNVneMXMFfoMa5qdngCiQxry5RW2d5
0n2BBSQQ8DUJ9ErIPxW78C6uWScpYyJFf+1Rk9xidPU6aABYzHwCtJV4hGo/GTGH
3B6Tn5mI2foYapNQqoOV+kSJYWY//qQ/tyuM/wr/XpdWMwlw0GMJq1bpoXxcu4AN
JT0rmBgJEVcaXGB3MGaPHbDLvb3+GQ5xwsbtFv2FyS0cIT0R5lj0JuZd2vsJdebW
uGRsFozehQsU13sddTklS/OBAu7wFiK/rM2KwL3tVWfXCxR27PUWPbnjqSCTBRZy
5OG9JMZBSpkbo2ptOv4eUl219Wvc48IjHvxJwS4zJTqg1oH4Ajdpl+Fld60zPqmJ
7R+a1Vk5NoFsksxTMCGUulG2fd6ha5keGIyOAfsKif5wRvMDw3ccpNWlEtqF3rSK
AdUIY2Oqb54dcH0uF77j1A6UjxTxBgud4hzc6H71APtu4lTcqZ2D1XB5tsa0TooK
RfaNyedO5KvDNlzm8H4NQoXwFmzEPuyRma+N/hDhk5HIhLAsyB7LZOkXx80B8tWs
XHWN7zBaS1g99fu7X/BlTnWM5aMig+BFlYOlU3R4Tmrd7nW79BbA8JJtFVECHI0R
xI9IGEKpAjcXqRQtTykLSHGLSiEDSl0Vv52c/7aLmYjvpTqNTN7tgY60+aizET9S
YRqsx4Gh1cBTRFagspfV5A8Bfop2FLM5XJ5wllA0yGFl3AIt0VT3wfI9rIakw1OV
5hYe5nHBbFq0OhAJo2wgASSQwGgzrjVsZ3/vT+76QHhEU7QlqdJw4Leo6V/oSnRS
FwstuYDkaRbc/SQqCw2Xaq36IrqERHzXA85m9EPyT2/UMY1S3fxYjdz3YnKA9A9Q
FpWE1BXX3GR7FWPA3VQ4pGvpxqN4WZRuP6AOrwk7rffHAGMiJ9qVp43bP7Mrzv8w
0++oPT+YrPF2KLbGWPfulfiu9cmXla1+5Byi0lOHyW8dOjIbjxOkfVc1GVkz5yO+
jFvLeTix7wDd7iEDUyZQhfiRvKHf0HMyqPamjHB029Q4b5+W/oekfK8Hx+wtDIF5
85inokGSOXaJxdnw/fDrv2XUHUXOpMfvVRmUIWiCkB2gi3y2RuXu3K2UxAKQ22V4
ABXJBXYFf0kgjtotnwnMXLJWE5cu4JL6mcWVy+mrcKVh4y1bY7rEIZ3YUgjBYsdZ
d+GUEVuC85VyKbE46bheFpcIhpMrASImlywcd18oXA5B+iJsszufDekcOMNluo81
GeEv+kWpJBP1+/The0iwe1ZL/IwQAnmKiSoYy7Wcat9k5GZi2lxlbfNfkonrQoZC
SP+VaZ6u1C2nqdEXDDR1NHfjpFjpdc75oKYhhuvkXkPdgxhn2ZUYujklBdxBAFqk
k7vL0ZWCIZiDpTHLzHiZD824yu3eGvcis6Zmzc+0TawunKx9/dxLo3+OvBaMbFnW
9dcpfnG0THD991LAKDhnCdxInU4/4R/KiDJspU5AEefDVOEXS4/0v9ZHUerebb9e
svYIK71Ir7uIvpiK2SteRn3a1VqdX8i5aA8q0zkS3QcLHgW0PiwUyhgWJW5DB9v2
/G4Sy843lC4ywwn/Ls4g7jnqVZ0Nw/WSasuzcQK5KHY14p+JYxgEmyrOFMXdBkRU
S0/dNutbGdOlrbUmZe93pP1mk8QSo7FV9+9tkUIa+juzvAsH7/DWHKEX8IqbtmpP
ht74SNbT9sZpaxIGWmE42uQwq4BDc13syqAvggmTqLXeOdHwfFoIHW5hmUR73xWv
5sr+Uvx/SesInDDzsbrHCA3v6tQJeLJOnHMmPMWGgCAZERZkJuD+lSXGrDyEg217
ZmLG47wRwRQ5iPmf93NvQnAiDF5D1AjRkF9CnWDMzwTCDIIygybJDwZ4ioQ6iYL6
Rca+TIsnID8uiO79G/MiXxxNCXNunH1y/yW0YZDSkdTm8UlMVJca1wDhC3IqYi5E
T5FS2dRpxnAd5QP1YnSFXTpmRmJb/Bb52nrXymVG7wcGg4y99KOAGTmhSaebC8zX
fJFex2x6NGAJi8Ka7B0YO+ck+1u42hheDFzcdKnw9WodpIsVmSroafnRnlDuWLMg
b8YYnH4ey/iACiXfyRPj5bc7HQYV4DCFzpRFRJy39JxvHLGr1xct36lkBu5ze68V
wu3XtTDOgwKs6sdU78rGF8WMEEsQ5w0ZXhrI8FegTbKBvj/ngacjp4XXk6efPZki
bHsLlMIrHDhK2BY0+L7fRsUGdQrBZsOdF+Nz6HWTfNnyh5vruo3Ml49Ib6k6GwzP
sIbpPPoNOwGTviVqtl9AY2zVUZG2puUAwBimdqaQzzuCo4ReHAtRwhly6ThneIL6
YhnnLWz0Fk/aoK9n/1PvfzHRvJ0kDxTC2+2e/BfgbQimZv7Pac+BE/tVUIA7a/xf
BKAVrXuzMn94eXZ+Wr25niY0Y0LrrG1nVbeOZOTJYgOW9975AAwaGqYOkdfvxbmO
79s10xpyx+CVkP4TA+tPt7dI7LjQSyS1GTLJRk1B3ME7/K9HiY4xFkHiYcb8GgPt
t9h1FXBfJJdYQST81ECVPpULgJK3ymZxqOsSzEjhgV8xo7uWPAIu4IVarTitTQNS
WAYrVA4ADPykpkJwJ4QmNl0xZ7WXm2JGUNcL/0MlBdAU0OEons5brZGhWyAGzki0
1g/4HE0z+fFVVrrDCzCHa3lrnwTb9AVcvSEMrZwxL4SAbMA4ETp+PBqiWeXCMdtA
uNRm8Z0POmNVTnYlq7a/BW9EknRnAdD+1HJ1As0qelee18L15PQEGBF4nQxeGvzW
o4FWSCHP/Vyz0wZ0kiel8aD2JqNyxCAyrwBt32ZezZnrRGtX6seYhaGpxXKt4Qiy
qalGTwWIqxvMqrrI667CDQAdWvInaFoNayqaiS9Tt8WaNCaagE29JEs/EN6sq6gn
15X8xHTG9okO3eE3ik1Q7wsRg57s5Jds0Lj3KVURPMBugMGzR+5VfR2njxHF1fd0
SPprohwqqYt4AAL9axZodSBY0jeQaDxgTydxT2i+rxlBnYXeJ3rsTTICLQ9R8zpq
ko85j4YG5OqIRBukpv5FoCkt0+oMTN5rTOBwvRC9Q/BFQLWZmnqLMz4n8deqYmSs
fnMrXXmhjPSAoyhvja6t4SFGVNRb/okuauX4EJ9JAYdPkughncQyw9WWCqBeA9m0
+l7CiszsYWFleuogyGf9KfKkr4bbcigxwtf7DpqhJK+M8rAGzNZ9MdyryOtcPMqs
yxGq4Odr2WQpe2+iX1AfjqDZ6bA13POtMljs0kd+furhpUYGehJoH5CuGBXZi3Bc
hoLNKX0f5+rBsOWgkmW9rR5USvwM3Ni5FC0fSsjv90g/ddynHNYWys7N5iQcctrA
TDzNg5E9pUUYOjEK6G9iC+M64NCYmT2+S0o2Ixu80vugVkBo38FVuPrDVX43dG2+
rB778+9jM3fz2dOW6jQk3df9qmfLdWQ0qw7U7tZicfgAct7VWUmofc3TBQNmaTo2
LvzdzQSw2s4zAeYWqbwxGeYKTSwUL3LP+IiJ6SHM6Fl4gQLmRV/ePH5b/W+axuUa
5GHLf/ys1O8BjH48Z9LiG4PzWNJ3cVJ4z6iYf37PVbrRBndCH2tUumeU+qCw4lKQ
Opx7/3+0emEFDvaWV7/85Cil9jRWkKrYLB3aPtAqVFXaWCZHF564XEQjOEdvVNkW
8XPlKDzFDjRcTs6lsC3u/fAAYUkeyrkewvK0TmcXVPOKT6ggkMFnoWM1oX+Ix//S
yTqGKq8SUOrtAkkOkOhGQcjTt9bPejVGBIDnU4Twr9lsnUKq5WEW7G78p20/vqqh
ujWqUHnobelYoOTA/jFztPItVGU5OgeizGMvY4YHJG+1IVxPSY7x/72+NKU9nPgY
Qo7SRhwqj12oFxwDKnpP077l8Z7Lg8nizDxJ/xmav4+MluaLBhB2aAjDpMOyfCBu
uQb3dw3WcFPhBZavMdpFIeDkMhwsZBEmH39cVN6Pb4ETlTOQe95rPI+3VTnyJI4p
m/gjUc5nX4vboW+C500fEjy8nnzV0P2am0Kvaa5baQ1SNlGAyTd8dRVZ92jsHAnt
345xioSQziraWxcQDp9N4c7IpW6wgqyRMaOBTwOSw6Ip2goyMj3ryHTOXubEk9AI
553hj4w+PuFFsGosckg6gUgobo3vWOERt1coNu/fNXsMw7z13Ie7mP68hhwvtws2
5jjBe/fPLLfM7PFsjHM9YWTZBGcsiwznrhTJbK0/7+uWwmUpISmfueLzmaCozIsf
Hc7GDpTsEtPi+q2htZiefrjKIDoadvCSvFS3WPyZX2wQg6qRW21CjXXFoMk+flOo
Zc9i+ciQc0xx3ouwgrwVS/5HfcbCMJso1f3xolvKhS+d21O2tBbYRXWOWMBoax9K
VeOkKy4gr7frtAXgaiDELXlui/ycVHNNDvc3ZMnlH8e08LjfGjWK7TAkD6f2UKvm
BDp94oW2IJUNz9rpEumDVm/d8bTvnZ9yLHpjg+dEg6fiNOMULmEvCKjtw8EguhN4
LLWPcf5Qan+qwC/51AE+mVUro3/mVRHZlSP1OUpgfsUbfRXaOMr0IUO1HpKGAqs0
5XrBffEO9Vod/lLGEeRppksmHgENkN9r0Zxp9N06+itZE4IqX+O0SC551yD/veva
p7XWxA7KiIT/pcvrsiac0VevyQLc4fYe1WqLpvmgHs/MVn2dbw0VOj/Tb+8gIRvo
L775w2I0V9wyiNtMvsNsxz8nJk+HnTASUjs8QfNoTQqYcPSPi4esB6B9+5m+jXgG
+GUV51Ij2kMkzpldLuDoLomemsHkr+TrSVQMxqVvdPY/quEVD2rbBIm48S/ZiDpZ
rD/S1OHfhli0bqXAO6yi9p01Cg9n/0obKDWaNEulhF8YwQSObnhW4wfDMgROpm/q
W/NX0WHredJ9kYwm1a5PX2UBN0/TsG9awBA/HQzl2Ib/yfDkuVGilxgIYIuV4AxK
BQoG/iIq3+5RHB5z7aUfLgpOtKQX1E0s5sY7FEngwtlxcpLluXQSN4n7Y7/SMgbK
4+KY3pzDjr0MMrx4FK7D1H1qDvbePPRcuIG/nHOsbKaReRu/QjbZBNwOq7QM+qAY
UeBMotc6EK3NW+y4MO0OeeUiTp3GCOpbrojCEGFlqesrJ/Se/NlZfQdI0XIjCm1V
Qr/Rf10ULqsVx/Op7EqkDfLz2SoMOy/EzxwEbw73RxhTxpk1n/S0GjJ/CnmnulWM
PDnsDAE+/9Mgkv2SZ04dO9xGCBJCd5O9Wwao/Ch6KQqLBD+VCvVi/9kvwXGC7BVC
AJrCKwZqa7V+MECiJ1BCNRo23mvBdZtlJG6AtG8B8ofar0OfWRvTigoszHxn9mpn
h8Vo5xr0cQxsZNqkgBpAf/91ZJ0tI/S2diZk/VWFgLVkwxQXHf45WJi8IB6Wr2jJ
vJ0c1kNHr9Z855qT7sYFwRm0DEMEhTx+zJaRKwjFhZxcQ9tl1rlEcYHsLkfnjb/f
kOUIcNod9WV8M0lcdazqr9b5bOYJsZzsMp1KPooFm1FCYOErsGCgso7xLfGPjMFV
tKVZjwMWkrTBsnRpXI7bk1VhFv4UqAqVNANHBesv/dFMDZ6JnKev6DZjhV+RntCd
vHThGo2MLrkt5nkTgAu1S16/6/M+e//8TL2XbQSkb3RTNq4G8lktDN/3QfQKcekr
eiWS5ZZcGXyYXIiEhJhEa35S8Ta4iJmoxyv9XnZ+8UrCowMg9HxGT8qz7QfnZl8o
qB2euF68r/U/IjaTErGasCMLq5xTVCvviVmrezXpgwZg5ZErggJ2z46wU88OHhyw
DWufzMnlSZlD9X9nCPBPZaF3I5qqfKbtiLlR5/UnpOGWPfv7j9V0SFtFYYjUjbgs
dWgETtp+pJCQfogSF+BhOw74nrpq90hrh3AibvOox4oIVCsU8wNENMSYTY6kimfg
anE1F5fTFrubllPse3FYP9myVUuXLdaBpLWfoMQ++3D2jQgKx0F3iNFRjXBHiIBw
7oYLYzo6sirzLzN81IkpRlUxwJ8mFp6GpnOvuyTVd2RAkQZJWwvkrMNaqHil8+sm
rq16KVh3kSNF/kRshsBrxarpPfTYL5MT6O+0agDeeOG+PayA/E7Kq11jJYdcJn6M
QGRIIRBVyBg1cE5G4A4ZQkP5mAhH7pzsgxK6/hpFy/NXBx0sVjOQOqcNsVdqF4hI
xG8oT1iYKOG6HvOt1CkH3VbnA+Yl7ezNLq734h19HAq8RqldVfs8F+3Y5S8As5rd
p9mVQzg+61YLnf9u7Vv2RWZ+0PL06oUojYEYCXiZcAUF6Zgb8aTiYUIhhh3bEsbG
/oQNgTXy40KEmYctZIjCzHPXwfic/LcLK8qQtd+FX9U1fGO83y2DFVzHy4Q3glih
G5H3XFvyo1wziyBpl6RxxHVqiPduU77QwZITPLKOLJoSSmsTvzkXYl9VeN+5Q3/F
phQZTnNdihF60DCQxgr0ab6T0W07p1i6pjTffnBugiKDSCqXDStEF0RGdScJAdqp
GpxxuwS6nv9jqZzA5lTctU3u62ayJYDgZ8uoVbds6p/HFns+bhRmtPAfUVYPGLC2
Ok/PB1ZmcirWviNz0+kC6A==
`pragma protect end_protected
