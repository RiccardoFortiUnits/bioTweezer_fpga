// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
AM18TWeDmy3ahRGqcP432YEtFqABKmF8wzFq8/WTyQrJIo8YVkCMBHCDSF8+HrBuGLK5kDZtK2Es
8KKSi6Ffnbdtpp+j2N/IXnvkEd7JdEtI9hEPb9q9hIm6q0nkQyLFffQcoLUaKLZnNcFphKpzsEbL
RZ0RwBxbQJHH1nMCRVZwPQlxX/eGy+jIpC9cYDzh8BJ0f78ocVeoEiuPxdYd+IWk55RpJZa2hUbr
RGHQEk5VWo77GcgowyLh4xs3//ydJduZWJks2wSunMO1MzFZ2ljDlii2mcKk7CkOF12X9XAGy8E3
8COdgECXrlE4L1XnsTRoj48UHvB843pnfr0aEg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 21216)
/hU2ZU7CECF+4VUvhtDjySAoHkzeR2n/iiEaLWDks+5IBYgfg88mIZqOsmr7vIHRwVjCFd6QH+rH
JdwLE6EA0kShF2XaW0uRWQkR9XG7jNAk2Mclv7n2AW686OKFUZ1wg7McfejlKEbmYRfYfSLv4LC1
RF7OoFwGOdvUncQDNf4cmr12cP7A2lqsSj+ho9BBps055oDd6YMYkUzdVE0oqTROgxxC1mEsGfTg
+oA62o8/vI4tV6N11PQWWkNbd6/i9PmWkrYgFBwlbPmEDdVE0DEAg9e6La4n9G4wBVP624yM3vt9
Tchm9JDTpn0Feu79xLjIPoT6zksVFJAk3r6rIJpzMf0QNFKyYgERbp25cWLPTIytENZblnkAOz90
Nxf7Y3CnEet/Sc567ACjvkP7tVx2N1i4jVMTFueQeYPRoA7iwbcUxBD96q8ETZEP5eDMy9UCYyx+
EIu6tSCij3MIdiQLbp6eKiFWQ0xVUvNCZwDDZC+FymPT5STMEpKdxRE3yBVpe0bDFYij8F9SidGx
2wVlRulbuo5RPymS7M+rz/RReHRo54KDXUISRJN90nY/N3nstDFNJ2a8ueTZoPtfSpTNMCg/2QYI
toQl4MrDw1eI8Hm35npW0SrlM30+L6QX4be6O6BToTuODbA1p3hokC6Fn5dh9r9OKZqMkGjzfO0t
E7IJZrKQojqZ5fjc6JghN/3IirAff5PBaJBtdhBd1caX0+1CE3XXtD2tXQ2G1bW9sf4UPIRkEkuW
HHMBtSp1CgDRoJmTCAWmMaVzw7iFoYdZU9HF8ApLnrHPMmh6fIHudY2mNqY3wkfZuqp/8in//BvF
iLksApAUTOYLLBZWX6sT4iwlLZn/KFCDpNWA2G61AYf4p7uHoHEDfTk1GamLULXD4EbdXpursT4q
NxwBYl87krAR7tz9G2hV3p538m4zR4xqJyB//K0LP7JEEkBfU0jv1SYTjK5ZtorwKU06bfA4jmIW
yS4ONIzk8wnfu3XH1GBFAmzyhKg2+B9GBMAJ6zaG00nZEqtDWzlgZans6eb1gYfDZ/svLbyxjDDe
9p4b+5H62v2/3e+JgwoA5mJeFmuWOwPhOcDTmxqX2MovQOAJTFuH1qqsCOIasfCbxJu6LCfDq0hK
GIdszfvdszIr/913CXQvHCdzXz5pGBv54CJgSYQVRJopz2eofAbvaqvEY23hAKJaYnvz0AI8ikMJ
i3Y7Blo25e7IiWsbRhLsLACNzOJwn13rM+OjeDEZi9zTXmYeA9eNeUPFAW9MqFJD9LTn6E+I4jx1
PrI1YZ1zmo+mYN97vnjlugwy1ld+iB9eIKzk5QcRZrzWlBKZHNzVSnqbgBQsSIQYNYvA3VLTcrD+
U50EEVQo36sUfjP+88TcBB2ZBw4e9vV4Zi8ex6j1bwJzzL4QQvt1VCJaNYoXTveDwSGKPUQBj1C5
ramTUNNV1sveYuvfYMx4qWTTx2zk1WRvk3gezOXTOFt0+7zEoCQe8SjRDQy8/8lRRIVHjCoU5pH7
x9Qir62y5O+qLFgeWa95SI6oyANk4YbrUvm39s6ar9HTcM2kQFf3miKPgiwfvUJXSmEPUACIY/ty
4Cm+0lVf+T7N4eFEBEpyXVLjLswFsIIZfvurCAnqvPlXkBdPeoJt39nwB2C/mkUl/nBBIUrK8M+V
kcpJMIDMMT6FXqoh51GfakNPr7wzIHnStW5BLC634p6rndFdmTs8M4OCXXbZ8MmXBEQ6QH8mWf3i
FAY2SecdPVKkq8U4EcC2l4fSCnEsFU97OJliGubKXqqcyVhkgKF+AghmbNsLPLue3hzHMOFP14NO
zeIv0UGcU2uKpLuFP6IKmtYavDYqQcbK3LYqBwepRUVBznWpjLF42xCJNJnqkBcx4+qVlgrqAe1d
l/kUNTsGcmMjVucYnWp0+v22dppuknE5HMLhsQPIkEdolwOCp/KCKeYEtK3eF5UAT7IwQK2gVCDY
/5ul8Qc6n2YwC24crMOCsS2Rrf8bVtYN2YGzmKQDrGRmTzC0T5XWHBo//dKORYw1IPV9WRvzTpQm
KyMZSkcq/4SuUZJzXdpKWvD7kbN3TH56y1dZS0BIHZTSm2tN0Y5Z0vZG94p8jsCUcHZdfjr1lqI9
y4vS70QgWZuJZm+TjUPpOMuTuZsK6Z5oI6EB3srKIl+vayIG69SjHzXlNqkheGtkFumiq9QsfXro
2HWYOAsoyDXcZgSV0/SznSjXbTrCazwcNVaazC+LvsAK8feGAllIkqEwRaysk2DoNv0hLDLeYrcj
ynw/UYcHyrGKqhJGCgiab/VfJjAEnC1Akj8nw7RlqR34MB7+1lVwho/LD/109ejgBil8rID8jfD2
2vqzqQ86sIlPiR+2DNBbxxnA7B+gYGhH6PMB6llVQPouxc8GOKi0BoSP3qKA4BeALbCKvmizn5RI
umashQMQSwVokfcSP2G4de+DGb6jWD9NdZmuO23fRZCYXDE8gmJ1R5jaXuk5LR1nR5hdunsirB71
oZ/advVG1jXRIw2Vb/lmCJsgIwT36FwIVrfQmDVELR+wHIPFS9iXg+FN43yRqjwrBiu4X4POzuDO
hsX+zSwxPwJAm/lB5qwdj9XazMbXu9qUpQHCJI2ZXstKKeEUN4wXW5PvxK1jcg415SWflmODQA89
uHE2+flX04WUEya1PjARd+ybA5mRwNnZHS18elJAjqxdDmIhhP0qmMwutbeQuP4p7k2Zn0a1aTGa
bl5T3KUdOh45L8O8G1RU3BgERxbumIdJkwT4BYT5vT5LwpSj7BLJn1ZQ99ZjZeg5XylbEL+aUxQy
bQMlaL0epIGOuxtXxSpzYeYO9yzqJic0WGy9z0wQdHQp/Yu7HRUErnKth1R8xUuzlH2VPTvNllRs
A7olXlxexdzE5vLSHhhOYMijdIqkCvWccC9FfbnCl71wiNaB3/EANzzlRBEF2GubnB+7NMeBi9SU
/DVC9883ewik+3PfHeFb7gjv8iAdi08pKk37m3lU0zX43ZY8nQmLQ78+zM4nac+Tmaq1I4fnKJ56
uW2CPe8r5D0ck9qgISMPBsD73DbqN9LXsmIW/pwP60pWHll/l8tmLHrdtZeqCyQMORfLq6EAkpxH
aPn7GpUAp94b945miHaHyMDJnS6Xd1SpkEfYwH21H2k1/cHA9UQYCZrTonbfDOMbTGPerjrEz2xK
tiN+/4+NKW/FYFsTnGC+yeqkYOgPFbkviYa8Kwmuk7b8aG6bXEfPeQdi78mkCT/3K/jjMLaAztgs
GlzeI/bL5A8Er0gows/eirFBFaXu6pNcAXbK3Z7kea7/mubmMetAlIq/c/5N6FsOG6U3aVEUbjaX
PKGoDyg1UR8Nd5yphJ44bXv3DLYXRd3f89EmIZRAWX9fYJZ/YJLlWiiB11Fb1fIBrtcofoJxAwVY
txezRGTB68SNLKByWCnpo2O2465Tt+kTxp59erPzx7zybVrohhPFYb2EzNnV/aFpSW+YM+bAG1Z4
3B4WEL3jKng13BiLCtsP7Av0coEWM6mzvSO91160nMZDjQ7XuM59TTBg84VshiBJAdc2jiXbUrlf
ZNaVHPRP0892CFpQ5vT147FM0zPvRU5VGYbOCzze2pCi0o5ChcCdSzvF5Me+Wx+gg0QyV9obOTYp
5ji8Yw4YTB6Ev1uhl8Dm2WTuvbhk+5VMCmNKRv2zs21l0TG0GUDrZ4KuZhHcyFiPfmWeCbakb4Ep
fNilKdowu/xamCUt81ipnJSYbj6ho771kIw7jqCiRWEoLiEnGPdTMFnjrIxiPePMI60kEiy5hY/u
CaBZD3lkrogeQN9EyT3geHXl4d/anA1Ba+JLJHH10yNW/pUaF5ze4t+Wr0maiIRxfDyyc34Zzkz5
Txf+48J12az0uPSUcy5zfwXKuxz5IqPhM8Kq8U+fAXIPznPvJoHwkBUvl9B6UBVzpMjVk+RZjOpO
imSvmHkI4OBawLs7K2IZn5SgNAhWLnU3OVYgyhGEhIuUf2tN1RAaQauXmQ2oFh2mYt1TkO7lTXY8
SLVdoIDRHgDP7NoRppIKperUPBMeQ2Gp1LscLypbJwQr32ZIZRp0lwM8Jjm32eYK0+yO70FBaU9F
qe8r3Gqt8J/14KLhAR/5ZR93f/45sO0TABbZW8gnFOYZMPLJyyTBK35cMtGE5nWCeG09jLcO4iXc
TPvARltcB+vN4eSeN/xomnLrXnThforPOQxZaNhsslsWhCZckjXWHMq83Y/rZBAiJBLRa/j/Ku+K
xwGeHj+8OxrsjrbqI0xyZG9HChvlWw/SD9Z/V4OLFW/8oN8vgsnaGywsAU+jrbJtFALVOZ1Olx+m
g6DpgIibdcrPd2qFVAhJL2GGQmlj56NRQ3eEUYg08BeaiviApnp3xHdDggDxACPbODfVoJ2/ov0N
cWFRoGRzBDZbCBZgU2wNheOMIjh44WqshkFAs4bKlfbtW/sIqQw+8P4m8DEOMtHsQa/JcboyzXDt
Lp54y/8qYRYFL7tXbvFUJwzSQRU9hE/e05t1KNMqsPZVQKuz5BKOrWhah+rDNGoPRDUH44lJ/9G5
SEiTz1Hsy/jjGCccEiVmiM3Pj50Skp+F0IwsE2lQlVKghndJyI9xfa7Wa2ToXlRQeD0iuw0IiK5o
WzWH7AMllZNA6Gd4NcAm5HVCjk6OHMUYyX3grNUcLoXt0U1lJdafHmGuim/oFYjRoWJRGXNqbqTB
hm2lxvISu3YR0UAWLpC4f3seX8v2kgNOvHUWmDUMw2QlGFHHDq7hfvCZKyq9L9jI7IN9v31c4g8y
Raf7aaquxoQyZVdtHXVt3sD0+ujBQX58z2khFMhmYkVevliraVlmzrKYxi7T07TGs7FTN/VveBY7
BNRMBZbeXNWtFwHjUXTiEnaq26SiCuF+028+Hwi98j6XSeSYxx7+QzVge1qlCw5DMXTOiiHRO9V0
QQcDgdJjDqQ0SJd4hs9BXOBYJ/63Enc92L021WK4cTW9VzquGFwVYysC5e4iZ1btG0A8NljrF8Qi
xK1gGrR+gWAZyURcC+rpBz4XBPGSOMBB8zzTFi+Jv6Irp/0T/kBJIqXyqMxILxmxC2PG8kUzRQ2n
hPfWxZ1WxweND44f1lsfN5SNbjoiTPu4RMFaXCbHhYHp400D0ekzY2wRGBIiTI06WcflMHYVdYtZ
qtx1ujD5dbLfpYYzAdN+g9WRjKl4BSKBu2v2fiPDIENfVzB9FxRY0XNRyUJTTYv70Hymb/fw0S3x
ouU8pqt2ycuGCv6VPWDcFN2Q+OZZyAns8eoHcumphgMxYUCvhWUPWI0Nn60JnE13PuOUhFeZf7rk
zneira0f1cCCgsfd9DmTa/9QyoIJnOfFH82tjrfaCi1V2S429EXAo1MPIYfFj6D9hLaqOu+xcTfi
liBvWIlt8oKm6mNwf/xAchZCNTJ0gvU7s6J9ZuTJrw+Ou7j+CoStoQ22q/qTh+5jm39AhBOxzrLX
KQ92YdIhY2i+U6RfGxNAii1lPmbwvsOACwAB2GfLT3OEENR907z5E1nDrvT/NFbFXyQK7jkMzyj3
EFxD5mgdIreafD1pP1qe/uQO3T9WWFgQy6RGYTtGvfthX0qX99ffkV3itxyG1NShaz3XTG2KYAIN
6NiJQBMp4E3i4UZTjes/iHxwdV31S6dQSvJhAoh0dqxVw3ifSUBIiCBtleHcMTld/YKSQIwmVteZ
scf0UjQ7BrOF2u8cDwX9+QXKtLdiU2j01dDSVhYHYyWpip1Pyf3tz94lY5POauMnA2PrLTpfQ8Dj
bLOcmiw9Hf7I7mnTkkI5Nfz0X7zQ2va3shnEUeDQ7I+pscVBtrIv2BFwWd69SWkqvRnu7d78n//Q
g6744eCoH7Z/TsQ9UGVyfjBKdsCcow/2UK8H3N0kl1fjbm0oAjNt5ypdBg7X1CIpB6Ns6KjkJ68D
v4A77cdwhzrYc0trCx7xhxUmbsvHJg7WgWFLzi+fXd00Igh+/zz2YLJ47ExvUoHqsE6OZqWvzsEQ
+j5zggRqPyluaQdDIqXWs7BuxHUJreOGNHMb1qpPRKwTAjB46V3K3ayuGhQhyvvwXh4S7tEhwW/S
g4/DT/rTlznpWfBucKaj+ZZq16vP7XkRitqFq34vGE2oZpG3qhSAC5i9lLgj89RcY2cfiToMob7f
Ffkd7iUk3t6Ew0QE7nOXLi/D9JRsZJaxjDvjbflKzcktS+uUKYKqJZCebEDygazYo1yU+pZfgVfF
h5+llcMUT9/N/TzBZUkzoQO2f8vKJkD6LIo1323anCZgt4LJ+sEYfnnCby6BoL18WIH/yoNyC5tC
PMQ2ScerWJ3mtPOLDo5Mqy+WDkrwyXLC+Pa5VF6i+WsiajWyqEeZHZL6g1K0putiqPNo0tauZun9
RHlCYmzTYURGwG2QUQfjCW1oBS0r2b9xy/raVw/R1/G0tm07/HBnM+EHcY6H53TMjJxkkkxyK05L
gvHMgBe8KOjfEEhTeSuaHRq0qqWnnOR/O0PGbcW2pwkm0ZgRWLhdBGv0PXIZk9aBjH7JuuCW1jdV
GpPZmzvEsghnGwUy1+/t5EuaHHnZ7rVUuZ7FwoJPT0pmHFZI7oS6N4BGgGgrmo7EhZuuATMdtRN6
jasB7wch2SDr+z6u8AbCrSbwmZEmtDrvHREB/eUzduaDtfVQQKwY+OejeysJ7o49NjmWef7JtJ6n
zMkZXEdElrU65lN51o4vczp+lHTJ+OsNR4nr1BYpTfJD32TbHKRWdRNjG8SVtZzllypiJfQ5R5xY
xug58b9VpA2E2rzRUlEOhRiJGlQSMf/jbQj9T+4IroOxjYROrTsS8o1p378A46cr+8Wt7eavky15
9vg+5dzrqfKeeOkiI97vIoQPj6WOKzHjWLeDpdumVevb3OYkofOAu5s+SLLKV3F5eHCBhJma33/5
r6p5zV9NKBFsuoSdTKDvmk3tkMov2bOLKBQ1O5rW0Xw/Kh+Hmze+uju4sjXMFTgb9C7Yy/l+OIsG
EiPkmKaeII1p0sTekdlAahYxhtz27C4prbjtEDZnc/CzSbNowbO8wbxWcA7VlFz4nCCaurQhWVw6
/bWNvIHzwwh7C9Q+JFA8bVad5fzYE49d24BfY0zdO4g+pl0bAnk2aeQOSygVwCPBTtWkAJMlySBL
9v2w0KduYAJMbZr5mfMHdMK5Jm193STbQxQQJRJwKrTK0KHmXn5Lx5+cGmTCeGSeUulHLaHDyevO
nLWRmV47VBg33nju18aLkujmIEq9XDX3LBl4XmDkF5KdE3gRqwpvgzc1NAp7fzFkQmF+v/c7XyK9
crON5IIPvdDJft8xnjjKnT/8YvtvREMHkeYZnlGzuGjHurOjamN1x1fpNe2XWJ+YBU/gjLd/BzZM
ZXFOpVCkxN+Cz0UJNrNkOF7ZYuaV4isNlr5f9y9BPfQE0IpUF1vhmSsiOGxL51nWZlUd8N4x/XNX
IaWJJtXEHilkg2RgqQ2k8rFJNG647MKg9pul2SOIy+5w1LozjuA/bSsKSFMAnXkXGCq3xTmg23Y4
Ex+XC7ha0T7KE/Sg0I+idtdNBZfiyt2RpZ4MHTg5Pe64XClaE/bat+9vyH8OV8r1tw2MO2m4SQcy
fREpyfDHDbsLYV3PVj1L6hqKFpc1u81UtnjKQRra8Nwpps7eJvCR8FQbGiWFcsKWC5a6WFiBduEz
f18fXDqM6uyMRIi6v0NqmpXrqWnuUk5mT6NU7Dv8W93qH5Apdvp2+zuKJr+mcpWgkMHZ+oSvdK76
/sQ1wzSsst93+OOmUeHKfHDIkn9q/KSVCfmWIiOTOhh4R+b37qxqhxjyt6wi1tCdDtVls3Pi38eV
s88F+3L+thVUmk0FW6jQC2PHZefcGUzc866+t9FpQCM9p6F/tkLSF6/uqxlZxxQbq03gtNeFYD8J
F0I/sIKqHiI4OyInF7J+2Npg/gXPVbBpIPcqR9D2w8qcYODsZFHE80ccTD0A5Gvesl5If2rfTmcq
/066OUuAz966Q2zqnlHAJ2rBRJ0UIMbYYMjsSG7/w+vc20lvccaDSE28p8unikTyQD+m/6tdjHW/
vQre1Z8O85exs2sc7f6q6oLrrXLQHRKfV99oSenw+s5K3xqdXPQ8OCaIfWfwek+0O7HTe1quwGyL
lxaNi5Suv2aJ+8cZo81bijQVZhQmF91DL9u6b5AHe9y2E2bnErXa6Rw284++D8lI+TTTRhIAx9TI
aCbEmTHh8Rj8HJqBqqLLJMHeBu7Cz07aeozu57JMMDIL43WKhBaQLFfnAFRqWnceQnkYlBoX0EV8
SnsNoSlTOKc57GJNf+dg8eeByp/b04Aiv3dYazsG1q5S8osHmO8guSFBOJEipYgRTZHtB6VVjyEX
roeMRvzT+cVIa/091aRpUjpX6Uj5s4HnWV8Rht8aDcY7wjy4+eV8NsLggg2WhG5yP1VvkiCZB7UF
DExPAguvr+NlfvqzpBx8EMOakrVgf7Gzg5j9ERBQ3EZoOrLUdDN2NAGi9R0V6GIvbV96sLGdsEtb
3YxMqd9UCe1gMs0uxAg7qMBLWnrj3g5sh/haLO5BJsnt98lJEELLLNnzo/Hv2kgrZ7CilkJgNgKP
l8JK0BeeekrVwYn3FtpgIntGKkLSFNpMe8j26yKg1QA+rTeUPSU7yCr5EK+XmK6Gh53f4jOnK+tE
4KM7BBgRxnMS6mDEIkOxPoIPnE8gbLVxxxmVJ2nQ+2DhOdb7ko+7XOH/JUBpCARMZPsLkq5P9L2M
l8uLF65MtgdoFtMEknt71+xSmFL/PF+FTlRSGttSSdGZJKn1ymTJFNVVZtHQFP3nmIST9cRQAW9r
0Uwpho4pmo+XI93V9+v1/2jGzd20LqsDrf2fjl5akYiZ/q4mthWe162EPWQzoyrIE59j93UKPPVt
wCM0NNVmNcBYrP+/xpkDWx13o3G0Tp63g8VqsY4A/Hfjdcf2acOsaqd2pPL16+NxfP1ZIUd0S8xi
9alIdbXfYN+wHF6i16BkPXhbs5cKxvCnAdF5aN3IbHIdgXxLeI3I27Fl4tqSycK6HViiNzD1xg7s
aIId8hZlJaNE3cxZ/R+seXWkYQYvnaclgVgVWwbLD/GmeXcUOakXNxvF9qn5tAm1sn4YldcKJqQm
6WryovGmownghGGkX+8BD9kHq7teVc1haFA7p8wRohuE2iLL+jh55oWMyOmjRVD0QOR+nQZm/yii
8NLkaxDJEIpPicHlJfZI39zOcSRMHBzv3TSTLfiwd/1Fyj/HwKUV8XNtVqMuvWKcXEx94rMEos3I
LTmZsfsdth5Ug1AQhjiPbBWnT+GqY5DnlDBYdbEJPhFLI5McH5qa1xlRY9+e9Lu8HpuohyQp3G5T
4rcxP4U/x4Jiv6m7jwdcM28XiKk39uMJcP7pPBdsN9sIFZzdj5b5gBEZY7DqkYbtoR7z76mbahCb
BjZmVYTPLQJA3T/MzcgI85/i7jqfazg1xsHskFHhW64TrUkQZJyPcDSvFKHZ5TnMFafyGIiboEF0
8/bR3sVC5Ug9FYYFdJT64W9kybCrP8xgmg02U44qtYtvRCdKUb9afBa/RpGTSZc+yinAyVi8szii
hpV7Wv+6BCQHrx7oxIy8S2fGAwXQFJ/QfLeQ4srQ6gShsHdAknqyOuNXao8A8Dk2hsmudykdO8JR
S2hpkTZE9F/JmPKWaYnSDpBa0cmu0LTUfcHjPElzZFMTAOmim/wEyHU6iismQ5hYvQrn+tBvJAp8
+lrhbtHkZpaDnOTiDEO6khl/gQOTz7s6pstZDskcrZj9+dd5ARRvtG3ltLBP/JV4SCjMJxqwAOky
L+o5xI3vk2+YpXSI+1KMfWWJXXjEJN9cznFsxTqTi18sIklKjX1exEloYjmFiMVKfLYeQbhInoOp
wYdUSyRnsc90PDR+PuOKLe1kzeJdKB7Y/ORi3g3e2+THehcEuMROw35Rpcaoj7e79m1opN8Ro9l3
q7+0HD94uFK1zki5dAzra6r+c4+LxWCTOGLqS8zNehc6RI/cc0cV2UJ8/MhjddjE2U8ETmwDpla6
OsIpHf66pAdpVxhMXkEhRjgRnJ9ld2b6xe+DgKPNRgHz+wVzuCOhHb2Rnja88GT6CtWgU5D0e0Dq
rLtpfyw37nxudQ0hDmr+243tGzU+G9NOy1dBfAxRcU5pVLSm4AtEXhQmHNwR1uimPMFn6Fjaqk+g
/1r5Z/se1ui/mUa6dM8M/OANo5XKvjdv39nKZ9/FQjsMSoH/Y3pBX61/KpG2nNnhIUxisnu4RkO9
8kXBTIddMt2J61bgsbTvssXH5oqhA5nXTrqtMEIo+Q8U3mGYu+TwkpTXL44TEnJn1V9gRZC4AoyR
5x8jWaD7lfXLdDxCJ26N3EZvIW/MnpMSZSNjEK7c8VnC5NMHYQjYskEd0OuXxD7JtgZBoeh14piZ
nT+heGAVV1mQCnZ328cKoOJ4hUqxuCZ71EoK86/aRD2fCcDwkpCuKRafTk6wSWOQsvYVTZTi7U1f
NgRr9tDGI712SjsI2GabN7MYrpdfuv7mHnz2tETz6jujtcayJ2szMtZQGsq4AdKK+zl28SCmJv4U
WvSWZGU5c9pIuNpk5v5WpOSr4u+vGNu+ovuzCvGz3klZLPpBeRL8NhqSANutL8CRPTNepEI86AW3
yMVA5ja9F2OBq0OHF9x8JmnVV7jH1rZZFWayHczhNYB8tj7wsJ87alJTOjCuoYkkqrdfbGhFme9W
CphoUWkgn06pkP936bouAkjx3+QHOdqoJtab9rQZBqmz9lWdP1YDUgaxRbAzwLcvT5cLLz8WGa57
XyCI8tvi2tX1NLrAScYCMHsijJwWK9ykHX7y897hX4PI1a29on390IbCtGJc3Em9GQAOXqyegms6
3c+DTTlEyCDrZ/CU/sIZeUk7exTzi8d50ivkjRfgmic+L30E1XRZxg0L8EamqMU2HsDnzXv6dnh5
sO33DSvr5XNvI5pWzmJpGmIRzjDyc/a6lk+iyKKFrugvsQuliDwFV6h8iNUZNJVAn3crrIjcgu+B
y8zLmWGejuEYHXeSIUc3JcXqYdItOk2kDkOL+pS4pUPcZQw2b7c9UR8dMhabcNVvWJpwdhSvgsJG
7adU+mYDttLIzcDHKBUFTTbT4YZv+8opcpUrlikMtI3oMvud/9/M8yXVARVkLJ9QLf1TvPT8K4yM
CRO6U25dy899AJ8zlo0cYvZFzZJ2nWkL2Hxb6CcroeiXn9wnNn5wIODnl/1kLWKju+H+osZgrF2+
Q6L5LetBF4WUW01jsLeiqbrnldSj1F6UzOvc1PkHJBNZjm0kF8sGUSkleTjjoXyBtoohE1VxT2z1
17fghclCfZfH7jz/+WjqAa2K0i+hyyit4Bz/14atWBuhgLSfLEKsZ79pPe3n6YnNG2sfUZHPm6jb
Kp2aYB2bYh6dLsItNIDB0oMz4HoaQWbwEtNjn1RzrbtTYdpG5QwiJ1CT7uG52d5aE7+wyMwDQmi5
AjCo2ydCjdqqU799N9GhIwCXmAdY9zqSRzP2EpiEm2C75syIb8ZLM7zWXkqz8fRzwUPTM562w8qj
al4diPGlfU9PfaTrpTRtNIq4pqiHvnwIKyo/m0l8QZqkwwj54NKYGG+b2jhKjcwQ+CeedziMR9KX
9FAN55QI15RyK1r4/gtKVG2SVHdBZgnidNNyuq748l6S4MLTN7s1XypVly/6A7wUm23EFt9gpavj
8rEmV+ZE9W8TZ278+ii398wY2nX4Yz/X9YFnCzDLP7WAY5P7kXCIvQy8RZLEeJ4w2H0TDRgbsb1r
rqHtcCioTRA9GA/uwWIUj1kWiCy4wLScbi/sXCtfad/z3xZvQnVuv2GUyTnuDncl+dxz1P+cMRRv
tuMGglXb7L2xSdTTGkMsEDo04GfDZLORWhSmtGOr7E1q0WteEdueKMXfgEwlBSTmhtMR26VDhrhe
rnaZ79d4lieERDKDj/zj0x+PKg1zg4Kzpu2vqCIONk5jc1CvBT5VhVjgxxqimLqlB5Tm14QHJt4V
xu/nxzbmKx+P6TlS7H8Gj5TJ2zBHM8wI/VDsXWz14mt97ugQNqRAVhX1u0HqTGIRv1kz4f9mj1f0
CkadJwva5D6/jatcXS/zf+LbnMMUeZdBqFPlpjV8d97jU4VrPWId/XovZ9aRVjDxKjAsHh2zPs1y
Pdn7unN6RvoGGSuqji5cWLthvUDdpPeAkPiLjWYxlp2htWam1sKDliAq+MvLdNlh2BH8Q5bPXCTQ
ak/5eROoPRPpJAaC8w8O7VFqQdDgcJPTxlPmHA95GzqlecndgadaOzipgElTMrs2Apk3xR1aZNKp
MQjX5aR82ceh/Hxw7FEtP/1O/Cniy9NLrHOOciQgq4x0GY2GjyxOz+l/TCxbwx3RIYgtBbsAM98e
H35mJfn2yyhNGepW2kw07h43oOjjrTXVzl5A+OJEQxLPi87G3jBzVl1nZqK07jtRtFOy3VvYB405
TKdl0SWggtCZJqYF1FhzXwo93tSNcXZGJ4ElshVjupOIIKHQyyJ7XVvichaoei8DTZ2doVnTikDR
+dFDRUqyyXPwnAUdm1safuPQv8F00v9LC8bxsN/PX/fw2jedKu0DLVkMOEjXAc41E3jXhynB5HB9
o8JhpK8DCGMeFoGWfl12/0McH4CURIJmvXBY3eVIGA+mM52ikyCptr4yKBnzVHwEspqXgNdLyH3J
1y02Ecil6sJ/Sv9CBgxGfRG6N+Z6oqNskXQ4IUb9tjzdJd2Eh22Z7rp04S7XirWXorkIXgUR6SQ8
fAegPDAAqSr5fx1mlNDVDxeMb6ogUjNEoHnNN+G4WTeCD5b/Ltn11IcM8/UH3lfrBu+Zt9rvKw1j
C0ugEWjD7kDJyKemQD6ckQaYuLSijcgpFCGRwPMSaB0UYx/9PPZ6Dk8Wl3iKxWx4f6pEUZLv/eVL
nIvsiHDVB/6iD32XdsoKNFuht7wt5GkJ7nnS4LRoVYg4HQipviQwxf9Zq0EEG2y9ZN9PrSnggiRr
Np3WvTV3i/o+Rny8jXOsXsYH9KZiasrEhpwf1ypGSztVo6U04p/tCwEZwnrGBENdHbZ7GTGw2rc/
7PYkmB3JWnep8Nv56wU9aLTwV8WM0CSMQ5T5M6od5u6mnYasHrYunFCO5PbIUo8YDAuSuKldnlI8
hHYvymm2cJtB9XPQJ4z8Zki8TsIaFgb3CfM7MGPK4B+xOsRCf09zYcOOwY6q4/c/BApxokDfhZUF
/k9Wjj3ukn8Ku9r5rme/37ABVefdUXWjOhnrtvvd/zjxMggZdC69c6ShKyOLiBNC/twvVxWfRU5Y
xrKbdTtX+tY05OH9wlAysu3JOn0P2ValFEiadFmPBWzSrlHMb8tF165pqBbCUxKg6C2fsp1fE8kL
P8Ss3DGuUOniEHkSP+uK8VT0PXZGkNOnBaKoY71MgW13rYJbP6IzwE/qiwuqnjUrQM3WepzRbnEH
MIzFuxv9E7WNfKFw+ItR2GV4tpbc4rH1nU0C9qb6OAOUrD39imT8nzEkBrvwc6S99oNpiJ2Vee6W
1LM/DOMqcfn+goQCQm6qHPk3oHGvHGa2CJBXDIYpuC/DHKJEf2L5SkU99n7JZ6hBbQtZIc8Dyp4P
a40jQoixILu2mob4uZlRjQOifQEinsZblNMqdz1JegnWHYCsyvCgHvXA4J4KbRh5AQNkxOuDa9TC
gTV3Sqrx8or1kKJV34Ag2y/JVuLwbb1Mnzh8dcgvj5KRSAb9BqQITId0f/G6aj9N6+YYgLolOs2w
RbxsYubA5wb0CAtyP4svFsbM7fyd8z6aiKT1yqNbizv3QCdleBtUnZKNQVwb/KLjamFowE60WTOG
uqCeEHpF7flsdCWoy9LN69SAOEnMF31qqqNt9Rt0sJEo7dLLCiYptzIrVZmjpT9txksBdoCcukHk
Ym6liExl1hVrt67ZdVD1NrrpFgNIU5IT0WTw+h9Bn69Mxzk6K3s8H1gnu5GAoeB1jQzGCszoDcbm
p1vLXS6ZLiDqOEFWhSvWAnensOQE/TcHRzlkMmRSXDhXp2WrWYOZC7prc6M+6PRVytFMIaImKxm8
45HQbA3kPmK0rv6EGQgcJNoVLbkm0/wKp/D6ECAQ6iOtTg38PdH/v3SOtSfpiWtNqEp7ufm2LAXN
wHblQrfORnfSdZS6RwNetooBbg/fUzGtwvUT4SfEeYlGHyqWj5UqXb124xPuDuJQS2piOM8tikb5
nkpScIg1uCUeCWCJjcM5D2t+GPNRU7PLZ7fKC/+zkQWP6DCxo4/YOt5zThHyC9ohezwZFzjw4adn
0zbl/iiRF2WrEtaKnOqEyB7VZ/E2UoT/ql72iUHjr+h2rppwZtcUBEhyQseq46b+kGq3FzyuBCtt
mQHIAnuSq6aStobIzuRyQoj54UsqBQ7w33DybkaIwLiBFrmSwUjFde4Zarmk0wm9PBlqwr0K7SMT
+LCgW0M8hN9R3l2Bk+ry5kueHgjEyV/00yX54j61+8Nc0dVsAuxLdhgmgAXTtSPZAIpwMskh9z+9
aM5eLzxyGUndpq5SU9qxQ+OeJPmYJjvxQw/R4Orm7LxJibDtZGTzlEil3T2RBl9fSZxLLmIeIQN2
QCMWhrofEGvW+n/prlfYj1dv+SM7Jgv2oXgHcFOvQBq12hk+uuQg3xWz2YJM6s/0t9cYhhxo+52y
EgMKJw55C5A4DUn772d423QOoFBEjk5jhFzqWKyXeoJ5DNv/J+ooO+8gbZq0IIfVmrbpxVbPRVSc
59fSchKCffc2ZaqZYpMDkxVp0lS/nRpE/YBuXPAyD2is/n6AkuKJM13ZsKWZzdFnNUENObHHi6Ea
Ff4tHU+gal3fVs9JC7NhQcWtgoK7YAOS+KLb+MyVcOQqqc+CZUcIK1z7f1SNH8xZ8qQ7OlgDzKs3
6PNjbeXnJKHmnocgU/oDvy+S1susJIxNS0FWV+r14Tb1M9Z5xSrGXfrFfi47onB/9+TxdobsBHEu
WGg77oNtBgeRZpnNzw9A/bETKjyN6pIXm58wFirJvQwk4tnYPIR9hwUGAPR7uRcXtfwL0cMBm4rn
20BWuAVe4g0JPt21rAB/oK6jFhjrCBDf3ehfFOigi8Gqp7xg+mxhgoH4rHXt/nKxeVrO2dtwfu6W
Ggezka1+N3YYlRBOGrApqSdfQ6jG6oESO1ZAfREIPKnx08v8vbG7qO98UFhSYYnfTK2rdJC4Urgv
On34lxzzRjRLp+7lRqbm48uSYkUsoB8TOQNIqcJuiPDejKZPu+vT4CcwiJL+dbvBRXX5mtzP1zdR
m4TplCEgb87mCM/ugI+7DspaeewdgYcd1fVr+e0wdWg8GerXLTK2ZOSolj2tqesoyr8FeaXoGquU
6IRvQfWmcGjwse9PpuvrfVA25JEJnL9KZ5HA8Y4TsdaTydeOxB/ECbzt7V1bgIDRHpjtnvlXicDm
6GVuuMYcPtMWxRECJcxOsqhT86Qy9kwMQKbGegO5JKx8pj9c6YiKSr4wdOzULYMeVooGJBPlumbW
qUi54sWgUPtjdJew3d4zpuUgyZwVN5C7N8DaHLNMvNWAoYm/ooKJnJWmBqx3g97Sf4H03HBKEGId
SPl42+GGbLEogEiUeyy2sPqgxYnJN4dK6spXSXmJoaTAASae3OeZtEMTBqXxpCQ4SZIYZBqn2lpt
rYnTvOnjwTfKzL7yIeH5KTRPqCqstBli/QmjYxLH8phrY/N/xHP6oE3Ae05u2LfHV1U+Gtyy4JCf
XjGPpW93ax1mzLi4qeJEczowR4GxsZwD0dxrytvltYyAYiS9PFlPumy/1oCn1ZnWedPWOpXEFVpw
E5jEAlh2PNikdARGJYGtfgMr3I/p41rDuVUCBWeBTlrBhlGHwIbDEI85zkcz9FpGdeYIoVvR8g5K
66v9F9M9NKWubosx2ddtiLN0+eiiSxhPt9Xa1S9Ox/8MGmDwjeTQeuQOueqlnP5NsYVJXjacIaXa
CKjw3gLFdy7lGyzzjbSM97R3bBKP39J155eIkE8SCwfdQkCeCexVogXrKGrJmIaKhedXmmwYV1vn
Q07cFkogmxvpBfzHsFRvvfuraWzML1cnChOaMw7yjUJ4V5SuDaHlGs6y79WXR0bE1PMYT+pueqz5
vNxCNsbP9nn1Cnk9+OCjIpeNR5SggzTascdYQkyJLMCXw6pcCQY7szhoaDzj+wkG5yqK48wIA4Bh
yFAM9P2sspladYIci5M3DzNwCd8+LOmY7rRIQ/Rwe0jytJxVuP5zE7PAle9o59sjuyrlc5y0acrW
9B+rtFjY6yR0OXtsQ/RIB4xtokFCoTDtuUKZuOcqFy42qtQAG2mFy592YQJzzumrMfaeJXkwm8W0
4JDlTJWk++tj+hCY7eeOTeUoJWTnzjo93WMwJfdOChEAw0SdxbDk1YRqv2KDezWaR9+oHRAgl8Qk
PBllGRnM1r/yeG+0nJVSgwxdNt/zkqWYVYWXOjqi9rByab/B/wLoLlV4y+/E/fxRJOR7INYblDKx
e9GCKtVgVfPQ85atbxUXWc8uX+izeNeYq56jjnzOAhImk9qfHGqUkeQ2OIiFrOyxXW5luy+AyYgX
MUWcbLzIvbvpSr1qT+hIPMF3HggmNzLeh+aVARAKUaVn13FpWCUdvpmrYZISFpBAtLe1rJ04QKM0
AtEok1Pg+vdLMCpMz78b2gTVahim8YCCZs+6zitm6DqbsTSaniOy93k+0GzH9izKGEUq4ruxSgwR
5AKT8Xqb+BU9rne3KkHo09JaEkBTTqHKo+RvyuVYYGDfOnPvIc3FOkRsBId1QInApTXy99G0fpaV
2BqqYc7zci8z75OZNy/Cg1NYHQ4N1hKY2p0u9r5+flFZUDn5Fuu12jyEcpRTVOYkMwO/TnUXGcsn
xTWCG+yTUpR60iZ2RM3vhHbWtVLYkuasqwaSsO4jshSSLZ2AqFjvdVLDD4JoSUP/2B/JWcbWiuFT
KwlS16iJCs1kMZHduMLk3BbT30x2VFzQDeIu7M3HLj0pzJ23AvbAMHKeHoV66p4Jfe7ERYcxFYt7
daPboIQTpf2h3w2VE74PH8aTEST0dHpsVJ31rYSr+MTG3uYrwbzTI2PZBYZAMoEaBAu/kGJhLIcb
HuDkn6JkQaLPqSxkUmlQ5w9VD6GDpuv8SEBu/mzEYX2A6ZEcUUKUOdq1o/m1L+I4wThY/KPPA/OU
L6+Q25iU5UMCVWp+yvIyq3F5NU7rz45VqIeeb/tVb+uKofklT3JdApcp61WneK9xN0qRdJdz6Sbb
n69XdPNQ6ZFRt41KMkqtgMybl7relbmQc6T4nGHnnbN50c4Far5VQz8lr+R5uGHlM1ouCm7JadeN
xKLUAV+U+jb6bVTyNvrv47M0oYQvOrLYEvhokMl+0UT9QvTJNfP+EFGZiL9/gy/Hbqz3W3ceHMBo
ftCocAJMVh5D65JXO9oTgnTmaejE8uP4YA1M7UacJBkqGIhOTEGtbw2i39i4+lyC19zEcWXzznn1
zwAYdh1uYbnOda3iMuUWZ7pCnQL+Zo3tm31lwnvXIMFRQpdKkJnTnfpEcX4WPTD8EyTtUcjLS22n
Ov2OuVhH3dn8QVs406u7GaybfZg+/e0TC7WUwqhm+1VqRM5LAda5fPg65YxRGHOTAZLB1jF+CL/O
LtKoGBdhMSyi4M3dYbex15tGp5qzca9R5YFxg+Kkee1B2sLzXDcIHeSJSayHNRmahVcEgeDF6kwM
QjRACW+nAvjyaDtA3N3btfgPbrPr/fzMXyyhYsi2aVH/tfvSEAYtjNkJastkWphyRVP9bzaed8ST
OL3oOPMcbmJo1+zxBOQ1QgHn+S4hhZHYfTh8ImCizoxF27KJbNT31SLm7MIBCJ1a+5Kza4++l+ua
dmKbLwnCKqUi9+WKTKgVWAZUlj9mH1j+QlSaTkqyzAeWHl/e9APNeXATf498gtt0Qpo1wOZl7rP8
vAU72mb9BKaknL3A6yc1dbZ9A6lcVCjqSY8LGx81B0eG9gFC8QMBLY3HaMHD7r3czyG+5hUqKUU2
cn0THlLYl/7Namm9/Zz6lKgat1H7BsLxe/HdEyaYp+JocCK1hMgQ7JjBCEufFZvuxCKzVASqomBc
xgbadcBgwAK/gRMhfKmU3RBrQlcWOCc7pbZ5XKfsjDk2C/oSDrR57LlGtnYUkNoRO6dyz3B5gUwD
DnwpAFB5kliUEeqdfKWtQzu3KZ3qzPEOLYi+SKavYIiaMfyY8AeHwR22OklNXhHZqFjegKz046Vp
KH89SfqK/5oSo4IBmNMNkuyCq+xrjeFtN3WGlQaHCFawVIUIyD3HNBXvuDHXiDQYRP4C9g7aNy7S
FTOG5dIcOEet+dHD51a52cyhtrgbRe6PW0bIHbF2tHlIPeWOHqrZ+39Ho8+GbqzwGWBTHTEwoxNt
JfM1hoymrxiLEnkwY8BI+/8WyWMjnqiyboXan1CzqACpxKZUelWZItIE3I1Pm1dpD9kjqKasllqE
gJZOdMoIUPIuYZM2HLYphuHY3rv90BsCGLiTi85HU3JAQYMiZn3ABjjSLGHGFcmZTU2rLJA4ynqX
hxg/SqAOoxD8l9JrVekx8LdXwTnTNIu8DD1JXJbHBOU+2QG8zRQclhZzRLu0nf8WCqxq7quFie8U
IwfLsdBo+rT+jSoBzAPDYc5IGSN1wk0qIdMTaBeDA+uk8yhbKqb0QPwNGW+vscCG9aCbupLfEQ3n
5u5MvBdS+/hn2hlRhFnMRLC7qzJA/sZomhXI/L7335/DuL1EVKQCMaYo1VrzoCliLTgEp95eMPNY
581EGtTZbPS7Ks9s1d6u3bqOM8/aPxpIr8ImpM9TqZCTYfMrUdOI2j9E9Sy1K9icYNpYy3hJpY5k
nKgIJFteC37na2PRP+BEzIyUQw4H8txMzvo2JSdy6aiIi0OYVa2gAUAbs9WTyTzCFwidRiYh9FgD
uMOTG0l7JT9yvGcpMIou0sAMOK8OG2OzZZdW56R/oQ5Rq6BX/JULQQbenpPk3G/5LLZ+TEhqW88Z
UdDb0KYH7Df789QPK7A7cPnSj1lRmcfCmyWYFC6L1VTgheDDeBrfmO20mnTgm2hZBD94o4h1+fjm
bkBmbIv6eq7/ZAIK6/9zFR1Dr8WAU9VCBscCYpZLTH6rvd4l/1f3fNE++Ws59EfBDQ07T9SRJmXh
h7eTwnWDl84mxCa6YlEG/GbkoFl9wXB++JS4HjkpVyLlDf5zUKzjpTtHEojkfut4VmhHVZGjqn7S
bjlaRa6+dElyC9bWa/OIXWxYXaTbJifG3TNoZMauiJNjdEjxkVnJCraJYFQSiAn0AMEFb7YB6nTm
q+uTPT7hzGeeXoTolarcMmk2lNHAJFxHUD6253xs1ufv8x2diyNg3NDpSLNFkTALVanGeDBu/ABP
6YgLcczeZ7GgxA+ILLkK2uEXQd2VoVNhCFKDpr5n7aYTP/RybeDUEbx/ZOZzO7PidaAbBAqhO7lb
ejlF/22ISZ5Qk1GfDI/QLXlf5rA4P5Tr7/wfSXiFmNBdPrZ+EGMcFWSeC03URsBkXmakqxT6PJRa
XNlGWqBR4cT1N1SpSs7pOvd43W/PqK07jOfrYx99cB1Zfd66dhupP1cWjmLgL5QFzL3YtN24Mh3B
Q20Mhkrt0nqfaiUgi4c3Onh5waJzJnfXoQbSnXUJVS97+lnGKHoxa16+SFt3QgUDdj6R8DnvSOU3
IanZdFZkdaQKx0NmFMEqNaTHFGNXVhlDBb3Az3iwLw10JdIBmxMuP4K2ZX41a+dkHpX2Ihq9YUaM
QHeACN3NMRTM/VhjMj8M0jqcG7FSv7eQA3aO7ZganV/Y0wC84ZjMIJYCbDBQZyFqEC8DfCXQAruq
GNIjg6Lk0b2nZiDj9ZI1OUHnsB4KS/Jl7jGL55JW02vVCuk4hpnIyBoR/AiBLOezyUgDIchBq71r
b4I1KUS7DE9uIbC7kDmCVgDAHb0jBZJqaNJnsWJvHVhq1T4Ce7RJmyne4MDjBV0TXgp0NHHCSwSR
UXKmm9VGCHv7vkBirrZqDSdfxomogoiwXr47lSfbBqan6ZCQStchtxEC2pBn/OIUclOgn8P2TdtD
JUd/+t8lSRLlGAD8w5o75mOmGw66QeYx+3+wIx/4Un1frnH7gBpjILbA4CKszCsg8EFj6FifyYXj
vT0uTjIsiqub2xODuILJl4kqnrt2QNQhey6YznnceDhxJb8uue161UowWTKxlav8EsuPNPIyQ3qJ
8zAlq/ZTN7Oh6mK0Jfh+dZiZZnqMnI3356IjXmVLLZjYrnu/TbFmxqpJ25sQ/2lvQfiusozmm44K
8DHOjUPiT6nYpxn9ElhEvl+yU8qcHnVrMYSCR8mO1ITIjdy192THgQ1b8JBNJjGhJaKRItSRT8Hy
NOmYSakTEEle5Eg2auxq630sS+cOTROJg3v8a+VSRGJGA9gkGFM+fjIXFrKjrGaKnIYuHWuVbq9d
f0mXGaQjMDzv3O+grJeH0gGO9AWQJAvtyCqvNsTA+9NKBWn3VcU8GCwm/if0UBRQd2+/8wWxlh94
mcNyT/bIPwzXxIlnrmVe/QaioSyYNdwxaIjE1ewPn6ULWchlPROz/42UoO04oVjBylN6/hJlmw0i
Ew9gyJtqBkhncZr6cTVNosY4c+jchFTSmRoS3VgUSyACMFNacY6LGyR7g1lhQSZU7ky7GwzjWpTx
jF2nlDof6ZQylDFQsQuDeCcQ4QNUuom2EoZg1H9S23vl5l3mQw3yFmVLgstZnecf9/95OM8TJb9d
QmEfTYchobHTxoblYPIXgu/rcSW3h5n/J/FcotKF8zEFqKu9KAHLNBHJs2ZuX/sBuoU2kqPorP3M
53iqHkk0/2F9O9ZxQtqM+QPK0nXoxZDmWlsCRLvNS9M3ERgQ4Gt8UzBtGkDHNacMWjxihpwy2BQK
5ZDqDgSFD1rTzc+dWYy2j3WCr8d/4vs5mKGFZu6ODVFj/BwhwrQmIJb7Ig6wKIWWZjWUQszalUCY
SaMzaSJITlrQ4cQRZnZWfJ4L+jHMpubUbqeAmoV9kavDJEhdUw9OvKQiT4nsH1/XUIPS3If73/Kj
na/wIta8QMOI6kAO5RLQYfwdbQykjg5iyDtBM0R9cG0hgU6h21MaAV8JZWwhF3ywgcOvd7pubDr6
6OsXzUgie0kCyMi+kPRm9yP2wDXb8uIJyXEIhgTK8qoOMX1ZdIHTIC6EU0HrUtfnLqcW1rNOMitS
WeMn5S9CGdSSvyOHxmiGFDaBol/HB+jeAQWGwSqC6wkyKzun2iOLKTeixSDPsCwHlJceyXzWev1+
/cDMVL+lDim2bYUz9DG10KbRLUWlYAMaLCEZkcFRtaL1kAGCGDmzW11zGyYbACvmxzFt0S86J71I
8qfgddQM/3IVtAo/W6bde7Gagvhr+rHwl9pXv/j7J54eHiXQTnUOVyMrEoatMTnaYSWV4eq7u2Pb
M9j4gY1mk6XNl63FQFxb6fdtq3ZBnaBmfpMDeWQfIX2aBQ+wv4AXAaRRjrCeRSjulPFoMl5/69MA
sSWuxTYCdmoQDAqNIyY84XbYWC5qGoG9NDt+2FGnNuxV0AdPWCdl73xfVvWORWahW2pV2aUH0nZZ
724VBjJDzWW4VQDmTnVgnNL2ZEM5i5PROi3rVC7AcwCCtY9nzAK/Kj2ZkFu8GKUYat5NJ8Ihvwyh
LcUDhl0IpLlEoeT7h1Mh+h37TiUkoIceTBcgcDH7h1w+unigOdX2mpzc8USrWZqziOeebQbkhumU
roay5CzZ0qUNThWbBETpjf4nAsO/RfLJ4cpVekwcBzPlmLeJBHPRXAMetkjUJ9BzM9N/hrqxQ0D5
1JFuK6pDdHsRl9AKn9T5p3nvm5Ug5TIrYTJxA6WtCk8LxiF0ryoybbxu0W2J7neoC6wYS6lR93hx
L2oGivZib++shZ/5o2QHYu25SOcK7Ytp9/WPjda5jBTX3A7vuyUKo8PNh58PF34WJeeBq9gOsBcD
7ocuclmRT4FPwux0iCrjz7N5Mvy3Ddlc9KEdxV5BjNBG35AMrZeJYf+MrRggQvcuKCf8AFbitg/V
flFr5NXskNspubHQhPVh/fi0R64HQIlycDTs3UI4H//vaDfPUAlZYYszHbgvzs6MqewrkO919CmY
HMC6BUwNNdNL5AZe3tsRc4QPWVrRUErh0ZrvsKQtxWUIVMFg+z4MN0O5AEAcMu+swhpgRoE/bMWz
bY3xjPh5W3kA+46tzC/xda2g8wfeRxBl84zKlAl4JGjS5zg0mJB2qqYtF8D8rNPn36cZawnjNdD4
cx5aZ2RpLr18y6Rvp8mdh2nFABQ/gPGXGffanbKiBknXzosA/EkfbTK3OkK3sDso93EKHfBHVZja
UiID/5q+nkO0tQACOsxNkYJ5t1w/gsSIQKPsEQCLkkRz4wdg7VbUPph6Aa3RvECllIvOOMcKTU7J
UugYnlx94jVqDIZpJ3l0Esmyr2U3QJfOkgGMQrdRdDcCKxEL9/NFQhpFafpUSD/F7dLUQ4y+xLPK
FXAJXCvXmgw+/6a5pnqELxhq0VO7toHLd+PU7jDXhMm6SvBMejfLhf7T81ffxJ3ZexuxbE2dPF6E
RIv7ErnbQn1McSnl0EG0u6SKV9E7Stp+eS2yQf2DWHju1PGASeAcEb4trFAHDkSgChnQaNBwxUMH
NMboEwjOWUbVx08efsZypNhiSmezE3lt3Koavx+OewsdwtJ8TgkVy8thgJxx2Z0ojSdval+LEQDV
3Jo6TfuIu+bROblRVWLfBKVgGT1b66u2/5pIQ/JUCQo3rPOf3eSlag4VO/Hta5qHDp5yxx1SOHgK
fInofD811GRLDQc797EMNwxFaBMiRDeIBq10meLQvxmVvsMU7tMHrnDkzbLCSL5TetLk5lKMWDk3
WY0emdpetDl3zxeSuUlWkbvK2pMTUVSNiV7crMwpfdGsUTZUt1kXAhZZQjU7Vjg1YwabsrKLtLqc
1696LjIhfLVnDHSu65sMN6KE0s4hAKdZz57t/SHplV89xGk774g0ZVCmKrgWfFx/92dcoPgkHPNI
+boY/2PVkCxvBJiGTWG0sLJMpnOKQrj+Wha6Blswze3AQI9PDpJXWO4/DhTzJIlxeSAhoqvVq1ah
4sOHreVT69EUOkd4s1u1lBSN/lKFcbLIm2bbKsU+dmiB+a14ykyA7visD3y50TTAqt9pQ+Mj7ALe
BcDygdmvgoUBoKZf/mUzzWbg+KydZQDdtlEktR8uDOJA515lgkdXkP2OvUWyazHf6YePes5Dd38A
/hHOD+w9ADHXmemb+QiNFVVplDxQ4LMLyZhjjUMJ0thIenvA+5Q8mD0Zxv+0l9cXeyZd5c+XqxdV
tJTIdcL4cEdW/fnOazZ/ThQvy2b6HdFTpq53UtS79uuf79tO9hGKn7PZEBNhd7UKiRfPKZDiH5av
Oaf0aL7ZmbsUScmGWtcVtDF2brwuyOk/78yihbcyiY2HMimEabI977g41RaroHE0p19tjf6MT2PK
moSDLYhBFpXzqtKdY0kSS57Gl3KfCedjt9GjyxONZjKt7NvrPtNUT4f2qks/GPtFcUtFDHKfgIj8
B0l6IuVGI5xFqce1ZonBD9/lDTKNjkxTDAufCQ6MLz5LAI8J1gk4wAVMQ8aI/rHWBtnA+Z0liwiB
sDwPJy5YeSZbqjUh1/9YaxDnU/VWQ4TRqBQNm8TqQRb1uoaDiRLMIQT4nqvsWDehm4ilv11S7oc9
L/vCCfUqHtKdJ88krj6cWyEulYx5CDCbo5La+QMCSwXu4aXox0ziOBkoVF0peylbRhUwLGHjdwOp
Rnr5xWqZNWXLCBcvsEklBfUwNie+bll1n7wo2/hCMysGMiuwG0ucFxO3k25SdOPxj7TtJ9JhzpRD
aS1FmUZgZpv8mKbnQg9t50UjzbgXpU5ydIgQP/jxxM29wIgdXqV+r4hQSf/nqGVk+jkNkh9rs1hS
i2DyC2mkC5EMT2NuW46xTSn9mQteX/YOkgj/4XIIV5F7uRXqvPBIqcu0fYkF7xa4Vts/zV+qsgio
BVxKtE0SneqHE5m8lj2cjzpXXf+Be9cUbSoY+C6lg5pD9OcQ9AbfHiWIxRPgivrO6MALZHs1Uv7F
PydXDHnRVImu93VITtdImPbasfnNaCaSKURXnNacCnqoZQc75YZ6JTptr2OvWsETdboxYq4W8Exj
sbFGz/kAZGgzUAFP3aJ9fjCcpLbr8ihGt7iXX0cqg3Xxyn/arIH/zQfx18VqUnjXBoiICHtYl0Hr
ZABjU3bSzIZb97UQqYIw9A2MakKmeo2bQbd8//j0c1L/+fndgWbf1/S8EsJbMlLFLpNmyHya0bgQ
ZgHS6g8ZiKwev/t9WyvWKXtstEc09P9piZk4OqdZkMm3lb9WZwTHWl1nUI+ETOYPvKTuxXZVVbm/
i3+wUSYpoiPDb5ErZworeBbKJAuDoR8N8x8bg8AdAkMdRWdNr13CKeSfQPQPj1K2aeOTu7H9/Zv4
fvA3lTWj5y3YxLiXoDEEspwy6T4SWeDI2oKdvTzEYkbVyBYMaNXWuyblc49qetsWqLuD1FGppZbU
PBXIF/sjD/hut/NzF9gSqp4mJACZ7s6MMugMaazzstamJf1/I+nwRppoUI/JApx5qfncUvW+pvO4
vWsOYfjJHA2/Hldh7Fh8kApAvJrUhMdkrgHndVrZf2OMDuVOb2Hzb9FNOX41rVseGxGclU2+J4uP
fVxU+kS5Yy8I3UiE2pK/ar5sw4CRk1qKkm4X5YuDL8wyr3uxblh/FGokutMcmhQcI5JVHvamLOyJ
3wHvcMczFZMNGngVjH5xgpRZ4KIaxEE31Caw4c6lEBMDLYtcJVleqgdDBA5gANERJisDq9A3p7m+
rK4Dt+b/q0TU1SgJTeY6FvX52tCpx9W5aHpsIK2VuntiQpTLRdPj54OVCDLUoaxje0gEejDNa/gi
HGS7w2qQk8psg5RGO+ZVEEv0FG6gk8sv3RnKWkmUvToEU3kbU4uKayZ0pwayPZP0aQxbdhO7nMiM
okStoFI24AiIbRlYyV06FTrIvBPz3cYTlvnPjWHVFqlsZw9hqqRk7nYgOGUwDLWgUS4Znzy4kpYu
btY8MHHsPEy+8k4WFTDS3bEoM/va3RNy8s0kYb+pfZmTP7KtlJe2GeuHJwlvH3dXvVZhTdAhsyqQ
Y/L5jbafVjuvD68Z9qqqr+AuA6qBShtIdaVsdcC48VoWf0Zwjz4e7FozPP9pkUuhTmrTSly/IcL6
ny8HJx60s9jDO16U+aS9cB4ZCssLjO+6BfaRI71K9nqu3sLI68hGF3suhEzsFuZ1Y+kXnqyawa/X
vUFtY82nuiSUI1msOej3+Y/Q9rUtCnFfKPwc1PQUWY/HU7c0as6yVg9+uPDXqrWb2oH//2h8clki
t8+0kTCjja9AsiLo+MIoLc3Nvp6RRZwUniXL8ggcSuJM8cqrUGZN7VpOji7d5LlH1myCkTy6p9G3
f8jfRS0r+toiFBcMRJ8/Facugc/bkZc2gMzvNFkswE9VE1M8/i7e5C8jUjI6g7kRJhQGwvJ61Zk+
rri6Tq80l3+1N4nBtkkV1Ex2X/N/eZf2W3JgeNA63G8vz7c8luVNiMgUwcDTEY8iVCrhZroPolA6
//syNHzUQ6uWSUuBnqeOIoJ4xYD5/iQECTjYUibLj2nhfzlTK+aeOZkn+khyWgOhxHMC0OjGSupo
dwOBOhSqsA5Cti2MHfg1UhsQdgO4TEYyeFQGrVbKXrx8U2tZYb3dlj85pmX15h5TDGw0CVhFbUas
VMLInp6oHoYsxi9IsxHZGi5vI/1qIOD2df+1CKYq+GrBdVE913UEQ8twfIUaEYmhIf6nBiZLhHHw
x1Js4oQZhmEGwCogAeqhjAUHPxKozjfUKirmuAC1v6yuh1GU0aAm9W0l7jTT0Ngjjn5jVhABCCBN
e6Z5ashKazVn8sw+PRhy1OYSNGbecOJ9A2WuUa1ZaJPl5gz+gEO3IjI/yCSfeG6wudlzfk+28Yrf
MksNTZUDieGtD0egK5BKxkxz9gCD4Kk8a/+jTIf+z3jskWvhxHSZYjgY997AUX59f0/e8M8f6YCn
rFol/eIo3gXG8XB2lihsVi5SfRdRxqPPDrStlrRrmsnmbmh6gG7HTOBqau+of3KYyKLG8x/VEbnh
lJxZ3hZo9qb1NKX3Im4WoaSj2uEfV5qFeez3Rji9pk16W7Afps5FV47Pur6+BbrQZ2JXwye97pXT
Dk76jgX4c0n7fkf4lxVFAVXEXkV6bpkrShpqN/tzfk3srxMIdQC7PA7NbmaxAQ6HQ8p1YGDlwICa
0zgc2KNnfwff39dttl+4C81LSO3Rq/qunnrXZpQeprlgPOkBtinINeuWK4xj3xWVkWguQyKcX7UD
d5Z/bUBA2nhcHY5l6j7zL1mJ5tvCtzgl8TpuXGTnfGGFBfEZHYySTnnM8mlg+BAHdqT/3dlaIMbR
CT/VWLKUVjztXmsgQG7j//UoM9KfgXM1NXq837vHBp3ttqeHPHaNWfHIRSksrPTe33S6xCMP3duz
aJvtZIh8A3bb0U4yej32Ec1Gyexq7ueK0DcBdINoDytr9BOa6+Un8X8pEl0M954Z9523FWMp9mOd
h2f8S9nPbZUUwLEjnjQKMNNeMXygw4adjAVxvmNyQrJVHsDqiFLcKe2P8QyEfkJMhVG85u5ZUDKj
hDOHM6/QrcktwNzwJXa6ak0KR2DZt5WNiucF7QvSpzsDma7DUxCtMdmfAngJvE0v8ASkS9Gs9nxL
WRtHejqtKhVoJquZf6j07HlPGWwKxFxgTq0OGlL5qMpF4G7T0zL/WoKKtMsfRvoW3neY/tWqiZgA
oZSOGETYNTuW31XazBc11efWX/jqj6cyqLLrNMwUNpI23hGJN/EKY7c5o69tqnWTsk4NaY00KfC9
i1q2NLNXEwxS1oCAAhu5lXLAFHHZKc1vnEP3CyVCARqr9xDpNHsr9nXUES6Uooh0uUjZosS3gajq
90e+hZHNCrNX+Cm4Jh2hbR/dyIsOUQsI+w5ll0y/dAKShvW1ErwrV8iUwEPtIv91x9tRCGv5k3IT
OJK547VARO+oq5i6UNUcK5ccSva+fviZP4hTuT07C/MT8s90thC9cX7AIMncYb2QTampsfBU8cdH
+czrCm+jIVvE6SIzvLmVtyyRxWabVEVP0bp+mCskbkt9bk3hMxLcw6Igew8qkW38CozTTc7JFf7c
w91EgpfLG/Y2HuJjDDG7tLKs0ljQs+FnQf16YoWvJOFz4iVKg4dF2qasGVRYguyfX7HZa1HViDbG
OB09tYMRKlivDwr86Gat8LZo1uiFT5TZMCqkk8cHsLf1H+D9vc8mvlRt5sxfnEafF49UGjl3a07B
Dtq5/Lz3I7RYp00d4OShNaOxznE37kMY/rQyp8Xp8ct9wndMkxyS6+YLLMIKlRSPe+SY9tPFy7tY
4oFeB7kGRZYiUjby5b7XLWwK3Du+VBONlaXCfOEYKXB1+8t2S6pbRNt8/HKNoJojgABetdf+l9bv
ZyxvHeAPJIejwAJ1ofoVLVGL2h4F/maF2pS2tqIWferOKFZJjbMBzxAfALdF3Ev3YlwB4RfnlDm8
M8zGG9AOv7JJ3mw4gIg7WwUZy4foxHDSfPcmaA5+1syp+iaxuGGEoW87gXqxrNBC/5/TKAy/7pkU
A/wxMucti647I652NGbdSCVTt2kWsHGNRpxUf40WoM1VLKiBBAZvmuMaFA6SBFZ8EOgm7Y3Y2bOI
ddxmTzXMpDEyUVfB/8C2iw81L4vJLy+QiXkjKmvzFTRHBJvM+nfXXYLlvsx8AvFOG2KrJYlWjkoQ
6AUUSgO8OWxSkQ931OEQmtoiDrsQ2s9FEAImL7AjHk/KLjCe8c8nv9uRThzQpc8IbLU03MGPNv7v
szcNBeAAvwIMtfyUk8K4/mFwH9pDywXZMUCxtCvI9dZk8t0y29gPgUx480ffWV4j1pZDF7iV4xoM
yTmhYSeGb6lTed80eRPuWH/oa5xyDeGQRGs7hqhzLDnosUoxa4VpmX3eFn5eSeTWxlKyZpBawZtk
s62veJAiB5RXHsz1sglwqg0uqnzmR1a3QUCBO7Eet3odjp6zXAXHZuhkbohug2fAMhWF1FqchZEo
cqeMT90EQ9AwIPvOKxUUbU5HFvnvDkXHuwsoVXX5ZTGsSmdIsHpntEmk0JdgIrYh8zwaBJwwDq5M
4cnErAA/e/AFZJ79gYd/m+AlPAuKEBYVdTJ5leRyctTOaXgcjOVQKSkBLoy2xRa94ajaL9CwVqXL
+gcXSmCfEPh0TmWr
`pragma protect end_protected
