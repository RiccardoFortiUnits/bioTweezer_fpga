`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RP+1Hi1ssKCrBN4Ygz1VsEPDoEcZr1klVUfsqvbuc5RTfvklO5JZ+n1lykNRPfBg
RBrUH4vnj4aJJdEx0mo4kOJWgTk7lgI9YkKbmbS/Kbr33mRqvJVDaypeB1rvCS4Z
7rNnUnoJk3duo41kt/0nmig57pziX/mB64KSJ3i2ojM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57744)
AtV5078eUTbG1NvIx8gaRalqauycawvep6BYIt0ITXhrD5TVhTVFOeudqcCKsjj0
KblPlenqIwbFsJElsvJInqukteq/E0+8w8kEDIF8yUGRCy30LVCTG0LJ5NLgxxfq
yrYYpq3Xl2dZtneCYs1BsUAdbPDEYC0qk7F+C4HI7/2F2UsjlxMBvyBLgK4dFMVB
Olai6zZaR6mXaLAucdK/WkJOPqUrLnxtqy/RofKYozgnuDvaWX1DAk3gCQGj8fZC
JJLC0Z2ZKYs6OrPxh1upRi0Rh068NQNuc99Z4ZzzditY4x/duVtqLNiYZsgY5c0s
K0VidEVqW7zlYxArF2iimM8UIjQAcH3kwOQmLo3ijUX/YtdrlhJCibSQv19/JR/y
ZqyWi4gW0HWzVbF2ktR/bwy4vZf6thPGhHhlLRyu+ZU0rqwnZ7Y8sPXUy0NT9jtm
2sOuicD+LWcrgwi5IconQ//KWaCjNVRFgToNo1Dq2xFhDZ2WghHu1TfW5qZpQ6gd
vqwXTIKOdBUyO4wXP7G3TOrjpzfrzScexaUKQIYKJhub+LEbxm07DjqdbJM5wRYV
9UcXNdT8Il9AwITOxok5GxFYSn/vaI5y9PdbUIhn3Lm8untXH+tRw4N+OKvWunOA
fd4XCdWUseMZ214NBXQsPMVC/XOr9uQH7OomBZwkY9anARGNFAWin/+NwNAzVM3Q
STfjKoBhV/pvmYFJB7GFv2V2aLjTjfv0gj5wAABhfrrRbWTR1V3NZvqxEO8P/06x
4Gy3fHrgw/fqalvw8v7jafuiluB29CJ75rLwnPZvp2JCcgWdyOr0Y+MV2A0VEM+e
tKl0Fp6oHbZdU6jfRYUHgg1vSfKVFS1RUqwq4+GMeR06Vb1eGycdrozu353ef2TD
Ezqpd/IqEzH3TOiLMwowOjONtEVAUE92g+XmolQlBNeC1t0OWwn2kYTEWG9WHHHd
M8jvqG/khWng+3FBy8wMeCnaRriMRSN8rkOp3FfwrOsm/iS47TR1fJWziMa+Ix1Q
LVV5GJYgqVoZRu0VoKabVQHPsh5quQNOq2Jk9vb44SW4f4m7GkF2GLJfw9XoGjuZ
YHAxjzBxjoTVLzEFQtUtY3iwjHo4z96BJdiesZ/fJr53/y/hwLkrTLCbkWBUT6bl
HW/Y15kcF9s9SvvyU8So/bqwlM7knfcI5M+E/QAv71qmWjsLG/jXiXixgJfqdHhH
Y6coaZPKqoT0Qy6xZ7z+BT+Qyoyu5EK3QvSP5ueSsatgo3XAnuwnqhBCZJFXoLzZ
ZZutXxmMdhGKqbBhnefKfFsRYEridB946a/d/GVesnJU177MnCRHA76iyqPJUgcJ
PRVYpsqQNANjElnxPkCRMGX5gFVpdfXpbcT+3KVVj7xH/4XJ2W0V0Oy/3AjJ1g5g
h2vqUevQkNJW3nsX0oZGy+fBRfZL6vYhaaNB7PPmYNR391emj6mgwMGsDyERQ/UB
L6e4hst2V0WU/UDHLSAYNA93FS3V1Om8DRv5GgTYkJYNNSLJ1jt5gjUQ1KNmc9rs
USrkluKJ0rf422t9jpwbz1y9I+7iMr+x6SOH3YKF6gBUYhthEpFmNyPIfIY4+ETM
1T+FADoXqX2Avov3pG1u9PG7IbSYaYygjIMPQTL4EVmniDLjg1Wc6l0fAifjMYF5
6DEPh3MFlo1V/0B9/B91SrxneR/XgthP8nAbsYnYDwlT90OfD30RRV/EPtmU1oXv
PxLflgpRMApEhSMIBXXLrKi9toGA/oKhImX33SkMU4SNWupvfsm3H9A4BePct3xO
v5bJGFDWYIf6cP5f/5RMHs4L/nNP4cl8NiMI01w//3W4a2xoHm77Nmxk3QNOYtuZ
YMNii6/tu80oBg7YaHE/onsSHH1bpHa7lIpI26e3lhPjiM2klOify8vdET/ahUol
899511Xe1/u13P9cQv/djYK7G/2psPlMy/UmQuV1ocaEcTHjCW45eYDaUOtsJDZa
Gh6fUAS+NhjY862mDVbS6S9HTzxTQgiIANyqXBteVl9dPFFSHM5y+obLvKnMiwnX
0l6pfLUuv3OXe5hkDVcLX7yj1SU9yYql7ol/hCgmmgm3h9Nyo/XSsDC7SsiIgLvE
dZORJuxsHTfh/C1rc04LkvrAjg2hKK88feulqjcJ3ZGPPue5HUFRq532iCoHUD1X
OjfRlcVhhUfhv0Z/os5EK3zIsHI8j3iPqIdHES5Aeb5e5vH1bjZ6ots5h8/ImKq9
1bT11jO9hB6AZzIyxmDpg1QyVrpa7o7LDYug7spbXqPiJYuDbnZo1ysLCDd5cHDq
Mujh08b0ruqs4MeVPsFy3ECCCMBJZeyoVdZ6b654feQbnn5+qM1jU1bf6YFXKVvo
Wn2Zv9nGfO0fDzZKiTR7CWTE42DLUKpy7Nv9se/WnfPPPHmEerSi4szF/uzYI5E3
K5fkQxTa1Ay6VEuaFHkT8XCa9clQzwPonU/zGsX1wjAh+Ze8KMTsdnowPSxTFy8U
tdyqeauVqMDmmLUbfHPkVnbyys2QBLMXBRvhvWVKn4HNq2W6Q+x++21MX3jAWoA3
zcQuPMhx12gz2i/SUdNBb2q2ELKnfihgyhhFftQwR/XOQ/bUc+Zussjlapq1dFvn
LDwWQx+aSD4VrUSLqU/WxzpB0yKCJy5kM6HwZo54+GXDrBtNS41eAhaVfWDlCV7P
V5P3ISR79EBQLnzLwaQqZQU011E3ViAyilZ+xDJEnqr07hUmXIuxFqtHiekbi/aG
SvSSl+mvhA5XTSPvJfog0NUTzior8dt6kcmoRKX3UPBq64GzsMBR8vysd8c4AKlY
d253Yx18O/lNS5j57lkM47xANBxEJEvVl6StM56b/3+7ycWpYgI9769+ReQXYr02
EUZrH74h5b/1fiOcVWuyUTzjj7qzaNPSvjrNmpJprtQrjaFUL+y14noWk2Ogpr+t
c/d8wLYiw79MwQlTHaxNRONxMrJj/8Nfn3S5u+uZPAchJe/UKEcqDDnYlVdmYSoL
4WG5DC035cWXfZPO67xwhOGU1yhN/THJo4XYGJ+ItKkyBNSJ/pBod7hod6ucunEN
+Eo+5A/WU2RCqpaUonck7NTCSqndpCSfdUEJgxtDZfTUQ7xmxSUZ9DhTmwF+lfg6
lFUxL8yGw730c/YZJdhLbIH6PK9KJimrf0KRBF/I9fmu1Ba6cZlgDGtBZFmodt9+
sj9k3OcqmRMakXNbuLFZQO113gGGq799X+Tvvlo3Uxar7XzIa+0I+EWjQtgLqON5
6OOTdNSp+/0+akyIVey8OxK8EtTzwFlvWiUuSamHLwM3qggL1XftODYHMmsm+B1j
bChCDPjjlTnH0GNrvIr8uVEvp/HeRy6KkMlqxvPddOaVYh8ReXwbxFmJNu2mT4Xv
o2R1d1u2i2Pei2sUdof4DWKgIFQj0NpiC+bR9wo2/S9kQUg3GUlUOZMcrvRd+Xcl
/X4EfcF4Dt+v/E06msrwxdD66+jHj37UgrBpNZdpvrHoclhYpmB7gPT6IG4kzjSZ
GavWkTWTweo4V/bvCsujQvxeBdgn7i0X1O5UC2x29FGig745Qwnyd7cDQz82krEv
Phve/nrZIVgPOqaJ6PdG7tpR6Td/fu8U+lpOKZtA0+WqrzsMjKDBh6btkgWkvf3M
7h1al/RfiF30NwmtSClPUNaQLsWKE5XV94S3qEw5Wg+ZV7v3Pum1JGvRbrwUiq9D
bHQpDHk32Kpj+dXUIpfeefDwWnyfjDBY5hWbxz5XczgzVUc2ioQavQsydxPegCrI
g4tlrcSG6PSEc0ds+Rl4L1gLrjIooTJ3HL+CLVLNUc3oZhxeuq1uNnDwQPcQS24b
BkJZ36fcerhGE+fOE7iJPbAom8py97t/pm/gTatnuicz8m0Mo3Ao+Ea+rzgBaWaa
0C1rYNd5fgDlKtgW2uIFe9wLf96s3V6QvJfk0GF88n7O/Mic5g88XLKgxn1xBFwW
3Zh0+NPIkfTMyz/z9UvzqYHjpCGULSHdfahMvcVPWjPMz1NDSJaDxkN6dLkqZTOm
2QjidYFkwocurcEzqksVwqDTcOeQZrB0S1BwSyrbVlqQQItmGf9YMArncS3RIME6
u/b52gTjJbT2CO4sm893wWJvF/cuqha79WaR+VNzFlJc25Uvhc2OeV3q21CYj/QI
OwsswOPGaKSnXs7HBqRUgUgGVyru8N5Ebtbp8VvVFU4CzYt+0oo1wOB8wY3GiavP
M7MGRSxJS77hdovKdPm7pbxRpR/X6E6CPwBdPtUwOOZAmPRZb+Mn/PVOJZFqwI8e
an4Aby70mrogz4AaEkcrMbTp8ed7Kfn53XOVdRDWRnTr2pBfPgepQg1S/WmyZqz5
YJ3mrsxLOicY9bntZlEThTTuKvwBV4Hlkg2Ei/YtHjcbDOiLSYvY4stO1djguyAb
E/Yu6kFmfi7jURRy+vGnisVDSnnDKwbHKRpmkF2XA90IXQpFGNQFQ6uaDU9tchOH
T0W2rdlZhVJjjKy8V5VL0EoK76B1Fq8yovkp5iVvrHhSznxNwQpXVXPneZ6ZBBzf
zLlrHfd6kqwWwui9r8dNIIP+1De0CMoGDG6xmE59LQaT/1fxCBO7EvrCyVaxqdGr
o+6BDvvtQId0BCQwZqWBCjVFqUEuHQn9ujw5sTpZGUfmKAPA8ZGylbFyitUUc7OC
Dcw0zmpVL+DbOOQTfSUX5uxMgfTH2xJxL8Gik2Tj7x5kHnJ6lQdtJpLmq0Nkd8XE
kCzwR7o9AxgwhGCWrS5rHY0RPxRV7jy7wcXV22XGxV7gCLxuX4ABAK1CzXo0intv
DDzp4OyApsVdfiEsK9FfURwmSp4LKvFV2xHUKGGOCpsqaP2ofkoz7pHNvfuNlZ+P
xOR61NUHaPz4/9RShx5zHvJTuRtYEKT4aDDLEH4jiK/kkwdKnltVQeZAGurVvTlg
VQWu7UmKnrkZP6XgBwn0bDqFFky6LzIRWJt9QzFrg0JzdHgmG6xWrodSyjRCHmYY
5qRosyXVW2tXTEv74+8wN3ZUtWkztKI5wyvt5ni1w0RLDC/BQUyShhyD0LEVDOUF
GfR4w/9x36KoJdhS1P4dhg/YbHMpBVZY69ibeY68z/jo2LMr/rzjPLF7gIdbMGtS
XanZ/3DiMIVEaT2HDQnSHYu7axT9Rb/PZ6xmxPDqIQIPjWQ4FbGQQd5ZKfO/7j3b
KnYJTKKPhQDFQQiC6JFw+EfTExaWa7xRS8QMcQOU8XJTaeO7/FOY2ji+rcB5FFiA
dHOOI/EpcyQg/Iktp+7ugihEG0S3rd/5iPdlidEXqJ+Y0xt1IaasMi7nxrkuNb6o
9uhVEZ7CeKUgj7UljYjRefXfKdAwj/f63OTe/3g2IOHpyUFJZTIiNZU2CGhGC04N
PXMwbDZ+iXUfTyKBxrS3aphI/vpydYGp+2xN3NSRnp/OYHYVV/piAWrqliu8WYTt
qEAMHoYjnmkDVuJXYZM2TaiOKqi3j2wXGSDOfyX/3rxGeNhmeu6Oe/f/qNsLEg3s
ec2Z6P05v3O0PUB9EBR7TP/R9eAqrfEaCNN8k+DqUpZslqbnTbj6phx2AsSO4UHo
71cMtNuKWZzO4jD+dSwLzPfyDcvlo5IM86Ud4c63uwcAFS3uEXuJdG1bLBmEJtHD
lxcGElu5d1Ag3DUzzEW+GY4OyCHUeYSCnI/0ahF6SS56uU0McCJMxJHsI2KstTkm
I7vVT2KlQ+ShcBJ3HCV7RcZkPUKcbkb6jrxJtDLte2qlxkQjYA87GgHFBqNV7HjW
1AP1zGp/o5+9Fgqmj+MgIhFDk6Tvrl5xJ918a99E6qXn3P+Or2/9JT+B6WaTUu3+
Bx+i+1Y0d/7PbofMigbweRox7hrNKhGysnGL6xB1uGHhVENu9jfHPXxDV4Ibs288
NZDvaMSYx/TyxTlkc3gwzR+LmDY2EwU9ErtZFZxYW4K8Wyz80aQq3vXjqq++VN9r
sr4ZTgcMbtdrehr6orpR6mBcCDV7Y/uupVt4ZS6GpFPJz2V7A1RmzFVfd+pz51LS
Rh7rblSNY1ugfJ1ndTe+EVFmUWlLdfVD3AakebgLG5Y54AT5Sq9B9Dh4gTwYYg0i
9Dw8MK9xTCtA26sAMhmdhjjpUrO+qmst6biq8BJkl4cmeto/j3zY7J754KAHkaIq
Cbzs8apkA8e6jC+nAVc8RqdnQh9Ynq9GhPMSa/O//9ECXQQ6BnNN4ZnTXqPo9i3Z
mu8HzafndEHWbp6nIYSmCKsVZB8ZMv2ERkk11/+3MGytoHDNAnk6qer4RkxoZyQZ
C6wVhVhkRqsR5SviZZb3akYhYmAAPn+vmKw5eMXRMpTGmMixOwyrOP9lw4kQfI5p
kj0Exbk7Hm7P+GHZWA/KTWOe94fIbqi4XXmYU1AFqBmb+iAZgQ6nw25GZoztH+R4
4zZ+5km6Gt/bl7KO2zlysLBMZ/h6s2BD3RddGINe239/U7fipl3wY5SqlJkpOvij
7Y/8mCP7LHIW7+1ieJESPXLep5CiYGaQjy/xFbwGfbz0hnT4/GOaLXKb5aOfEA5n
nlsktQS5nYorJrvraHyzOx3PbUrTlQKldsiV2jXwqWuhvpADqd+TPwn9QFi0cVp1
kvg9a6piRil9pDPBQfY9LS/0CEpAGcd6olo8BMSiTX9u45y9J4Kvir0Ah8NQnkNI
s/D/9XhvLkNfkjxxqSprUYouyt4Rm4RSVtaI+kMcIiw1VIUGFzSFmYu5PF/9KVZh
BWZBOH7xUhAp/8ZNIziUFGgRMUIzviqPiTQ+QVJHjtTpkacc/ooZ7obFIr0qr6z3
LDhc85f3QPEzi7MeuGCMTHoLRbiR3/v7MCg5Jdkx18/yiUCOcoUNN90nxkVYp36q
DnhOmO2DxYbMGJk3zNri24IxkyFL/o4XKoCIsncKSBRB1GLEfCkLDgQFsDqsjjF7
bb5/OB40UD9rHxaNUAyfyihTnHMzQyVdb78IDgHHTs7NkfPotvJQnQFqxWNS4x2B
GAsv9vTICj9wO8a5b5u8LCPcCpzvpEJSdx8CcodkAj54Sfo02OlW6x84DVDEdzgg
/EOFD/W8JxBMJ0KqyVqc6IgTRe2xk+1HLR1xzrE0mU4XMNRlNIOneH6zLVjX+gCI
zmZikpjzhdhnCKcC1MgiHmiIR2iUkmbTZKb6qHUAWqVMka9tJOuvxLiPtozvdHTS
sJR4L99mXzHQq8las4J8SJ6thWjsi9EnetALHRkAZRfMkg7NZYXJCoMiwvgMF3Q7
qSn/bETZ6A43BpptOhqVKbnzX/L0etuoFC7x6bi0mKFdw2dUOtFWdBQC0yQqWhiF
ii7Goa5nY4I2mJCNF97AIM7ckbYZ5IMoImzsUl79roQfUbx9jXSbPb825js3xKCA
88BfH7K8fshMKpwGJDDBNaFHYJ7kkoQDmfqklrGSNlJsn1bdNiTvVlvdEOCF0Z/K
z21qbXkaE41oUDfIuq0S4/Gse4oFVhS79T66Wg9DgAHM9nPNtcoO40grOdVTmYAt
L8KZoqUR85rt1S8EuyyHx+0sA1QGLtFxl2GV7QUb8QqSGnNc1BhuLI8JzBCzlDMI
NkqwhhFr/tN4TeenVq25XPG7gCFK79Pp1etKJR9oVjDfgiUSMBD0Rq3nETKpfuw7
yxBly4pYuC12igVMrQlU8pgJvZJV4fqT3JXi2UiO2GO72xNzwSa/ZR2MYdYKmFMr
fPtRfQ9mdX+wDm6Md/dmQ0H0mUjtBZStSnYXgJkUUxQaBQpLIom25/zjeF/gjmKv
QrEBu9c8fCbO1INBzU5+AUqDfsHW/KnfS/wQKAK0rcPAaBhU1pby5Xd6se9m81kT
iYOeKa42vUjSLY6qhBigGuvJJwLHMWV5YjCEUbUKDbPw5925pATSchKhmQOAee3o
37Ggkdr+G+NPxEEs7x/KUM5agN+KMMtQSVvBV951ocaKmP2yxgVml2DNitCQejhE
60mjq3UYYySwUx0aFLFRlZyprvgbBNiAErtb2W7QyDBVwB5guO85KV+i+z78MsO9
PDjxcc1RIjlHKZ6/sSxrwSFplAbnYfSxj9bxorzvwtoygyAW7xphScTlFw2uSVR5
DdPRvOHqUhqb5H+9C3wKM3b+I8RCBkc3x2jYfN2tWQf4cQKH6bV1YAhgGDiWZBjH
XAOfmtM600/oYhhSEIOYWG5fTN8QjbBg7A3oXjdLgvZLR3Hd1yijllih2LEg4NGm
NdXeSDSq5BPgO1kAtGhg96UNC19VdFmeZfv6QZ1zfhtEyKbHWLDQ29Kr83Gyx7GE
QMxxh5K9RvfR1M50imQoJICl73Dp/1zybOH7ipKsLXS+o0SFRojr+DQZxK78Ys7g
Hyheaj9EIqTBWlUyyHSSj9X4QFu1iPTTovDd4XRNEConrew8dXpf3koqKqPFxJHz
GiZ/+tQopZRz5YphVnriFFJtNWRHcAb8fafR3pkzpcctQk3j2ufFykdc2upFQe1a
l48j/Yw2+wwroil6r0uUHihwJpyF+xIwgfnBkDgrTs8dnMhvA/GOIccb+6eWruJb
AqPHT71LQFgy6dmzh4Gr+hNCP7366sXoHqfnLLQtRtF8GwsaCYcdmS6qbgc02csw
gWQABOP1kzwNqhL7PRrciU10DH6tfP/EOXaEF51YyxwoOff/3q6U2EVD0Bu4EW8H
239daQb/C5M6UOCMNAyNO2MW6L0K46nZhzVLL6ghR3zmjA7AzQgu0LC/EMVMXxQV
vRRowHbDBqIHRL/928zVLY8iI89mKcvU13wXLKAK5/pGmeBATXUtjNGNes6kcYjl
nhqoLsreIZCe+6aeeAugW9/HJIyazSqwieHQyga4eIhltCD199gLRVQ7tZ7eY3Da
GBgSUS2cVz0V5Q+Mb7ebDSFhkQvGZtJNM1CUUdJ+QC5/YL+ARLPVDnB5BYKoURGd
BsEEF1cClKHkX8rD/ImB9ARoWaEwNuRAO8zkQYyaeaFbVnRytnVQ95PBaceP1Q81
tkOHxiQFNFG+8wACVgNh7STR2JGyEDfOuhm+D+VtzZqm22qxDmjVpFPFnjQpDmPB
DqTdMfES6NoJG0MfqoAGCVA38/AzuJ/SSz6qBErdoeN/DyfE49JPq+wbRtWBHNmm
z9ZINNmLHkZbPY4/8uXISvoS3ZpcLYDI3VYKVKpmQiyG88kAiAAnP/bkdw54CYx4
2Ox3uJAuTGfcRam0lEHtJqqlI5U6Tb7c2QGmq2nrNC0IsULvqfa5i8Wq5J6do7GB
Qb6uxm3nTjVzgfWa+K9S8nyNsLBxqstvpWB6DbAObdYGzEGDEYbsmQBXxnCA2TXt
UCT3rNlpuFn6IPJcvrkcQw8gFKxQfghwG090FEiX5TQx9voee/8In+RhxdACTarS
YBTJuBz6W7JwK9boPaIgEPLX9Sf9y4LcYnWLoWY364KPwGDPyzu6LC6YHI5dxIkj
XBg9bPAyqz9oGsSh7209ywy0GArkEYje5yqNyaDWSze5/Qw5NXRL9ddht0nz9ASL
lxoS1WIEyAiklW1cpBS9c8j9Xv/O2UlR9RKxxYZPxCX6K6vkdMswW8Ow4TyHQczV
/NkXMdVLoA6sHeivdBO/euGZkJUpZYYFr3tSC7L6Fjw+ESK0Z9fNQgpIVdBUH1qj
ZdnA5j845mmW3c/cP2mBAQ3DUIi/iTW0WLHFzy0FWp72XA2HDZNtD5olG0MOT/kP
CKhJGawgF3UFtOPES5tFkv9eZrhlmswCqoszrJejG4rb5u82ejrplOP+A30PrV1F
VkQug3vuB5bF0AF5UhICm+dm9/XQOZl/9xZEgRi9XScPOq17u+U5g+63rtlHaHAA
FGNKgrhwLsR6AglT0sc5zQ4w5YxE5Bsm4JfwrhSzGWOKmvwPpdoCwZXRG8pA5kgd
784kZbXFKxgIbtvsrwKz+eLogWCRYpyK8nFw9aYuwFdIhjX749N82Y8fYtEoSF0Q
D+5u695CGyd62Tu6IPyM6LhQrtpdneAtMyE0eBT9j13QZ5E5RscI0WVq7/2wMnWc
T/md/ybhg2WY73Lk/G/ed4eLaAmoH7OqY89eoznHdUQdcLxim1gAqv9lAFZLGb2U
eOnJn349voI1fkRKmrd1TP2ejvuD9FbBqzZZYmGmiXJnct7RpIRXVlzXccjyy9FE
o3RL8/sxvvGSBdgi4tklrqXCkHsnqYbyQ6PvYYpjU3iBLzxSR7YGARWVJbFXyiaw
+cHixSzbBbgORmlCeGCH1akzgu3R7Poi3cL345FrT6NBbHyyJsxH5dazRGKlDaYA
fvXgWl4WwT/FOWMe/h5kYLmY8kOk5VxDFphhgUUwSp0MS0y3s9V6XtGkTCnBiycy
atV2qf8UuYI8q4oMhkYk2UmNJm9rM67q/TecTrrnm/IaUcKPFNP6WimkZ4s3k8CS
517HykIgm7BvbmHlQn6jmfVn5LPViZLu98JOiCaKlUXz72KL2EjWXaD+uI6uOcyl
gZsKA1UyFue42U8MyAHAv3HDW37B20wZzAUNGJFEfbFoX9tZfgmqoKX8qeD5ChX3
T+3DEW+Rq4yzLskP7DlJew6+7GbgUCxcXKbUc06X7qvvmV7/ji9nm+75ODV8yFZA
zKz+pelm9pM6oGQYjtK4jcros5W+Mj9ePbT28e7Vm3O2SpqMLLqMxpVewUYS4193
ErGHa4JFNNyiUPMCRi9dumw6YsL6Vp218LI5nOPNpdnyNKAgb6uWzyQ4VPCoA9sL
b+QV9h9rhYYhwCViG3dIPiYmZ2ZwTGm/0xp/42f2PQtOzogaGHiI8SL8+IpQFyOD
gDMsoe2YRGUV6hktHNofDMFG0azxsfGmm17ZEZuqhJ52/O2gaKmKUfhn7B6uuK7u
9gunQBdiapPnThNcv01Q5Gxdy/agYbjjgXV/UgfOFXPTpaj9RLwXv07fMZTRQ4Ti
MQjw+tsJZnNBeJTAIkqaVHukwiSNh3ANMH5PPa9D6QPCyuyf60SkRNeaSgtdQvTs
BoHCp+vVIQavAVQwm99ixfszYtd9922mlBHVgbX1x8cuir+r+hXC006M7k+qmpRk
G3HKm25eIrkivXbn+UbZ6tQ63eScVwFN14OqwTwB1NndRxP10wXJAUGkWfqtGZct
mAx4fg/bLfFNTMdcdzl8SCiRPgfPO8B0JqtYRihuhEBGdJGxRetMcS+47L3iKKO9
SpwGGcQ5b+fDPSVQpDLxyIueUIYwmiu3FyRnsHZvSHcamGERaPalZvXL7WfBomU1
vjp4uJLEO45ct1nk5MHfpNnGt4/SSUN3sqj/pTVDljxbQBPMsggj8/s/4mXFKbgY
SZAF8RjT2skcLexDqZ+VpzOuSDVxQWY+9ffsIzcWd5MYfvdBNbDhbTiwGZnjEffT
jd7UBmXXaHegeH5JG/oBBO4jX4lvbQRLnz6GNmwQTJvH+Zlu4Y/aUIK2H3H/EcEt
e5rnBgisVY12+rPAwZG8J3wiwEfRxanh5FY7VkeYxJT9uPrr0LfRpaWyqj3cNzqD
C5krvHk6i56vrL3bcOnezJT7EaFyzzMNjPy7Neg/1+uJGi9q1iawSzmtHeibBI6p
5mx9rxy+gGw6maMajEU7B8ILEhFoTqYB3ouTqJgxrdeIU1eTvy05hRFcPrLKYU5E
GpNQ/fK310dXMHyxQXXXkpjQQsweOFJ/EA3LhjxFzmERNtAes+PXZheW30pJ9HeD
y1B7yztpgp8zTktS/ynqBLFcHA/iUD1Y0Tw7/DQZtiZglo64cS3Je7wX0fahOR1L
pnfi2WnEILRO2IQe55D8v0N/PRz4uEsadv4KgNF0QtKWFD8skcNYyALN8BdHaF+z
coMGaEEmQlZr3ArkVZcdL1gMZLciezZdbrv35H3Vua81a9CWl/ZhT8sYlTyqjffa
vbfxDpXZ2JvbYyA8+OuyZ/1+xgunjXCI6TeC2Dci6/Wgb222HwOOzpWMdFZtJ/dT
TVq17qginpwoJMkjtBD7uVEEM7T2jVQTw1WHLzx4rmogc4pADo2DxrW8a+S75i5d
IEY8VI4JGe+9UEcJOZefKW67r0kGWrbhbQpL+f1flvbNiGHq7o3WHUcb4blAsgYR
LdiKCOG8UV80gKlZs6MEV9QVhBh6YIY+mcuxzA/+nLnI4lDgCyQ2XVX5foLo6hZp
bQGf0M3xzU2JviWwuDAry3P/J45GgR7na8nflcrIvim/6z2O/+UZclwaG+OjIeOm
Iv5LmOlQKepXu2nkIotFeFCTecfMojoGUv6bP8jaHiY/Yca/qnhNlWVX9gmW9jfr
eifHSENhUuRIJbyo7TcM1N3U2uAwSPKt+amttEwq/XcBBVnWgmEl41iVeyR4rqRX
nNKoHxH0MBQHIB8IQXm188v2g1hX7Gz2jn5y35wjNtlfMYq3ZgOHI2X56IJrwt4e
ohlBtRPefWTmlq3bDnOQjSYFp//AuuqdBkWYFPaJnkmb9CkokkNytzU58Hu9ELzV
pzjotuhjeQ+e9Hlwhd6bbBCwqFMk4ADDeBxmTnmpVrdCnMLkI80NnQggdrddLecv
kUczt75h0NIVcBUXz5/DUpt7PqacWFiZZ9cwg6tXVBjrnHUFT9C3KBlnQVEd+m/b
XDJVfIEpuEc+aF2brtO75rOdplqbInZIbV6D699Ppqbi1jAEPPHD01gCQtMo3rDc
TDObZIf3LEsWm4oOKbdHqyGpHeE5D2xRoM2pSUrfZb7X7H7Q+MNyXD79rCBhS4iP
ntksMGWSrqJuOCf5YCbHZuBIKXRMj8+hUBHe6WVNhwK8ABCc2sbc4+KfL7La0dcH
xc9S96XjQGIuWHa+scyQJBnVGe9F85Qyhky2huNGJTGHw+WAaIQkSqi6LWaRlnXo
ZWPTN28fqvxGwJqGiMnaJyFtMGufZdGKrC9vzLQzJOhCWL4Qn8nmUGS8pfWOMgEg
IgRNRqv7IqHsfGmLglTPhIqa/Hz1pTO3DbUqOhID61EMtcJ32//njnSBHrrgBCB9
q+528BtDh8ZhwPo0m8s+Cva1DGEB9LfIkTj9XbbcFz7gFMYoOLW6tO+M0K0TYxjg
4UaukFI+Nb/wBfEsC7djCD8He349dhwOq27xJhLZW4o9M/V5CKuynOXHTdRorUU1
PFBsmO6B2QTNkU7pZhMQaz06SYcVQ0XtOsGyrIMzpIVR291XHLNPUMPTOE2TvV+d
TKe0ra6Gff7wgEx9ErFXUMqG/NGvZu3TjDN5NiRk0xgv7ijOUHM7987uJWk79MjE
LLtbSX6u5Kq0mZ3IWr4G1dJiPfo8Wt/7gPHesB3EqiMGkJjSEn4CpskFIq6ES2ri
9qn0mFKEVajDe1hePtUxFY6mqvdxaOfhXqUjiEj5qZFNb/kkemAXfVrNzz4mAqn0
FQGOcRPwnNcVazaESXTM5dEz7z/j5QW8w26RyOctrCK+24QYousPwvB0vz3dM58g
5ZMMpNWkDBZKoC6B9lkx15+wJ6ciseuv6+1hXEuANIMws5PBL6QTo6MreFjfXOBu
M5GnrnWYWs1Y2aP9BA6m4dMx6pymQ9CdxQkC8XeVKHRAKxDchVJMnL6XD4UmNj7N
NC16L2oqy3vHkZT/PvflT+Ve7lQqgoq88f+262IOSnzmR8YTGPiMUZqNHr0KDHDO
AXxdSbEMKZ2bPgtJ59MlZK5RnavPLatUaWJ9flxanSsYBnjJAJhpxqwAYRMHaSbu
0TXgn6xVPTfMzVVdrgqpEZMHTzknGT4HAmPXSBj4HfdTfRbnSsMTYm+AFyonrxHy
detIuYLn7bemD+AxBuQJQUQVJd/qZW3lv/18zN1QrGgikrKibJrIdO663OYiTDzh
8Ds0ccqYsPCdhF45GDtOrSxYZCsuHr6hQJ9+OHwCdrpgP4KVQcKyz3CWHfKneHOc
g6RrQh6j4RZv2INQd5PwVlkFc1EMYJBMIllno98tFCBMladXI8+3EXXfn9r7GpWN
mrpjXXvV3qq81T+PLH8QHaPAffelpM8GTLfQwhDT6kdwpkkDP+Y0saqauXJoBfMW
v/20uv/VpNkmoqxyEH4QQqvVao3zz0jwWva6nDGKkxdxoUHaubXicBraUhwcnJRF
AvV6R8fn0jisHrWV96L6DDITCM9Ebhn/LTkv7it03VRytkVZrynz7Nr0CtRvYiEP
ccge+F8VBDJLYEaOWIJZuTcjtsw7LKzB5TJURsPMQIhi+b+G9UCXMpm8aAWmlV++
Xs9bMvC6v2VJdhkl49ZTomCyWkdMDgoCPCcX3eVQfO29b6PKfNtCVyeOLCsMGJGE
dq5AWJ10XSZSAcsYnjUJXGGUz4lHPOKuCUKBLAUMcOud8JqmwGdA8eJkjpSXe7CH
zhEB24l55W5xoMeUnNuKRHgLGCuZIbnxiKybIm308NC2bBHMj43FskNvYUU9VQxd
P+MC8CzY7s3KK/hGS4+qGfL+QJdzKx7e0dPkBcEViEocjqV4Rm0Kb15b8wdwerqc
dmVEIprSPLBjj3GkTByVAnA+oICUwX2vvkOe7qEuk1Rf5SC91abC3zB46yVcMraT
qOWM8jRwwbUbrNvFWT/NtBD8kmK9V7Jxv+DJLgWH0Lkoc0tA7YHVT8UaWq0FHO/a
eZePewCTjQPFZHxhaTfsG7jBJ01A3MJ/HK5Ie+kwrCIJxLoDzj33vSgZw4h7sCUl
IN4SxiMbu/4az+5ftGUr6AcZsDutl/DtWn40uQMpQaUpifUen05z4y4sJ6kzS//S
UJBP6OWkL1QLKobKgZmGJQv2Dz2wKg2lLLi0xo4/lKksfi5X1OOXxdMmDEl8alH1
Obww4yIaYzoBRn+otemBsQxh0KQ595e5ZOUeQ7FUU3LzKcK3Zm/EXgcVvB96OBhk
g/nmVg3+208lAbLBfZSE7gjvkW5xAQIeR1UTTReuCyaBXdhI1l0xvoefhlUJWZhs
LY/R9ygTSM5m3c9op8n2RyQpFp7BsLZUNiSn7c54TGuUAQ32+DwV/uj7ZK5ht7O4
pd3L50AjUdCYYk8FWZovZQFdVY1RcWPGI3+SsccKdKoEk+kRGA2zW5hb1BYZgSjk
V51Tk/IMkjMoFkXMxXjd7vcHX4Elgddaxc35krPl3gAodY2XxNpwhOJ5CzUbz20t
Sl0pxZLOj9B5BFDu53mefWFs3EeHqB0lJtWhqgcrgIJd5DpW5pV1ZMa3SVA6f0e2
ANwAadmwklJ6U9hP2vNOANEtAURrJ2sPCFKhSpBTTbgPVKH8klGOA4fj1PAymFuO
gE4LRhIwkun9Xg/g7zxPHvmt5PhN8ztA26CAE+b2+B43kXUrMwkqZY8W3dOAaDg8
QTROsth82RN8k+iyztUVgcwVgJYwrmNkJ2/94+c6z2191kCHvQxmCgcTsrkm7luC
AuiTnYZm9b4bPj1uKI6Gf+62gglpjfLVodzIYNVejlTZyqZrN3u3yHJB8MbXEejT
e6XsemwBMLCgS/4EQyFVXJQ8D0j5aggyDQjIwSto3SpafAlRBM8YUH63pbdaORU7
P+pcsh7TBJyoU9EnCGWAA4CE12fWk5werTWbsx4Gu0G8qRKuBwspWf9jVmsCLwu1
A1k6LXUYUYboE2IgZCudELKXbSISqzN24QhU3NYNKhexQk9SGW/xwJ3Exo079w5j
3oBhA3TStSvkRuiCn1d/cNS2uRYj9RobfRVbHKJ7RYPP/5ljTOtIO1gbbpnzDRVG
o703V7IqT2uUHWQurtiQpLnPN+Z15FqJ11S6pUarb015NnqN5DLCBHtm/bktJMMq
QGqnF5fpzdK0yDN4aRKM83lhSCZrMxetKK3nPU8qRvWniqMP8HqU3+CHJkllQKia
e1VDW6w9vV9meXdaYC+yHbZLS7jDhxGYdbbZdez1RK7mDc/+R3uf/8BfKjQgEQjG
FpUbRHz2vlP48Yj+WZez3Dtg6EMS764aTHhO1rhqYyaiUs/K6A7/SxTJ9xUcLRm6
KyssYUA8/ACYgRwPyhjeS5UQDLdHEepSYdwJRbNixcO9ymQjsuFvK8Loh/PjH1oW
YRb4ICPBo6gbfu+2kyUnAXQ6wbB87Mdod9jxyeJu1zWP4eXjqP51wxJq4aDUA8nu
hibv5UDRotUj00+9AyDt9LGSjcMuxMdDknbZCeVF8DsrxsQQPlO9mIhO23l/OtwM
PtUugMS6zJ975zop5V0Myqx4s+59JUXBSbllRLl6EeNCR0d/CwyTNqNnV5gHZQzI
eRvh7ehzOjH0iC2X51D2n+ZrLHVS3yB8N0d6c/bjWSxgcYUCONZZTo3aJ9wbSkCN
wnl7tsYhzAB7O4/SQrZKk5QpkuF5BBqCMuTbqxfs0i5x8ULxIhPart0KpdDAa27v
BffxesBLL6QyCDITfPIFG+3i/LwBqzfC16PPe5+Nbk7LZ3ssgnxd3V5laonxWGGo
Pj1hCILTlWPfWfSRI0ea4Fakf1oxDCF6xUE8VCTZSiODnhytARUoiO9PerZoRfac
+8jC6ZfMiVkDKVtRwMf6OHqyzEpC2E1gBybNFE1hk9ZXJ5RjXcJL9QFZn1NqVtJr
tOw9ztKMYP5txe8yt2HWzImEhTEfpocI9oNt0xNry0v+uCbk44Wudbc3a8k33/by
mzpD9kyd13VQeWE0hrKFP5/mZ0F5pv+nSpYZrfoANEBA+sensCYVXzz/HhEaek3f
DrHdY5/IPuIpvfMjD/X1qmlVblNR8xtAAdxLBSs3nYYCUENWUzqwBDG2UDaoW3M+
9zVn9EyVjAfIIrnD0sof6EpIXs8UoYY5UUCA+/yedh3XWDBLUGOYFcGRrLCrg2rP
+EYDbLV3WBVWSfiCV5Tn9c9EjGKPMkn28bMfGezq9Bu0cEuhflTBpSQUsO70GVMO
/K1+DZW10o2L+5OveB6nSQsdLRiD0MUzXYknwfZ/v8EfyQnFszjLIG3oKSUfMgja
6WehLujjrXWS3uBYd4dZj9mdr+VDnMYNK2lV9Bsb9DFRqEHmFKEMc1sqzKOqiAag
cRFjSp2Le0l9RWFrPQbKWKbRSiuRVfhYmeV/A1YjoMLhb79Ro2oFhkZDEAjrWIJQ
hZxUA8nzFUJMIDTmkXWhat81PzdadlF+7VNgckCDzl9hl91/2/lDaO7K3OFSQunL
OtYKTcIsS10yn0SgcbKEfopV2JoFHXeuyVjBOQh8z1rHA3C5z2Qk9r+r60jxS9v1
QQy9X9yK6gKYtyJT6/jOGq2FxlLuxxOEBjY8lxHuZeMJuJGeRxp2XMY9zqj73WlR
lRdBbyxlJLHaPVFiFIJ3CuVoeB1s1RWn3PH7QzNXgR7Q3hYF7dUmjfXPZFue2YvO
FakzwcQ0kiPTRL5pUJMA1gqCW2e+GxegqAOXgWenlEfyBuGxGDvVI4tn6pI6P8Hg
iaUTyC+hhkVIoXv7ZB/TLXhQ0eAaiUzVVuXxmgp6tAdI8XRtFFaMx+iLDjc9lG3G
SfJOft9DXfe9pB8DMcDrUP+iEQBPg+GWZd0WpDtWDGr0SiCiFbIs7igpqol3DFpc
rm+hTYjd3Uiyke7MkDzKcDgUHfxFJPp4XjYK9tJdSDfzp5DXMdSGSyRgOA8DysfM
FFEcW0RFewHgoxabsJIKuAsmKNqojmN37CoKPRo4bUZV5v1CsrWVdAxUt+hFc1Qd
EMJnBx4sb/9KSn61d/Po/HlqLnepZ+AVfHU7IxLv9DYHKsLqib2qtwzUKrrSJ3aj
3hhC6zvxYi1tUkzTFxxpWs44ruZyoTEGHYJTuvLNSQ4gPe6sQSvcfwUHZfh4K6w2
ugTn9qLF8iRnNzRm4/ivcEnl+A1ZrYYXpW24FRX1nmJlxGlqqSM7iIsrGthmVwm9
YCqh1YAYdr4RGkD0rL5VipqoRLPBpivzqxNBB8K4l/4RSLccWHW2Nas7bb2wi8pY
7rfG94QBJizMw6PzHq7jZRRxdVHjpwdWhgI14IfckfMTUpwxqPoGshndiqcln9Ad
6pyeHs3nFz9ZZy/W0nsrRE50mM3x3Jrjrm/g9l+i775jKH1MogYI55UzAzPDeIXw
/PQvle+mAAX1lyFPbXmmYdKmVLutUNbjCUE2ndqio07M04yAD7AwtZnI8okvEQgH
cjDQO6rUJOWgqUVOJt1vX50Mxpu3mJULCbglVNZXVlG6jXSRctErc0zbkrmc1cI6
iqg4DdTaAM28iLlgOIhufvoy5IKW6lYZgHR73I3mUydYf/E7DrsOSEeYr3h/uF+t
Ssh4JkcAqacwGiM3/wG6NIa6ZqsKXwJeu78nH5U6o5EpAk6Cyo19ddZpw4NHb3A7
V0DgZe6M5il3ySNyKiZmmtmd2/QtE1GjFidyMvndYaHYzxTx7cx0sfxLVopehCZU
uUQLRN7dtZCRMdE0/8ks2zkyYtSKN5cscP325B7SsvKYi2Td5NS85+HT/GnjpA2j
0cKQikXbkp/DK4m8EMb3DQwBfiPlg6zQoY7fpjQJ28Bu/jTNFgJWz6ba3x6qxhKM
0hyPYJxSRx/HdbFu40TZbwcFW6+Vp62Cu5iOnpNgTOTexRjlA8AmQj0g5sIuWu0E
fMlIvwWWETPxppXN84Ipg3VBjzaxOoNCkL/48fSn9YuHoHygk7FJmyt8sd9d8ims
V9qIeITx529s/Uc30OWkWjTmdf66lWevdhqIkFRJqEgHdrAFS8PXb2cUQ6yFwXjW
oZBIG5XFXCc8rqOOCI/e4zE4BLPJxyv88KVI+0MQYTaSvgM27HBo4ntJSCdWz3ry
jHtVUxv6ubKlRZDMN0rIbmFkxbpnK0kkPREo0gDLHOrt6qZaLenxyHTRKR800Gmv
u20imgG+Qy08u5/fn8kCrRzzfQmPtFn3QRLYKCf7H+Csl6RLWnA9+iOJ8TxDa7qr
WxeArVvqlE3/rLPBrVfIEKVBv1NNLAFaPRcE5tW3bPzHTbcOfCVMngK6IG8baMRT
NHkcwj0GGnLUCsKzm87zCveHnCdRx3uNxHji0hI5gSKITq7dXSwWlmDjJ7omWvIX
0lE/TvNKTc12ECO2eVnJyEsrb7BmfO5E2Jcd6AGoXt9dY+nTzorT5jUGL2Y2YW9p
IqiR9kY5UttxCtyBXcCaaDmWKHZoShK49Hp5JJor96uFKaAzUJd6wM6AuDwQDNjw
rWsfoZ7BMaqooA0y2zlc/deUJAu2CdOrDmSiHn3Opwr8n4RAOW44e681k/fzJWyq
7oi4vErvuovLW6njiuk7VG4sTV8rO/5BOE/HEcshoDr7lOqw5a9sdehrDl7o4o4I
YA9jlfMEWOtlZ4ORoDUWgb5g4vy2YyrDDrexVWvuRANvfDPuxLCTkTa51hz0/HHx
cPAiM6KjCc+hMzDNUE+23hCKaWsqz7whDJsaNEcgGzb3+F7qfSrhjVQqoD1/8Le1
8s1Q4K0YA95YtPQBtFtAPGp+ZrZ9hhji9O+e0my5sL8wD7lDBovRCFcZAHU6P5xO
X9NS9QbyPDS52HFBZvemWJakCQdeOA/vV2QGlAppfKL1cOULcSxKdLA+4iWVMz2T
Cq5QZ8mDP0fXFevrmbyzu2avmtYAmv+HLa9+Pn84P9rlROTzWE2Nhuj2jD8z5TA9
pDNKePPfdrpILGkjWGDNLHP/yMUNTxt9Vi1IJ/k1KQfWTgP6/ldhfSxEWETV1fTB
Us8Hzq9tmBUVhR4qEsIshu5R/W6Ibh9gLSeMv05omTODyq1DL/KRG8fOm4b+/a29
thKv8dx7IQidD4bN6NjFfY7LXqOWMQYc+QisGwVvWCLIHCHFwJvhbOp/4N5VZmT3
/mKo3+u2P1LvFIhNMsoITgBxhR5QL7drxRESPx9LPtAXVKtZauPqe49i2iUkC1Nr
sDpowe2pZ5RuXWteL7J2qQ0KuQebcSpX5MYK2BhnD4S6PB376eDAdqKNoi+3GETC
F2s12Zzm5B+DrLYlOBWE3SqSUHXt/a/MG886WbVV/62pTTRWSPW4WX/jx+164uah
l9xC3DjocehTGmXwXG56HUXfZEL6rv6RSIgW6M4mBOEiAzNbGgrPfYdPX9UC1pxf
s3nGPByy0NgKWxdkyyqniF59sV5P2sgvZicWignzG/C9LUzPH3aqB7qWurRbe52k
+OE7Qyu/Zz01A83QmldpBGLqFGuZ3hZPO533LYnKAbR/FNn9BNZMAbcOLu4rbjbk
uLwvqr+yHOuJBHvak+pj6aewcx+s5/wrfsk+YflDi2fcKsteXZbXKQaN23pjfz+Q
tMgL5HkfeuRRr74rOAPKnceJunwhSyWgCOtrrmjftmmY8sfx/6eWfqkGTAYLvYKk
c8QW1teqmZ/G313XXoVgYG3Ij5yLWhveRjSEOwZTH4gwQwnCo0Xv9SW66tKfiDK7
U66Cqm5nREaGWzHA95bVFrdwzrFb/zeMxusCvsd0Ek2Leq2pYa4w+kDR8MshBqGa
UWWMYrL/HmidPJUIJMpqm3N6NiXIUSkjAs/34lWuTwbMb91g89z39X9qbR2OubiH
liAJZb8/l1uZD9wk47glChcSbIx6l+MHaMWy0MnpGCzfpxL/5NsIuCXv9iDN5H0T
co+k3jBEVubX8rdphFS9ui80SGCY05RMMfT61p08lBa+Z+GMmWeBr/KLwx0EuLBV
wizKYvpkC2E1c+6CR7zWuZOO4lm3/uvz7+9XCJVKOgxUdW18vq70Nf6wl9B6VFiK
cAEC5o8u9AkF9p8yuMfGcRtrCtMtrrouTwQSIR/1kX9ba/t1J+MSlPyYm1hwC609
vsC0szuL3LttotP9WtsVXXEzh9gfzQHTk/k42eCWd2glIGg2uw05T6+xYqC0BG0O
XH9OwfNr9kwxKQD4DaQtfAZpGv/KGjjnPm73PDhscHXUi4AJSga6fqtn/k8FyaHc
bM5lsQFZ6+Xo7R1Dkc+/CRjPO2+R/5bTAonH68ZpyxYPHNZm2oDXcehRcv21HTs6
ONj4Xqbq9fUk0d6+IFrDxpaCMzuM00d0RwB+WelQVzUpxUDH8OtCgzg5Ij8FsH3a
LJAjEU7Rq5+F2vm2j/htc2I6vA651yOMPhJWWfT7R6W83frB+lhlcLc4mF799Q1H
FKWIVkgwYd5XlWUDaqCSnK6gpdW8wfx+aYMRV/ShPV8bsh6VQnII03xdmJKH3iVZ
AQj8AiVuvDglVhw+CTb9bhAkQDfFW9RdoEwd+xLiOflkXWkd/6tYcUY5d3389d/K
owXNH4Bh0kpHcZdg/rB/Py1ZghLw3alojhoOO/C+mDqM3Nvh+twwPuEEzFX/ufec
ievuZu+vow8GHSQ30QGGExf6E+PVNEPGINyHhPKFGbx3sp9HW3ywUrt3ChonJBJB
C1a29A7TArG+teAdOa+2eK8vif0+ZSrom7cwboVAzeXBolV5k3dpNKNrakq87n67
pJfp2jFfS2zD5/2x+sXz0f9zBSdaNVGz9sPLPN5ayei/aXIkdOLinHdi4SsypT73
Gmikw1DGtVXzNOkGBnXcTzrClb8HTNnD9yYkGMcSTZHoyi3cK4ivFUaVQ8etRcHa
D92bx1OYLyd/8Lwh1RhSV82D3xnUfFk49oWz+3PP0YBQvy6i84Qr3ScwEkynB/wW
FSDP89hUo1amOQT2nVX2kzXhjJ2GzEOsxtF9cQdbm2QZGYl1PkBBvh0rM6avY7Ls
yhKSzI4HnH0/Lrc/Fsjs2A6WMUpDWy6vWVb7Yqm2Yfc6KqDmQSutR4LPjH6BDfiE
M7ybHsok4gGow7XLhWbv2cN+WGvo0zgi8Szqv6Ylrg1w5P9H6xpFn/t5ZvIdt5Q1
znRll1sVoDiynQWCIvNIM9aCyJftzDuGp6X+l/VeNUstJup+N17PX63Z8Is/3fWa
mx5HOIyW3P7oVXBHW7YHEX9o7jHBfKD3tNriYk+kfgufGcsMFu2O16bZ7Gwr5v/+
KRuzXTzWEhOVhoyxOoiFSeqlpEw0Q92Ew6xetn1ynBNidpMiJls0VIPLPw7D68kQ
nR3BkHISk/wLpvu/Iq32DJlZ20eQGsJqTF/kOiyIp1XH83NLktPEkBSkbc9XgpDS
z2EHMgQ0bH9mthq1xyGjEQsFKxoQXRooMx6SDk1c85HcTPxHHb68+TNeppTJP1hX
xOiLu9ciwOgaClMFD9FTGbYqw9MAhQCVy6jH9TJLhcD1s/piC9cKXZBfm2a4+2M6
Sj6kfJM5lhJ5Te+JMYvUJJY2rUgZafTnK55NxbAfXG/YxLaHqZsROgfCXxl9gBEP
Rdorgu69AyVPkqWgUY6QNMRFPYmf+U8igSNLfMWFQivFOdNv8BcFcto7eDZF7lNN
kho93fCECTeZG/XF2KTt6cVELaUh2zPb4W9JyvDnmJOc6lbMWv2WSEGVQsl/tmqx
zy5Ib0bTJWIi3AXYLdxRl//dWbEfdc4AggwMdDVUm5iyqEU0fL8kdlWlT1TzpEkF
Sy9kzz2Ue0WiBMnl3VZnP04wfC7pbMKuYbtLIA2uddhVwk3D7UQplOwrDEdWwEFk
Op9SWbnQZHNg5jlcWD7DVXv6BAlgQE3zTaYJhG+FmAo0to/t6xTyYv5HaSoK9Jds
YglEDWBtFw5cd8wu3rj6V8tVZjKjUBmBjnrT9TLt78b0ZRP1aWQvAe25yLP6ptah
zXFjjwWYitH8ydxraNr/hrvBCcDhWqgD4OaiokcwdkpgszO5kW9rnDIKyQeV2wM0
WbUJzhnmICu4wTdXcWW53+qC6LrIJaXa/J72604B1iXFDyiBuCZzDgTokkttHfse
zhxpQaYyZSIIE4yjal5dJ/q5PZf17lLAsZgpGxpHrRuTqvaax9GXiviM9RpHZ6Hb
QuGiR/Hq+CXeTyY7QT8VQyGyOzB6s30E7wzlE5OfSGZ5X8o7jlod/9EBNsK3jGSg
A7Aqx7PaoEtDuB2cgxBfqW3KHMsTnHFeyiBU4ziA4PttUTG6K6IMVktj8+DChVIZ
0qNK3rjKwLqaY2bD2Yksr5mR6p17QftTHiYyU8YkGHufBiC8Aob6wHRaX2faXoMs
/XQVYWo5nuWUYFv58Tslw9fzyHOaT4C+k8k7IYUHH6b6uKyashtB0RZGH8TkoR8u
vudtOzSud+bcCj88sYNe8VPj0jNHsq8zqXjEp7QZmH2NhHooY+hWVdC+ROS2PqC1
ecF1Rd0QmX3uW2DGPXgHCmqwNi3s9rMIox0YGYAo08As192mTHbZbJZSasBptuhC
FRqtOxMC1ROw7V1+AdwL1YAf0dbmiXOou3IRnFduMjC4JPut3TP1udSeZ7AR4eE4
8kjIU6nXMpo0xbU/fWjU8q2HOrYHjytqBeKA2alMdeGh9e9M19IybhDSO8kzctbI
hRpUG/m4ssAyUnUWASEUrpYE4GxcHnwbKAQ8mm/87uXNIToC1NXclnnS3FKc4Tw+
m85w+hkzYkMV0CA1Liex2SiXrOWHnbIi5Is7B+6igBaf6ZNpXWQdByLBuf3oDwzQ
J+9GJNz+zP26okQXP2XJiq/3mPIIsoHiskDcqJemine3F/ic6gsT2R1sDQtlGmCk
5qy5rRqf/HukZt8xDjMG4+PE/rQ+O0mRd+tYoXy/sN6bGog/a1yLJe312ha/Vm5g
yUu7RbM7OGBX1vUrnDf1ikVBZxXviZ42U1EI4jIf6gaW2r8SjmaBDg0Q0I2oOrc6
NUTcUV884SmM+UWo5P2AHCin3KHVaSkkcQ4sIsxV0xxcc457ac21qNsiS3gowqoe
SuUjRtbdml2fHt6mtatWK4Qq6jHMKp2A/tVV+/bqWb61xiloK3qh6QiP1gEPKZ1b
0mjIi54Y1s7bzngBP1W428E4xFOiMhQPDpM3P0bzAaCvqz0wkAJy6RjVTalHXa+s
AZUVDQ+PxlT39qIA+/Kzp97h7TIjzmpMzftNTG9q+WuIKpue2F2/49Xmm7nrh0Zs
PaOu5ajMbqvA6xS0zZ8Uew5B+2OAKZraE9BLzRUbxhTWw/nqr1qUVMKqFhSjdR/S
VTRbu0JSsdo3Ag4HfucYbFEvbp+gTT4vMgCSzUpCWkiPSJ384KRyu5D7xoFAhtYs
He7QQKmvqOhyTQ66GsfJSM56tz0fC43yTwWD5OFtfXEtX9gXa+fMZSsyxf9iuVle
HFw6V2v4g2qgbFwxOXipJ+gn8lqL7GsY/Fl3LQz16dWnBmXMGkOqaOvcRD1yOuvD
u4kJQgWTn6bx0A0pLXg5IjEUvF1r4n6n2Q3/NMxNgBuTl616T9+OcD+I7LDdLLJ2
xgbFNRepjAvbYbd0ua1i3CV3PJH9J+nyCTb/Sq2XVQhAxAjQypLngJ/2EN/mBqbL
g21QNOxbrTzca8JPdNVQNi+Prn8SnJWKx5wqzNajGVDUl3VyRheEofj9dk3e9V7S
2eVDHXjjqBHEDiLh+CXmkcIkz0zM6eQc3ESQaWIa8Jlj4gXDQ2vtzwuyKewGwDrG
aI264bL1L/P175xlX0RQl6edNOiBI6yAz1j6Ko0QR7ks84/d2x+GZZW7tbW6zw3Y
hJZyM+HvQHeA7QuowStYIDGjtfJWlOt00223ZIOAg1PMmNKWytP9aBiUnCiUqJc0
seLsNwrTBE3qCm/35MCIjsW4qCXSq4M9hqg46eXkTN03IBYeEmQlkhs/n2D/WxP6
uoXypWyj+t/2urjf/AS8GmtAKapSto0X+SZ5qHJ5/rrk//tgMp/s5/nwEuD1qMur
dAmJjbjpMWDkbz63qPjbkTQbX0CnGtF0muAm5XbTQG8L5kpg2CsXlGAYtqd7gMwN
rCGTooi8Ll24CHnoGTe9SKxaRE3CQE1wY3ZrjWRqXWt7TnWYxXAaz1zOi5OYbCH+
mBsR8CAezq96neTcKPZItUt0FnmBbsa/JMh8z4cSobKn1MeCxM051KdvFCUVUTkZ
KHekkLRZ6kc8v50/ZVfCSXHc2SNQYv3R0/5lPuivXTvJneeFSZgnnF9P3fiovqaj
2kRyL6qR+0c0UgDAhQoPBu0Gh3y8uHKWPw4JH+ciadheVMdRd06ny7SVLwGLmMrU
Kp5Q6wctsj2974ZIiMjOUFTz8HAGsXBp995ZQgj5jvM7IoQVBATzNapuOt6zsNqF
Qzsd+w6b9kVWYPxUIFIuxbbNnG2Z1Z/8w5iyCpdkCbT8aM1AxaCe6f8WtXQvV0YZ
3ZTIIo4lW2Wx26U1vUQGF2tO7EH0cQXV53GI/oE4+FNrnNIXFIOZb5qH9JCByNe0
95rGn9nHVyVkqNr0expVumNa2VqAcSPr2YI+yQkARlR7MWgI3PrcSKGkj06kUG7o
n8ufFyEiASij5HfWcU1xYefcixPtnHXb8Q0eXs0yfo6glH2GgIxwOJi1EqXkNCxf
4GopxiM2nXunb2DY0JM+ucI/wea0lMhTCo2R2C7xy3EGVQAu0BYpDsoyrh6b4f+U
bwmJlPnsPH67i2R8RPpgXZuZ6TmR4CHxJVCCj4P1dma8Qx0astlxF7nuUWgf996q
NYx31oIt2KhjhW1IJMXP9eOywIyyCI7rrfyx69pik+WUVYXmx7k5pSqo+rALbIbe
54/8WU2FotaYGqsnvgBBQxEXZ1cPI1COHir0bFR9/n2q7yMypudZHizo0CQwvnrD
uFvscLgmuZwV1GTTpIFK5wh1t/ASqdDJSoXjl6vCoe+C5ACoUqsp7r9jzcVO2Ip4
MBebc5EAeFqjddMMirbtMttLZ3QPQtc9dtZm47P5R/dNYuf02AHfjkkLRQ8tYjbd
C4UvdflEGY8imvWA3xb2P+O4NK9y5zALWjFQFkFy3NVCfWsKQAgGtKTsLDYpGoR0
8JTpbIfYRKkMbYqD68XlONHKpW5oNvS9zvfv+gofyYYN+UYZalTR1q3bNOkHywfK
/Twb4y83zbF+oPxtXGa8hm5clOK2L4cxXBw7WroVrTA5m+0RLcPnBBScsH+1J6Rt
ZG2yqsNfjDvQF633YsNhy2DzDgX7Fl1FV/feYaOGVvxghEkxipNqaA+2Wx8YuST3
I727muiGYbqmkhKtFyb5KdQ6AVbCUcDvoTuv9+WK15mviqdkPcAGEBzxbL+Us51G
+63RlCie/9EymK/sn+GJQiQ4LsU5UXONu9DJBs4Jd7hs+DdynKuzXhz9Ir0B3Fw4
nSKk6vUnhmPXwnds4IoOHhze4fyHXGfzM8zUlkJvh/CJnw154k9jX2h4ITZ9IqIE
YC3Wz2tP9NQ+Za7fzuxFRt27Cq19/iKZJvZSPBfx2nc7zqMIR/V2A9E+hU8I8wFl
HGRx0x1wMuddF0xBm73JrsAqUhYImuLVv4jEM3jOBNRb2SMn/3pU0xWQozj0cFOA
zjEbimdb8CKsQlgcbjx24eTqUyCQauqc1xLH/mvDk/5se4Kt4Q1G6tIeydfIIoYF
TbKpzjQkAu/BrppLLKWZkL4jOhXs6yCIk8/DuUn3uck7FdKJcxAayWf6XKjwJ3tC
RMw7YlWE+a50OtVIpTJMZ6MUA35qWkcv2/k7gNlirhjcxzjqMh7JIJrFq5OB6zLl
PRcKTkCdx7wAgr/RTfzTgD7WGRQTYiY55GbR+U94h81hEAoRwGRmMTtU3k+KkIg9
P3xQUBY2eD8In0xlTIOQbuLM+HiX7YpvGpKy0YpwrMZbwlGO2SxPp+/8TlTz1rfV
9jj8+j7SDm7EFbK8aelrLNXPb1aDhLbmFoYpIHscneutXDfP+eqJcfH3x04Hp5jF
S4/pLPwFLYJj07huaL8loY9d2r+EuIF/atLE1KmXvTtqMzQgs+4/eoEjPescXHha
6Hv8I9lWWU0Xz6R84Y5zZB8TLq8D9h9rzP0Y3cEBv4x9QgqGhiUhAgT4du3TC6/o
GfbeQjjwO8tOXB+qpXv3R+5oXOFEpHCvH7BHwO9VaMG/VO3RxUGU/HPhkS0dDGHD
EBmE/5s0Rz7BOYnZWLs6u39GZEXWxm0y1iShJT9c0N7ToreBYtB+t1C5FN2cdncQ
DwwDmWQNrQpfISPpWY8+TWJcIuoM8JqpwMuqzkEmLLNHkGsgJKh5jHnzvdTwujmk
HRyBL5n7Eaqo3uhO3IhHTMedRlQZ8sxe5V/p0RiK0TO3OjaX2CFufWoX/UCcnLdX
YEp44MJWRYqpwi6lguiab8FzueyA+OKKqogZ2RUCkGHoUAexZvsoeZJ0FzPV0PYR
9x1oqns/5OSUoDrrmHhbqRUrT6SEiBKXXJXZW/Pvr9zsbg5tCtpuIxBnUipdssBv
N9TRD1qevkUG4OT6HlRDsk56vUUmrczT+45ciRVw+wp6ngzMVSgNU0EGjvoN58Am
e4zPcWF1w2Vim3Fg5ucTlUbVhc1sma51gQwNvlOZOTTuq5IuVAvbX9xVbKsDm2S+
BGFt/XCevO51ez9cWeGDkD3tmq64dx2jOxeDa76LTjgNihll2mnfmgdqd6tDWPkI
aY2ajCOnPQxYwPXfW0QIKuJOCqltWq+IW+Wcuu39oTzsMKuK8oxh2QJPJKC8BkHU
h2ZsRFXji5Q+sYJHv5vqQmJoG8fDrXRJhshvJrZQsjfw5bBOdVHVQfI4nCEiWumz
NdbKLQY3SRNDcZwetdbSzgbH50HKxeSLvaP3Mm0jHqUA7uhTlbkay/6sNsmC2xKu
kcHJglD7s7G/83bVCJwbYyk8i7THX9jcSzSeDn8sB07adBDP8enjRKJdaCN73GtJ
0NlmFzYCZvdO5Vtm4ABL4Hj4T0LIUmR9yXKLrwQLIUjkYaPivnVzs4+w3FQRf/Ps
M2QmHzm8HIWXe8jONorawmrjAI97j4cD+o3UfKqjS/vJuBKm4e1FKfLZz5LxgxNR
bBxpGvMQBkd1BN04g4V06GZ0qyjseZzP+eK9J2GcWiwH5opiUOVPlDShycHbdjGt
7H19kMscfmBIG0X9Y5P5TQV8HDcU3zNcKbpEBXIpk5hhH0JMa2Y/03xQyvfMmJQr
4NIb6qXHZ/qdbb7vbug5uAVyLPqazJ+oSrGK+f6Twgu1v0dSmj1OLDk0TsX9zIdo
h8NKGYzO2h74KzfgIDNLJJ7D9T1Iekd+TWVijPK5AzQj0EJZFGSEeM89AL+3p1/Q
JhokAPKiTAE2FPudGmZ9GdE97vDEt/23W99CjpgMALzBzYGTR19aYBT3voXOizcA
okktn5bHqIWbGlFIFRISWcrPCwGw15eNFA3TJao+B9xG2R01sqLzkB2+xOImZxzU
Shf1i2JlCDn8OamWhBygqn1aBuIs+0ZQmMI9PZoiUx9MN1aCeAxCU1cifGTxhEAe
Yxhm7tfSqD8BTnsgO5wdlTa9IEPeIIVXUrHPDRwAiq17CYalXg7UURPYi2quUmJF
cxdW19O/8fv3QuubEJ8v8NvUv5YR36TDh2RugwheEGfRK8nZQZVarwds2CYiPwW3
a+P/0cTGoa0zk0AvvCiUsgb6FZkoywDNgGIh0oIBixF4PIPWB4XeC+69dJr4RnfY
eXTGPhuBAxPoLgAJQ8gB6tj3hpuRs8MQt6q6T2B8R9d9GWd8n8fuR/M3u6q4Em2z
MwoqRV2eOO5DYJVlClZz8ZJrbdhbWI8LCzt80Vf7Z/e7vmtcIzvQWZPWXcCIHeEn
wHM0lwqXlqyJKe11nM5IqYf8SrsK9B/nVveJQ13zNTt1lKQ5nAU0RMqw57WZOPnE
ifXLT2dXczCavlxMT01cQ31ta9ccNIdHd9h9MXR6nE2YtT6g5Lj39zI+tTg7HXS0
QOa2lYU40AV0gr/RiL1bW6c7eCtwCZIHQi9KnUrMCEWE6uO9ytAgpdpagk/66iqm
jmKggXcNyZUH/Io9dRALtDcVcg0wcF74K2xBrWtCyIYelZbqLAB9SAG5qI9NGseQ
Z0hb7hlVyuYt1lLO76Bvr40dxwESUUtB5aLerkAyNCz34jwf5o1AotaJ7jlE+Qsc
7RPl2Fe7uI75tFBzu5DwDC9PzrmA+huRr4FE2/zOkNLEc9FpRN9L87jkabiK2pI7
8GEYjt9I+CZh6Hx50KLBFPXKe08m3edex0f8kl09kWE+y8dDX8qJPE9VE/9VvcXd
mElJCxYbdqXfpHkDkYdvEI4EL5DT6lti/DkpUMBmj896CyxFhUSrDmvSfv1dDg1N
GdpMu6anvsoYOG/JQoTrtI+Y1vXwK7TpXugJebWpuz+cKlU9nlx9PnIC56bOvIe0
VlHmMMr1tVoTXYZsm13NFdujSjcEFhiVx4ZA4gU6x8QD+AVDA1Mm83UWcbaf0NLa
1bGiG33ljT13rstOQ3D9xN2uJHC5LUri2jpsRBcbSwaZ/HD4OFnetLKWf241HC6z
gaR2Py8PH4q8I/HQFiggr8oUfX5SYqVdllXp6gaF6QCRlyTnD/jf7yBdmlcxJX5r
+wM6W/7mA9dtBnB5Ni0fmx3CHc1zng59t9Yi5J/q5MsE1+gVn+bBz9cmsEuADfPu
n7bRX2YxxWH1Ws578uBJG12UwvJea8aX4t22TdISnKYD089P0ooaJKAl+PxfyfAp
LCRBJf8vDBMGMghZBW9AaqeXqsWeaFJS14SkC8aZrOviD/c+kHJIr5pVs4y7bb7r
cYQ7QExFE4+xnNkqTbEp1qgLtA2I8zpe7IjuCzXMw/0wDoSTjCgcoDbvfjVHyuyS
qs1VvnI2R3NdMMkhanL1ja6fMo019fKHPprSn6Hsh1XewMuo6wMb+73VcWo1kEa8
dNbJYbrWB/S5mH8aUIicXwQFZGu+MUM0OBjlLcSqKm6PzW3rW5tc02WWoIEybOn/
P6nVCAKCo9HIMJGlr4ZcvXD31a/+0GAUPqzFkK6zLglXtQisos/fJSjhR321xzA+
z9TaNmuB+/0ME8qKPZ5YDAQaf6f28P0N7hfaYb4wUMm/fEuvP4GNto1+Q4Z8hlrr
hEt6K0DGWqkGXQ1usLYnJaCP+HHd0Km2oIsqZfU7rI96LPIAW74FB7PD/U/1zt34
WV0EunSup562Rxl1eSaCvlSq6hDnj1vJX6ua7ThMJRD7iuvxDYGuPqkCQFxkhJdU
0P/r4kqI24pcZdimp6LSLqXszjsGYvgCs4prMnoa39/MbI85XRri3YhA9pCVPHy7
681BY8A+mOFIhXBLmCKgr/3Rxvag2fhXJ/atVODhBkuASO672lS6obZQyhdazUTK
dpmvyz5ILxvKVQUApOBNONOmj3bytpRMWzZADoHqRCmgMUNbIJo8IP2Y21w2PN0Q
LJ8OKixSQHvRkZpBpc3KNxCCYsLtbkYazv0a4vSDoNEpB6U/pQ912GDBHyYrECJD
PUr5iYooMwPPbg1u52QmKWJUgstEMPJeip7R7kIMGS+kjsZrYc8ceaG5vLUFwwNa
v1fN5PtHOMWh2+2t54HNTECoB5HTx0mbnTzxP2PCdkN5bfZ33exi5RMex6wtlNdh
gqS+GXGE+RHNufr5JvRwFrdpMioKen8//THG3KSyAVKoK+OCie2M1fauR8mhh3lI
OLc6vKytn/uik3rhmDIkdxQoSgj/vBM95JZ1ch4KGipQOBPYklivQuCEhtKd11AJ
cy1oUd3hPmcUWJreNsgkCcK1xyssppwIb5uJT3bc140cB76r3Cgy7kDaY+eRhXlN
68zfmd4KvJEj34UXM8FulD7i+D+3OPWskFLoaEsG1ZmA7gUZpg7idfgZRJMxCwwt
Nn8o3nmDuRtF29M3kF2HK51+/gru5udbmPpkUJPJRMO9WnkFK5JDy51RC+HxWZb7
0vCI/O1mVLokuQbdNU56gomVjZVTfKmxqrYBN/7yPfRrazvAwCiCLC2/hm5VwTj+
HskoXHHefZd8QQ7/drccAnsnwFPI2O3xs0Lfq/poFptarvutAGlS+GzYXuAh6++O
96YsTSoWvldYwQsb29HiOqHpar7Q8nCG+ErlWY4dR7UJFjslGiU2v+VVlyaDf8i8
m7RpxEM5GrgCMTNSRhr/8w4Xb676MBKIcVqo1fDoCcxHoKEFuqNbFx2iEl3pNxBK
Jcc34NvtgQoANpQmstxEpqEhGdRfE9JopgGLbaU7nR+Z46U7w8lLVaStTXTo/FXb
tep5clcE/fguErm05tN4Yj8KlDpWzHyoOSLTc1C+ZcHgH67BbpjDNAsaLxtL7osN
YSUZvGWFDCqwlKxRxU2WflcXxvJA7BZiqCn0lIqJ4C7pRX9zjhks/DoO6SFNL9Lj
It1z9LjwU4FI0LiM2LYJ1VxtE4W749nN9906bHTGmCR8yGcsiB4I82EXJP7RELmN
TShuH92RCoagr313+0N8iFjPa2Nmn43e48prOr/boL8nvyW6r+Xmm7VG+6aPqHMa
RxxUSP6ZK3LQaCdOIpODfXBYmDwu5pBqBxSbL0Q5zJz05VPj/NQ6rNNMpLe7uz5D
LvaVGIK3pwrsBLKd6J3LL9DCgJUP/VtpLb3zMn5u7ATbExvA0ZPofYhzia2SQAc8
kbme4LwjrhelAXvgEagFED4L/hMhFxjxCByJ0ypBPy73GOzTKs8Y4z7x5Ny7fEaZ
7C3hBcXFCeGE6RE3A9fjw7+EK3DfNMBFVIO+iCDlyp15UbVMNtSMzolZ/xAQcHVK
LTk0w5dCQNfGegD3/VCJnT12V5MrZDj7ytOA9Ak8L95VXbYClBTwQllqGQSd2SiJ
uLSxrCvmJeAV27YTqTetF0toWec6hGkr3xgpbO4wuxymjoBAWK6GVy2Y8GxTS+6p
6Hn7rAll9kW0/s2QJI1mn461wWPfgaUkkzO61ZTXBClJH/4nD5sUjHrKluqo6RlV
WFHddukhtpWE7XeH44s1Od7MqkIDjLqgS4QEPnchEmjhTNO22XESjeSZZCU9BE2f
jiizvi4qTNrOHDxuFBJHkKXkewaU/2w/efK1rfv6snWHxwyeYygIKHimHJ81Q7PR
JrZhMmF9dmjtAwkJ1t3PtJRIGH1sO21gulTj09qgvd/XL3SDaghqO9Ahej1xlJVa
eU8Iu+Xt2V3a6YuqzDmSpkFuwTW9sPsLRgjBQIPG5VkQ7KsjPZQaHzR4vFcADWPT
BXunECTMQ6uaJZlofqaVbaemJbYJ86cAve3173wh5G3yqsOfnHXfwSOpsW6QCO+e
m4QEa4JqPlDJu3x+LpyD+/MDPvNfCPDFL2w32zSB7tF9XanRlUvZ6mh/Mk9f0s18
XwxYorG0ZXRacl6gaCjsdBvucPwyIRGuQGo6B6rS9yMRdapRUx8gMOHOUn+pRJJa
aG6otW3xy8huq/rQJ8UjGeUK6sqJgSm56g6SGRbHwcb+ryLyoN0Ut0p2X1vV3YSx
GlFFq+tBN6ZedC5+CbZAR83w6DlSkx59MrLpHADSb7kweX69rcVFiCmDmim0KdpR
9n2qTI9SzFDnZwe+IMoRp+4kYAjq4a63/S4/ifklzDZJ8cSwIPSqzeyofTUv7Kt9
FBnQZwz/xVLLmusZqT1Q8r9QGgJ2SCStICPyOtJ6I3LZ8RAMVEkFtqWhfzjM4ii2
j491celaesOq4laQYCLVJs0lr+sAkxmUiqjucXO9OliSgyhI2Mxgag0ydUwu/uNY
9E9o+eSIy4Gnqy5yMQhgG1aWzwjaOaJxpa51fLIvgNZ4ObfvXljaC6fDi82Ie3ep
wlve2PUzgNTzseEmyWt+UCy2b7z1me9HL4pM76bxOpi1yhTT5u/2HokDa//uM4q2
OVt5M3X0AjbbnGcn4/LuCG6k5xfkf+4dOopKGId96qzz90WvJfft5zd77W60/5lR
eZuFmrU+w9jMKtOt82j75x7Fh4MtxzQFVhjPMT6v7wZXFPCoibJpMnAMCwHkEEcb
woO82YfdTuLTn3cH44WOym9blgNi0BOnkeArssJHK09ucBISEpyfqm0pFT4SacXj
v9QsPKs9bf4XcOzgPUI5sYmaNRg5XN8pBcZZwc5xshsFbpRyE655ONhbLJh34aHy
5eK6Dy1L9g8eChCuIwbmdrNhdzclgtnKoY01RKvwhh2TcBmDFROsZiUeC9x2Af2v
8Cce97iTpEADugmpFfRxK8zbBofOpTaJxff5hsDtkGOggwj50WMSp/6mGxAeLObZ
4omx5IaoC1ppuumayqyoJOwO5milV33j2MqsVMuirW+Fpi286zYcReP9BV7tNciA
TEpuUB9Vsof1fSTMC362DStMNAJAmud024NLvvBOVrd9QBO8Ct7qS0+hUOg4D8fy
4YyE79/kPdBVehjX0penrMemj7DFrZHLGvCqTLe+oAl9uDLXavehbM+xI21WEOKZ
pM5FaN+EWkazw4Rc3ekZK2jgBhgytpAfbGOTlhWGIU/tZxvwvuHRKWL06h2JJk1g
BkKHk21UWhfiZHSSQ5WPnVlPlZfLw80GVckeWtqvKxrjnibBU3MN/D6xS3jy25wn
A0XZeMn8mOEPj33FVC8NyahjmrXIc77IpsJTUGfUAfXLLCFasNGgjR1/YqkKEO4a
euxY/RCCqG9ztHcvUzLWm1kyfjCcnN6b/dn6lZjzgZ7wlqzqgCujiQEoGIBqLGrU
HGDRCAlKtylH0fLOpmKdi9f3aLCMC7MQWPTXztdXB49zYRLLTDVlsm2PEpc/dmNG
cS85aKcGX0PP5HLJYnSLrKbFaHkU9NzttvyZXRnuqtncL/HSQb4rPeaCotXT1pb9
kq6TgpuzUbtlIIk7334ATJBUStSaFgGbwVvAq2yZCERDIaXsZSEOSb9Tyi0Ekhtp
J+IFkQ6zvFRXf/o6imoqWFjq40B7K2OzGf725+u/ExGHSJXdcVwiKrGnxHHE8kbN
vYGvNSkRB7udAtO0DNVSDfOoET+JnLxht//h2DkEycnCoIEZK5Fmqe/h+WhRJ2gT
0VcDQIN05Vt666F7a8C8aFexg96PDoy0p9UQC/KRl4vr8hV/Qu9c+OydeOnaNtmf
4OtPb4MuVhGfdHP4jEM16W3PT+5z7KVVfSntrYHLeKkA+S294QsUK3vYWvklIzly
DTlnQ9a1JQsOV/NBkEtv5B/GWtnykfeWbWrW18XoZzBOh+w37lOkGCpU1f4zNXKw
tspHgFriClr7P+LYYqZyyDID5VuUFllPwI8y7hoXbdggBLgf+tlpzMQnJ6KZr0yk
wkqDr9fVH+HYFCvhMOYVlH9k/2evt5HwK+6iJJRngobTDF6eQMgycJoFnrJlMduc
WdrRO2cjYh7mm9HiEEU311AAI4j8HcYpMz0WnoDna+bX7atHzG8Tb//coyiFhT3+
o36pGVDizMCNvQhih9hbDKIC2igW4SOa0pBmnDNlnuvmQiXE4Yr0VNcjtKSsuWWA
HaPRyeTglJhe1XZ/ikRLYK/uudosUvCM2wpJQn71lZFHAl+uF76U7gXUuL1Pnqpz
D3aNp2SqW0rzW1BU3DdevGRYDS55ODOQ9iAMmfYjNIoimbypJvyk1rJd/u+nh61A
hXcgmvyV8nA9VaWvrwyQx7KA2SbOImAgjpbL0JW44r4Rd91xNpfTkeJPfGqDw3a2
vBUgtcJJPSNe84ALHTvLS3JjXRHdqC5XkjOVOdtO09SGcurwdj5fdqcSJ3Gf3swS
7lRUQfm6UvUfaDLE8SJ8wcbLdV1dGFkRDaSRS6LHrs/h8IU635fdBcrztlY3ooI7
rEuH5dbqy1XAG1TfaFsgzW1SfmDRFlg3x2EU3sM/1prALMeilyXjDxzzIDGz+mus
1vgAzjA1r8/xOSmhZqetA3bo60801jEytf1sO54T+3xtvFQw1QMlgtBGah6/MEL+
g6jSWX5TZfrAD4SudvGotC2q0bCCricZhjqVnsvkkIZnZrPP53ubvizfmet3go8Z
oRavdZ4u6dL7CwHUkLVD1hVFZ1REHy21KiQ2hwXiivVmZsmNuJ+fPliIqrU3/59w
Od32zrWCOGLB+V2gjifc0rTKPLgr/aojFq2OzrOfVZezhAHNAENslLdX3gnJrPWA
Dj4foKDiMlO8sZMy0Hfan6YW94Rx6A6wec7IdNEekJd6/hAFfu4JJwvX2kBn8SoH
WMgfqHjE4Th4XV8Bqsc1OX9XWKNEn0G4A6wmq5rQIZuUHS1aUfXWB0++QbnKKorz
d6UxPMP2+/3+NekrLLJeXfqSF03xbx9Ro8ic+3GOCoJ7fbxwSxpEMxrNP84jVSOg
w8S0fZfSVyETqXSv9jBBVTb7JLnrqr6qkyLWrk/nIUfyLQCY0vtFIB1T4oO6LCjj
G2NzAghfjZ6Mi/VzzEOhCkJ8l941xp52YzCd1P5pkrhoqbL0zBCiLUkeQbybebYl
EPe3F3TBnd87iLfyzblZOpo4YJfgVkE1pBSTU9N0kQ434GEXcFWHKU3264L6jMvu
VeLtwLyC8PLb80/Qic7ftfaZOs4L3zIRD0MO/LFrODHT3DiIhIbLxAutEpgs2wgg
3OlpfFAKE0o80ESR1hh+QQRZO6Rql15peVp0H1+AYxW4aPtx5u+7yVlR30Roq/F+
w3Uip6v3jOg9R4DYpChrazZcV0Vfoed1z0JYoEqiwwuj8S/uHcRsST7xN9O/fGSn
eAhCpY/Nm7+LGFYM8+LQUKF2Ygv96K3Sl20l4SXTJHi5Ghb4Bdtxoag77ve6sF9U
gSx7/F+kY/ox8/4qcZCu63BD/IPZYegCq9Ke+J/F6aD7uNVR0KuemO+XeHUFPvsX
EqtvuUHBOYZcvHW2nKVLw76zNDNBQd3JlYFLiEjrreCm1XT/lxnlsejKUl0p3xTL
Ikkw+3yWZmgzz2EcdXJw9QmGW6hILC9Ulzd0utoD/fFvpK4+7kZuc4tTvzsqrPe7
SdY5+rx0pD4O8HtJmCNF1E64rEFlAj0zCRsaOu8rOQCDBX6UHcoVKbBxkYdgHmFF
2Xf//od6XxexWFSBafwEtLd/+pcK26yDIDgRfUJe8Myl4ze2OVmfHqo5jQWx/fOE
aK9nEm9dOWo/TPyk85g8EemqlxMjCSS3aYhYSu0RVcHDFxKJuCvYAIJMi+dEloPV
tUp+kkP/MDylcIVgCrQl5zmVSnoWI8mXFTrjlorGJLf5QdWtC0wsUigBUlOBuV0c
Z9ND7xYBLAO6bLIAv8on8jeoFqzfwmc7rhhj5H+d7V2c+/Czhr+qsnik6ufPMKm8
5E6Lk8Vf58+TjCrnbC1TIkJ2t632s1CCmbKf/2EMEG5PT+PhvEd/UG0dQfiqYiwg
RRLLWkLDm14K7FTd5UpCy/nsI/PR1N0Tnn/rES9aX6w6IwqK4WwcUyveuM5dUVMk
hZDdAs5rhZB3nx6qi8Xyqa7tasoFvh/uMw17zT+C8J1aXub4miiR5AqWe8XvYLCL
VN/jahhiMOY4SVsu9LaaczkMbvgiDH4YerWvrLMr0ZnJwQOpN7FQS/uf4BzSVRQQ
J6nn4G/i47vwuObAEVTH/W/ZMTHSdOu4nxNm3nweAmbL09IsALdb12+7f1BEUjYz
L/Ta3QelfK7/G/wtwp+YgDr2IrS+qeyGph+ikN1gUmgtCzNdtIA/gfUlZcNcsuFf
chGZV70zXflgq+oQeJsdGRMgXRx9YCtNGhaCamLYt+9g66XqNCC5MI67I/05GCl3
iLvyOmXcJGlLLpytrR7PAizmimreNAOmjzcma78SiECIOcR7gAEd19TQrx9aH8rf
lpcBjjzWTLSLd5OEECzneoxNU9XXN9OGINuyLVWqflaSgK75lY/YLnyzO3bEOIuG
pqOh8VtWi0LbG+/9cS19notzPUOTay8VVXTrJjj/G+c+wjA2SAzgkbW8Fq4zlYG+
99Vjpeh+6YNFe1cUGLSqY/ywwhhcjTuMcSfiL/aRQDjTaF1AoFGSQ6TbeKZG5TOi
avYNWkKzkDxQV9LG3xK7M5ktADnhlkkBtv33jmm+7VTG9CLH8REnu2BAWP9yEyJO
B+YJ00mgy1ZvEslv7PPD4xDJmfqZDvZRVAMHGaYApH8J08rVmkelXTdz26qOB3V3
QAumJBczwOu1h9CZrnmjhYQ+2hyQ5CvJiMGIWCyltDqihL8++U+ZlpMUdZsxtoF0
rpAYiRJb8QJ9kpze/qgh9e9h5RCezhW6vADdw22+qI41i0JG0ibtYEKNPHBeVNIa
14NQcD0+O2zkKQFxyTgbMblQvpdrQplA5idzSjvegsLD5xDKz1s5MRIBsGGnV3Kx
QcG9TO2W/Z8yB+L7hLoher6Bss1zUCFGCQAtHL+DMhrZQsUE21wjW7CPOOkcsdaA
wLeFHEg2+Yo1aMHHYNPPKNST79rXQJ2SHjajvf7GTolF4p5pLvMY/++kC3mFpg6N
v1TJ7oivrWrNRVIr6OrharK6YEj4SWE3z1JUo1ybg8Kt1MJ8VeffuERfxD/8HYPO
gYQQZpmwSD0WpaP0SOngkPRNe5oTfGKEpsWDpiR/hguAs+ipWJ7PFUIBckNU7lOb
udHECgIkf8jCp2vU+FdUM2yObLUz0hw8m5R/hMhmbIqzWU6/IYZCOZqnYOMybBrN
+FLV8rEETmhDtKxycFXG4Z+RDtZeQF3sSBB8MCzx3b/Kgi5+g2cl8Km82zTYQJjf
QtMWV+RSlPNp1FnxqGD/30sETtwljU1o72zrhBRQL9BSIedlLJ8tykGHhOyLGAoC
oDMpCPzraaxydZpPU0AWwqujYHW0MFsphRUSiQ9fb9r8Y6ibRpmYISrZTNlr4ryk
lnnezkUJ3dtd9cIh1DuCKLSqC7MtuWNwnQuTW97jEQ61bAgQezwPy/izBitKeUpd
BzBYsv5lePDgxNNpOu9B9B8jXrLBz0K+KQ0hcWMnvEUNjV8/LiDZE31o7i3HQMtv
zL9e9NXKJX65hxWA2SbiMoAN03nKKyFv+bU+iSCWJsi0tWnT55wpuHOhWQfYd1gZ
s9h4oVHSK0pAmEMLptxH/wrFxFOPS2Req/3l6/NBYYCpkqGmht/joEjhKh8c7D0m
mSiDw85zBeli7FrAYM2e6ucNk2O9fI/L8RIyctLj8JOdatjBt+oBb0xMudnVTUuc
P5EdPwGg3cWEhXv7VaUQ7yabk1wvbNT2rTtAxh6YSd+FNtGnNBv/SNFPSeitfKLc
ZcvFMeGgEcyhnFxX61y4J4+KeX11kCMyntLd0Ks8dwRaDrdKZxN/13BHXzwkWQyA
z3QcpcAYLDHmIGliiSNtE+HrteYj5NxoQAU+2NRZxirIDMEHvhyBViQ3xJS91PkT
7nMH+IlsFRkmhjjWFTZTDGK1e2G5pyd0FXAqcpq5UqgxS9lB5qnVXhk2ZIFQBiN5
6x8nAM6SF3QVZCy6YQchLLS6NGPoorZJdV2QPJ3qYDCFgq+0tfalco/0v6uTy2SZ
21wVM9cCp35y2vLA6nAXSZFXKd0VcENzmfcQHfbfOJH0tO9pMhAHeist89lSHNnv
676Ydp0Px85Yl84BE2rshSoZogzOuw8DiO+8yHuK0tj9NNRnQ4FzrmBW+pkGpQ/T
gBcO/lpGa1vhPcbnMbtFAohrBb4i11oz08Bezd4Ki/dTCyYSz7IjVVpy3UKO6ZrP
e9z0IRT8MjVO45bH9msENU6vGxJcDbNER9h5qvERI6fpPk5b15dRgYE10xFic+Yi
ryO10w6lq0lUoQF2s6+3l/65xZpJjdmr9g6Mwrym9xNQyFX/7mxgQ2VjFRXFR2lV
z/WTZJMvB63yM9svidVIXhwX1tIe1tSd82ATKhkm3U+fjnljp5p6HAtGkkQa9K54
Mo59Nl3CkLEWjJxg3MjOvUnr4Y0ehtFDgdU6HenHDmvlNVT3AILRIO3cJ+igyeTj
0Evt9PBJmz+HhovERZGUbu44sOZNv3Vmjs7PL3MalmSJ/roLusu3u1UY3ZAZuxI8
hPzwYPl7Qyi+yMorCErAF2bxV3785D4XPAcSEss5NDgA93GjeWmpXh38pXOExjZ7
MrGSIvbu6E/3bTmujuhvzooLmPFpIPqmGo+XaAfVXM8qZht4cFn/DPVybfHx5+wP
wfRQPeopLQiqDJC/Ae/TfirbQM0DOZYD/NIWeEs6gvqI24Jx5RbgH1DOwUKj/cus
SK/6gWLyHxhoAJRwpT2BdLri9Obm7tc3I1uJIJfw0Fcu1nGisMMJYsKyIqm6Itkw
MzqviEeSGBwPEUVVq9OPrnatUeWCMFGvHBpIkZGdgkelZ+li4tLAXsYzJjGNKpov
6XRUo7AwKDKgdEKf6MDMvNqR2cj8OQcEDfBHg0z+qNF1ermvgIeLdTSCv2ZTCe3v
Zd6JAG/66RKKycfZCtccBtOpL4EbJ408FNqbslWQIGN1i7hREqXJC9NQiKYRiKQ0
NxWdWSASEYWLZnOxdN+N9rgmRXvTOLhOz4UuygknfKWhHBVRpFFrRemi5HWH5zsB
6zz9YSwVRUD+OkpWDQtsgsUm3wGIw9Gndjwm8kvgm2wn7d9ANNSTKnXBu5ktdyj6
v+Xa0GATqmhRhaUDKAUn6yxEIwSoFtvjqmXwfFAw9ALs0AqDk4XEdUI3u5uHG8pQ
F07UQJENnExD+cuhR/UOWQwvaGH2WtWe6e3Asris1TXl/bV4NjGLWE3VmmuruaAj
lNLuukaRgnCy3HY8x5gWoTevrVg20mj3uG6teboQjJzga/ElPpdZLCjQyVSzbSCl
X0MJ2Lp5+JEg0JiPKqFUmEkQnTWSdGfnbC/Qx/DHtPPwjn+bX80GDkkpo81K515p
MUN2ZGfg4dGhQqG5ry6CMvPDQ/der/1dr2YidS9M8Sd17Xi0ID3pWvwkbEHDaub2
evUeGENMJ9RQoy8eeahtGbb/HqKhUMpcGM9BsPhy+VUCEr0huLmpiQhVXlo+xVdv
He0JofbObyD9/TZzQLTpp9fL9RB1tSP4oPJKvAQaZqexNYmUiejxyXCzqZlPb5P4
5tpR3Byn9/lWsu1TeHkPfHadBqr3wwl/XgfYiuL/FO1Vuen+4iFd2tJ70Z1/4dY4
cYfg/zv2r+YpT8vvhenVXvkSO2gBiU6GcPVzroBiFuX8cwede2VEYC7raO/Osj7p
NFmJKJ5jJ4MCOVXEoLl2JP2KEh/os9gMrPm40rpkSXvfhG1CeLaMOdlOmzGB1W6a
UrEqJbMMBr9e9Agx0J4PyKOp/xlSm6PodmIAC4YQq+TiSETOK5ikSNSow5GPuf3V
NaZwafAZyb1GTqEZxaefeEc7gJCdD2sTTxNQK6XoEI1aR3MoKzlxgr4LsKm8eE9l
rMSlyLeEWTPLvbuX7fsDGt+wOHROgY3PldHQZdVPvOlryGNb05Q/Z8oaAHKsyxRH
1WKTf0vZwzGyyS8PxBLaab0VObeKIFxCIIS5fh01Pe1LoCF0cpSitodE4DIgwXVe
O2aEINU5o4ZfP+dKf5OEVowZhuJMioDmKnqdgCWt+qtUz1lbz2VorwqjEveAe3yJ
CGxcBQQcnsmhso4fvfWpAlEN9qld+7llA9+ztLbXrdROMLEFUpZy2D/egJ6KBjU7
5WnJK5KPAZjlbf9Qq2Uv/zQm36PLtbHoM/aBcXDaDNGJ466Jg1ggjAv8EgS1qJyY
lgqSqA71ycF/vi+ZdAKy/BBKjfDcTD3q5YwXm5SPKGCtlKDqpNQzSZw4nHfqvzwW
cE4LXCG1L5Uk8ghY2sIOdjNw10yYCW9197nfVvGX0JgBJx8LCoC2ASeAhWQmMWFb
QccoyjgRRAk3JSPDdMaZuJJzbqUTsw7jeOksUooR28GbwiCBlEgbEhpHggSihe6B
sq0KCqtbmDOFh5rjruqLf5ewBtBbeny+SyhErhKjVngH8YCzxA7xjI4bpumn5bdn
YHh/OzDPixsBbv2zE/rgESSzltAujTS17/ABMHIB1aIPepDa5ohdyU/EMtqVIXg5
BvP+ATthgezt3oVAoCIfcZmWQzxvnRXHEc118pBRi86C20xQKvk6OhRZaKBeuiRX
omiNUKf4dLS1OdKk4axXX0cIKLew+4OY8tKka8dAki//Skv1OHcqtVQbhg9fyRoh
8pABvPe+9fHXLu84sHioo1m2WL4WvndBNF6+vdu3jttAMNo/3LezQdtqE06npi4T
kcZnTxoZQ09VXhNWE/V2FEgfNQLvK5O/0aGwEtU9jHuj0O9JH4xp4Cjxw0ks4nK+
SusUhBnXqSmm9OnzOjIBPaZaTbKxRJlcF47CIq6BSOA7MlVfNtSRIiBiugGn+KaM
Eynblxe3EgqnFPc6fl2rZVgDYMXMYdwu+d1hTSDz4f7ROUOOrXRdt780XgoNoMqZ
jlvskWTx6I7S0cxj3q4LXIiavK26G2X7FVTT4aukR6q4C0tJpdm6JwZQrQfafwWF
MjvsqfDREY1e3v3LyGybSi1hkhRkMeeCKJUTH3O2Z3Lb2EoBm/L0bRHEAQdOSoSH
cxQyFICjYKbSz0Z7tpgIxwNPgHdvdYnKkAfNfIVcgt3cgr75S9cafY9aXFPxkyj7
PJNkRzm9iiHNW808k6dDQ7IJTirJ+E27gXk8iAmULinepqo8dWbe32J2XzQM9Rjx
KsosuZX3nkBzEu/irrpi2vd9sMYxFY59D8aGCk+X7N3DdvscTbPBizNYimhZXjtO
0KduO3HmzHYKKy9Wbrb5WqfYGUpUuq3hVEuCFv+BRP5/SxUkxIAnbjmHHMX5B4Kt
EIi0AxMoqJkMa6F4kZvPDRLDiQzR903vHQlXrbqqsJWW3+ArSVHI2edceGr1ZO9s
fXXTJTs8VWKQ2nmcJblhnAneQ9f2A8W2Ch9ODt/X/93MuJgpdaU7DbWPmqTfw3sg
urwGe+mAo359EDCBlHoknHQG3p1nQft9idTKUIGeiZjnTDwrKmNeDgrefRpRYDYE
WGxhXwX+UC2CO8czbU9yK00hPpJwEztZKJfNzIxmj4NjKU5phupBUPdTCxJWwNHL
QA5eLgK0U4jAZ8r83nthMYoCiXCTXCXyc12FdG4vQY9t2m/7Ok79t6qQODSR+cFi
dgeN/71113koz01zE+kkPRc78d+zebnuBsPly3HiNbOS4/+qz3wkU8vhigFkfqYK
5oBbnNq6Dv2gF9sCSyqQKvsrh33rP2uZG+zHH3zbgV2h1VuTKtGFVB/5v8WUVFXC
yYoxgwZSxyVY7bRKpkAVGEXQSfuqIM+fCRvdp+rCc+VxLuPsYnEIYFI+ul+o3+h4
A5+l9yxr4feZqf2vAPSEDrCl1zoyx+iFvGyca5Z+Z5bxVWQcdm/WRFlgtVHJRiL1
XssQa45oTWnaFQKnTl/nTzRlPCifPmmS5Dz/xiD9j+kGYlX61/rSppLGT1VOT8bU
Ue6fZy9JrOu+8WSJRE0x0tQqzGiSAZVM/n0F1wL9bWyLS+TNL2PpHOMt31yn3ta1
Yg9ybgoUieX184/m7XeWpZM05lHAxYLrjqpZPTtABXPf0cGch0Y+m4Vrgwh2aKaz
bufM5D4fzPz1x41ykqSEJU3uje3zNMXNcOEZU1lG7Vyilc0L2BA/KAde5kx7jaSa
mufVrFhWQZn0UO1Ipxc7nhjyZFFp2Ye/5y6heS4f5UtIhMblH94QvRxUGBZy1hH9
I4uWhVmNadC3PPyvG2E3Mbt/EYkFOPh73P3tz73Fv2PavfsGGGLle8ocIMX0DdIc
eB9Y7czxp3WGdlFbLYAotQBZCWLDdrGyyT2Htx3zYiSxlY3Xa4ewUmV8FAMbybza
SAX7f9xiIr592KTxWrMvuB47zp22qk82qBR/tPH0/3CGzuZ47zwQNRyd44svE+Ar
cZ/B4Ug/jAr9xm1dO5TqWLe9LkxkBoVIUg1gfp/L8gVFLriyVCLC37dWXMV1JLVA
qHXTHNEj1DcPALM0kl5klIbbBQ0Mc4J8ztB37TP5OOjKI3FbFzseYNGd7Ma3tIqR
XpKGAltcHSp57KiGw1kGdOFkcP73rgxdcfYn2aDW/lYEPmSPnsySgF3P/dXIrWc0
0ovE7N3UVflc9xkcFFgYM8Ncz/cAn4bfkyNDVoYIayByj4PEJl3U4wgVBbtPDcvm
T7wlmrMTOrkZwv8BUd2y79lGSShBpiZS1c+WVzGxpTLcX9AQbgJ+qF0qagoKOmXF
KeKUb+R+pgr1bDioCZn7fyU0MUxbQNrknyK5WsKCm7Yv7B3Jvx9Ar6F7vp3wjy2f
xm0Sc/uPtzzGc+d0zht2TwsQs2OYR5wbJEe//IBQb0prahfZNofu/PFO2zgH8LBj
H32pXcdHq6t4/IuYIQ4RbPpNlg5mjosZL7lxuLXFBK1MHgSgvBLXCy3SiSbkIzsE
K4iXs5pL9VHwLhuGvehqUpasLVuD6b1hgMC85dnqvDRYdB5nV6m+GarPIqxiFmW8
UwztLi9WrvKCbGSnbjqwXiZkum6jxzhjvqv6Bqg6oOy84V95bpyXpehrGg5lhWGi
1FyJWkAdHbZi4GJvyXm4rZ10xy9OIEb3/4ct5aSKVfiuEgaCCLqeffm+jFCe7FU1
a3q7HV0sKX8IK0TV92MXYb4OhVPs0mCqg90Duwe4H25R44qE854DFjSXUtyL/FJQ
2hrqdcL/O+cQ/TjqPT8GhcIvnQ22PgS3ttynN2MjOpZ4riSrtq4Hrw4HuVoZwU3o
Siz/4w3HeSTfH6J57U8o1RouyGdrb2GZI/8VpyYupIrXedwuP1EYJWekZ88zzX0F
paOKrzdOXavFQFvNdgwhx42/37sU5msfMqV6TyLABSKhjhDK7DG98xNg2QU6dFU0
qM4o76/8yEvUng7oMNK1Cc1+sURsEIqfSAPvsFyOzWt5XXo0wARbrbd+yU6c+UH1
NjdjrRJR3bhYYq+oxnRtpSqW7zuCR1OiuGgTfp5OQNWGXnOLIYQvp6sSD3FxogjW
Sk960kNFnTxHzkCIen7J7eAM/NR3j7ELEBmHqb1L5Bhtu1M+t/m+V4nd1p2a7v1M
lggpJB2TM5SKFtO8THYXnBLajli+UncUyxJ68i1JuxfLvE9ZRqyxHif3p2poVEKp
5Td3cfY9/I9IzX1ze46TsE+NtNdKf45p2m1zmgByM9+UAUcw4niwGLNJbEF2DbWM
kmt+1bABAtnifao7Q6/wn6S792djRyEBSILf+6joYjWWzNYjdrnF4mQCMXK30FfP
f0ER0Z/7kEKBjCT7srOLmHAOca25ozJSc1IyOMVgushhd18YPKCKfm3VFE2cmn6d
Exi+IDjm76mQ4ubRIv6jorZpDPXauis9+DY4/jTH3fmcHOsbE7aG6ziHKbZPkVlZ
774mrjGhUbcJaplRQ0C0HHsNLbhwx1e5oCun5OGWjq6zI+v9ej/DTfR3PQa+yt5U
HihhQuxxbU1kDGQJ8oi0vN+r+7rdjrPmCSJgQUbWFfeVCrquLP162n0Q/5d+/j4L
viMMImQiq9J7uTcygeflDjE3/NmqcsS/zOgLzbfjKvGQ9js9WaSn0Wp0iwsA4EtF
DxWMOJwUUAWmqmItjTR2qMFh2myuMhKJQmHV4+V/o3JB9GD3BlnHSV/Z66+TWtT8
XVn9zGbMJVosQ6jR/FxBSa30znx5oLBrI8cHPZvEN41tEDCRF0q5zJZKN01XC0Hk
BuvMO3riMAI8qIVV4N1A7uv3uIdzARVTzX2tSx0R1EsyWDfl+rpdoLMlCzauhm96
25bfWKht4et+fdGgeCQrYFyYJCed1VwmX1dxB1Uiw2VzSB0BsBWqZyn3dVmgNH7m
asfSouHU2dRF03RxDyCZkMtyuyrxoUmJhhW7frQ7NbkYQSsGXcrK91E3n6QC9YCn
YLGQ1dnERDHfcqXuejb743WbwUk9I+rPg7vIN2j7x3rxBVx/fo/7YAHZFRMKaSUz
PTKGJfYdPXG4Nz6377kZH1LyfsEuhkMnlvB58wzVY9XayCyXJhPVoicBF8Z6EGcC
e3wtmWTC4hAur2IiCzg4rNtexvU86HfSp+6oAKp1FAIMZpmszAR5fxlmwkitTQ4P
LcgtnAGJTYJZlleya407jxpTL7rLwZ5B1FOlf3O5RAHuor65H5v0xtMBJIwBehux
3YZB5ar0Ck2RX8qnF9x6kn6C/bOorx0HJi7CjL5950i2W61XCUwJdFDIIQboOoYO
tk0wRKQ6oIMNEVTpSa0sHnV9v+FJjHPIIpxpu7Nag73TFzQm7y/jO/nC1aaixzSo
1gDtRZDki+0zB5+J7RR/U548JQH5xYbx72Dum048ksPr8eBJSTvnb+fS8FlhQPPy
nur+nXjoR4ffqKCDJdqGEsFLWtUFbvIXPTu4dq7+HZXYnxGg2U9wkqwZnlgMsbYB
fFhngtvffvuuD/QRoqQgySI16uhodcNQu6gNFf8U/uaQk8WXYVH2T/o+UcaLwBb7
GjP3XCODsQt82K2nYf7LB0rgiOoTAt2Qr47cOjKfym4UJx/kh9Z/oP5rKcyDUjif
aLZyD1bSrgE/BfhElWWMPTAd+w4Yh1q4xwKulEgHLZ1i5FzBSh+OXV6q1aU9T3AY
f4PVDcwaG6TCYK5L9oP96Q3AljwqKYG6zsiNYE6mE5+aqUxv8BhtvNTJ+yTd6H1v
jx+xZ+F8Bv8lxX4cAc3eyikDAPhdLHMZ6j0DBYlL8IOmf9ZzT8LZupzYBV5h07Kb
VtAhl+QPtvOpjf1uLkFWTkhMhKQpVeSahbmfFefvfR1hh0hPEMiOPVBOz4qfSiFL
TZNBVc0wWs9zxh9neQh4ZJycv7E9vmCGflIY5GhkYG7Qb/Xco6fxO9e2tm2nH3oN
CXTs/wLGi4J8ywoUoetYzx1gL4LMzejewNZGeW7CRihmGsxB/qdKQPztYafBZYTQ
n26pj2HDBZY5HPSQ7gLxN3aTZD9eCpdm4+iEIUMrbZObxHP2PZKDPMKIq+E1W+Tq
enAArZ3y5QZTKwBfvdyxUHi240XplNQja8OZrx5ZIW2VETZzff0vSJ8D1gKrBDuR
xud/VDHUvG4zxxIAtMXDFOrRFYkouUBTi1yrjr5Sygc1ytseUIVMmjFdRQdsAxt7
QZzjBKJW6quQSGmE8ZtkLwKj1+CiyAyJdrLMoed9LrUz5iFzzAFZ/7wc9mKFsRhs
xh8m7JcLTi+GB84pWJSrx8NvsC1c1nGboBrolY2zLJJoHB8mauL9315ecvFBQasN
CLzvaOQFpjU0/zp8yB+IUsjEF0PZv++SMfWHiQgHhjgLRA3UgJG6083247cxhj5R
DQMn69F4od1IY9rl35kvwCbLTq0JLeOFkN/rRKZnm7rLemHpmDsPtkAmrDHHtyI6
OetUVhfk55wJkefO8LA19KeZg5L3ePHU499sksWyNW40+7Eag1H+NU9Rb6IN6rBU
7PKSKC1IYeFZF5G4W/RVaQHzgJ5hvDteGKG/H26zys/XQvm/0cWQlMt/6je+PeA4
Wldv2QWFtjTy827uya7WLw1gehsJyNim1+giaZucDt0EAXE78zg2C6+PMfiI6lX+
ZRpBDCdWmEUSjwmsb614uv5sLtHR/Vxdqpw608cpIVKojNjz8TLMosrXxl0Jj45w
yYJrFUqbQ/3hupkFVWluBIxyhPyXw9VrdsLNJY4EVJv/CxSW6BMggNmV3EBbEcCR
c+oVz4qD1hQp0Haxp97b/CsnrMistnf7JuWagWqqMBue1/xVqEFhGh72x534Hrbw
p+UuQZU54AT1VEAS8yBFmOrcYlr9dC2B2fuTLrNXZEJoFoD5+jfba3jyeYNFUGlb
1u+dLksgNCDgnVNIqve+AX6GzZ97KxKko3hrC00nUCKhoimpi92Cs8vfV0bs/4lR
TCvJxhmSgSBLd9R29BptLmsN2R2lHrzd21ByeO06fch6y7b3PwYa56JKrh9HpXAs
8hiWdd2TyIofapXpz354SmKLJtySMmeBiG6FRG8p3Dg7Bq50CNR9S9DhWw85L2/g
LrPZjlIsE28gUyxnybOeVyIJqMKQODYW2Sl6xgb7V/Gf7AzWCS1PaCqouKn/tjXX
5hmxtSeY6yuRAK6TlLKgvH07RODoM4twKzvd+OvZ8q05LncroJ5hALyOo+tJ1jRk
lA7YVXXmDlDUMa1UIpCKylQO7mz878xobXEELrfD8YX6+BEBJCbXO4IiErTDhulA
BQYpB8qCc9g+WnjUrH6b/26TEJ6v+HDs7h2N4xvi8syHmYKbHgx56V2Dj3DY6Po0
IVUPyx66RZxwr4UFzCTLJp45/gNGEXsLkNL73LspwNK/qGNZEPXr5uRm94ML9Aaw
rCAAqlSjfu/c1mvRSUjld/br/GrVliZ34BHQPHGmAvf7aFDAMrZ9r6N3Df3JrKok
ocOuOLbNqFZlc9oieJVBWdYR4uykBHQ8CBfcQC1YEAam0geA54EKpya+U8nbsSs0
G6g3NKsJuVV3tNbQrzw7RosH2vxTJqjIrDe9YK8AL9meK9W5xwxEOKpQiH32f+8c
BcWt7FRHOWA/kBoy0F4PIOfK3tpX/pXaCDjvVM0IE7DkWvioe17qMZ4FBe7vGRUY
rxbGJ4vEQ0KguymxCQwq0Aim7ncmIQ599JYRKP5zeTSWxLASDC77DR6tbAR9bVHH
QVU2wNmmgxRofOIBSq0wpwmXQ+QXMHYl3dvrXKsvEYzau2Wp1/zFmRZWlcRf+Wr9
ijBgEJoXu8va53Zz6dRyZXdExfQFwn47UkQDY5Hl33mzZepesrAPw5xSBkdWuc+W
QNw2rKu0c+JTO6HCvqv9qknMsOGbsLAboRbK0N/YMJseTYYECYHTzNLHv5Gxu2bN
d6yWXfhghCV4JcYzznwW3maRUxeVrvhv1E/UPCL5CDhnXddzoz71YbO5+5W/Z5H+
mtXFVsGwYqG0xPmfS6J7StIMd4fyLnEonT5qLqXW+lVZ8aSi8UOCgpu9FJTBt3vL
/TdMnkLQ7zL5GIQyaZ4S4BVNFO4YTvbbBvNwqa2N1MksDL+Guat8mtYXqFnVLT80
3PFFJ5LW0lvTGOmNLShB4ECmnu1LLJOGD/WOBAqF3FJxUNt3k7hx+bVQJdByLecT
yqxZpE7LDE1cwFhHE6P+FOg5hAOULjG5XRv6Q3m1dhtoOuBeNcykTBnTPrLtN7AD
U1t1+xNQ3xnBAyMaylwq9o88RmjYvFphz+jwmh4x1cNaW6MdKr+UusKqPDWHSUjb
XJc4GbhTF4eTq9MAgTYW6RdXg2JyWzyqrGrKGiUhaaPSX5U7+8iyHN5rA8KceZPM
MeGreQ49v458Zj15VLTjP/zPmtM3i/pHArHRb4ZNN9oOL60tG1ex/ciTm1etf0qu
np2noWuJZo7oYOoBtz/j6G6N6u9lbMRWJ6Y6rMmOrSpxfWgPse37lzstLvNuq1py
6kXVoGpTEp2FFevhW7kl0HuNRqAcwxiI+X0MUcKgK09Ek4a9zk1ClDLrWRfIpGxG
KOfRKnLA/M/zMioE3BL5If/1OFbuVadoMTn8ohAPL4Hp2Xw5v2zMkwmsNvVxiyG1
YtX0FZ3e0NDs6wbCm7RY/aIffvyfZJNqnl1cwOLWJVpEmm/PniIBvmIo0ojIeiis
ItKVFVshDovnxp8YGQkgvroruOQXOK7wPBN8yUAk8KuTUkIxoHGBSLTk8Gxy9r/a
nwSC1D8iviJUtxZ3akp57lC1AMvlu4360vgdsHUHOLEyrtLHgk25XmU5IibzdH3Q
2NJM98BrpDIA3QCvbr1bvsN4WuoxzzUCy8SEX4+PbBqU6AVEozMqqe+OabmZlF/U
8jHZ+BZJB2g7FsNJn9EhbftM+2c52VjDb2QWcS4L9r1DlIpv6aWZUbTsJGLnkXEV
3zFoDrZisuWgPfgxHQ+NQ+9H8tzp1MAPf/xk/JV1G7WFqk3I+HdGQUZKVdJUIXTn
lVWAmJnsXctI4r1l0lrlCJjtOxbiS/jaDiEtAKUhE2o5ApThbhcgdzR56k3M2fH6
BcPKCdtFkRNPi+cpNyJpveVavP7b35NWFEYDs0rXpi8SkQX23Nrh4zWvcnw/CVIb
Gw7JPr0KUJ3Yl11aiktRu5UpUNKTLEPFB7IkguSPVGcui12W41bcdGEnK98zZwSa
Nr83Q6D+BgsQZ9E3XO58aXRd2UGk1oiYIZMtYvQsDin3TdI7mPEJheRE35wnBjrR
y5LUrkYlPovnGjidHVJC1lTt9zLc7LckhZqIf012TyiyGy9TEssbrx7jwUHRJSo0
thiWXpT804XZl8XCV4bNGGhDDZOcs/Hp3ko/N/mVANWuQ0MUkgy21bQmxo+Mgr+E
4SjpCiI9iV8YPpvhgN+iPLxAZT4Ew+RUTIVoPTWJY1+U6wz6X/7w3t99XVozMxQB
0U250EyuSNHLu+2nlZJrxVX0wjAh+1d0oQefGwkXKqCUm6QN+hWqGJHrzdyNpEhv
tBDF2aFadHexYLfBIWRkuP/5g6/yic9moPrDt+2EJztzuZ187qGF136AHNSydFL2
h1cfC5d2C5YgIK5nSOtDc80aRe01W1VB26nMaFNU5CJFBkX+HWUwhQ6YIlBLQqUs
dwYkSIhBXKBuX22/kVPtPLerl0ZwGLVBhEFqA3PCgaPuE6kFjlgk4Oy1dauPi0j7
pQ0CDye+mgVUaVVFRBSxyAS6hI8zrpG00Ks1DEIXVUoyr22MTc7SVQjvYe7oxehk
eYs4nPRbjUfyuA7fvPOE7ezHzlD9VpQ2O/xGksWWaaYHxcChe3n0O66dLJRBN7vM
0UnGvN2OXZMNnHrn/6+3wsGhM0VRPVrI/2r0+RWehxua29v034PMovoK1PUudT2C
VuTC3HYHy+ugL9okXCWh4AhA/JzCmL5qsainChMejqOFkJfju1L9KjyfUSjUZPST
kINY87gNcFgn6RZevnetfvGzStj2UjwxD7VNS982jMJVWdY0X8EgaGyz61KniPTy
KMMSL29nA5RK3oqTXTJiUdAqRNzCuwDKfGljW2SLzy9dq1R8Aqjq94Cry2x4jcii
3QeULHKkqwmeaZTXYasA/Q0/C0o4HtP4ex1vt+YOUhO3jZ2XcwWUjvHheyssDMOm
lbHaj3xKqliJuIQkhgOa73W8Pd+5Xa2Ou6rWZ2Z2atyK3VX5lflA7/jPmmIG65M4
U1LI9e8/TpaUElDEOsnHUSN3ZLJQTuLN8MLiMIDbexb0hV0hYWETJmIa9D+vzPHy
rJhU9SGYBZ+YUMju99XaziARr6sMiYzUBHRINTV4QsRWI95y7bj1Opa/Ys2xV1Vg
K7Rr0yBSamZ87WRRVymI+9RrESwO5P911RhkJfY+I0g3C6EuoDJnR348iAGWCgWy
rRk+jXn3glEE/ImVLPGWN5nOrcgyvHPjgDQ30BKYMIANeZYEa3z0+le5lmNJfhd5
Md+oYL1BAdo5pR22YdMg6tVUfaebGD2t0NvM0PNIILqfQmDXK3Q9YpwZM8c+gMD1
fk9UsLWj2IInZCsoKm3HkkqNBj0PTlRsjqZogmA/GO993qbDJRiL4+Q+/DDwLLWD
sWhbT9aJbg0wdPL2iH4MyQ1+JiUcAzO2uZRuvCU8DEFuPF03TvT9+8jIzcDSqS4F
plqoTbHIYargZ2lRyP30pUafOZAK4fMYJ33LD/5tJitjSBv0fWBuhJrGtWN8TQbo
qK4kjgYVbF5exuZoeeQD/c1d/y40gd2KK59K7DSDFTS+KLE6MokWC9Ix3TxRG1uU
8IqHxSr74epQ+OHR+jAcu+NPbgVEAvm1Ir+rK7O5sV8QXuKEoU3H6Nf8tUKqNkqG
qG3MEszLmdmvIPDVnB2cQMNQ652WIGCUKSFKrH64wyEijow0w1Cok5HLQCWvaR1W
0e2+lg49R89ilbOsEdbY1TW5KsGYyjSp52OuqSn3SLaC0S5WLDSiUuTJqHPsG4V7
4H62ImAC6rFFQC6k0kav+oEfoLxVjo5L+hyOjcwXVHNPBcH80nliQOEch2lNwQye
AX+l3RBIVDh9B6xlQA+4KluNWCnLf+uDMYD0/DE3JzK7/IqqXxNBUET43G7Qxn3X
WmCqPRvpOejgBoXgwgPwuGfwXNL4BZUoWWvo9eQsq2tXf2JNuKdtpFJaED7UgImG
1aBuNV2GNkOJ23NAjAyiuTBpRQxthF5YeCCwZPjjNEtMRCiuR3xacehjEoTE65jb
7najth9ivNbwkJZY0iOITZV8hwg5q3GiUOUc3bpCELIEz2wMLiKVeY85W2cwKgLb
ER+AJqoepWhSAdRbBsySA98TI5WiDUrLDdmGrKA6kHm3KzCy+cASnzRj6CGGFVu0
CCcIrvjmqiedcGDczaoxHUdYOBWIjujaU9nPaQtkCWqbhB/qY6/KpXZQntq+XUsb
/uWr3ak2JwparC3USjluJTwoZAh/bCKXMiPrG2p5qk6fDQsLKfKp9OMKpytuQlXh
WcY/BOQpC4Z1Wr3Fsi3xzhQdDZyRc+fV/u3UUq/IKSBqoln0k9v3BOdxJGMdWZSD
imXP9oS/7nLS85w4uunb8ix1Wcd1tDLb3RH01pLt6EIaTaRoqxTwJkt2FMRFumLM
10N/ekbauTI6FoKoDD9qmY6CQiT49KTvYzVNwB9HAr3qMXJYcCo6lNdbEWTSgCyo
LGU+PX2TZqtyUE+3X7we/2jinE8a+/es3v7lAWWZ9ywl960dMhNYnjUE0MrYaTeG
35xJi6Td4Y3KTnTvKmIgtHM8hv+EUCKknj5qRc4Eyh7k9PKUlRx8E6ma5M5tl5oI
4VqP2xuSKfndvGrtDGVo/4nqNLZAFKqVNLpdRroO1CB/KtCbglYUIwt1+fP/4zef
1Eu4hIlt08PA7RzMYMEsMnlNcCpuf57RQtCFOmzH7Cu8OIV58Nfp6ZiO27kDBred
oQBwZbww9wWNDUUniHc1vB9fV+8qJA4vGv59jeXgJ7QjpvIMAoDc9gcKe4mgMVSe
Vqbh+hck4REGC8CoZV9B+xL2Q4xqQGFnBE3+Xm8tPfR0stGY8Un6w2DzdKbZsdCg
konNBBj+FY8ivukCkL62UvQ8osVrW90p3HFB8FEjlxPegn+sicC3E2ot2YzPtW57
wL1E53WTRnfHaeH5CjByPEPPlHSLALbNlAsfYfu3G026TrffdUb7r8Z1ukMfNDGb
K3mN3CzM8eICW/2oqrS6NmTIa7jpVnJ9ni5LfhURP8Kqj9lMXJCPm45xW1NxUWKw
nqnr6T0YJzAtM3oEJ6JyufHjTgGUcxZqoWc/PORLA7hAQ8XJqCCnUoGBr7O7Ddns
IQTYKXCwYSVRHBWHjP2jb9lCR5+spHyqCdBWfy7yVZKvAXX7wcwL6jFjRmpAw/Qy
zPqv0Zx6MOwed4wdD1ndiY6dlQLSATqyE41ha5kv6IxCevwyb1WqZ1T4Tsix4Nai
9KhBUAcIhHczoagRMrL2CotgkuZPJ8FBEXJQ5UHcLf9rD4XECjW3SksJkwm4NaFV
YlqOh0Yxiq6H1BjhH+uct3XlnHMeS1Le6LwXqkWToOrAAjIcKZ83Ks1keF6RaMnO
42w+b9K7eEYGet+5oSbjzJuI/aCJFG7ZeQZ5RGXi0x00Ar70CVuNBmUmaq9Idaq8
PP/NaH1z7GObhcpWI9L6IhQbNgZ2emJYfK8CdVvxoGOGsfJlrtFY8p7IIoTZeI5m
P4eyyVsoIRPrvtR7iJAaFe/RrYrJVUIPtwJTmrxsUbaK5M9HdN2gOkguA/dwD855
tmfXfEerNzdNK1bfxu7FkYOzjWChheIbWN5y/4uq/ythnQwU+HvbS7SN2dZF6baP
OxDw6ll+HZCsXhcu8aSSxa8n96c3Yu1CE7L15k1Td0GxsnSmNzZNXTloFh9zpqJx
s4w9e/DMmXeok4SqU5NFrZKCxP3ANmJbJB6q8T/e/G3mlO8JEKYKm5o0QSdyuCpr
9WU+DGInpykigcVat59RWHWC+FBw6jYx9PYLN3jS9Hhz/3R1lota27XWXkHnT1z+
kQ53dIVevvUOV9ft7K4ojBtP/gu0gwDCSLR9I4On7c5bp5esokgdoS1JNJ0rsHVx
gJCBiBOx+fkDBleS0CPRGwsXELTCIkpyPUww3vP/NoHR1aLq0vPVQsH2bQwnFDiS
lYkr0oVdZl+E7FWemtt8jY2aVLmEpHav+XXBxWuEP5mkE+TTJ4rpK52ei7FCjs8u
brpK4xS61AtZNQqpGRFSamVqXNGRlijsXchmmfvy/i/+fgkEj64i0CWHeqthLihq
pLR480vAs6xe7P4z7Nf6+vXfdIBRvN7y2x1Tlavg5kcCQ3vCB/emuVOontiPALUg
LxnQajIQRqRo9j7vA8DnpLRDZXKjirgzuS8qMYSY1EOJ8GDEmLecMYFwo3mcfMBU
aLFHCT7FumG4mH62N6Bt1YLw7xkNOMAS1soTMZEKuv1HH96nkhQiv4uLpkuOnrL4
kGMt6kCPK/T8tHRtfzGvIgic3SoRlQNS9EhFiGl3AWWioDw2Xy/ZlJMYU7JupaFL
hcR4f2n7+sD08+YU+GS52ywSEI56/vXcrFzUqYZjoMEmQHgtS1Gw7jDJGD4MG68B
EXZcEjRxdmolk0GDGRhUBnfEj23/x5OQkHkC9B9CszvBuQoXQzFZ59QFBJWtTwMx
nJJkXcb3CrZ8t4CWB1VPIGmOBKX5LyCNYNLPSxiObtRYvJz62zJV3UwirfXeof+A
o4/R0Nf2i7Ldl71J4mLZEMwbdkvYKjYJqnIlpJu2G0/k/427ICWx/LtsBr9MMYxb
cxZ59UvW+V7hqbaNvZvpKdFrXIB2Ua0xC6q7i1n/ALZPZHLo7E8ckFvH149hz1VB
m16Buf9Ene4AS6TjdTjoa6lhtb5ahaTIkGH1YHLY8MKOjQX3GcoA89b3BHyNGRP0
3hJwB0C+kc1+hLgmVf8XF8GUBdQgjqMnyQ1QdtsZ+MWUL35Gv9e9mXbfB4ZCVMwH
3NzFSvOTwHzjYEIAaLz/UECdQTt88UbPjsGyNiA3kS1LjH3/8qVONABmlN1vvPdt
8XedZCeJrrLrvRYWHTsXCJaGMfvU5Cu/f25P9wHMCAiNU2YiA4Y1yuoOprVH8OEH
zuAnf/+Rzbh4l/4Xymp5YVLSZmeqPTibaHqGEUK/IgPEM72cCHPgH6C2NtM4b/Wi
NV2vmOYWw2L0xt/5aqGM6witAujhwrwvpk4ml82rIto6tIsMg7EG7G8YUDxClPfi
RnF9BEa2A8C73k58g86C7YPaq9H5T2MvfhpoB0h2j8Gxb5HXVcdAL9ozxtvxb3Cc
iPAtXoHPI6XES/vgv01zVRWLFT2AQM/Ox5ICqBcXPDEljrceRcMTbp5gLZO6drXl
PdqjbiYtQzDJUdu22RhHbYJQP3Lvq/4Y2/N+1RWSelFS2PV1aHcBCSZUhWeIE5p3
bXVYOzqT233kPvZfyFcIiCEwhL8lEhZ8b09s9VE9rgC3mvevS1dV7da/pvRBt61n
Ht/BRx+kc9vduPs5fCFj0SRkcU6Z1Y8SnSD3cdCVmy18rG0aNZzZJY2OSLLY9NvC
PR/xWekc3cTiMifXAdecJNgqylCh1yzxCecOyNU/mLETikfcfm6Zc88FnYi3uUER
IaIbMDlofRO0PSzLaRbA00cCdogCXnPE80Np59AF4qYcmReY5hfOhlQuCJ+P26UJ
1/SY7t1O/jxl6bJsffWLKJC1bbUWcYlYZ99nBRx4XoPZbTINKizHtzZ5NiLze/UQ
CEmcsNXQ9spssFI2DSTCwpzCMSktRtP8BRuzZBGjnM9IU4z4aPvY3XWOrT850Y01
GvH4oYReLyiGhP8VG1qJolDSOlB+VACRCJrI387DrJ7oTjNMFYALrvfMNFaQ0a8B
38cdPKlCFta2xlEFWPgkaZsCPVRlQfTzpewahFK3FKtyJsYYiRyXLt1IDQvt9Lfl
HvmkrYM1S2JjL9PXLKqAkgsxxJkxPcQEKKk6N8aBxWpUmdzUHODE5kOrBf05SyR2
vkNTmv9sMaCz7zwJR4lmPNrl1pQwkm/IVFMeWY/hBM2vUzXIRaIu+qShbgmrK9Ll
mQitzNs2RTGkKOu7cWt5D1rbdB76O55rhJJ89t7MQVL2K5r3gBOxGOpoZySYYWzS
rsv9ZSbK+zbRoUa8FYyGiz3hsADNUxwVPaYGJ/A5KD1ZCYCsYOztsFyZMIhDIldD
7mkqSaOhOET+wuyJJywQjDw8iwegRD6DVhM4vS+Icd94b8i5DoQUOIVIjlNik9Ui
/Wqn1vlXJIMRwPmLGQegmaofghK1PeH0eMdmecPlDHHJno9Bck0Ovx6Ue71jkg5r
sySU0NXJypxUm89BnxjlnkIvgTHGHcOxo7Nkq20AfxVVkdwYoRASBFoN+yGNfKLr
7cn9miS1rR9o/BW2UTxZolzY5VBTXnFybSZU6haGHi5cBv06wRIdcg3bKWIPLspU
sd1p5QNFyk3KVn2ZDbguJu9Cvrx6jU9sl6Xeej7FLUHlupS2vyW7xPiLi8C7sezK
MTWcC8768NQsR3k0TQdcshTPOQR3WGfOV+kPg+/WyuflmLXm25PMw/bHAIf6l5W1
ALPo+exT1ErKI6FBZIziaV9xN5cSTTvA+Zpr/NnKsl0IwDQtCbnlpmBwMztjEaGv
EAXL8xsSowZ06zUUU3GtgBFdtBmOQyO0MpPMnS6B1yclf48MWK9b4Ps+AYQUIvrv
aPIlPv57eZDEQ6J9esOwjbG8/rt/e2UXqCW45/ua7OFYJHnjWlu9iJT4LVtqIvYg
3sx+PoLA6bCfP0yNf48j0gvI1fEHjolU8qs9Yjs9BeVk844FIK8/lCZGN0iqLkuh
Fl/jAkDwcLjFuZU0o2RIoZLHPwGAmtxL5tO92NQHCC3pXiQYYP4Ccbnuytz3JFB8
M6S19hsY7BE5vNxgUFTOMQXOGsgqhaS6s7zENKT7hwBO9VrQJiBhke9xrnCMemfC
c+AENJhS88sEPj0s+svNyQmLdNiR1UePHSW24/no9KXshWI030cmJt/2Q/F0FcYO
0LdHfkpxsviYcTTKLNUcc7cqC7uRRzzBq5qeU8F0T/tkaEbJHPqw+4XzwDZtXhsv
Geblm+V4jBw17NeUYYFRlhG544DP0MHDjWG4Ym2mzgKlEjt6vZIlBN7wUHKfKP1z
W2Abt3cZVcsWipikYPSFpqg5zw/qDkNvQdh/h84ZiWggiBXUpWSsbJthQz76tBSk
fBgg0rSQ/csjVInUK9ZoRTfLaorD2Uyh0d64KsiqDUFrzVnKW6JWFVGeocd4/C6i
XjB8WODtpcvZipA5BDPy9/xvR36GsajOVfsE3d8w5YKn11anEUMu7cjPVN/iS3+s
EURiz1/rVPqaMkynDqsCEZcQtbmRVWbP3zLceKQwC0MEkZOe8K3UebbkrAIRGGLZ
cxj3X/VlpLCQU5MZiemN/wJWhcYbCcn4QWJaoVZlGQfznbind/jXkP92G/ez9mAU
LS97mXaQzIOgHRndZMQCuMUOy9H8EOlsmE8HoiEw9CcKUx61c3Fp6F14uiV8S7GC
vfAh4ppQxqIRDrnjxqhTz6t11YSrMzeZl6tFd7F7PYP6uh9qGs9SNJUICKnzM57f
sDY5Opmi6U1q2yu9xjIRGeLC8b1fmQEaJsmVg1hCk7Yx//Jqw94mb22qMKMsWht5
CRJd7iIr5m8zWLNvF7V44vQUYUWX/6Pf1udQVxMDTfH+LYOcwxx4FCw8UoanOda+
qe6TUyPGxndQYYjckBYUsLsb89rgvO6eD2wF5SdQTm72FjRuvGYudM0px1yTU8/c
2TED1xF6xpV6fgkosjUWpUJCX7SQH5HJQtngakvCqHMpLHThL3pzXyrIJTTNd5DH
L26IIPojlFkQW5NAi+m7Tzof2B8Vq+Iq4SXPpPDFMAeIritO5Gp/UqqYJWiFThTO
cgzUKZ+aeafqmPbhsG254HViIAd4X6eWCqVG/czo/5sll3QgsoC0EB8zkDJhIQ9H
w2mtkBaCOA+iBKPH6Kp4Y4w5PxtC5NQWZ4EmRlkNorJGbNkMZlWjXqugnVpVM4kp
aSa1R2z4SMJkIvMaJjP8c9W/NYXfvdaPzpKTYQHJ2DLr5NHRnrTP1P06VlSOXf+f
HPB/qBrIPxDMKzPgdpLklP8V+GRCQ5WWfeFcDFxuuxh/PFGdTzQJDN77SbXx7KKE
4Nj3pOiCSGLyO3kRQ7yCE6uEFWFok+9DS9Pq63pIXZiJK2B20s4JFH5dXTkZV/H7
5nyI4O8+1wGDUHtAhDzyEeGSzt/U/AT3H9EpzdZM0I/Dww3lb68QGr/U73qOp+Tb
JYwoGN0OpFv/jiV7c3Gn6AmOacPGbftpGod7e+UkEkhhrL2RbABb7Z254x+r+WGt
AsjwH+BQRtoQbvdHZXaqruMy/0fjMBwrLjjqtLGllCyTy0CFRJzPLOHNLtxySlNg
vvLiC19P5KCapVZZEb/3cIY11BXVy+xaooxm0vDzNQDXIwmacA8AI0v0V6T5ZCQP
Z5pJYISw1OtlQRxt81m3qjfHZNrEmAl1Kbzbc+6qhThopAKs2vHEyfBmUgA/iQrR
jJv7k15FMlGRfd3U0fl5MJiOeVxqhvEkGGjvfZlF6hxCSCXMoDDjQAZeA2IKFYwm
AAP7b7Ln7ZXqfAWKpnkJdmWGmFG4j/2LFuB/th3rHuufDenpJEvlom5qbj4fppNk
wLKy1iqG92aH6SF/ryvxkyzDZDiaRwngAYZQQDC8LExwPVuaN7LNUx9PGu0TioMU
iEAPE8IPEIdqXTniOIsAD2hE5Cy+go6L4HhsPhIvZuIv53ho/F4SdK+yEQ7ZHRsD
uL1o8Z8EpJ6P118GiAoumX8+veAQLfkHXVIQRdvKOs5c9BjJu8vRrjIonLZoz5Cv
s3Ht0r+5zqoR6KYSd0ey6A1uYXW7UHzASB2/I/Fcberhjne3T/DCUDLaNveqb3ur
Yg2zoY2d/lxeEFEoLur8fnQ+9s+fuLnKThJInTSr8gXMhRGv/XrL1SZRnxD1Tux+
VRCZX2koJ94ig9Jzsr9emmeO8DkObi+8hjl09avkL7enrRF1YmFQ2WXimDCt4FTk
qxsSP3+EmItlUlprQBae6Z50V45SwMr+imydo21FiIc7OiXVVGlHbPSv5gFYLF2P
dYnbuPaqsy/ZQ18/pNiJYxJkiDTeZRCxMCaTMHp/7NRXNhEUrVv1GiY9R5rXT7vK
cfq6nXHcDMriZxLoAJts9JxfbZ0/dEVax0PLqf0Gt7bNA+aWFU+4l+K0bxy3s6mu
R1Et9HK8Hk/jF2rGDj+CScqhe8KfTyG0pZFZuoxmjUg4UyIwkAZ9djA6I03tpiHO
oEgf1yzfhKSDcqsnaingGv/65RJLPlKrihkOOQS+kscGEIDNlRn/cPanvudQBTeL
+48Usk+hy3l2COkF6tBksYWvppXtjsdvlKirkNdlxiamHmDtVHgbD8rSSATFH99R
s0JKVKhU7AeMiE0Vga5LyUu9X8gbvcp2v6DYpoT57Ub9yErC3Nk5KWnd8mXG8y3Y
LyAMvjva420KBwQk04Mk4M3rJDsyb9X4MT9QTrc/0tivoyS5oOsMc3ZEn0PydC4M
XozqSyUNH8+XeV5H58LbH0XcHIti1af4fyJGqCwA94vOMxDxHNNUmAqM3nqfYim0
y3t7BQJW7U4XmK4MkRueW4zztQLtWsZNOUI5f9vz1qB1dCTBV7FrylDht/6zTrji
rMUiHIZJALgfof934d5i7DFFq5RUmCOhalZj8q0jJmjEHMOa7AcR1rgvcIlxZbww
C37T1HLo5xED9G+sGBk3nG42WabGfNejMNt/dcu/PpluA13LY2tDcHsbTbT2ZYC2
4ooK8P5BWM8HYNupaoStc27ou8ceVQVyQlRxkfYTMzQySW7Vcek1oU2I+MspKXZL
P5CusccEluQIUqEA2QC4npEXxAXeigUNV+Jlxmci5rsQNfWpo6Te8BrvxgjvYwQP
dvez47Gc2RxA56QUFPiszwDPbdtTY1jZrQc8EmAsXPYfimRYvdCvu65JKqVJXf3r
/gaenYo100ZmDqBYdKGUPcPhEqUX+zubSISJ3aGCQ8oA4EN6o7y24ml4EZb2q5el
UDk38oWRfTHqHsU6yMoMqAq30ZvfFVvd49GOWRaBkDJZbyPPBRnkbOMnkHjhTnlz
tuW+woE5D1vG4rFUKnmEY7+qsylP1CFAHL7/6qEajsf3Dj6x7kfMGZBqYw/z50po
55RRS5tYo9I7Te4rFXtu6DB9Rs2jvKKLIF5pNG+5SR5HH5EcYDiLOr7+zTBQJy7I
cH2Kit1xwslsOVUy5xeVPrf183elH4oQkPnZ1Q8v4SZofChVM1A0MdMbwE4qB/Zi
P7GrIOYgx10dZb88LiSUgKZ2Ye9u5jgArhgKs8c5i3ay9Lr1qj/bUFRc502cpcW5
KsaHMc1JFk34GWaU4HttnfaSob7ol9E6wrYHHmYF5t/RfBuT3+gTHCSztKSofPLI
BllEzehnac0uIPg/u49Pp2vve0YQPROoWUiCi/T4er2noAin3x8JJet3bQKAIZDU
p+WGLM21JV/04x3KW02FGd7t6/buGfvROY6muIND2wQP/+PiyB5588pHKML5z6ZH
r/AwVW9zVDFInrSQAOMV2DapmndiKVPH0CE6DYauUHAqtNde7y6vMKp+7zimZiEm
CoBxY3IzVvoRUU/76+pjkbdTFPamH/LnHl7vEFNA1+lNmGq2suNtmsJTZgiMzX2I
5xA6l2Hq2IFW4dDMitOvJkDehsNcAV4LRmt7kMJ0MFjnk7GHr0iC7Z2fMQjgOqlc
Sby45n0QVqeP9cSUS3+QjcKEfaNfs/OrdmovkO3vWIbNhO+dO+qFl/MHTv9On/Qk
2U/NEhMk9ligT9CraeoVv8fi43LdUw5IUbeHiR6qp5M4KEPOYFapJSg2ukflD1EJ
igmlfz6kEmDUMR48Tap6mP92NxkQOuJfe6tUbocnLH9/5+8o37dF33oQC+dSasJq
LSydCKow5Y6JXt+j/AxLkKbPNmp149DOJ8kH0zxLtZsE1PlDwfToBGcR3R3WW1jr
KomCEoZBGJcacqkd+ylZbV6aGDj5RRFt7RvHWp0I5m2X3rRob8upxSWAnc7sY3wt
dAHC33idhZTydNNz2OOeg75u7WbSkZI4+yTJrCab1serSLrAREZw9lHF+Voa+d1e
3lj6Bmsl07naYJfDyfOXBAFoIj/LYtTJRPvPq5B9bDgDbxlF5rrTqEyq4hxVv2wO
k6JDKBrAIcSpin84N+dKT57wc4ZXdeHDoLeS3kB6ehsUQbdQLYdEHrQS7nXdQSJp
BF3kwAMblKi5umFEtFuvhOdS7E1689npry2KRlV/y60TpyaRfL+9D4ZeNJclowrc
BzYLmO74Osd1WlhQp39orbIAJuPDYfVnh9X54VJR3kacPx2JaeLwLgk7b/li3l2e
B8UXntpqwy1mgVX1e3yAT8UHyW1VFqGc+BM+o13kp1trTSY9XS8uNVMwOg2AqWy9
M64utYLG3MVPftL9kN0HHIpBruwFeHz4ba3d4XHGo4c/ANNxunu20BHN7nyVEK7z
RjZhOHsu2Y1jPWSQb4IbkDGXlZ8FJgTL4xUxxopcPLNeITMSCaTYBkLdGXygE26C
Hm2O1WYtmYiqTSZubbNgX20GNj2tsdS3S1RFpBiOW2yOInUYub5Ut4ork79+ovXp
jFIDMUpvhNs2X4OfyKPOtQ7VdkBAuaRFwthpeQwf/g3DfXKD3jYVUAjBVKEYqi8P
ODgV5sljEwJhx6xOu2mkIfmPtBK2bDOj8aia+3GsblJR31wUkCbMFlvIh/Kl0/0S
dJud00mdJg5Tx40cAxmAC74H7mD0EF5qgaILptvvocpL4VPdfQGL054JFDBlMPcp
QzrvDKhhqkGfdUFX92r9x6fd5B1T3r7onOOfCWoZbB2Asiu0SALUbH3tQ8iYuLDf
WwjyIWY/jO7cGqbB8NYhD0lG70f6EDLEWGQYYMppGAw3RfkA12vxUf6vWAgItAyl
arWI5bfYc6zKWqFRTcs7nskb/2NE5fwLObLqPwrW+7m3jy7NIop/xUZQ2rLws/YH
ytoF88W7TO7kOVEysyagmS1xa6ZOFUbzhCiijsGGAbaxKh57f+v8nzlgW+J8T/FF
AZZ7ih9882Ahx5DRC3Eilr9SiCb/s4jR67Ew6QrDGr3FoOQjzU9uUiZN/rv9Z1ca
qgTTQ7qHwv0h5vsZ40e/eAbrX1hR6YuPyVHaTBOWDZx4la3jGwsj+v18YlmxlYVX
tK7iNUr5jM8JMvaeDReXD9cdOfVsCCcX/v43KBADO3EW9mHcFQwkr3vmge2a7x+3
pyQ6qa52JIeJQ1DDZ/RHYJqVZW8d3B+8X0Crv4Ya/9wICo83rjnG/NvddfQ4JQ9W
+ZzS+uUUErq1zljiWnBItPwYabywjBXn94qE7SidzbQj42xJfHRkW0zIfX3ojhzQ
v0PBY7vGo9qUFHoXMOGP9pW0UGRFabWjuN5DPUO69p0Utpiu7kY+g8jfNhZ58Ry0
dqhN7olzlHTdryUdZwddLx8znwlYB8MV5DUaNazc6LSb4GqvkwRzitEWx0g1z0eT
OjFhf0806WUqHwF3rZegctOPyKsT2P0IXgOUb1UasHpa17PzseM7DP2c4cW9QA7B
EQ+REPpqMmDe6amPeP/0fb82Bav7QlxomVAoBMEelgFXyXxTkowpAdRGCbqdI1h3
41viyxq9Vg4mXV2HTjeitU6Xsnm7BdWzIL01Lw8FjWzlZqznLuIUv/GDMvCFqA1c
7WnoRgpAaihrHNZ6cD63pNqLNP3AQ4uOvLoy2TvwUPFG9I9joGLwQ7EU4tQEfWOg
GPWlgDF4SzHOUurRuz/8SwPFiVZT32juDyEiLfnVcS5EYRJP1TJ9pnzFpUPE5r50
4m+JB0mvj7IK9zCoSsC2QGOaJobEAHhltxarfu6fLwbXvCkJopxwj3wxoBT+DUys
fpzfy0TF1Cw14Mcr7zN5lywl5SdJYhva782FqFaxfFWaZ+wq63tDyekkXwFTn4W4
DZjAQF7r1WNEDRo8OwMUO8mGO9lJePpQslLgyetJK6vRv0EE2T15RXISjWYA+viE
Tmn9af6EjmZqna6GejRrsnyXbTaZKC/gxZPYniOWSx1MuIAClw71XYPS80VfamV/
kMSicveZ447wsAmuTZrxOc8OlkWg6kAdiBwLVFidNq6kOrym3xV/ChfOQKQSchdE
JJrviYS+d8fSmopN76wsoVkapx0lpHwrQ5PwWvzsBK2nKUzw5cC79loE0DTBU9+m
LDSPZ2x58gFHtxOLYpdRUzDY8TBaZUg/PkfIe2ay1v7VbLtCA0mk005nSeWa+XWk
E+AIM6hwKAnnJFGF0yz4+BkuNKWaP4Zz5Zve8oRItQYwkeiuvjL/iZuA1xSgL0Ay
Rbzh9XmwmPHyO3AQFKZbFyXCB2NXZmCya/y7hl5hjAp9YBOWWcknFjiBOtwcWXIh
JmF1Fd4nM1KZr1f4mnaVJY4p67SkIkQzIi5DC6AcDeWVaFPo7Q59IcuL+/dg+884
kYWa/CltTayA1QojPD6n2CcGsvSo+wfiuTTfW2owli3D5UcZHbBao3jEgN1ohIaO
H/rJ0cZTryEwpCE34aTN7o+UPZVlN/od+jEITA5cZbK1tBmrlveHP3Iz70juzf6B
/JOjYkVeG046wlD9jnNwV5Du2UwrY7GGuf3UqMibhAREabrU2BRB+FMab++ppP4X
28VegSemjIQyftVocIZGjy0BDK1PJrY9KOCLiLzOQ7Y3+vl808yn3pp25e5vz0eQ
VVUwfo01Nzv2lHh/7lltWOdy2i1suo7fwt+nfMrpPzA6TfSYDSVsIR+0A2wq3giy
VS+lfUm7sScn0G4xlG3czGRfSXRgyTejKEOu9buXXqtlvaAZqM3LO+fPYjyoMjZf
dcgGb1ex56C0HdHeHF2Fbh6PksQpAYEjwSxov9TxJCW79+u2BLA3prpz/pKMJ4n2
pcXualV67u17rkHB7nnPKUq5dGQiwmrJaVxHdTfFzdaWZx7eqkK8/83Hj6laUgsJ
UWdKx3GcdB9zo1U1yDf8i3grQqYdLzWgYwQWpBzX0e7/kC6pr8RxJ+RI6E0+OYWH
HPEwGvBLi8K2t2x72j9FcOvPxRwuKjO3hVy4cfpXXzSxyXmwTRwhFrZ6VT83qB/h
fUiNgE4/MzSRmlvOBdLI0SycpWWqquHX4WiDww8UcuQ91FEoD9+1DbDwLdfXBFCn
V6ej2PwADWv99QnZ5hKTz3Kp0mwcVxh8SiB65oLOZk777yWnJUAy83DT3G9HYLZ2
C432mL5vb+UGn4YtZdoE0pHtqX/mOizuue6RGxMC304john75kL8dZf0BLsvq+H9
tJxlskbI2LADI0ieqxRW79rfpDvFLSAQ7xWQ7DLT8pXbYxmFRUoZguVjQ2obEv4a
klARaDq3o8vL2rV2F//iZyu6VX3sYC8o33HaszIBru7fufgMzdXKHA9FLgdt88vI
hmGccYdEKqHQJ9Mt0P42nDobthQHGfnu1cSiK5NchB5DzEteRtfNVji20y05N3sB
YrZYs66e9DWJaaHb4KNhueWZ0RjtNCmZ17TISVMxQXMNuVj2QXrLK+2dR7mrbi40
fslQEJ1uq7FnWc3NhiywhVVx2a+FsI+EqACIh67VWwm/ZCxEN+GFw2W/lEj4H8Rq
i8ubTV2UxsHRmv9bY7JHoai84ZmxhpNLcyHUZCDL7UiI7/dHw2fq6TTBRc4XpXk3
dh+SbCGCCuAtnbS47vsyX5gr6LP9dbvuPaSREzaCJT07Hih+jWY3mGQfe7l5sEbf
aEYGx3jhW7fybcA6fHWpC+esvxsIUIlDt54Y1E3qWJ8LnHPIy5mWesHOjc/4RDbR
YwFolQKfX+GMpA3go4B5BGQ65HjQMoDV9U79U4vgkKkABunCb5Tt6xnBQ4cCWtOj
CHKa3IJAj9FeUet3Cy7ByJigrERjm9RsGlquxdqgZeWcpBOWF56qDkywYKnSeLrR
s+uleof9q+2/E+lTTmYxWYANVeucu8+1MYX1OLJvVSrXKxCn/5/BoujhtlFXcyD0
2sEuL6Budhl0enf0E78dBTxgyPt6Ac5klZAVkbynMHUS6bYiNt3tl8sigG5FFJ2k
Hq41MpsqPPY/cbrM9EUwZNYrSrQwEDETMSj3cug5bMEaziEWa79CLg5hxEUiC+19
LGLVxA502kGDY1kz4rtUuY/qZqk4X2PVavQvBSZi60zLlQODnGeCBVcS6k2uUHnb
m91MB9O2zP+evtZxGIB0al88kVDGimIEfpKjwdVAe7qMKtEwAwMZFSn/3kbvvT2C
Ju0tE1Qpm6PujKTk/Wf3uNhdy24QQx4cCYQwFmcPU0HQ4vmfVtXt/v566URgxWf3
4R40Ozhnwa83Q/UrIIQrL4P+WLtupTzNgFDDtRpWzccFYo5w6kxdesy8f5k17Tzv
+ds3EAcvRZcWfTgDdBPqHAElMyPwNVLa2zgwJ83Tr84hYJYOEZhXXu18M18/GiHj
BPcp01/10iNrO2lNy55Y3Q8C6WW5WirciU7T08dj1Zc+eX/6jUcm5FQFE9PqYW8G
PHsZGKBMq/i0n/Tvcw3V3c3iAbiN4WLFdiT/toWDRY8ZaZ2GUsalMUGcqb12IZbq
8nIwKvVFPNl9EvQY63EokuOtV5QbRmCq/MPptJc9FEeyLr/YEHt0t0r4wQz37inh
SNDD/LLQGYl4KiDyI6QZlXqWVC/UlVo9XK2U+73uLL5YuWiqjExei5I2wDnO25mS
VYD3hJcx6vGTtLdQECImMX8ufTuQe7F9pE8/weOj8soqn1XzsTa+HergBmjvtGzL
BgWo+WyyglR2hk9YERpmKuBJrZG/tyi8YsrCR+uS2G/4nNmnlnyGF9RSac3MJyt2
QLeGz/6P8GPoaZR6BkGNovw66z9LsVMzUP1I/WazaL1ih5rx3gm+AfFrNqBjOKpF
EREQUE+LcrWFKRE0VuKiZe4H4vT5tj1pOUWOdGGCv6bt8uLwOZz16xGxZiAPnzCZ
O7SINhSDWqRyZJFF9sYThpAuaY/cxa/I1wV8xvmqGa+MXLDLEoGABTThzXMoeU7J
VScBe/TzIyoGocTvedqHH08lA244Z+eehSqrqwo/yFsSrwjBXt3V85kTz3fpoGfL
CcOIWjqtqnei3O7+SjRX47Erk1QsFtUU2U5TttHHmLxFhsdPcf0h7G0mA4jlbNyj
CtPm/62z5qKbGvt4JyyRbxYKA56HL+uadsxoLEUd/8nrII7p1cSPkKwhr0xkb7Fk
C25LGgMI6dS3KnZwvIdFd/I3VHANSeqjHIWjIj5zWiYsZSTb1ibHHa3HWrA9Nc5/
TbTS+hYgTYlruq24WAidIss9lZwl8qiMWyvFbuxzgxp4aXLstHnH2b4oMy42EHbo
td0+mdTZ6tpE0FvuYuDiK5t6/QTzSAyjztQZ4WHC1jRQMpzayP3BI+rllMcbcNP5
Bc12ekkbO4LrxBdj+remCB4P6cJlmhsmjoXUwWD5Mv4TXq0xWozYBtr6yCLHYNzm
81oVvMn77+KPMb6joH8lyNZ7nLg0+fQ5vLALDJa9N8Pd5EZDbEN6BqyRBImLhH0f
izaVCFvcusTsnesCag8fOSgUsXPH9aT+i44Mt6UY8Bq7rzjQF3MwNtmVqHxCN6Kw
MUGEjAXl3ybzgg/ev5+ebgrkMHSvosWIHL8f21L4pd1g8KIPBHXdNOoKm0vXbCFa
2rBphBkhsMUviy64FKbSsEZ7O92nLmBxzw4olemNMG+qAnZ1cB8QtOp5gbbheTOH
PWPRgSB/4oxBRcD/vseLNDOE1dg0v4Ch81JmGgi6UcIQH/s4IUgteZ9CGay9LhMd
Gsv3+BccU8GSNqqyWPJvuOwXN+QyAF4pJ+ozRD2Ag5Ih9upsMkLwIrLn5Bu2cICK
0PfXA7+AVCvUoGY8UByILZef6CzGJAm3azP3DEWeF89WewyOk+AWF9RJszbJzxnV
zDRywBWAtA+BrHQhHCsxmcmU5FZEn6UF8nkbXn5a15sWADqjLQP2NjlTpM/3xale
aq9c3aTGqvyesP5OPnnWD0ub5NywqkQIqN3YGWNlDsWA3M4a+2Rb5MIEgnf+Bshi
iZeSzFrWEMiHE7UHjLkS8Qgc2eI7wF0K0fU+RX9jeNc/sesA5zJvvgRrgOoJEHR1
ljafgZZN7VfSORcCTJnBn7sP/rCm1OGJa320qPO1qR6oNx6+6zv7+lbel2ve+Y+c
U6bmo7B0VWCk3Vya92HTVtUwGYRg4v2dNLeRW1qwRj6zuO5ah/NKAT3G8bQ13mwJ
2M8yno2TcsKsX6UZAey82o60+ktSq9i0L0NWZFvm5WzufDa4obtiCEGF/6fptWyB
a5KHVAaTj6V5AX9nm+y7KDiiRqhqpIaJFPLNxSkGfDf5WgO4x5WJ03WIrEKMz3Lb
D+N29GUpTbuYQ9CkJxntcHzvsbf+wHNVMr/zuE1xl8Zrw8QXWllfj1TRNNVH/Xbz
tAwKT9+GCEIOR1YErC1GWQfo4YJK1GAL8RVT9CcPv0XlTKEGFSQzhdrx1xdvrq9Z
rWc/TfIE9M0uSP3Aw4TVkVUTOGXfAl9mV4vTdZdRncjiUkyWA7K9tfy/FGUqviw/
AReqwByWiZwjLv9jKW9LKhH601oLUI+VZg5/Y0h5k5P3zLe2W4GiHn08s4+CA5CG
cQeryKcXAKdq9OK+eR3iuN8j17RqVvhgK/GdnEh0zOz+WmWJXAyU621Rf3G9V7Xz
kxijjPB4XxsFLYd5mgp1by+NbAumLuIcUFqBizCw7I/wGv25QEXoWnuseiZfOmvJ
vbE0pE+0VuMLSGtjyzvoL4GyQHhJ7iwzj8wt9FxIRW0Bf8xeiQBgy5UBgrKehpsX
NMnlqwV8mdMfTHx3UVZjC9VAN2bKJZW4zPmPVkEY3g7OUIoyinmIzhUpFlSiBozt
cz3jusx7tcHU0fz0bBpsYxsQTaI30aB+cunsMATlpyTPLfbbYm1EIHGeMu+jiPOf
irQ9ZQnkGX3gbMs34EL7v7bGkKg8gR9VLkRhn1fvIr0CiPZeLaAC8X816iiO/Uey
8sXHVkTw9BU/jOTC7ddEiq4hvl1/2A+6RAh+1UR1PJtx1kOdIA9TedhovbkPsQUe
oVviLTUyKH0d7d5Znc4uJQSV+jAq/HyVufITaN69UWik4d/omGdTInBHK3dp86eE
32sbXINxvJ92GXOT1Wl568v5Hl7hNzI8wG1ipLKYsu4wa2HlT153xIbUZN6ZlczZ
ODpievqkVca7tFyNiMcIHpLOGszYlFcD5eYra+LPixAVwPqsTme0kOjR3rzu6VgB
LJP5E+BWcZoHYuAJHrekrbEzFJa+fJVTVg35ZeK+/IUoV7rbl+Ay75lLMZvH/zm5
F2hhTUX9g6ZWERKwjdWfwrlqVlyyt9Q+8yPUjsypONfgHfqm4N5b+giyiV5F71Hc
515SQPj6juSWDM8WX3oOPHU9ha5sVczj8GUGVkbJ18MYFwv+vqB1ZkY1JdUjggTu
WJupS2LHOzVLhOgv0WRhq1q2yafrbn4ynT2OJ+qMCDYXYUpB/ilnmH5iBzeTOxpN
mOgxDZKQ91rkhy2tcN4ZGybadMp9e0yW4fkiK7nl/i0ZXu961qI1sQujP+CZ0CHv
SSZLvJIODkBpFj1Ig0+gemBnMfISECeUYxJpOF/eLcGse/pbfQUOOMbXT9zFGR2y
cznfVl6Odme8ajH3MDwjNTXJr0vPAmDgxa5EUZTYwQqxKY9m4ht21BB5WrA2PdQr
VB6xdtSI5ycPVnnNnNiYbsO5+8cbmQio3+kISP9L0QjUNqoiENzXklhghPwMSvpQ
uomr1y+XhthKy7Y+cLmpfMpMJCJnkGw9r0v7rPBPEkgGR30ZBIBFlbgjRHIlncGa
K7kqjuFQa9OzT+9ZHiO7FsPRxVp/JepUHJDBHYMN4DZu2AKXcCvGeBbkTeVWPEGy
Fp/mNnC1bTTOnFzRLEx/HE8eThF0YwizXPz+qmU/9bIQXgzD8Q3Zf51YfodPBA2K
ZKBBH3+vBeBVVs9zIzJx04yZ+iA5Y5upsNOw4fvttTTL7hnnoqoG/Cnk7lh6mBTU
4y6HRruy5og1v81dM3AVXmeENKZMORTr3ntrb1uIUSXH6UQDHLYCEp3/aalH4K1N
lJLoevpX2lQBHjiof+Og9dJ5QAxE9B3ZDaCwFzCuANuIMPCm1NzW2TQ7wtKTWgQ7
RoHzsDx8ZJOEKrs+qCYJ77nJU1CHbgyKESUISWVAGWADGOXBg/ZV57/eLIRNDeeU
5bydnTFWNl0LvCKy0wm+KaEBLMMiAt1ziso1Qn3PIZADfWkSgV/WxEoQgit+hwYd
qu4HCnruEJBqOE84kAxuW+gAVJcylphgAW2TsX7W8TuIvZrB02bxhx3qdwQPl4N7
BEtbx7H6QqLSTw1BdFo6+2ZN76XrUyfbAcKc0r6FTv+zr+JGKkeLJjXt6errNGPv
dzzX9Va2O/7gFJtVyFBwje8DljIGSnhyKnYT115HqoaJriEWiu6/afymoSqdq8bC
dIfAJWq2kyV8XZVGaTnWOduPfsMJdd7iFjiaPFYUORM997ISuIs1aDfopHSW6jdW
1UnEayLHk8Zt+RWi3zkumHMfkyt8oHdPRle029aXqq6RHm9Las6fye4kugyTv6sB
NK6XMdmDrpaa2ifcYzi1/feteMEEnG9AU6mpclawRMe71u+GRVaBc1FWG5iZW7xC
/Wc6C3zcSZqEp1XhmweKFxgLr7ayYLQz47f5zzge4gwKnU5+eqYEx5vJ//JksaMU
6gv8l5olZtXU2FxjdlTxx4ynwzdQ5roYeTFHhw12kXEGcGLHhQRfol5CQn3tsLj2
J20ZrgVK5cfT1wLmwLSxvhHai09k+Fg2TBcHkHafqUrqG5GqgHnYjwNfN3okusWU
9OpEFFQyH/gXmeFCXkKbYrElAvSOpfnka/4n7TBpN6MeIlYyd62PSaROBWbPR7hO
TnbOjf4UhO3+fG7S76n4O6pKFk2CSCMQ4LpQffPCV2v/k7YTG2UiRoxZS1LF0Dda
4wcFMM6E8oDCYxKDZJny7KZr9nDjvWIMzivsIlRkELbtkAo2lZw5Xnb8j+KzQvKX
RXBaK0J9VgTrdsGz+CXWXocqmQArvDfP2Yo+b6USofLqQExsV1njV2PbzZ2JjUzC
ls69awt99m8uUFEg9ZZvN9Y1HGWxXb466Q20IjWU1PGnk2kCkKjdCgeCUrbKq/L5
kiEOUSFZJ6nJPlY6kWBz5N8Gg6+UwFLdY3yo3qGTdKw9iqNnZTKSzr1gFJ1Qx78N
62HWJrVGoVwdwi1YTyAv1yutejjBH6x4ztjeJl6i9wUaq2PlfIOQAJZye2u98Tpn
kM9tqanbIsWzlWo6JnwRTe2IxuVf/Vjnnyo1VIED5Bzr14JX9U0dq2GvFIl8eQhV
ogARtWMk0sfPMa4EXqTFLN1K+n6rwrBUkok4ub5BfaAlKhID22h9z4TWMQiPqJvP
HnBD5JkvYUjDpy6J5IK6JsxdU77wU5sixuAdBLog3NMg8I5UxmeqMboPVl/7UY4q
EuMJShw4eaaJLjVAerG3YoG4aFpOT/xnUhDOb5cEfIL+u4N9tAhdKAp+EwXa0jQ1
1JGHsukLbyGHFKB53t7Ezg0ZKNuqsvhyDJqWq5FsgjBijIXn8UZBQ+EwxZ7ycmHf
kBDs3J2DuwotPiI8AN/OPLt+w7Jt2Q9V7eR2L+utFVc9trYUYGmUqh/RijbaZWRw
gM+jXAqGtjUPmtpM11o+6iLKy6+q8fVt+CMA1rdz+AWO79R2Ewb2fi53tq9q2dOI
PMjM2WboHyZhtNlpSg1ruKbovoXWl1KbxvcfkvIOG2rzOa0tjd4NBH1mncau+i0D
3gdbzQ+4MNJI7rgHpFMEcE7pnWgnJ5i8+LOUvfEuwpfaEEwby7R47TVX4gtxIFQ3
/ygA8oKlJuQLUUiBf8CJMvuFLZgdGFrHdCWrsdRjUtorjIGtvObZnrLaJaJiISpK
csTvb26CZwb+WlDJm+M9AbxF59Z03WzTtVe5l0dekiIJkCwU9BGBmuP+/4J0KJdq
Or3DcOKlzHPA/yOoDvb3BdW8NukoIj7jLBajHBswjklb0DMCbn/VJsJOToo4Drvl
w3M5qlI9jisfaNbTzM4bY/uzI+UAK5/Dv3/Mli0Mwcf1b0Bw9oawIpIuwDOh+Lfc
HYi4LNDw7hRkaZb6XLuM7ww3lGaK6jJwqQsz5UuTk95BSTwNkg68rO7VCfaIprdv
V+uJiqqI/iigdDhByerzuGS5NNs12PXccCOfBCazfNbvWT4rgTJQ0Az+g0/0bgVS
aKvDLUS1nK3JYbtcbIdiLrIkhvl4dgDFpn/0hE8t2UzCnOwqCOh+WoPa3J33Zr1j
02IcMJ/LHLBEJggZvdYbJbvtn7RQrJIObKjujmazfid9WgH1HkHfH7P4G+GOF8MY
THZH70VRtYH0NDBQ0AVp2Hubamq+zlzxSFP40WTxPuNS71CvTwXXVJVbKBULjsBS
3rMTwuOMZM2gkIOc30OolamgomoKQ2D5BxaPYPds/tcu0W8TP+qhDgv5YU3xZGj+
Kv9tQSBOTM1fz+Z8fJxhTrST6ehmmHePQsONhSQQdlTjkzCQzymOzWiQCmOj0iWh
7fDCc0xaqQL0cpVCW8kvkxhFxZSefGQPqZEf+9r6vTXztX4zr+j1RpaNgvfk+heG
MrXJY2OIiUz+ZOvYzD80QDGJDOl+Gw4/0XAXPYB94XY8LSx197TKNIYXnVsUE9tB
GOEZ/VigcIDtoi64XSYu9Sa/YddvrU0dn+HVT1CDS1DmD/rAHsBRrrrl8NfUWRG3
EAT/2ZISv5eY5qXVp5entbF8TzOv6JGr58zXwaFgNHFBeYdWdwAlm/qWTZQWGyxa
We15uL5XOfp9VqUnO0MH++W2usr1kuYj1eB1DUlK0VkpQFE36oTlkS/Kd6HcRAbv
11GiKAVWE9gpgYmJuGBVJOyBX5cCDiL5eupGaD43T5AVQrvYfxFm0Q5+tGe5OTi0
63pwMVJ7u3Gmxw74aM6FwrhIBJ9+pjtNqwpvpVWwqdDGdqpWJ4tmI3l+BTFrxMiv
R6TY6r36dfSDBMVgB28PAk3My8qZavYoZZhmjKCF0InM+zsLO4uNtCtN1wp3Vdml
Z9DSIDNOnzBXvOsLWoMMiXpK9n4yS646IiYrvAX7SKvbs0rz0jcANOqpRKuLZPJ0
tOC0/2RXObHu2sqhlSiNSsny0448ECD8pIYG0VWIMgKQ5Lj6GlWhfxMba2RtVXsI
XyG9BsyL9CpCUP0cls7o8GkUABjvH6OPr4RHQ36K9W9XfYn2J2U1i6FLDAvigabu
jfdlVVSsiHzhzPuuli6Xe7w4t6AuFiDeDJpuYmL5I3T43WPhOaKUSt+zLuPJvUS8
MuFtpa11UrwETteX1OaV7YkKj/Vh9ycgDQibL0vB7KUFLnEnWWuRFeDtydF28hHN
oC7zyh4FPLCVqAxGqfHdhYuOH+Hok+db8BIdhsfYlA1oY+WoFxu43wDZAJz67RK3
Wrz++Dimdi661hj5aZNOzYPR5otwbGfM3HQZzSbRNbkjGK5YMN+UkIYYs+DQty8T
yC7ZZVNinW7ozheeh/J9L0P6jmU/NjflMyxhIlm2NXam5/RfU5/A6liSj7deOJrf
zuxpop2nWzBYfxxAby23PN1ul+ucnzpbc+ZZljwfXgCf7q8QsLOoVHi36MAcIKcN
Qd5nATb3fTwesnKGGQFykZR9+WKrBGvgKK8Y3MEP70cIh1nsyehGexW3TdKteerp
hhqIw0+YG/GPLB8VqywB0jXYuOnI+ZjYad0sQOCES8JQKMxcqjkQ0n7WBwx54ied
4VfPF9iwOG7aDU5tIFN7HFlWGtQ+/EMC/q3j835cQjamEQSN60KuOK+6D8oeJV34
86kMVNJzMxNCJOY0V7fNAaJkFiESM2jlaYY8pRq1gfVEEclpD9pjCn4MNVWbERy6
DexzFDdk+rYvnUnKfQRPqSrmQKVKrlHaVBwBWyAeAEQk8mlyzacwzKBW9JU4lnIg
vtmQWpnfo1I1CJ8go83gUF9qRagDSfoavdmQQTSIPGOfvJeCep5z2BOcVKexl8Nc
1dPFquE81zcfVDagD+6KNGNX7LfVgn0gTY525ugju8VEaeP5Nb1EKS2bOA6C+cQ8
9dDzxYgXsVAtthE0GTIwec96XzqvEJPuKZW8F12MEdzU1WOqqKMdMGJa+EvKMx7B
Qmw/ZqqJYdT3RiviGQ3kUYB0aisrvagdV0cwjdo1qTAfB1BurBUalKKfkBAMqzmg
NlzEos3YQ5dVvJxv19e7T/hnxKPvF87HCTixvE2sq2iT50ZYjBdyW7MVhP840lHD
rQnN3rxsb1DueN7V04sX1x/cydlpfdhHj64bQdvw8ApuY8CV9a3LicbFOXjHHVER
pbjr3MYN7kLhcnv3RFDa8C2Afjr+VzulGp+3VaIwh+k2fG5C7euFWgywAFcUPEfk
0q3SAOXmK3WiD3yo0IH6cTX9sFS+oYY5N765krbqJdbokCUuEsxDCOQZXak14tGy
ZpAqjhAFseRy8l8XvFENN+A4dIaCDPYqcutS6MiGVYmDnXDH0LhJ28/ZBYZwpwoy
M7sDPms1qJHn4mZZCSbhIOgi6gMiJD0nnwOyqbpkLY5PLUnJ9jOUve+TzKwB9EYg
SgVDJrA0oSoBrYZmUfJwhxkiVMWCBuX9eN0Xxr05raM030NQQxWYdDotbu3Y15/u
mHvK9foOSD5IYMKz3hiSHMz/NfZPisaOvIRS+oObOTLkOiipH8Ym3GDoGEJWsyCw
VtJyhfdL3cmVcgKc95Mr+NIqUZu1ulyeHsa7lwGm42J0jB/mt4AEA4c0vWCDVzfj
WwVgEnSOOdY4ovDC8hEvJEZuhLQn5z+dcFaw4Um0N6yeM4o2ioUc945qr0cqcaJi
NXI7zaXQagFMSJYuxXWIBcAxUjfAbqn/i8taE8h68mCHNsIGzwBfklZwfcgb89Tz
KjJNhD7z5UsCj4SjrvDWhO65wUWl58mwrit1TYwqZsp9vKCbkuFVmy+jpTrz4Joo
fCTT0wAPTnTThYYhJgpHxd4uJePjQPzq0ex+4MBW8wlPJQP+83/VZi23U0PgqLeT
3llnFjNoikDBC/jTEXv160NLaNGcHlsOu0bLrhPNbBvRTG87tpEbdnL4cp9os4J4
D7V56BIO+UeinzlmLvM5a+jztYOnqA2GIZZ4ltMBwOSU5oyitqah2ut4NsCMQPMS
gimF7B7ZmZuPpAtIZRnwVJDE1Tbfzfv/5//VjlqLMa7v+0xEVvLixN5S/s7nwq6T
M1eVRNM9Zhwnj3CHJ7sda4k9k/WRWsBwC88BVBpk7x+rLzyOHbIGyg60pmEB0XWD
H8hx7PZX0f3LZPlzsirOQ9Mzl6ymqNiNaJuWCdKJM+2U4lLUySkZdpiZQUaGbwj0
WIZeMcxoIs4rgzG97sHNw+hfWONMtYZOZS/NBywtjhIlJ8tEkBkWYn4qQxTAuJ88
FILqYet3oMHgLnzwARkwO17YDBI8bJASlwPpzBUC7KJGilvX+PY4TM20Ey2ODjrj
7vfjnUEwrPr/valofX/+BIEZmp2PnsTYjyaDEoUs9srz2Ev75HvFaeXtlPdxcNjk
B3GjhyYQmWJkQjCJ6oXKIoRtD2Kc/YoM6QFfoOtgjxx9YYsMKq7aaTWgjqzT8GH+
JdmN2NA69rMuAU40g9ZVDpJNCJ0ZbKqRyMkai2DIV5qQbVUoC8lz1brQris/3HHP
lFURFwKmulklLH2BqdPMRoGRgW0auoRZtYpXTWJJ/2DPI9hGGXGYl4aTav0rv0Qs
zCN6xPPKEtT0hJspGxoq615YgVtoSsItRvmI3g/DLsDSScY97M6hN38ubxu/cGX2
wATRXoli6yHokjUmy+Y6UnhiTleiQ/X+kiL7KQbsOigSs21o9RpNnr92JzkbnIpB
qDbBivRHIN3vV2UVfd56SACCNc6Yqd4JB3zxSinV5VgRZOIVzrtPUYVvyioAJStG
D54C4SwkLOzu5vgjbY2SvNwYmsydWlj3n95hmm/RXQfvl1Y4+HwgMnRND96vhDQf
D7oO+k3vkAKXIMQGyQWOXbAvU806fhryN+EzI8u4AKqpDQmwHAF1W7FRi0oUnezH
GaxmY2Pr0w/uJPIjsfIWFm0MsOKST1U56dRLcI1zLH16FEn5wOeCH5C8siZJg6FX
c8BJRqdxtS1skU/kEyFLY3DqVxQWfNr0busWQQLpHOYmsTTgA9GWNEbAcbSq3oJW
VacwLJrU72fLCRKRZt1mwY17yQ+/6eY3EZhVjD+07jytAbtxvDxZGSHFThY3xysH
D4sRzHrH9a5ATHeLnqE/LKoR73qWMxDGSZRyMjseRXQ+a/qQuPVj/aVEhMkwUJF1
NMol8nPcNuRKoP2BE1TqRd+RDgDDzc/Aus3kcRjz9RFxA2KGWEwpBWA+GnlHzUHp
uDZvxqEO/sSGerRveRn1tCqE4B8iZCRlXVYuQuk/rDpi6KvrHgoOQQdIrriPV0eY
F4ew5dMpGGp8DLCkXnyI2SvxXvivLxIYMDpBbCyB8PmUyhfnLV6jqrZQhoIioNRZ
7LqDf5zmwILdvMQatl/CCys2591lHZUW6p2nCnQikQGu3reWc80O7Gy0NRTlPV80
bmtK3weKzuU3U+BpbpZRaOVfk87kP8k1G0XqLCRLPD856JCTJ20aZiOrL6da+zt0
lpJpHEQpmfeFETbgExgmLH1naqlkcvIDLV2yn+rEJvtsm1EMOz0/4Qi2WZhc4CbF
7oUweWPvb6bdiDjAuWto79oJ4RTVP14I0odNSQy0v7PoEW5ju42oesY1mtY5vrzL
Xf0O92IL5uGFc1StvOxELDgoGtnPqO9LXXObJ7AbNTSv51goRqXsrVrjEii7UsQE
mWlZoHl8rZ/ju1/FTcTlJ2vtx/ThOuMVWrmp7k+0soQucZIr1mDpCvzM9o5UVQ6k
W0YU6ks/PbVm7+HvzWOTzMRF/EPevv8UcPGpSnkjMW16oNuWDMaL6XrfXUzrZ+zq
VBgDvwJoB0WF1z5W/m5yozguEzMN8OczNaEfTIPoBo0CoWxnOzRaZ9H6Goft5eE6
1+94JsvAd3ipEP3pcoyqVhWDMdYzqo2nJQ/ueZ/up2zoppfNrmAhIQNHRlDIqL4z
4HIR37g/GblbzmJ051+AM8pYeWJQzKsVFoL7pgUJSpBKqmTHo7/gOSF1eqI70NBQ
P01g6gzGrPtaaA5x8xJtRMvCZ3FnhvW7ulVD5aCgQ3FbkYqGVinh+Iie0ChuIp2H
FED6z7MNA9eQhdqgIoZ5l8CFuLTD6Zr97bz2KMfrur5eIn+Urx/NVCGTmDPAm/Hv
q6koA2N7syf17LAGZg95AcD9xiaQg+oCAXe000FGKWB3kHLC8usZ/KYmk0JEL0AB
7HqZvJsYYW8CDjCFJaq932De5XIKu/V0lQ/feUGH6VKkqLVAeUqe2Vf8ajysEOkt
WyYacRw8uKDxBedHZ7JuWUPx73FLqHGk4RLflw1i4ZEwxSFEMA577cuGO3aGpwAJ
j5NgZwy2u2tZ7+8+zVpeg4hzDG40jN1CrzWvUvkDLodTCigI6gU2jh8X9sikDRve
sPqGe6KT2PHtSY8wonaBriOGVGc+DWucoZEm9apIJrJAXsfY/3u7ILigZMVoTud3
EkhGxiBOHKFj+qT7gd0bXFo84aLDuHpEZgsgdLleA/cG6hLTcb0fQi8mRBeh83yU
245AZ0QSffAUU29XDjJrAWL7rBXFv0VjgcU4Yh4hGdv6Qu6OdX/yPF0ncIIFqcbB
H7WmLoh1jMx20SN34sakS5a6bVhQL3g3UYqxUDM7qs1zxGCOH8UWG25J/9HdhOYN
DAdh+/7Vlzu+TkCZi94tQLnAk59se44wz5WKgLfp+h5mckB1W9M5tzSxEQQxDo5t
A+4md4Xr/DKiCYGBnh+XygULDfhngLlO33reXCn1q4QOeNyN7e0vdJxB0Y8vRapU
4sjX6J6eHxFkhtgI4LVVvt9NUTa22IVS+CRLSdPgBjMMIKtAPKrqNXKPbML5OayQ
hVhyup776APssIEtRDgr8HobPu3kA/tzhFpwiAcdwYoVrclTG+lyUvn2B1AgK7Dv
YmU9CV2gkQEfPeV6DfEp54dQcsudXtGwdgr++IoWt9iLX4alinZy9VPoQaCtvXs5
QWl/aqqtqJ4vYZ1g6h93ub6JXDsIsjwuH5gl6w0j9Pl9LxgeAO8IvONwwFC1adQ7
es7iO1YnFa/RrHGxXb+VMl7PJuadxJysfGtt5Qjicc210+MmKh/j4TMIFL3Nv3I5
Mr6MQlYH9lNA+WSUras/qpW1x3ZLCkNU//Qdpi4hP4kCIk8mIWDrYXHD/obemmcW
ocCCVM1B/ddTADFRQyOzGW4qzhxpywDPeWVm1ygHpNLQR/B94Lj+uKH059SiBswQ
KnH5oElz97hJeeQ1Ko/WxImtHy+MvzXScIhdKLUu4zC+G/VRHTpsn7OtBIDvgUEh
BUWDiNs27+69554vArxXaoWK5DCMFplkv+YAsjZhCI7hRBs64JiL5RzzNk8+Aa8s
nY5EA5FZcZBA+F5wY6VRMQG0sALU6siFSEOxzc2IG1q1u8cdkKR5FGmmU6605yxI
/QLdUXx02F5jz1qePm8kRHIy+lao5QhRBk+Z9xalxfYkiod7/ZcLgAhqk1TRSzsC
a1mmqv1WgfKussgIzulD4tUlAS99x56rrD4LXfZfcH61xc8pup3fbStwV1cKiwfK
pc3NGQtVML8RTRVsiYPQSmgaSGo+Xk8YonHYSLzzXAypwWIJcsevoy+OeZf7WNzw
zHfirtPi/L8YKgmAL40bJVPhPcW8VTRE3VWn7r7RUCy+2JMPADHxJQAU9sqr18w8
IbXgbBK7JJx30N4aNVudHP0hd0YyStLQzDf4/lLFmw40fcSc1M8e8dssHstLCGGz
ZdsP6hUbuY/vAkjKK4udFJU2SIoQk/sNlNvb168OP31wAJVkE9DZP3dLHOKq3bbA
fQOWiHZsAz+WpcofJ6Kvh2Bxg2CuM5a7wl8EoCHPt/rX90cT4YEDzhtPBNerMSlz
NNoLu6lhA+HIxGAy7U7i4kWL/EDdk1WCUMs35dZ6sT9Axeu0Pv8INHbDw4TquplF
Q58m808Sxv9hPbc/p1H++NFYZBkQ2NEGDvZOYc0cShpgXVoyK7MAp0BettJScrR1
vBkPVpUWUhIf+uInkEaZAWKVAhb39sFbrAzfZREdAFncokDtgOaWR0mWJdeZoQFO
v+Vtxm/3+XehrzHesgyuP/mgwVRnmQngmEiDF5S15VgNrUFZHidxz29lW5deEu4p
h63vEzgIbmrEuq8W3kv+l6Ten1tME5wNxXDn8ZmIiwwb/xXfPhpxgCCHkkmyl9//
/9DLFiPxMsOHFHCjhlNvL3O79UMqnQZjkkVVxGauKGYat6XF3yC77r9w2ld0SelM
9oX0kk6aL3IPbSXMr8zAMaaOYqOALIZl3OCaTVZQvfXX0lUG438JIlKLdGQr5dEr
LR7T059XoFWUiDtQxuMT1aE/5j2ugHRhVL37nA/JbmYdHzpql86rsA3iZcyGtK/6
`pragma protect end_protected
