-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xgLfVrunq+Q8zwwMbtornPgist8U6FRY9Cjrf56aIOMWMu3fZ049EhR+pcEDV2JWv+QwrlY6YWX0
+BjHm/bXuweNv4kXSWAzIxMGvcQmZViJYcJOfuguf0qDqwo3N4Axp5211cEZl0CRRoHWM/WyAuyx
l3CdOF6Yw4ijyzHOW/WlfIaDSNLFDMyJUs/b+vY0arhvkkzpK0FI/7tO4ebJbNfsF4ZSORKZQw+Q
pBO3kVBz6rhHIXHWyVz+aiy8VeW9+lVRmYRebOeSJNeWr5vfrgvIvzlvrLhjAwRxMNmF7janssR0
PcwznXtLZ84ZH2cX9ZndknQi3mz1ytnDeGy6eg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5328)
`protect data_block
Z8WhNWZsBowbC1aaZqhhkdkXAaM0qxr+GNYPaPiN9eItaWjewExoQYfPmcXPXUA2LR/oXkWKZ/gp
Ta+YEXcWmmMqPBP6SSeg7efYFAgJEZ/GZCJ4/CBqPXqAeBKDXiysw5ATJ5pe0svJnmCxhdv3jxV8
s2v/XLbggTmBp5aEYCgwyyYmLjaiu7EhDm2e4eKYjvIx6Yrqchj2DlHHmNb6y7tETNrIxXSx3F5N
7Z12JNrSlvnU9sRgmW93UeSUsO/AqWBUsXuptYirZtuxWRQcjT3go3v5IcnnuMaUuW/Dm28RrHEb
ge6Q/cnNHupM+USEWQd6d4htMGB8k5uQZfJH62fevLrmz4Q9IWvpavfEhT2ow5pmbNmlIyZ8S+sY
6sNQdMirqdc5tl8kBoKfiT7OOMVtRBBccrOBCCG5DtsVb6ctjty3G+xQwfrP2lgDZuOhKsTcynlJ
9d03uzLu2mhvRSuA/hJmchNB6QlO2P9nWsn8H5AIP1YknF+6yRyUvPmXULxteoIbNbrrT3whoUGN
e7G9L8myuNThIOR7TGkuxXcPx7lMNVEGPjG3oxN5PJ+To6/3nbQeA8mRec+AYD32ohpxI3PV85pB
QdnfnTspNEJXJGUC9mAW2IwHorg72F1YnIlyhZpyyeJEEgN8Jh13tYLQN+wDm+0VR7PhUWk1z6WI
Uk+S6f34qqTdA+AXDPmtlM2EMKOzQNFK0HQWDw3+om9svBKMOu/Av7wa4oUDi0xT1x32bl+5tNeS
ObK503mM7ov+ObztRD/p31a2gFuewikmMFkpcN1M4MkqOZIgygrrfxB9/exkyOK97Npt5e0Lwub1
ueU6tuzCKoTps23db/LqAzqlcT/PWJ1+Ow+zV0feFWkxKD9xW74uzlEJSXUNfCVnJ29Rx4cM91wr
HGLvOuYTfKhwk4DbAeZNJwxIaIMssT3P1xsJjr5TtuEUJYhhHTwD56rXJD+SRHi+8cJDCvP+BXBv
7td5K9i5zSFQXLH6RYRdz4inT2rK7LOXxqPAHgiUt9mNaiExYMGlByOqV7J2+IA8qZ4cQfkxzavc
8pFfhl0GEPtfK4GYqjR/K7SebbAQJVHPDkdZcV/I7ivxfxA+9Nc07l47GavZk4ccSlif2j0+8GqY
/bqwBYWCho1uL3D47Qh5rujsA6uNIDc/RSgYBGBXLkU6fjsRdUj3WjZr2pwX6osh/Zb5p1MhKTTf
/9C6XJGeTGwYe9psUzw3NcLQmOFVXctNAUiLPLi92Iw15P79di4wv8CIRv3fHjVfhpAZHNWl7d3R
l/IEPja1Rjf3bOPn06UY3q2GPP2CFKN3lp/ZRJEBnBilE2Df2uCCBRq6dLKgn0bE5WiPITFM2JE8
uXKXuVE5YhrJLXdWh1cnKWEPOChEDdvd+uOcTrxMBCXqJNcDy6v4L9scgXtxkUUIOYa3Y25obQBK
RD0R1h5psFSmq7kwOVzVKqmk/sFF7mXIRMVb2XRXPvSj1aQCFbb09SpM/Mq9zseD1I2Tm3Q/AmwX
JFGGJklNgES5p9qS5a/KUnuueqLDJjx4kqMfigr6LjJPbX6DEMEZWVrZukCwyyowgmSBfhOEW0Lh
eWUDqxTFLDC831TtT2LEvrLziPK8u3kqJbYgVfTGttHv6DPrwGs9tiOPrKfOMhfkTSVVAtFxIpnu
3Y2MnvP8Ve1GhiUTur+UIxWqZ6QaIeDSK/Z36kKXvCMrm/pRBSUYIoL/hrUtYAOgCIS97nbH1hZI
p4tcVRXHprnUbERRB3L6SLy11gDn+RAVpvXOMP88xLhHcH4TNJkVCw44SAfJkB7Fpg0zP2wpscIl
M6RcPOev0/uAMb8bA+71NJziMEMy04JlF0VsCPPdcS8ciGHremm0PpwIKySw7Gy7VbqMHvw/soKU
oDwHVGxfEYQO5MHxly76P4uql5i94penD+jtdN96vAOqeD/VkY1vuJ5ewer/83DS+hk3Qx+4iHn9
hgceeNGJZ+Gzo4rMUg7/QNiFktIY2Mt9PSlJRQo1qHLMSrKOHFrSGr4N1TXA/0jkA9oLaXQRm1oq
c4OsrdgWfaaxGG3LLLMyNIxJE7xaiIgwWDzajdAUOJHPpsBNb8BbxThQWtxfw+CFUmIVEsjDUkTV
Z8dxlMwd2/t8S110slipVTQQZ120/RJ4TeJKo/wcBtLDgrD+GYBB0cftGFzj25hFOMFT63CFqYSd
xoLhr8H1vw+ioj9ilQ9z3OzPmj0Wxb/7tyMFfaEBuh59mpM8p8fBL/9VGtC82S3vLcy13xj2h1Vv
jmQPSLv/p863cqrRqLEYJ25XQJ0sNyNVGumlSvtQDpA+NHNUWZh2btsxkVmV5x2/pZBC74BBxAVy
e5ujiaRSPqMLR/YiwlkfDCm2by3d7dcXLtnyYjumBhMek3eG5vujsZzoYcPoHEGgoWNU1wMj9KHe
/MxVUPxsH9EWwDwrS8idQ1q5vtmmbpuwt0GaeftFztI8T+zV3wW8ntDflMKG1SA50VEXth7eItMV
sXjjfDRTbGcgIKZMXBh2P16l3Mqa348ucqsbEG9E5EYq5UrCm+OKHpms161X4Umhsoa7ZG4k/uz4
0oMGtTZ1SDHevxz/jE0Ovjcpzn3kYeppftmpAIm75Kfnj4B8WFUHRQyb9H8DDOrlB7kG3/cO5Ndy
Yf0KvKoErKubx19wZ7w0YnOvS3izVW5fAilWe70GkBeVTW206Kg087hL7bS6MiVvMA4YjT+k6eoU
x5wRYQ5+ZF2LKJyPXWj4MwNwGf0QHs6rRNrcIACekh/gxB6/gnsQrqq3MYOTaqvezlDF75ZVANej
YSava/BlF72I3MtUOaTXFMeJAQHXOdvXzfTGW85WMHhrN5zFIZ+9XSOGcSpIKbizcIUeVsDWvEnC
jOHtR67k5CixplPpBH3u08QzNCwbpILQHngb3wAdHZ4QOzZ3rJ3QacH6oIEGVx/Z6Io1VYrn5/5G
CGNGSB09SLFOvrU7UvAUkPmGDcUKDSEd15o7f0ws7kOgZr8+Pn6FszLrvbuFAR4XqeP1GqQGHQQ6
9VzL5S3jnVfPBgp3QaOjoLNGhcrzgO5exFn7FjXRf9GKsHxHZGODu315f3sURMbeKyqrVlsjAssu
yATG9/01rsOdukyUFZwTbU8zn3cZFgCdAD2nmxcz8NtB7QCWRgvPrvNAnBd8Q2joDKZeiCH/PRns
SHVU5c8Z80vxupLnJLMu1rhSlReMS1+ykleDLTecJ4aCtlo+7JA3d34TZbKhVpHzmo8vC8YYdSE+
b0nKZNNZCAtybLF+4Ki6zUIL20KWXFxKpyRla5l9neo6/zAbcDOQiiLn3cmzor6NEgygVl8mwTIj
p30YFyoB0hX3L8lJNonXh375A5Hpbz+zLG3zbE2q3jeUXuX9/MdZAnnvRGS7tfSqnUxYFMH2G9+U
8q9gG5W8KHP0PAGHAna2KxDdMtHoy3Ey5ij+EXIdOyWQNseDFMovJPtvC3GDnqGR6DolVnAcX2M8
d4csjtceiIaA8Uew6JAQ3ZMkw1V8JfXGbxO+YyvbTcqBN5VJnVCIEEHLGahNe4+A5L6RQ8pllVJC
TJ6quKTTkURSekG/84W0ayIUx5Q+zdc6853DSLA6kQh3BBi1sRzVP0pVN3TdDx1B3lmHOsghS9dL
9nVzKexf9IRjpgLQwKp1gIANx2RwrpU+V4yEJlQs72Fu4s0opa75eiOibM2j9lfMHLMXqYsQAH08
ApGohvaQ2euX+5tdz1hyiaRfQ+MrOogm98DS4Y605FREWZBV9yazKbMxaPuBCwIY+VknNjI8Ewdr
8JgbQ4MzbHOxKZiI8biV4gKKTMwA/8VaFEP4oN+atC6HPaFU4fAMbuP2vdLAEJx0TNkQ9GU76NtD
sPVpsiL5ocMfD8xPNNceNBl/9jp+jRbgnFoNh7wcMopD2t/zZI33m43yU3LJrxLSTSeYipI3OORI
XA5gNnAP/mX02YzKI8Tsh62dkMTw75WbE1bmStFui2tA7ZsqHqGK4gOsgiPUTRodDBOtlZSbs8U8
SXb11nNrlyupX5P2udGGoUHjcO2gxvJaB9Ye+mh2dyL48dpreJiXPABPFZp/Wc73BZTnRUx+4cHO
OvbZC/YbaJaJqO/E7CRm72oK0aHQ3aUUlSFh7PzDl1szY4ciPqVEJwGMP7xQClUz3ESn8xyuW+eG
2bGgInEG2poG5yst/wtdeN4RpEIhZU8ebgvFEp8QLLZSM8cUAfne1Zka5dhmBoNIO5fP0ZL4yN/p
0n1UnLIynWOtBpagwK6BOZ1j9Id9o6B5lI+wBkZthdimI1yg21jRtz3PUVj2VikCSJ6Ifi5LvJwl
19UAdSQZ4gJP/8gjhPtS+xSCCSKPaVXtmBuicnYVNcuWEcgMeL1Os0klotNEmwFiY3wIfOX/r4Bp
KqpnCzulJpxKHBknLPKT8wAjOQIiR1V3L3Tq1gymor+aLVpL1lnjjU5+XdykUlfvtgZwWcPTgRdA
z91q2ptTO6zXN9YWCzSceQPVxHN8cBIYXfYeLki7792pf0DknXmIUQMTqPCzsBzOm4JT+AoO7PA3
LjNXtUmvmEfeGotkO77lt8zVogsPIrjFQt2eHnJLIaK4i8xt8NMviM39aMnMz40Ct8Pnr2cOssGC
AQcN0NHr+RecztktaizxoZBZuYOWuv9hTfjjARtrxwq4krLxaJaB7r3cojAxmQURxONg6VgjDe/k
9A6kaPi5bqX4FCcLQOphRoCP6grRD0hhO4m+Rt720bgJefvbaL2ZqgMuHYP0jhdxAPyDGzcDeNgM
GDJWzClP7+bjjExIBWxjYb2WNGpeKIItpkNDWYPiyMX858+pEPd/az5FwgeMf7NRYbV5GrCWNoi6
HEcT6NgZVaAYwD37cS3PZtj2dPk+znhbHygRLA9Eh0gDszyo2sfROJaeoWG8bUTSQZwEECA1eUIk
0bbGdvv/3CdHt5vF/0ws4qhVQxu3rhU2DvxJ95vmd1MaeRK7xDx5Hi+rNEp8TqBKAwA8lCTK/jJi
DW6mZUn306w7TboYXEG0G+qyHfCtYUkusBed1a9Qitlmir8a7EJdmiWxaNolC+ehtK9IAZAoJQ6O
/GsKVZbuNVGnntMKXwjqrCx8taZbkFlNex7uUCdSCI6vmV+1zE/cONL0pCoXthASaxoipCi+govG
Bt85Lcjk4ALv04PUqPg8ldh0rE8QBOlF3oOwRFRUOIdBhT50kmHdVUxBxzCqpxl9TsdXWEOLQX9D
hOAdpM8TPjyHqM6GtreR8C+WrSdBXzCY9s10G1FgEOvh+MnEhoyjLCQsNPgZUkYS3NFtlHwdJb77
QYQkpnf7YOFBNXzjtBsoUgiR3YCqLZv20O3jKmyuK43NJUUvt0EKTZRXPp47wgUPyhTZoRNysZhM
RTGGNASEmWrErwRC59Dz9btZokH6q7h6KtYQxDBhFY4/o+lG2K7MB7uv8U4r7fXuEpm01nIBGcpU
IR+dQyYuFRzSViN4fJ1fisUO0U34v87KUMZN7ZmSICyZCH9gCvUXuFzfKUHNxHPTiQI5470rRXsG
a2C6lPAv+CAkJBOq6IP8Ifw8TamG25daRY6ny731iCQTKuYQLdhNCvFTdg2pAaYpiaFyyVj5W3Il
xUHqMEcBaPN6B+TwslwF3OEX0gjN1uEu8ekb+svrAa3RhFQxBhGr2Y5Zx55Qiz+VvdzTMcUQamyT
vye9Gy/4+GqGWTkafeETtUjX4FcLzaqCtuTZMDg95vgU0qGpcdV/uofzzYzIX6cu+3sdMduv945A
f6e6XP0tyuwGc5OdLtRxdFNiWZfJmbT00qa96HqsWkqCqVa6zNTlhmTFsQ7gOjucAYfUPg5QdieF
r6ivKvFJfCBsxeTJveEWGpW3sJHPuEhYAncWPrJm2rI6jFbrJxan9yObAyP/wtPckNv0HLJjn28h
4ba5tjUv2Wz5sh4oZp3dRh4BkCtcWhQL069NsrT80GkKZdUZ79JgbMzOvi1sH/W06ltk0v12qv/W
NKVdPlB7vO9yGvWGZ9SIG505LbR6TX8X8GRqpMKRQjYBLSuZ7qBbCYrECE9xDezpKFB+n/z+Jtkz
6ekLYa+lYg5+dlzxpvNRN5HQBkXNQjJdaLuyY0EZ+1Ws6fJ0sJX6ddzWGMKofje+7iXT/KhbSc0G
i/FPwM16f27Lo1plNm0t4r0YZC1tpmSqm2Fxl6gL2TJUZzcRCZxtkI6FNC2ek8EKGoPiz67TVnXx
cakH0q2/fbDlfyGYIZOBEEd1bvxNlm7qi56I4xfl3G9ip+zixrEILJeC6+eRwM3posAoYULNJDjd
xZXSBvDhCanic9gIiUpKsRpPpgaX/oraACl44aqdNgUqK4SKtnJeOYoSkZhGoMOu6zwzIafjZ5Qf
E/HXa7mlUDjpq+pItmlF112T559t13v6nBADb66uvG6sbSevaNwQ98hPD31rQnJUFJQL5G2oeWv0
d+BrKzPjuvh1uhQnzsPtljcP7pHJ9OyY8OiwUOKbKEnQAZhqiLT/X1xyhmBnygEUeMSMjJ8L8v6d
qBHSBDpyoxCztUPwkt/8UpAa2ltnnIiofQ9tDUbKyM+luYYPuN/mb2T26JQUqznTQf+7W1qiYLbQ
Kt5OpOVysVfxRLS7JEzHrtVK9rmFSikU9jV7UQqHVUArZRq/tJOQN190TlI92XeE1J+LtTbezAIP
ZrUni2TZ0NU6xgw8cZZlUtMfc+HtNxwO4YUc/SI3uVjD2Ld067cfB0OWtGL0e2DbltVt+12O+IV4
gKbn3lfCCwxIxiLxDAVtLOXPB2gcETHeDCXHWqi6lJJJVT55MQ6AjpW/z0X/a0QS9QLgvdBQLo5w
9Y4bei8Au3mG99k+pOrrTzuYfgPGTMR7pBPmbmi2kd2/IrHtM2/M6eaIhkq9Yhcnl3oHXjT9xBlO
TZQbMFyq1p9A+qSmbwFKzqKIcgiAZX/Td7fUwaRDv3nmzeZT3Zj5G3K/T3HOqcdclMPNAzg6viaL
cLxydboe3b860uhsSt9JA4pbybd82UNMDRM1U8Eh5iSA1Jp0LVyIAHMV4pukAjlsM05n8sQBKMYa
dv+Bc69gT2ZqTkJJUjLr1HD2VZkeswxcjIET
`protect end_protected
