`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D74oyTD2nrNox5W2wItO0G7PYLqKcnf5NFimHWPTEd64mvFA6jZB/Ebup1v1ygp6
+7ypA5F0IBSN6wzLSd/CM39TsHwb6UjBc1rVsk44MjWNvgg8Wu/IO8aV1ZORHu6a
MLz6klGVya5sqrPuabz8sFo6vjkN+vur0Kgt5a4EQIg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8256)
Xx8x6BmXkW2AbOwZnhzONY8YWeIdnnRDmB18AC4Vn252u2HOTh8Tlr/VH5+Ey37W
OXnyRQlgw26jWfUoJaW/TT5ikl73PqMPOiRUuTk4gb+KhLm7BreWD+DalkLOIgVC
Pb7H490nlqFk2Bz0z/6w7NuxDgBrlyDBHbUerrURj0Be4x2Ks0FYLNWuZAT9aQA8
6GYTAwqzZ30133t1en2mdAmIhQK7XzfCJXU4OodgTrqd1PJnApa7dYsJX4WhMMEO
R8+qIzKW9Vr7U6i0y7/MuldC8qLibIGk160D9+LfPa31QTW6aZMt2Au2uao732B+
FaxgDIa0XHAt2+HeXTZ1fv2Sw9CCJPkQm+M37QQqyaZJiHhro6L96BITAq2rW5EK
S3+taVI3O5/cCLjpanNMo5FhM9BEYbzPNQYsBuUIrs/Dm1uACIyrWnEodbPE5OY+
Y3cCQMXb+6l1TEjJmagcQjwqTiSD5in47tyReonnLZyWCJEmpecbY3XP+rhi9V5c
QElqZ3viS4jCf5LFEyJAJ7Z5VcdSTUba+j73oyUaBqecD8wH4i26/vHrwhAHj1lZ
pS1FetTzA2N3R1iaURVlmpaSf6G0/eaxAfKd3wmejkQiEz2u88Ymch38XfGvdwAS
NJD4KNz2JNRTPUrLvO3hZ1eJsDA5qZ+XXlnaVn/VO3TAQOkh3CmbrOn6Aiy5r+Eo
A02ci2uW232JMZwhK5wTkBGUemKgE/0C7CW5VC4whL4OFpMfXVOcth8Nb86m+LBt
AuwRsXeCQfeimGVNirB7WLcIHQtxhugwMWxXS52Ndhc7haCxXCe8/+0G+CbDk4K2
daUvIUphDO3pfCYrVagOvELZEms5WOiI8dX+wrZtFwublvCBSc9y99mx/QVH1O2E
s8UJFN48UO0j3OvPIwXPZUhx7+9p05dTY5XQImsPN9CV9WMGLn/E67xN+LYl9++X
GsGipWwOftD7S0Uy4XirERXWN0QB+ajIDnGfYkchET77ypc7EUILPBcVeOHHINNt
Wt3570D6NOmazNbPmVScm5Cx59fALi9iE8ls+x2d90d+75SqqF6dOQnx2o5z9QRV
1ff1xCQ+Z+WDyzyWKiqRsiPAwxUn2x/5SVeDskW2dqC4SJyeVrxJJfo2cNArLUJM
rUL7JDuTvw9diT2ZAWd6ncjrP9JM3epEhuolHLxl/Ejb/WLASgLUd/YkQ9PzBbpy
aJYEmBwqqvwH78f5DNfLbjjjGOLTCPc/OSNVVsy3CMkHLGMAxCNdhUZ8TfbM2ipw
4LZjeSA1FQqFkyoZxXsvFrUpsl2imke6T9oWAldtx4aoMXEngPvQs59teEY3Cbc5
G+3Gi9otcqKoFjIxVwpnTrI6ki7cWikewtfIQ5XrZhZplT7bo8dWta4Ji9GKF6Xd
n+bx2Jf+qoPq/DlYvEBiQyIqVwgindCkv1nfQiFsPe3uRLjny7fCI26JaY+DLBCY
fWV2QeYu+CqpF0YHiYwvfRlAKgF/CmRK2rJ4eqQz1EfcaoDY7Hu7637h0YDYbcDH
0Dw6PSME4kOMfOKpi8UMexSUZVA7y6UV4oMhyA99bl09HjwUYAp4eTz3s2W9QC82
+y8jh79kbT8fGmv2wVqTB/JsCLhZaOCCEzHyldIr28nscvhe3KCC8cLvp7Mgcr4B
UCgv0VrzH7Oc15Lj5dc+igq9d59eerc06W0Ww+UU5GMqgdk6zERxntBZ0KMBKoFY
HOJxr19HcUVPnjbprlPbKqFl+3REirkX7ZVBUfIuFoLEyaEL2Qq9CKafVcJ7FxRe
j34AQ8Ip5ELpz8Cn75wyBUnCWADmnDdJgYPHK0wrJrm9GZHGJf3LrfG78bWkL4Cd
epNPXMOPU8XfRL5x73qiLso+CG0OP+auegQrGP+AJTPdobPv151fy699uRHUkle9
/CIr+du/WsthQbZVapYD/qJyyzc+EAvgEjOmf2pCCzQouMTCs2LLxiOCDCTq9KNt
WVSpca/7liOXsuUn/8dxjdHBDWBReBesx9wXrDzYBozEdFnIHnGf0wd4rVXlmWHs
bC1mW1bR82TZQ6+lTksptbnrqj+mNOWmaHQPwMuew11c7B5ptWrDj1nQyVjxxdNx
tEp6nkhn44I0l7dGrCHC7Uuhj0pKnYD/LGymgU+6ylhkVc5MMV7ayFEul0TJGv3k
EkgSn97H1ODCYFkWSnKrie6XKoq4KWRqGW4wwTrqXh20OlCoL/klzZuGW58AhtxB
0OtMq3Q9/pmyZ8YfKeCoeuW1fZyWbs+fxJao9WN7mJ/qQckWDkF/WC6V7QV02fpZ
gmFcq8KaZSXe0jGcPyW3RaUXY41zbS3ez3ZjrWDrjAtmEEKTeswpkevw3FZH2OFY
htklSuFqu+j3MXsBPbNpBm61y+IjiMEljspPUQKpVJGtBEo1F+8qjahbHacSMqJJ
gltDuLDKhZNjADwEFVjLkoDuFR/QGWbtRKAaUWG2z17dCW9zaAP9grQPLiMDfeo4
I3xj5AoTuSlshXJgFmZsiS+zQkSn0iZfI2Aqz4jde+aHiVOcHgxbtx2zZPUfy/OX
SrvoLCbVOM/gcZkn6APIV57wGh30RjBhy3wf+9HP0WIxzJiKnEcvL6mdXkUjqpxt
B/iJDVRZr5y/8MkUvx/NkpQVtSv03K0ezF3+HomenfFsKYpvO66E+AF3nUtredsm
/hY3KTJouh5nsA5sOtnSbtAlHXgwtR5OGzODbvg2HhwACs4nAme6ooxbv2W7ke8p
MULl+i7zB0QaiYCyZA6/INu8LtuyydmWY968lU1qY1fXCvlogDpO5fSlXN7MUCl5
DZobizNYP3aBDN5vr1xnkwprX2iKXQgmTmN+SpvNJq5r+d8Ji+U2/EIYdVCp+MZY
98lJpv+dIeZyCj/CC8xN0eBXD3wNfgOOxoNjqTlHti2xuJ8Y4wQzSMSAgz7FjoC+
wCg4BU0KUXGw4+5D4sltDOZhwzlLzhZJpYhpzI7p370/iLu40iX4JQnUADm4laCZ
K/qZPeoloU/Jj4tMuCuG3iD32JrMMCYDQWDLvtpDx6eLswdRzP8qo25KvcdqMxdB
rrgcps6oU0ONRbwL9lOVuwatL9iW3bsajrySJ8Q+KtaCeEpsqzkdXWq1eeWjz5mN
a1g+ufvRnr/KK6+DaAwA/r+V13HQ7cv6KT4692TRENQMI9HUeY9yC3G4HWJ5Lgby
6jShViJ1DC3BzMd40ufscGWX4Wsodo+vcikAWCUs5Q3VqYS1vIGEWYDFjVHjXVV2
eMJvr5TM/j58Megcl7pi8EjdmtkORPCztSs4KpoqPmvuso5hy/SNDIB0J73PEF0x
qc7G+jxLMurU8HiyQAW6eNzkiAybW008bsxlk/CyNEXrZCISTnHTGFTAcXBGz1BD
Sc+w/+R9HhTpQ7vxvZT3/cSVJRKef6bpv2zUMIQPqLemmzFXun1rBkZ/ba0Ub6+u
rFEzeOWGEC263715P9tlrrgc5gUwiPUHV2m7v+S9u3tg+IgLKeElhpwccfELxBQS
j/s1hBH0VOZ3pI7aWnszSIGMNtOa8Le/p5sxUEMPb5vliEdOoGIApe+Qbx2bx1Hd
RIovcBUMvaiaa2Y0UlnruoDpAu0cz8jQIrvHt37uJ71TBT6+I75b49X6nbcQXaTk
nYl2m3AcehvezrmPz7jCwFlR6cBjZmks27aniBtQedApowOcEBi9mKQCzKUQr9kn
ZnF2Xq+o+4o36duAOAKq55Sm2qSn+9i960qyxI5UpZTHLuUi5zqw6G5G4avTe6WK
9N9AuByvnpUTK5gTTiMNfy0v2zUPKdbMz+y45W29f+wR2fqBIssoG5rgLP47HFZc
baXOzC/HXVkhLHq7Mjjc1QbpdVx93F6ljU09LvByG6GQ2KX/oCjSR2pYF6cZXQb6
0K8ctC1axbuEj/+f8Jyhinwx0lJg48VcYbBTxw8gNLeS0vR15sJvRUEXX3ZvuNt1
jIeHx/ypW/DSVnyyZ+nMlGF6DCYXjQqkIJQVV57NtyvTIQ4cNVEmgLvXK94wrZHj
nsrjehe0UAsn/OQ2z0+Qgh6G9PLlxn4WCRu8B0sMvg6o4b0yioxhpL+MJwk8v6iI
Im/MWKmTeYw7nYUZuTcDdpSf/HZNUVqNoHfP0cWiH7zPKy30a/e+z03Imi5icSfo
XlguClua9HZ+TaOokiJmug5smdzqeeCf4H37xzldKf7us+QbtJrNkWSJfSoi+b9O
FKbrfKsyFCeVd9qd5VnqR/uRiZJ1Tj0XrQ0BI+4/C6pg0pR5A9+Xyax6PjbKCR8f
DPuA1VrAsNAM8JoojxrlfK0y9eKja5XDF0HzMi1Y6SNWIrA+0SeaoXuBFQeY9Xeq
efr/HYYFsiMdJbxh3UaYbE5Hu2GlNnIWaD983vJclEzG5WIEjG67W07uwt5HDuHc
oz2lsHtN5BRXIHDKr5K30pAOPar9ighp2/+1Vc2dAn9Kb8+I001jcVPUMDhaMlVG
4eVz1YVnNThJHLbCG07ZTumRcBwv+faaHAWSuNf36uVLGV1+Y5ZbcEIx2KEqc7S6
YyTcStKYJO8tgytblUz5sDH1UQDEfunD4lbziHqjGPbJsvAO9sAAqlHFLoaDOlMd
mjodXtB20uyDgZTmtLhkGuLh3pTn4ycvPSkoGp6Wl6REOmzdVA53BB91RpYn6fUR
cGoDbzoeLiSYLsfCMQDex8DJlDprdhl0MqEP+bUtT8aIT4KcZUWIlyrjHh5w5cT7
czGB4XlKIareE+b0x6YfAye6Ezn5WAoqmx3pj7FcojjOgKZy+nPGGiZhtmdzfHTG
K1/d6+/DCCBxTd7LsfWzB/QahT24KrNkVkYzjnIw2HpT7MfzBLkxm2xuzFz7mN1j
i2iR0CP92WK7dSiXMrDLauQnMtrFwonOngzmyN8yvKYRDrdVwbKZdwgfk15CkU6c
WaJLYKzZQ375fkmQAY4nhMbmYhiMv4fMlvyunzyQbHHLjAN3z0KZGOew1MWTgoIx
xsERQifE9j05OLTmuAZssZxL/heD5vMZaNghEztxsjLp2WcXFVzxQCVfSdzkUA7X
87+h6tTdsDYkhl4ZkXr9a/6vLhWrh7OnW6b/ynHCserehzxC7vh15FypC2iG4aoT
6llU6m2yitCAb9zSEbdihLoTrlTrt+n502taOEAo4LT9wXaLHyceRzWM5FZa2Xr8
rirfN98VYd6RTwpBgNCMqR469MvUqbwsxwYSUyAe74r3AZUoYV407H/D7Ugl3Sb7
5xzS4ryqRu+qmindBjzJYGC6gHLPERqfutsv9htaxsRouVcgsBuRITiDuGGzS0VI
0RnPJIHDOUUGp4JUfeW/F2OmMYKlTwaoeVAiYvlskhbTihjGE+4qg8h1Re7uZKFG
ASpDyz9xIaTmd720qCUovgGQ2dszZ8+4FulWAem9dc7XBh4saT7hIiofnfsqIO2Q
SeupnsPPpXaUGoCyHqJWmnU6vfH6Z3jjIH9hUkXospE6LGa1KAQqK0MlSUw5X85K
NGvPJMzKhDRdkWfA2C1uD6bmSChw5cLq0bcsPGabO+PKcpYv5XNjX5y5j6Ud3wF7
o/Ee3qKy+RnIUpPZRhHXsm0lvU1rmg7zhdpgu4bS9t6E9VX8heNeZnzKtIDUGb20
SB6PQCbjYiDSCiHxL0i2AbDfLxbjms8jTopB1j9v6Iouv7XQaaQl7skk+kfzVPWU
+i53PHpGPn/aYTwKYOdXw5c75axgxUW0np2zAwA752Zy/iud9b8DevoeZx/fquEw
hoPOEvxPg/tPM9vYEq+hPJqmgMNkaAHHWvdVrWE4/Mql0w+I7Kkq/RYlauvSfPdC
F9ftq4p4GsOuF+sRa1dBB2LZiDNhFtyyDUsd+WSdxZF+0yjOJ+k5y9Qw5ynWTyEl
gMTI1joWqD8ToyPyA6SyfGJBLxvvrksv91A12Xeis2Xd/BGZgpwv6usN4Ijpk65t
U6IzqdE2Kirf5yuIX7dfSWBf7hZBTcqtFbh905HHyI4gdK5GYrLBMEJzhwSoiUKB
XQ9w3M0wxBrcStknixGnphmlnwFSFc4te+6OrOsFZ3osS3N27iZaEhGVEUup1+uK
vh9qsuTe/1/yPVHp5MBTgLy7p3vsbwXh0PqXHbUHZKYZIluy6aQdF7MCyyDia5P8
XneD3rb/rklZVE/jrx4nofkLHQNDmhewkmr/bd8lRP6s9Rhc2Tc65h2sQuRXROAh
lp7XaCgo2tGZsOMQtORT+veJHdxMQ1Gp0BgvWhlDdWlxPbLKf+BwTUjd72Y7g6m2
1/s7AVTGyCKarOve370yM+mSWl5lXLFFJAePru9xxlov8Yvle9+U1NgpzzsAi652
qjY72b8nW1tzIValW/s4LINDGvQSnK90+PrJQ5sT61YXRWX2bfUJGTI89siwugXt
lJuLNVOlpCqKHOI0vEw7u4nw0fjEkJmoLUsFrs7f5sg1HqQWGASYT2jI4A5De16G
1GsTRx46RLgKuGOGnhO4GeUZH5xyt2GzzFTgQeMaPdLi2S3F/9BFdhKGrPiBN/eV
rQ+fB+PMaUUrsrwX+oW6UkOI13v8mNE1V3kqGEyxAkZC9R1mr8cLS/hF6HP9f3Ib
8rgjyj1n9W8q0J+1ku3XE8cp0FzE/ovHAXipWhr+G83yVkO2Nfm6yGc5VC84l8gh
OzlvFDMAqAWPAXs0799mpUpoiL0mkjVUXKQnVX/q9B77dl6GfEZPXwLSjYysrY/v
B7vi73f1AkCRpidcj0itS67Zw23HF299J8NjhgrNfQwa4Rn4g9soRl+G9+zg3EC9
1Yw01j7oya0tmtLKXmRmAsOsdPQ+auORUXBQNkN0cA44ySt8+msIAQwPNPOVqGpq
A9AOzDJ7UyEXAHP6uwRb0aiVqRNZliMvzAShuYkLgRRoZZqlFH9zoDMSBUmISi3h
xbwF+BWBMviaK9JC28uqKCo4I/G5P1y4ON8x63JmQxMuPpJf0pWLQM51/skf8AWH
rTpads/TxN6aHif42psLO7ZRsNExTraj5vQnrOkG7fpEeTKmQo9mNMYlJeHNkOoY
ciUm2/4z3B0uXXq1/ant4qL16VZbT1tzsCs8FUnec6MWjiZmhdLba8KRVIRV4rfM
CQ9vYedpYM3sKLB6lwGmRjh8A/xPY+qzJmI6wNf0G4LhPxwnnhiz0CYmdUeGTor0
loliWCIRkMcN0VMqCse9YzMuHFeDnH2ZPF53rVkSASlKyqSnfmneTqxgBAuVc2tE
8BYbzNasSr0JZ36jFcum93U764WyBzACuBfPEQoQKWpUhj3qcaoZMv+53S2BYyNQ
uvm+DnVhWOQaGOEv0GBEk/noeybAzV492cuPZT5nWafs0g+n16ecBz0PG3ZvgUJc
sGbFfIYR7FtOM8R1tg1bekiUb7YOl4rmWxEdkffEjjj7Xw05qDktw/MVlXVV9mqY
fP4bXzfgs5PQFzajVdpVeAaFq/fSdxXncFNKbXcr6MSI+gI6i2nYCoYrjvKOWHLf
QRcIZfC93VK4/ESZcbDHQmbjRxTdcsM52sz6kRGEy9ZQVU3nejBxgbXEoUn7YBHI
wJrrRw+wzJnnaI/tJQpBVm6PyB7M/dhddx4ejxO92KLg4qDf1zANI31dJD39g9U6
DIwbByZA4kEFEGe+a5FtQWg6VGq7ilEd5g4Sx7eUh3DqWn9EEWmKykyIMYKhLVqL
2TDY3auohtNUsBMNT89GB/fdP4T14XC1+YNfuTC+L15GZLTf+gA2njPaaBLe6jfa
AM1z6/xGyNvWjmxXmGP2ColKNUmrBSZBDPdfE9OryX29BFcWSjx3MYgSv9bjzJOj
kRz5qgC/O2FL/HmqmsoiLu119W4xuSMEXezBLLw6ELjW9FzHIJYOva18WWw3+E2d
9q9IZINSSnh/jbxwmzWAsLL2oPeZzGTrR0Q3+fh26QZkQrn9mYwIeeEaUAePZELX
tITqIGNIq5voUVALL/gCyppRypilzgkC91ss1HAI7StizLK0NIbItEfK6VC8eEkT
3sLGvMJ+i6RrvcKX/ryfjs0xdBR7Vnaj8KlUi7gujM98feSGKZJ+ryZ0aJOF9dxb
ZqP1nvjPyW7eLKpo2XX1ASnehRdwXHbK3Cdf+kv//q8Q1Q/4+vOEUkj/sR10jTcf
EFXiHGIqD14m44tnupfh+KJZqerIFrSYSncrn11wd9470hw5GZafVYvAwtA2t6kM
IeaV2oaUASBc7j8DXl8HDsWN8O9BTQD8j1MdHRqnYUOvyP/CRk3kgRj8FhIcZqeP
3W4bq0xG7sAUVI+i/KgVK3H8jzWMLefELaNy7lBRIrnwr9MkVL43ikKHpnJT3Dyp
/UJv/wzlmh5+IQGUi1M6dzD7kKThQiTvzJazp3ZkQOcJOUWSEhwxcG+Xvvmw0qcY
oMJYWZECVscS/Q2YlcWePDGqbpx8JICfshbJKp6PcNz0mGURff6tnnyNQyNNfceP
ZSOBd3NeH0xLY1Dt1N05kjxPQELBFiNTuluhiEG+rQ2lCvE2kaoFT/ukqqQkiODA
7poser4wr8K70Dk5VqPzDun1PjAApT1PmNBkTjVn+bhnQ9RR7QUmupUKq6Cp3gp/
UkdlA+tO62v9O2/xJdDVp1BUgmcvwIZKmzu6OE/Ll/UUtWgyLbxJ67Okxwcfk08L
XhZ7PU2V0e5iLBswY/A9vR6QLJOp9a4s36SLs/ftwUT7JSsnJg+pe1naFQjNXnEW
Bfd7PiUUQfRZ8zy5/3altbkAbkgGfceLOxgXuXXzNqV6duI/p6grMLuKv818JYL9
P5l3rktnCCzMOJ/shMFyAifqPAJpUCzCPy8JiaiXuX0xnM4myEPjkJvjcEPCIMvJ
qgNm/nqlGeZTDzv9xO8MkgvyKJcY+7gY97Xj0un1iF6ctvgbEGjlLX1Orhfjbv0c
KPjl0mWi41MW4YQru+GoSOD9LGJ4+vgi1NwQK4BcDVlbJYXBFto1rWvPlrgBxrzT
1iB2jA2eyTcHgl+vL7RNey1XKN12NlDBX9vtw/C1LcVIQtGmhdGedIDDxNz5LGK9
7KKIzrq19xsZtjN8hkNINXd1Oh91KY+YmiMefaCTJLz92O/nQGY8yr6y9aIXh7Ly
vs1T9DXrazEyxoMjY5rK0LUAXrROrC+eej/Kr7L2jIsO6opNHZ3027X41rrou1+b
1IZBtXWrpgs1FmtLIyvkXUmH3Km8bJ5WnHEG+dBKAT4NjLEIfBf+MrKnWEWt8+Wd
k84gDIoGzh7wGFJXtshXiclPh4yfRAHs8Ax2rwtJG4cKn/OD+qemnfzBBekmw+XI
1D7yRaqbMfMmXgiuRAI3IUbnNCqYlaTtuxhT94An3Drg6ovf0BlsFZTqPJqOJqVT
viVXBWmU8/FCXne3fxT58wNRbNcAZNUAnQXQkW3qjkmCeWHS9FxIxP2E8yJwv2J/
VL1fx+1xI9Blbw4bTmeMbDcg1M1v7qYVvGtFTs/NdZ7/ZVFpNY75kSFFLPf//IGV
uuKKZh+EPAfbq0IVJ0q8CwSO3uu7VogvYd0i691EQ0d64Fuz1gsf22Qui9j8mABN
4aQeWnY6s6niVYfXJlodPqY9fR9Wg6TcjaOnprK2XGq65nFw8jjvruZtIK2aN9gO
a+WZ4fQfba2h8fpdJIZNB5CzmesJB4wMcrl93IK8KCsZtjqV/sdyce2TCUVy/IVk
HG5hVy/wfMe9X0VT0+Y3Z2BbspqfSNpN6Q9hTDWRZH0jV0m2bBEfdAZYSDydFQbV
mVSXUPKn+SwOmHkHfE1gQN9UDmPhe4LA0iW2qga5vx2p/Y/gEM8ZNAbdalEMsBKB
2XVKqwzD8m90yNnUVb42X/e59r4ZaVmscnUaaW4S3qE20RR5B8of4oCqMI4n9Vvl
O6UawsseY3IQA2bxfjgEk0ttLC5jka5eji/VBOSWYfZUfdu23hxyi2RDLy0TSbhO
dLK5XYFZetzszKyInhY3uu11NhlEyZNixqYuzg2ej7vHPUFfzv/xjs3apXDc3Nhd
wQg3ReLR86r3/F1AAGMb7jcI1L+bygQ7V+hUgZ701xqTtjqXbC/DXetmsYNYr1/l
K4KjaugA7MCYVsgXeBu8S5KV0Px03L9Atf+LEOER4Iwu0sqJElcX/ff/9MgDLNPu
8AIqOBcRu2GNQvazvIXqbVG1AaWi8trZ8Xea77GiFtH8kFqSZcJd+IhQbaTQUUbF
J2kyhB4AUzplRf4Mlz6WZN9WldMLAu3+Rhzg/5w5PZ6dfMyqjNgV1Dg+ECH5s5u9
VAjeCGc9ZkK4vTirXVc4nUte4AEqkm4F9FWXguKoJOGDK1pbkmCHB0y12sRt2ttQ
ZFkYSfXXqIpT12fvPZtqZG8KxsYENX2nV8bjteBq79j2ZwlHFkA+LhbxwMJGATDN
MxOmREAnUSmgzbLvhjJt2Geb2QBhKqijXLN5l3BlwuUOnmHWDPj/cmVq7Xx+RFHT
g6rNrm5xFtmabKzcKSwagKynbxrSGFPl55n7MHy72NLXXG4suDsMjwsRlNUY7gi2
ZDdDLNXzJV4EWeG386a0j6dbClG14mfJtPDS13kc/rF8x2Tuma/u66XboZHCkix+
6JsIr3SWqflxsmC6DQZjlZc7QPJXA6GIdqObu1Rhe/j5fFX5AWq/V4LnEruvzHYo
EUlSz1ZSAgQrQi+MtDoZgsFj7dzR4r1TQ2K5LlSC47YpGGRnLcR6881dX6fdEXkF
sLXD1FP+r4DPlWCdWIZr+Eth5DejXue76tI6f9b5Ys6Dz7z+MbTa7BQVUR0ewMNy
YWvwbfxc2ct55NnyO+QyzWjIlbe2+P9jNh7SibChRJkNGGIUbxydR9lyVMd4TSMQ
OMZBzSzS+Xs2RILUczr2fBIP239n2anQKntOUkqDOijSEoLrhWD9BRF18EBqX+SW
APv/a1GCcGMauIMk2cbuMmtyKV9t3BgyISdNsiaxSCcSZmF7KPxu/tfOA4LZpjPR
DGv167qXeHFeoJMoB4SQ2MrvtowE4eFq52eIop67D6R1vBPTUt0Z/RQdfld3aKYi
`pragma protect end_protected
