`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cT4A3fvsRbW6vouSagkrPfuLHJQhcy5xwgGpM6/3q7Ss5Ng4fpJgpHBcHT1oPb2b
BfiUGG+pwALmha2INjIda44yRjxZuXUj3VnnE6NG3fSzW2Xzw1dPs874j8mceU20
Yj4lMJHDIQdndRs2b51geTfUl+oSWYbxMKY3Uco6D5I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3280)
0UNka/57w/DxRkuznU8y1PkffeG1fA6CI1GpZBbj1qF5cWrJz6fD1YD7GNxRf/94
aty8IJe/4NkzOUPka6soU/5kn/v+beeTZoN4HXI83hbmz3SSO5kfD4LPr5d0k4Dr
xyuVWDINn3Kfepy99FgLMZA3xGzAxS8Le8G3kGRRtFYQxrCbUW0yhD4e12bk2CcC
zELcM7cXMXi66ugbCr/HUVSvwpQAdr8N//rdQNMAHDlH4RJSCItX2WZMTI/Eg2bd
wMX2jd/6yZmfEltdZUgQe/coBjVDLeNCB+gPJI0Lqm130glxVI5Yqcw0UtF1Q428
oqXozXohZzTyRHnNq/soQmh6GHR9n8MfJGTBpuaKopKlLJkk/T1qDR7ttaYDtg68
wfzs/7mnI5oMV0+OKB5GsKagvkIh65vdLrLt75Afc+mmUpY8FunGHA1W3QNL35U9
jknIDAAsOrg5NmU/YNBDdT5ezTkboSE/9p1IcZhv+FBL4usEaeBW//gAu/goHKvr
G4petNBhNeL0X6tQ6Nkc9GmkBmnVrAZureshPLZz2VABhEizQc0XJklj5VR16DEv
3g4nD5Xb0y+snJurq3GF79zwGmjlJzhLlld9Eam/5FxtigFI2QVBNfAu+jnc1O0k
sAc3AsxU3Bs22EST4LcNFsA1sLhskbnktEn5Q8r9M73bnuLFhaex5pMXazutICzG
ze8jQer6c1rIGCOmq056jT7Kc5FMikEJ9QjAQ2hVySgzpU3TnoFS0TYdCuDOX5sV
k+z2K07eY+Fq/Uyq9OJvscYqF8IiwDDfUcenpLQVbpI3nxmNsQYSZaawhimZA1g3
paHZxOEmTEVOvzhEYrPI4KnFP22gJZSOoJLTIgUuVgXJg+EYpXMP2YpxAOr4vR9a
5unwrBsxxC4VaZvSN177gpLk2AGZU8lWxIB3Hv/lrvWkfHTHI2mhJuXngxeAsj5R
FFanGIOFCVxNDlT0kzQcYfHGR1PTGhX2FJy+GhmcqEIlC1dLcaGmPA0oCblxj3p+
zoiDHu2KqF+EHb5iEUCyMsRdVOAPqBROLuuYs6J0P9GcmKwyqjY3+9yAJP38K/Uq
GJ1cm0a82p9htb49/wYsDJahueMqq6zts2gAmqjXffrlAfldISkRqpl6qFiW6voT
mi0T30TmlBwusVdeIJ8UpwvNSv9PRXOCHPkokHfPlb66M9+DjysryWMFA8mr080d
dChDl5SFNA5GFvcLL12/cZB85gPeiLYDbIymebF1stv7GNogKRbQTzTGH48PbzgT
irqY5eDDsEyAgTq7wagiFNWN8mHYcygCd7SPS8W89mEEnNSfUDfePhJwcAyWs9Gl
tDaekI+5fBFBcHH9En9WMkGCYojbe7NmejSsojL0bcgPubGtDFGodUC2nX6TfW2K
ltVsTF1S7f9gLjSSB03DVq2TVSVXFDXbDdxW+QMJbHFWwijuX8xAhCsQ1JKoE+TP
IdkevHzVRUd/LDKBIn+OjRlc9M0zUNk/Q6UwVlXAn5s/YE0KmznpgGF7F8giME+z
4S0sIhRGXBF5JgHvpJetVGgYVfbimAUbw+WWr4XE3T+8XXCmL6u3ju9OPSdkGCkI
6G9MSyWgPgwAIHDt+WRue6dbLVC7ychDPGvx6JNrLV6PjdEVGxj7IpZSsu/FF2b6
Lub3/23x106fISTGnrDVkgujduLV00BQqB5wXYw2LB47i4i/4YD2CHnvX1i2PQyx
uWYpFDSJuBIKkqumfvBDXi6QWQSdOA6Ztkl4cCyQvAPT9aole/o6dmubX3BQ2e4v
xYhdxPvbn+FmLeNzrmY/UvvFPzwSCMsoB4sOawfo0LEMN86R+8GFEI7OWSHq9p5p
Z6nhW8J2cEWm5j4eoLmp2ePhPHFMrfew56B87lmBdDC48bYFc+Mq7zAqAxoxz5EA
NTHJNlEUrK/oWMmsq82XlmWjxNAi2+S8zhFccpbP7ugzJaTzpeFMBZqwZi5eBA0j
NUF4qzEpq0mAiI+g5Jg3dUxTddM1/CP8wB/qAGtXn8EjYvaeESYEuArfq0uT+KUF
4k7yhYVWYfDacx2j4bG/lUk92VO0zwC0LfC7EddOkCcVte7NI85CNkeHPM+XDrbc
brz01AaMnlpLaPVAznnTwnvaGBoJVRU8w+GMTfcTKDUoWvY6ya5ILY2FHajOR+FS
20UJTQnp06pxE0yLTHlbcOzsP7jMS5ew0Le+35LTWm/+QMpkXin5mcrEo/dip7fE
vipYhokwyAjWDTEGOmumMwYgUC6lCDMsTsYuAA3lgU9/JUAwCdHPSaQJaAuO9nK1
0Dro3ASBaoqVum8KBPYRlhv1L1ISiuRuwlhXVUtMvKOiuGjuWOx4VW+O+0LQ2Oki
PghLG+pkIDMJpBQ407QI9qpff65Pis2dMBfNzQoPuFi8ENRo6tqMEGazQV+45bou
mzevHn6dmgB3O3xxMuVv2ZeGAWojOhczCkto+KsTEOniHAvGrtsVkHT2pPq+LY6A
cI14+HmUN46Co7pTl9fxpu4ZUX0mXeI/RUQzz63TpBIXpINE/ljtSo3ywIJ1GPu6
cCxA+gaXVT6uzf1tUidKioaKdyWJYC5FKLZGRYc4LRt55vXzM5Gwyaze7OFu8LtT
Jqwf3NTH1G85vJeJNmAIm8y8tR01CT1deoIfQNlaflvl9DjR2c8dYh/XNZK8KHqK
OgPhsfSB5/wYku+Vwyt0PwjMsoS/kkUhh56HDeRp/4OwQpmu5zPW9tl57zil5H+Q
GB1nLCPdeku2VCsB2zVO3ctoPGR4rZYimrzQ7G7kYjj0QZqjZvTrt3WVaxt/Efgk
JRhjHb5LBaK+MfloQtbuVUxZHfHayVbksad+6qNGWOhh2UScS7NCEv+kAtORwIO4
XfyDc4lqaZJ3PrWF7OuSByhepmw5A5C6KPhf44sof37RC5UyIhnp8WyH7dtw6A+R
yF5tXnd+zwM0+jp1k3GRS8eDMvw0dRt/REs7yrw12Abvk2XPGlmpUhAqsf2qlln8
DeOl1z6Egp41sJZljOfQvOHQCiHlaOtPj++StA1ZVpxwkouyB8KXGno91EnUHXyx
RHmjz1t3vIY6x+VaQFSZZh+t4pi4Yd3CWZZT2kcDuNrCM9ZO8XPqxBjZjPqa9BfW
QVrcCV++BA2cl3+G4M1a/81Sv9k/tTQQhwzK+1xL5f4jS3LgkrJwxk9hKTqxNcKl
4TQkCfqQazSRRgNjtaF9I3jUtNx3SV7rE9sslNk3KnKIH2SCRHD0e8zwy9PBxwUU
zYdOgrlM37Vn23w7OQblrAwY1m/D3ezgcAe09FTHTCuoz+wGroC8rdPP0KFfGV90
0z0Dd4+rlUxRlUXSy3zhDjy5DodFozBfPICNq5Sz0tH+jP3zlne3B+ymeCiSbXkc
1dyKU/7Zdmbfu+5Za4NJUf8xp56Y7qFc5d2jxoVi+SDY0a8KDzALdhhNpma9UyD4
M+XAAZ3E0vFbFsadsbYAXox9XkkhJr33lcop33JMFZ5yMHbNh+LNli6u2XoRrTRH
2IQh79v+R+Olo5/7N9fAbI7sjdn0S5OTRP2GAOaE9BUPLVcbAhdzs5HVg6lW8nh6
kQQ0zUoyU1c3laO9ry52Rr5Eg2gv1xK8vR3DWnHrcZxlQERLSJri/SSssnh7LQ7K
xvBiezyRqGy0BRp0Spocp4iq3kTawJNZUM3fGlBjLG2P+IQmldctoB7Yw7mx3c8m
x4r445NYOsf6JyBjHZvxpiQ5Hb/Yx5fzQvTTqs1YlORKRt1Y/pfpQ00dAV3aBphN
vT1B87IdCJatEGNMLMcaIIoQljmxe90RGQLgEl7M1Pq0FOHUewXnhWnyEPFP0tEo
PVaR2KqN3bR9yNJHarGuldi0X0r0G9MXWS5CTVKDHghUwJR5EEDMInZesNhbagb+
QuS4uMOIW+Ib3O4Eoc/2f8Qds9urDkL1qsxPzk/x+IrRcZKUBU1vm+UgP0s2IOiG
1sGbvR/t3/V4DzCXIicjrAmS89mK4PwdnMVrmmE37YDhk6WOKiyIBlHR4gfRHJIf
kQoSSwAyfqIDT2xABUQbSI+do1KSy/ehzZfNhdrLf0kK+xbDmq3JCglsIaWP38/W
Z6a4myVciKRPi6MfgKweii5c/xSrklG5iw/z46ViYgC4bhlQx2HgOb1ySa5ebQVc
xCREnXs53zUxc0ojkOLjbaq1gO8W5ZzTqLOBejcWG/a9YUMCxHtD/sFfshgP2uPM
H6VEZt7G+W6V34ShJ7dkZRUJT13hwSPpoUoxgJ0wehpTVXVxwCoref6HYnGGj3Qw
yK4aXZ87IIUIPvLH1j+qQwbY87+td9J/b0exvdaWXR5Hni5ySjiz1cqTBWu+PZx1
Gt1rlkiaDg2mzkDLZXGckg==
`pragma protect end_protected
