`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ok8CwbYBAuFEZNRiM7LYzyxeODSmj9y3r8Pkxa9hqQBl2jGxB9suMP3oax5RsHBZ
uaF4hKz0lrMyOMXEchnxG6eCzqGepYaBshcpR3KdptEBSy1Pj/pK9WOHu1jNvGWo
XdiPmCzuCcQ3wXhlCJrU26sf4i0THJMzdLnKF0vdvLY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
zPwd5URK40Q9s+K3os58RQuenuKd7nCRs2qNqXS+m17dbygPOzchJ5E3D17aWqqY
kQZyQbyrB64t50lqoPvObygg85FQh7I+pR2ALSJmN/y2qseVedKFwiJa3hJLi0Fw
HD8DmOo26Vy2NCNfaYGT/+fO7UDLKt7lK9JuDg+ULRnmYQrXrvpIzfd7V4rMpFWc
gMX+2CGyxDu5s0hrnSXcQO+XI90v17bTnPsajgj9uFgCByaWjH51RQ9rDPapmQAw
9vPbD5RnB7kLgAwqQgK7NDTlFD4kdNJJcY9QONQvtvUqQKiIcAT6pxG2a/TYtPPp
bdZvcr3xdgLm+QjXzDkfdSUKaQYTZKmrLq5F01i6F0bAVQCrnKN7OI95+2SFcBpq
OqQY89GXwQztA0V2P9Q9uB+k6oezSQpxwnYa2CPVkol5WfgcXqYzVEM8stXS1LYd
bJITYQW1tHwMc5yBucprhM1oh7lL6Xi0oBtJAQSN0amSkxPYmv1WIjy2PMJaANZ8
jkqPNasdP1ETfRMddHUeKwnL3Tt669qip/Wh0Z+J7/2w5lg5pa5lgww90i2PvC9G
U4Z/WF6L+f4/pg1Kf55WY+5HhBBBd9DjTXre8C/cjBjyN5qsjN6MEK5FnvnDkecf
rhZHS45utSaM27mZSeW+m3VKIKrjBAnEFe3LDhV+Bw3qjqXJiZmYMhDndG1dWyaF
o/gvZYRXEsYzY3b7y69m6zNirFKq8KLKr/NBHhKWfTp1OaZ9HQlXgM/FQZeIIGZy
Y2Sco0MXYT2ByS03O4mms4yr7NejdZ377qAl/sbI0kAnoMVKyWVj/+cbrizmTo8B
rgU/WpXwv+wXUlR6QNvPSveJrx/90cbhZGZUAaHW19bbluP7SfEA2okYxAMCleQ0
6yRL2oSYwyckOFheqgYpE5WveoNtoCCgETXOF5G7eUReO8NtfwKI+jNS/xvYrC6V
kAzPbtVo5rILX8im59MkGl7sfF4gZMcbnY2Bu8PEbGStRxtBFalOgXFIxlqx1tDR
GHPa834wlwiI2J4COlYMY6h84wtW1d+3ABIk+qFjkvpvEHbkz0NdiHBcMlwGNkSo
97LsDfoYFZuAffzeII9KIr33pdUjjDyL4ELH50DRCjzfDRINhZRqdshS40lXDalA
s16/zj78Jkt0nTNKEn3h/eepyik9ISkjWdNjflHAoBf6z0259aVp/wotLh+RmdkD
L1qGa9iePH4Y3GGmsaR5aVLKK5by/Jio4a6Ef0x5p9Slw+6LfB4h43h91O8mIbaA
aygwqkZ1B5xG7ocaBXWTTrH6Cvujg2wB7e7rvI8M/t73tu7FxOnAgTBsNntFBeXu
p8W+nLnewkofbPe3QNXkLS1NSkw+cDrCAEFnfsS2Q28ZxFmZR/DWo7mZhvQCypZQ
C9ShuDp5BnPSxQ+9e08fRyJl3+7RzAjJncMBrnpAdDGaasd0iYEqwcaJN2S867jA
IEpXrRfdmF22oxb/Gfgix+Q7cc2tEZRME3/KYoyO017TM7xUQ6Uwi2h279ASa22K
LHO/bmg5qQF18MIUu1kz/rGOLgZDQQ//Oi8EL98OwVZS1ntLrrfkCQjWVNbK5wYt
Bc5WDHe6yDYhQbn9HOgCm4wjRZoEOeKr6gcbxhFw9ILJ+NDSPwylePQWW8sRB8wc
R1AuPakuVxraWDqd8WDuYomp7F00ozbhndANMv5/MpPMW98ubyCqy3Uf4CBFfwcy
SP+ngPxQ6M3cO/tBnL4d5cQcP4Y3Yw24su/5Rr6JcmmfPJMrO7ToIlUgCEist2Li
6FZjHRlhh1TQG5qE+96J1dffhHCZ3wW9wm4lySXJFWbD4YYwN2hzj2sq8AuH2T3d
lIkQGccVs0QfyCS+niOmV6x6OVDBk5nnGcaJFI+KfiZHZ0GEItOr+mE3YHbfKelp
H2MgQDsmg/JVwICiuzley35MawGecDIwTf1yza0oGpR8PA34p5WXrmDc7EJuALGK
XZc8fbIkfK2twJhL3OODuRjvBlJnWZSyIbJEInKgbVkz4Ez59yfVpEDU50qD/Doz
8SDixPLEhjcoAcU/OUTsbRZkQ0pnBb8Pu969M2QG5bOaQTNAeTPeBkq/fTSXRERu
tkwcVQm3N8PqPlyIAnaaNuaVYJrWQVq1as0C27HUpfZIMpC4C62Y8UON2I7IRHMq
iNiaSI+GakDQoeWQFK7IOIwGsh0ijeyrrFonT3bpGsCZIhREz1oikrVDRbtyYE/C
eW2ggdIFuBS43bg7Uw58wn/3g2f5Kz9AFIJKgp09Ttecnku62aoWu0yYEUIl5k6g
kSkLbpfBoRTDZk1gGy7m+NEkFbdTDB2bNNHTWXdFFDj7txM3MIG6Qa2Ko6Ed4oQi
iiCC8a3hu4RdX7FaPaTiEy6vrrmZLnH25VGscED95umIiEIVeDlfWGwH3Ahb8OlC
iDSY6ov6i7NOUbGKEQMYuX6jRF6To5ENwdajiDiAj6tSJwAu9fnHVwgfkARvIlhZ
IcAoOJFOO+Omv79USS8Stub6HrnSpxz1owZ3S8fiWQ8lP1PLcPDdfD/D1n5nRQXT
S7MBL+igvxgAOGmumTtZhhcYX0mx0ptQxs8aGT/vCr8Ra2M1k4nSvGCRJHk9+4Fl
rqj1TuzECHE+uQfbgHmZOAymmUfiNyX4Z+zywiF50Od86M2cEeswednh6y9o23x9
8MyJgDvFSfhFZ2G2RpcG3NbnXRGkP8n4H2eFgRwkOdgo7Py1L1PK1/NWYlTJipcZ
3aijCvzPxgxMpbCxSlQbxt0y0DUqQvr/LHbyO/VItO2A16BWa0q1OhOpyq58kSOB
mDcM5GQeUk6WD19//0JkFvUAQaA+ZgZLBHF7iU7RLWkTPBhMkOEklomGL1QN5CpB
qt+xBbYH3WIU5B3vV2/cXWLY5H6RNHR0r5yukmHzHu0RLJ37oJSXhgEfYYKfNg2K
xdz0Z7NMRAfQenBe8l1TD+IzOVAAWtxCDPa5voYYYJct9IDBcUSpykVfQEZLxLjC
gBA73PW8kwYRwPTx1g0Ew6EwIR9dfSf1HjGmUQfDGem6rwuioprdiRPVhb21YjSb
PJXh4e/z1KVbafCt/SD2O9XI2Ib1ex1Me21phLCmaZJlh1Boipnupqjo187yQX4X
`pragma protect end_protected
