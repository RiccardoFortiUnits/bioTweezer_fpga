-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
D1pY1/gY4juBoziza8YzQ/cO818lWLX/6Q5K0AkbnQ4YNEoB8LR+82ltCedCI0ERZ7INUJTxUi/6
7F3nNI/Vqy19Ge8WJkyWvwMFrG3/mJs5jAOfRwmrIm3l1qDzXRutmuUFGyTrIcxvEVAQL8+jRERL
Hpl9Wr+PTbsZTjur8HUutipFJmQ1l3sjYgC3QlH5OsPW0eHdRcsVIxWEKNlFIyGvKTXPBu4q9aoI
F7P46org5Ami6kss6l8F+eC7DhFziNN560lFmwIan0J/dg2J/gdA5ObdoC9//z2032T9cpru/Wen
7rdiI+Ga9qBYeIoWq11MSgOPwuC7xKMGqcOUXA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8048)
`protect data_block
xBXUuHy2038wg40H5OaJhWG8TeRe6Mk/ZiIF0XLP0VPvndWRH0JDueSf35IsgJU8qxsrp2wYFe+6
gLL2zaoSR8QaTvUXZWSAcH6nYmeBG5JCAEDZs98GenrBjR4AppeqS779m8EAEplT/32cm7PVSzIX
MUtGD96Oocs24Y7RZK84wD6ixb3WmQLG8vJrmiUe2g1QonShorILT40FG/OzDhHd4j31j2V1V1z9
IbsoLH0/0k01l2ozEM0pJZ0UNUyRtMDMtdVE0FgEnlhx6BsYJxc0of36I+2ALtPfoOFUXxTXveAR
ReLK2ThaGuHa1u50SWA50Ltw1rfiXJ6vTCtkzAztOUZGb8FsqGvyw02OZgSiQBvgN15b8+kFtCoC
iwKVsxv47V08sBo6ThyYWhALdzJQxr94cHciGglmh1wTt5+AWQoWYDW7HmKR+3Byi75ydJmEGfb+
8tTaHfnj2YsRgV02lsmQPRJO4zFhC6yi2kvsSz+NWI30723kRVO0TIERJjSiRVsXzCEyNkwgLhml
EBPleUbu09oJNTZjpW7IT8xVGDAThIoDfhiTF1zRhSFKk6T1957sVAQ4CoaPNyBqZMAVnaRS3hqO
Ie/bIA3Gzxpjsoe6kbfk2P5YWYCBLD9HAEfwPd0PkkBR6v281FOj+/AKKDd7crqzB92zuIaHPPYu
6BMKr2lNm2ILysO0tLMpioFUBL8qIw+enxqT8hlWvEQz7j0+TifeFPr3QdU1Y8g0lurHdkLDL+xp
oFZYJKVL5zAWLoWMdOE+cB7sN4Io7KpvDvzIaAbGuYvrFiO++2Wxl4u5jdkY3UI/aCz8WRpGXUhF
MOzD2tUnjZXCFkbG2M7zHI9gPJCl/Wj0P/ViGV4fC/QI67SwO/RmE66A5Outxyq5YRXGIMEdRjJ4
XPEREBM5yGe4Dswyv0Yz5E66bnBqruS+4rgDgkWVe3IVz2yKR2NJZaL89rTcR0hhh2cMepKZYC7n
nqE0Sw5zjnJBzxoLNsdEtWNQhhYoZkaEKaCNgZycFmZ8TMxsAG+nbgl04SiSo6KvJx9D6EScAmx5
+FpFM7laxeesNaRJKSYnnO/p1bpsBBxcNbqbHnEQgMeWfTo/7jPgOzekYM4EeqLZEnwhPbfsS9pE
ghC8Bo/BdnRBm82mjLBudZA7At+U3s+KsQyPusiV03V0sZW44Ee8nzSlqbCEl1YHwX7GqMyVcRnC
NmMg4OFjaMSV2504dE0MA+ljCvkKhKIpSfoE+L800rCk3icQpVgo9wQTTbhe6W5bUA+drG8ib7ea
kqk7sCflsbpBO7wJzqhpLuaOr74fZ01/6SU6FvgU7AOwPXdkFP2fmWczyRTjKikPaQnA06Yv1Gbt
B7+NUcNNWs8Pm/qOZfL5gXcQtzefaCvZPHBVjUPPwHND5w/bs9GVcyzkzJckYoM1JkhPt/+kMSyw
XLfKxCe9jXsVFcMktJudwItuukSPxWTU54z6nOCYsS96tv1tzyXoYQh7NUJx5lUwjN9tn62Q3pRR
KQNEhmMKyUYxz0F9JdlZX1/nRNpqhcZycfL7Gbsf5NfSh7nQFUDK6Fhw0Wlbm2RMbPFSgXS/q0QR
Y0Hjimio5vUh4Ba8EXrnU9xl6NTvbRJ88XkGfDF12MTYtImaApKYkij8/sK+I3BLFxIRF2WzVdFA
gEtEx8ead00ftgizaCI2Neaq9Ky50yAnzUZqdtoCWOqeKDzufbBr/CZMbMKZC/V8DqXJNGxUvbNz
cEby1VIIR8d5VoBMBVY23mXJQTyz8+LNwt8QYkAHeF/khPV7+IvgVxFlS92ne8nUlnSHcJ5Cl918
g0NqjqbZR8cS39NZeejaHjQ+WNx+OA1YW6O474+V4RWT1G80hIodYMZvcCWRdcibKgWBFt6OlZtz
cW+9apL3BTG5GVh7cs+oHydAP1fc8ZtHFU4398FZ3q8g6y4xRD+NQZ+vKQzKDQfmuSzV2X9xl2ZA
FL9Yr5g3L8URewcfw7Wsj1TE2vMjFG1JCybrd7vr/N1CGxVZQpn7JmcGwE+sTKtyRC5phOCzYKb6
O8Z4sS66wtrZL1CTEGWhfXUpVLP4o+DzKG3eiUzg20/HQCQTvwnGveC8lOfbNMc0SHkeUidAB1qn
hBbS8XPIOAu/k2QWM+uH5uIe6UN5MwYe1TTNsBCLVj0BCvBogVOSNxacb1OKwsO0uwow0cMTDmn7
+Wf143cvV0mVd/Sgbu4+IfQVvgIqQdLzU8LBMHDIG0d24KLM1nVIUwS1SUmwDHGu29dAklnmpWzR
ECdOiyW8KJgc8lXKuv2yRnfUgDcfsHdTsJBfhZkERv2CoA0A+Kb3K8JGA6Y4QBNR43DqwOetXWbo
FhH31afahHcjnGIaVpaIEUkdb/0d/t9dZbCMMJ7osaY0LZe6OhmWSYtSJsjqeu2XFtYtZveB6ZAS
QfVC/AbDAmZVZAJuHEvE/rWgJSsz0bZFU4WnrxoJIzOoM8PA9OMyTQuwMZVYJiQdWsLYb0j0Z4PL
qbKcwZGDrhX4DNhh9PlXWe+icZtNb+uUFKkJwBBunSlAcDgxqmg9PkzUtiI50d5ZTUFXdsyTiTXW
Fh9HMsWlypIOHny6FFCu+LuXs/Jka3kHCKzBuh/V30ltpmpy2CqQ7KV4epddoiWUR7/W2L5FkzmH
Iwt77psw4jWmP3vaFCjLa4LQSgjutXE5W2u/SWpjHD69Z7ZAH3Tfpigr/yYAgoWeGdO009W65Vi1
h5fHqNLdbT2qWF6qYEAYS7Ii/hAeYk7iBNHWRqTegqqsuPBya1Cco2GOQcit9RXphvxkR48wUKxE
M2meMBOc2HwCdL2EJbadjRLY+9EMGCMEvhFzEGUh17AjFkoOa3i7yTRMClgpS6vMzE9uMmGawti3
LZ/U33i0aAClPnABWyYwoRO5uff5szWMaKFBmL2W0u2/VoPpaFrAHdf9o0uaPYjvxLjSLOgRsFju
qMmM67keAxFByRPd4cnGsK5CNMWzR0cJBg9fTGtMtBNe7tiz4xrP6K8y17bQEjLDbhwhtt0sZ8zK
zqNst7C9znjQo4YTxGvj9/0LW3ZrPMLGfdPZ/hEQHT3XPHz0fixJ0Z+HFOPsnldW4KbOVWY1mPhm
ZmF5hB5+q85A21zPcbznNQqjL7lffDZ52214UyYHNtqNL3+peQ6bwECsjn1TTCPp2voUaMo3Ax0F
lAUxys/Uzc6+bLJFcs4vLqKW7+qlitUgZd/OIiaoRI4FIBNPoHyYA037rcmaLhZumKOcUDJzIRj4
fu0RM+/pZkIcrDJ/7cbktHJEy3IoEdsXgWeQ2duWt3m5e1AraETQXdSsRQa+YZ3eq4WkmVNKKSim
QfRZQFU2Y4AWBYfhElHncunqLLD4kghwOqgw0Sj13eTW3i6vSTt8l0C63ylOZUy7jiEoHr5AETN+
YSQK67EBqUO2JfCcUyzJpFXe0M/WNnGTQNihpfghJclR7yXFWAK53nT1SxBDPyt+SUG3oHelOwWY
2MW03US8RFgC1tFXNnjbdyLB/2Ixa4WLe/LXToU9msVszhtHkhrWVjWHJsN5ampMBdO75rJz/nDJ
JHcvBm/2uwUw/LVxLfpckfsvlQUrGb1I44OVqzuhSdlvHOZCOGJGSjQdw1iAtlejUc2fEXbYyHtn
FmwPPTgr6zNCswTqv2CwHzI4JCAop3JVl7xc/2nESIjq+PsADUUCtKkvpVmNiIm4mgfOYxWJWF5a
nJTyPmfua370C8f9iMErZboV9LTyFxOQmfS1Gx9dRTZ7unvKumWUjii7euEAQdhqRbDg2XI0KQX3
2IgSemEfGSVO6FpQXcUvDlhrNhXqwSbnP74hvw+P2mygUiMZXAaE4tfAZg6wXwPGy6gH0J4iRfAi
AotAt+nIYHr0nCyyl/QR5684s4emUtD28stXO49WCVbtUhyMzWZSrdsol3Z+6+lsg3BYSyDfCijx
/J0X4Iqqy7tYZyjqTwuzs6jg5s0woaEHWgm77ant3c36uWvJLNnDk/tHMSxHhT4HxPzT+tUST1zH
fIC/WSMeY+5RXJENaH7r0jF1ryuwRAapE179lMmrpyd78I3IGL2GlLIbeYqQm4dGpQv98W3Bphyw
DZ3j9yiotZ5gqjd3bJ61RLZ6cxnP22xvGckmFZVytUds62kdOe4aCON8hO1oZwLdFylWsIXCMRNr
CdqmEShmB4dgx7xMgkOmJw0ZojfDo/ljWJU3UgwLGHsyZcJLVghS2SeBjek/SuJQJytjHC30L1en
+LcY0DOTN0Ao1i3n/cYTSNHu8PJm+1fZivTtRtAx8+KqlsQwwQYSdxzy48RNbrVRJbCWDvvFPIIj
Ez31EcCixKVfNgPTfGdCIcmaPisRrtJDl2+yKHOlKDsE2d20S4nSi51Ij9kyGUyXVEVTzElFkGOa
LaisZhMgnyHIW0AFAY2jnB7Iln/9l0EMr0WffXF5/l6xRXw3RzyM3FlP0kdKLfYf3bHuy69u+3Lo
F7fobVYdFlKvLS+zJIbqudOLmW2s/Niesl1hMEEwZ+/85TpBcOLQRZJmf47IYORWm5a+iWRDXEy1
0EthdreofaAhMwUMakG3ItSa+3HZe/MzTynaa/wM0iAkySIU8AugJqXgD5BVUnTa5gW2d3Ryn9hn
su6vezFkKZP1Foi+c9I5KDlP6I0bytynVcHOE6m1Gp8EW3H1GpgvjgkUXRRAuP1WkTkRMJ8/ab7r
Miq/YV5nTjqNjKSO9a53b6X8CNeh96t2mtpcVH0g7FNyb8iKAIQnFGq1wy1R34WQIAgI0IAP82YN
OPDk4jyF/8mqyUGu+Z0x0jaEWjDFXTei86Lg0qkRfKQFFSYc2V9YlYnSbXWP/PCpxaC+PnKvcwuU
OXzktcUkZPMSeGspol9I/eO86QWsdlyImwKvp2+mZQ0wxURUeI17E8/zXHnixlcvrYJS/7VNXPkC
/vcSIsUND2m7f1fXWaTuk9JUXs1Jh0B5s1a/WeMB1n9HvCDMWIb3hAqLL6v7A8hUcrMxBxzrkdin
jFnumVgrcWibkZGqtRIJtSLG1upu/4p41FlgiwXgnxfI7PfCQzG/vr6ERFenOXloxqLqNSI8qVfj
lIlBiEDBjLwJhG7rnGnUpxE1zTNAWkXCwfKvXMsAOUbQS/ZR3bMMOmKCYTEWoPyatIA6dMEtqxiu
4WShxHnJg/VYwwdv3/ipupipQqcy/REaX/ucggJ0qDsBE5RfEbzECHhQh9pjzx6ONxV4J/pjahvE
CZbPejqIHtNX8gbyCGcSIEeS1+HBsq28JQCVP2SuqhrdpG3gHa9/ocOtlXJLJWeaE1nwp6DGXJfw
+X66JyEEnzpS6lBX5oswA4m7GQcDGydVW7jKJedg8jxeEV+WLwwDxaJic2jxoSsIFxM8hJ9gSS8S
LHjCl56YuEnft8GX2pRgtheBfWrGZYeQpN4figlz9v3B2gMgR/Dtpo5/xIt2AzFeM4aQARCSD8tc
UklklpVjy2tTYM7mjNE3IxJb3naty/DRojw6hPsw6u1XvIte1yYhHFcgWMmz7ve4ET1hk0ihvsf1
lSOnGoSuJQvUsrMgu+Qdvk3tChD7c3IgAY1ChMWqCvGtDf4pHWT+se9HDedMfpfkhBwnxwgUgQPW
KLASQc3EeScmsiVzw9ar8VzkvCyA8jerzx4ed45B8e/CKbGvRKIaLjMiJK1YqnsLnHC++lkQ5CNd
SEO1mjoB9zelAKXLFyOj0kr3NryYdLYYMmVCYuYhrs0IO9Cvri/kBIo+W3WlpP7S1z1y1Xr5m6jg
uol/yB36nniXISfY1e0CKyJNcB9NcRMijzKbnpHsSRP1o0kopeT9xIKk6rkVw/FFWjip1T/NvDZ9
JQydoMgLKgG0sgblTi8ojUM3vi4dRyXYyJTiVxpDo+zSNRIYaRquFSgKwpNpFznhr56/hoKxs3tB
0hXdxtowg7fTYpWSB6yf5PmkYcN/L1BCVMgSjif16KrHycN3/GW0ZKntlXIU/lRXbfULzrz8gyHj
NpYELJSK25SUujjCpnZy8RddhcEdCqRNrElW/zG7RguWMHhUgTGku7GzVYuxB3VtNN05K4Px+LOB
aVTeT0SWTrHTjgA6LKYl/zcqsYs1ofzeVKQOQAFf4yMH1BH2YkXT6JZG4tKfQOoDUlnSroDukV4T
3tOJ6N0CtGCB8EN6ulzCyGv62JKqDCIp1tXHcpSyBC//ev1NNZzcjtpo8zJ8AStkcCmg67X+Mr6Z
l4wnLSqTHtdKoTSwYPGJ/+lj19pVMkGU19pfy/xsPvTdDSFjwJGBdYKRo6tAa8mE8xg9o+oqs2FV
J3dQtSIheYmGNToLn6YOnzERmeCbUnQLWXTYuKrMN++g4CrRapZGV0eL9iGwpsNEjZQY1boqSUDN
0xyhSN08aiPaz2zYivgVbR4iovtnB+m3gW9OoK7kZzymPzS/SmhToLdOZZC2cAD+Msjv8xGDMMOw
T4SF8PLjtaRN9vi9vRwKhQUm5r2UJ7rIqETLjB9g1bHIM7lxsudzAhRULiGm/kHC3O8Wj/EFoiNE
PLm5qqi03ZkzUwyhPaUmmyoGjZ0LBmumR0g8JDrC0CBo+lrW9vs1EUCghN8zLxSE/+e5UABAeV6O
FcgAaC9PUvuamJXB3yNpec4FvCxhoBLellf90oBJ7QGgHt9FpwpDjaNhkphrrKlvK3iDsCOPVyYX
eTR1qHBh8ttNciRWvfhHml6E0O61UfUu1hZ320vkupkbM/TZODBjE6bjcP9llFckiPQKQGMzjE/C
hzsRY87YVTCAM3C8bM6BPoC1T6Pq+OAeNGWGA5FK/kyMRJtEBz1JhtIia/fYSLhUdm/jjdIRNtrv
LRkim2kQdSay5GVY4zGipaQfvNRRbB9qbUEBS6ARfZEBjR2M04+xLzsfKg74yw09iMDAvlVVqXcn
Cr44mJXQ+PlZ4oCRh7vsrxiN6WcAUhz6B4JQZ56DL7Q1hBLZjDpOr6nkLJXEGub5R6ecDGa8zcXX
vnhkQXaMeRr6LKJdy5IvoabL7KKPy9tW6NT9t0Vsi89riFn0oczS7UXclBTYSS4esDA8T/ZHK4+F
pN4vs/4wtIavtdt/teweafsVNi496ZkMBHOxcYgN2Xn1Ts/SkfEp7MNW5+eqhf47X+gQfrfF1aMG
eCdyPhi1jHT9vaCrfnoCmLu2LsRZXZBz9nna4QUmXSA/xmhcMmBk0fWCW1sc37Z2J+aqr2e17JPq
JFjACXQ0D99voRtTo/V0n88/TOiJTMIHAGKyXcDeZNDukW3jP1nVxsxg+T2M1Nl+Cneb13WE3E0H
OlSly71ZcU6qe94o3djSGZSkMFFU3IIHzPSj2uEu6awOwqlJt1R5P+0MZA7Sr5PAU/1XkQITaVh+
s5SieWDuKiEfYgRfCvLU0JrxV5/wPBb9I5WeSJLDOBhEj2NQXR0Uj0/ZRtPkPczCdkOIYYfkVGTi
dNnVOmCZKzWUiL94mWBDf1dV9DPTzdiOwLjJOzI5JDLVgodHj9kSj9Ey+T3bvjbEvD6Rg9w/tjGo
HkNAaUXrba29frcMS3lPgWIlseiz5JY2PpIyapOqi7SH+4zMnnXoMxNUULVSOqqyuBop0afkpLDk
7ko4QYaX3kIjlOD01NJ9HaXqkrefqSzOTXO/D74ypQgm5VFrw1FE6U+xCnC27H5I9swlceZNhTsN
/iEdwLlFQVfq6QhP0ve56MGhkcaM2H68L4F4en500fl+wU3GrjiJii1ZdL81ByV4ZzHfTHe2jM/7
P8AVsKJ1RICEcl6nCXbw8GAxVKPuS7zGGGUDenDjhxWA72L+ifx8UoQs0TF2ICqLuOKLiM5HQblp
n1WD18L50VY7rmSZ+G785rISts5wH2mO6bFdA0Us6k7vwoKe994WhIrQgLFYYQ6NFQgu0QIlwN+4
qLhNuCxc6Wk5Fy++yxdzNGjhQNGvgOVF507GSlTFZeBg02PeMtWRmNPuPiV0En/jgSvCgFJm2hqR
6wDLxPWETA5zzkXm1owBMEowkpW6MkG2XCm/FW/BT0dcifVfRAMN0NBUO222GeGn53xivYxM7bM/
8wrhmSfW+p2e2vQ1Jb+2UErTC71otQkXryKG+wNe2mLroxbiGsty94qeEf+9klpRSwUScufWlMcP
cXnYmeRacCM1TX4wgKeB9sDjQGON3Cu2TZ7Ex1UeT2RumK4J7PFSVEQ6A1qvwESUDvRiV8z+XqVx
7RUSKWVuu3tT02zV5nFyB25iXwZlX3GOvrA9l8TENy57GI+6UQ9M1Py2fMw8FRb1+Pa2hEFZfyB2
tD12AptivThYy7CZYygo6zV02xQ1ChdxS7uLe0AmkeB1027FPcUcu1/LUkZCH6gY6YTpKmYTOW4u
rpGbg58zf6tbqTnnRLxqi8kkO7F38uaGpb2cNqVDLTXvBxJWq+D8b8OiiHY/iWx6MPREqp+BjsYQ
fWgTb6AP/TrC692jsxoIELpLXTtFNFq8NXFl0tw6N5raE5WNZnJxmjs+POxUGaGOjTF8zbP9MHKY
MBVxD0A/s835hTmabFL8amWyLtTD68wf2EwRB+rVONru8ZMqkihrxllCfAfHgpS4Uyfb9C6t1zth
Bjf+EcnNVTz2ArE4ERtLJvfPchlJhvN4cJAcoLSqmqYCY3rOL+FU+uXfdzUY70HRyucgZHnaKHT1
iqecBW13HD259yEaJmj/gmdkwd3Hm5PifFw4M18Nh+1wRsHuUdaSMn4zKRZjcnlKjiq57NP5t3fp
HvLOznoeJkbwj5W98NxDYqARjm1QN4eaXJ3HQg0l8g9RbHd64lpohIRz+MSuw7zh/4mLrEynuJps
RCI1CSd7A5dcXKYj4WbsfueHOPeQ8RS3Lpqkxk+HjmMPFMuQohnPCwaL6Y594A5VmnMI2BTra49g
ewImNe+eKHi5XovUYBwUfANnxmQCFqMvgkwVgbi7S0ZHirRV7rvbN0aitq7AOoOCnocYD7mFkdXQ
buB9tiiZosqbutZuv2OfPgE1+Ro7LNgDCkfnP1sTX/9oyKKiadt+QA6cH4o0UL5uy0mVErhvWPIX
68GF6l4P9EWx9edrvhTBeDFuoxdSrlc4VBiKOVkAhdhOGbJiF58gW8EhWBTbMKAe8TwusYL073Th
OhAj6GPpydOQoNMpb+MOg61mFnaenSIg5hhMCtEjJ1bi4eHgTw9fkyHzvFbKDLqg77/w4udLIq+O
M2yzSMz7wlxAZoHQKENZNRv9LJJejFQisMq/aoCiMw0cZT5gdfmYl9aqoJw25Xh0yd1eYP0BCqDq
NuBNCj/4nty/CYmbOq9DigDfHPCJ6xZSyeiYjhQ//Jjztnj3OYUkEMdWhuMRex00StMw+ikbyqRA
jBKuEA6jMw/sb3B1Dz1fkmXm8ENDgfFvIIh9p7LMXPLWp4qYTeLo47G8HKRyiKN24qAdIFWYSOlj
TbAbRgCcU/K2eL+2Q4iDZlEmbCTEefRQahbzIdfpAL+ncMHHXH+9wgOY7GvhP7bVP7LwiMce8uSR
GRrlMEzv6XSGVkrNz2+JExHbUOsNbFTGAELKyGbJmWzk9OM0XXVJzti5NHz6JnUz1EndJEL8IP2Y
rYjFxpLpnKnItKGaxzdTWHuhlVIVML6ojeQedZvo8vQDuA0Ldrd/caf1gmdQc2ybMoPBNLcN2vGU
rmYAS2K35U8KaqwDKR3BCpMcELlhUMpfGgFTHC12CeEbyeTq2E76OhTBkczZEyKLptQJtC3TF67b
w++v3pCqyTPnetGFSHVQfFfYLmpHsVSSD047+y0f3t00W8u8jfLC6kLQk6ZzGIyMQs1DnhPQ+adg
2rn85pa4AuK9geT7VYVGT+QIWGq3DaDVwVEbrJhOhn5yYtNDmFBV7xNb+cvco4FvHtg4r/AbjT6/
aU9XBZubcTi1PvFJoRjNocf58iD59uDZl+5hTvdXluMv7qbf55lx1zOoK1oizjpuWl3V5+f1nA1Y
GQ0Uqfw7GzCKwWICrKeuu1mvn5sTzVVtzcNQsbSP0MxI8+aRzgWFlb54CIpoIyv4Pv4KFvDYT+ps
utoAoj904vYn9///EVh6jYmFld5SDKG7n/DJ6pY7VZCnnEVEpvvoB1KAUzo2NMLl7ETbvkDCT7nr
qLEpQVYLOyYR8CpNdFnO2NIqHfZQVB7nf1BdZ8Az7DZTT/GXHIX++7RoZNj6NJ/ER5jGKyCvHdV+
AVqtJ8i2Dyw2zoyXT85nZ6E4KzgAEgLTFLSIphQLCU1wgC/RrQhJ3tYSVNWsl9Ah79wtg7Qvt8es
PsGf/iP3XfEgbS6IuDiVh/EYoCRRhtn9lk09qK2NgPBo/GppH985zV7M4PZ9zw5NM1Tbe5g3gz7t
wij3KauDmW6df6+2yDMZKy/krmbpSXNDj1K7HCHI1Zo/nnJ13Kcjw+Lsu7JBCzL5dsmm4w+7Ezwg
oorOoGQJFjTjtRxzLv0p2ZmQbhuduCBR36r1DYKp+l+fWK3S7bqlYsBBS//hGMgJ8utVEGEiT80e
7v8i8r8Iskf42FO9WJeL71S2uQHNFQh1AcdkucnbuJr090GMYeVC+btC2pR8JhFxMJFmd+vw4+X2
1p9sX58FqgSPEjS+XpYYrr3Ze7t01CMoibksIGBuBlm9LfiPKAT0oZ9iIfLTvAoO4UD7UVBpCuy/
edCiGjgTXbRcELxbFf+dVvOX741nG81Pc/eZItSAeRIMW2yuTPowVI/fK5dJ5SKSK7mz+DS0Mfec
TkEj7FTqk/xiaCw=
`protect end_protected
