`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MghEvPKGx5G/p0lnu+uO5V1nHtK4AdvY4MzESfBdZhyGt6+bFa+XY+pc84JsY37L
8QZSG/PgUqeiI5+XaTyCG3i1yw21eKdWxKFYz1fW/iN085h5VdldCfsB1bqFL6xj
p7Q1AVIwM8YpFIPXaefdvbssIwK8UJuRqoYsnf+sTyg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4848)
+uSTGgTzaSUTP8Cm48CkTs8fDrwP22jBtWgRtpdDn5HRiRhE+jPENNdFrjmJdgv8
DKxhOn9Kn4s1F2CyIkzRmpdSx7NFHQ75Sh6NUKq7bd2BQHyIT7f9SxPXc/LItO2h
Rv5q6PGmnQPC0GnowNi4D0/6LLOIvDtTZrVtXWecNsp5zmhescTwbX6WxE0FzD39
LAvdsDUbg3IvBYaSqP7YOfpBmpvemEqx0NfN6j/mPC52N+wudNMrKks9sO5TJ9De
K5r40vCSNtl3CQ0OjSygOus6YGii16LEwpDlzGhQsH81JayJw5eM7q8AYpOXbGz6
YZsc7D/ycXHwwoAbIJmyFm6lAxd1PaFknwO5iSID64E+C012nzEyUUBhjsVJwO0i
2aZQvELKdlGex10bIMpoyRnqTepPF8c72AAlnyFZ/+Y5hyjIXljb+TWzy72cWS6i
7ydlfW0+HiPK7hRcU5FvU4vl5mHc8Yo3CUbdJ/QCDm4YYq4qwmOG0t7rahVydJTq
tztPZrdh5oryNFxf4viPMZcotCpd/djHK7f2j44mRAkga4kgR1VgucijwXIAC9tU
Ssp1Wd5So4/pD6Jx9b55bED6XtE+6Z7umu6GUgMdkgDQZdT2na9P9U2DNxjjlTxR
4j9ASSRL6ZvHy7jyWGxCnmg+tae7Lgig57lZAH6LWktnUZq/PmqBMwpri00DE4Ps
ObRKN6OzbFY8yVkYcX6nrmixicLzZoj+RNh25gTIj5H8O3g8ZMBgeRCUhOwoE5cd
hqsC4Uamo6KDqE63oH3gi7ipCRHahyIVmIGNKUMkkbzkrD/q1hE4DvpO/mNq82Jt
i8mmv5Mop389uNpyOt3D1U1SgAaxgSPYF74A1VrCGbj3SWpgmG+VeTYQ13aKHmU9
U9aJ3whZzfa56RFYqEvw7zi3V9YHxjqMlr/lD+oQfPoJaFvb/sepPJz+DeuVDuyd
fv2OY+EVrnMw2BrXceM4v1i0QnXjsH50ODmiw2edew6fT9E7A6voigJ7ss7+5mH5
/UtJc9g/dLYN2NOVlytJ+KlXtRMFBaBKnJ39NEEPv5iGfsejh+I0q0EoquhjO9ee
6RQyUmu1YMAh9uiV6G6WEiXADHWhuZ6wyrU6C0cIzx/R1tpvwnvoJuzXLij/ipG7
WZeqcFl/D7fxnP03cMFRVtdkRfGfzAW1TpnsUoCeGKAl0TSRvDXdw6PEoGX3zkVN
5jzLsFUrtx1Lta/m/HJmusVltl+npbnN+3gOQ4y/0LsfGzSvvOWQJUjbtCuS+aIu
Y3VRGsYwFtCItHv0BVwxXe2j3nNNXxk5KzTgYKWpLmE2myo6g2dVd+jdwhQ6SqCU
Orx/cCSX9hoWhP5zBboMzPmcmIS4WzvVqG/9VhXpld/yrTg8dmtog4ygR/0pFaOC
ru3t2SsvmAZdwH3bnqHfnsI3HceAmMDTa6W0CccV/z0uMaWAtd0FJOphoGF3Hxm7
oimM7U92aCtji/zb+Hh3eJ/HuI7tuv7uAquctfV09T6HD2+BwI1pl/1ZRdebNVSU
09gW6oLfahXlV3VFnZB6GAIkDuMveBvhE7f1C5F2K0PuKGSMtAIrCp4Fgp+n6L/z
7wyWS1MPFzAnFhKNKWL7p5XIjMkRyiLuCu5uP+1pP0CzVJHWZFiuQmcJ67AQWeUR
REInrb9Ym9xyUHqaFPjUszAoyQ8Syg8L0nS95qEBPVdeEQj8vawr9MsxSVR/U+Mu
7i4pJMVZaNEfvI/MJriCDDZmOcxRhIa7GG0P7vbWaNxDSC0a2jvP4X5CW0rYqAAm
oIzZy70pnRKc89FhXGJJT9pByBcWagYduM3vZHTe7hejSna4eXaj2EbPpKyGxfXG
fZWBzkVajpo0LtRhqHIF4Si+E+Rs+Rvh2YAVDKuz844s/WpRLU71w61nPcKKlX+s
YQA9iYwsLXa8dzYyIEq2a7AlardImB42rpKLibGM4yJz8pUhqpqnQowFO0jFmfrD
y+lbD1FeTBdI6OxjwXKigEN5P+JqCZ+GUlqs/xD9Tv/kiYdUaD16gfGNCORtQrBl
UrtQ7+Kq46EnRec+ibBe5WKNUhkaR1lRT0z8MbC2Eh8PBuaV6Q0VrK6c3OJFA9Qk
M+TmNUsNjCQwJ6Cb4drOVdjeVU/UAwKXmZRsZDPO+gFCQjbvzuvZfbPrbnQcCQy2
LLjSXEjBwafnLIGCgR5VS74106CWU2HxeWevyZuMPda7u3RPJ2lHGb7/p/Fg5ccE
TampnHM9S6pgU2MVfpOrY8B9/b51EylHGZv2XEMhuHE2bLT2jatgvqYfvUSZAFDO
K5ozw0EPwp94mLeQSlPxkjWAF8ZwdKyHlMLJP0/U97ToczZ1XEqMJhDZZM28BKAn
lEoQ3gDNCD4IjI6CpagZsXy1S+zgtm2KZPLiHevCacNzs7gB988nWx/T90IiZTHr
XmWSPtPaRCIEB44XnTOW2CstXlUOr/+7TC4Ey18eecJqb3voTL76kcAAkn7G1j4H
YqfCOry/V5KtZ1beHz37fEy8XFNbpqG6KVskHRGV4SkClgkkl+rZ4XWbj5mE9B3Q
oeEyY28++5Nk09JeKXIGlnB1cUPVjnjFgyyn9kODY6qFxBeLoN5+aDUf2x4QxcPS
hNfV5l5cZ5FpWQ+hxfbEI5xfZwp1mg0DgEZ6sNbil/7OrM/5aAfx4NOXI9m21H2s
l/TBaxnVxZMOMEAA6bEIaCdygIiMGCyLVaUwYidmzmopgYcLtxL57oxu+oeWyzfN
hrfXEF4f3jYP0b9PAmX+/lV4aeXWjbtJAkMIClZbNnOYLtJtVBewD6J2t3P1J+Ho
ifeEkf0o0si9gPSZWbHXuW2mG5xQ6fpev9Vf+UNx5JxgY+oPcgs1q1uMAuHAVgJ7
JMVO4rx0u6k7/F9EL5yEY6x1uv/ZPqCNu7d5TMwaD9T7BXn5OpV3PDGmmy6nwrGX
iXgNNmpWhlZWfKFQmF7gsoZt/mTrUZj1ELllLCYGe1mq8Tfkb9ASAloy/9LoFcCT
SCcfbE2prkT2CyheClAUIbaMTCZtNmZV7O0ToIhBQ7iA9OtGR7TvWNEy0YzAI8ec
rd9AWVxCAwbiJn0uGzxf6NHrJ/yatq9YurZBo4gsdc4rixbUN44bl5yd6b3+8d68
JhIlBoHe6kWvUN+hZWiQde/euUjUBxda4QTYtymoVppvyBsUJUOHIJWKHQTXi3CD
7YXWEpEgOTjpkFmZDUFqW+O2sZLwoliLceflhQ1mttXQoXw5WdY8WMjfBp86/Pwn
8+LNAJXlD+yGRlaAKWBK/E3JE1VzjgS+eMHD9gPBow1USh7UyXFK/8r4fonW0Anz
cJgG+2jdqvlPXzwF2qunZu7E7FOSOLkumwnJIT26q/w7NzLRWoc0RBCt8JYQR4cy
6okJU780kakeqrS7ZgUKp9y13Aia7vZzPh/evBS4DjP8KMtbE2P8K74iWICfJonW
qlvL88yRd6+DZKGGGqNIM8F5NCNZcdHjdn8Y56M+EX1Ykiq8DxXQE0ZNkYYkRtHE
/yGB+0KMHrMlfOkOsedFEUe/LODhBuee+1fT9FebXkXdDzZI0W3RCDn1Vf207LIP
xYSEC6tPREzc7JFYc6yTu4PYJlZS4s4b9QYcgt8cLYfWXrtlaHylexNCmepNYTGl
v4WIUvKhUmg0bMxVRM/MvCd/BAkH0aD2jd2qasnzV14hBegHI5lI9w6urw8xAY5j
pnfZ0Qy1YlDRvLND0j1HGu/VP72CcjqXncAPa7tVXXnsj2+P7FyB/adPBIV8idN9
cyTc2Z/xbhPvwYRZolkBGAsle7CiwT/20K+X3ggC4OmKVRnz6iyAkHrr5j1HE0LJ
Ag2PPyV/z0lfRgOwJx27NMqrPGP0gBW3tTh1i6M6AXW+0ixSzhr58+tpILA29SwT
p1/BQ/ErCScE5nD+wcFnFaiDjUpOFuvGqLmZ5Nz8UNVIZnyrna7TZZIKcg7+27nx
q1tp5NlZzGuntk/n1VGMEBvNkzDMhZPvLd+cU4/IQiDHqrBeIRIK8IGjPcQkUml/
p5kB7Fr/H0AV0pqy9Tjhk9b5ITveIVWzMQG9sMXEqgbC84mPrQOy5AF77bc3/3i2
fRrIg19BfSBhUGb1nSw3Dp5UrTlXUFOthGRhes1cx8W5Pynj/wy6wXxxyc+UNpDC
zaKPmSpfUiSJ0jROghDRHC4JRDJmLDDI4SdkWibNy2kS7t8QhEmvQi71VsD92VLa
cGZUrTXZjT1Sj0b6nPNw+ykrzi/QFxYGECaL37lbZVyC7Khe5CYFFZmjCbCHmsP+
0rBStlgwUnN7yRElljhGPz9dGoTkeKAyFNoq8VMHakD0slsKl4L5IRUBehmZzfWp
5vOUdmg/Jt3jU4RPSISj88Tl+Ka51uTVohy8WcWajBI2fbwZ0E5ux0+hZvyYpLw0
dZlizWahixhFa0pj3CqfEYE60B6DrZkiRjJbLDG6VT1JJmu5JpSD1MRRc6a84fSx
GxEnj9sbJU761uBBiQK1bB9uqFwLtGVUEASpR5uVaB2jDxWAhNS7vNp5U56Jx3Jd
+D7JXnAZG2n70bM8tkvFXek+G51rWpDP35JYXzKdFPKihQQqDMBlTOA4I3L/029l
SfPg7LPrWBIex33NX6bjpKa8aAHyk1USOQ2DzYDbMqMTcIhVR21DL6nazGuN8r4w
m1DI/4YfxJQHONkiGevWzyrpYmDFTDgRJhg6wcsWuQf9HDqAcc0g5Mfb2u7nNIY6
pXfEbj2tb+sCvcLWnFmLHAcGdIXcVOdpfsflUeDmOQ/+mrzwv838EJzrIbUvbYJS
n4aHksHSZh1K+M5n0UTM8MQ4LjgMjQbTVTlJv2WOT7WdF+HI4aIKdyxgbyDegH6r
b6ehg+hv5my+hOqsPbnJg8b7SQwolB4n2UixSzjBzGhxdITIvBMfktVsWmt8IB1h
epqVCIPytOlGhf5ZZoY1lN1BM2ZMwzXIqqHQpmxsneGfi9H4PSBlFVr49cx/1faE
IiqC2NqWkAOqJj/82UqEDM0VEUaVdcMFbQ23WCo+47LZxm1rpoS7uOw1kI1bwMOd
W9PWiEQa4IsceLwu8GXV48ynkJrEquaYiSXhuaJbUCgB1vbtm5xYT/lkF4cvK/l7
CBtxZZY1Bm4jYxYprzyOk9jhEg6rJ1MiAigOddjQLAg/nGVTXv1h79S3qRptjS3Q
Csjqp0OINU1pPNKmMArFYe/y3R7CrE4M27DgXawMvb/E7eU2YFu50Ig17pi7Vv0g
BN+yA5t53zwWdL3BUljR4mahFJi9P2jJaGbb00mWr4ZqmgEpKwMuhK0Ri/UvJWXu
tdvmZDF6BNYTA1AKTdu54i9JtFkPska8AAhz7XG09D86CKZwlpakz0ZQw6LuI6pV
8Yqa/Ax+h9ki+k2jdhc0bV4NZ5aYAgmG4y1imyk3qAAMuLlpROogBwW0RAjZxoAL
/OkOmOZ5ItJ/1snEHI6mf/YbnpnT4hVJ+9A5wxyQpFwBiM13GmardHKM1oSxmlk6
MX4vVk5bOMoNW9ONW5K+Q/OhBZVfA0hWERkHIgIdHZpGwpgUAZ8s6FErzN5oqmgN
+78dmIFauQjZgCMXRCGeWB0+AywZci9hWBzPeub7Hyj7xsiMAGfwKl3UNnDv3m5e
nEBOZvhQN9lZ8V+pZtEfJuZp1/emnBtlCg62dntjyLffEbQG5bqgNYelxYoDN+7b
tky6rnA/uKj5qCSe1dBmpgnftm+Aq4cI+UJrN8w34u0RKdqJbu2+ffNYZpLPwYer
nKKSHR4Mxk3fi4oPtU+AKCDsHdr4JM/2A2wjWehWa9VtHNAHrVamsBLTh/puhD42
7ZxTZ7Lvn7flEgk0lzp2WOP3/LEsfHvA+iO1Y18jaTdZtpH54zaiIq3WndbPq64X
83UIKjem6LqwRkSfD1nsX3oiVfQrAF/iimwRUmKRI+rFOTvEjB9bosON4oN6X9C0
aPC9R3FbrfZJbwg1aomgeHLYLzcnnZEVObHeIzvFsgzB2Fovi/Z53IejkeEdrIF7
tI3SVKMbE4vIH6nka8EHHEINDUFaFi3CMINWB/6Dg+w0+eN7F5q/udx+6CLrbjC0
ff61hlI/xlQIPIdLnseEXHFZJ+3U9T3iqEDeuurqNovJfPsWO5ctkDq/VHtWxsZG
ni78UlCJp0phhsPWG6Q2HSTYxYWJQyJVQo/8TY3EG3ISrdi+kbc2ItGtYqUbQJzC
5hn5F+PDx7uA7DDgs7QrGuGXdLWLm2tMPEo3h+Mp07hDGQr54O9DwJLVRROlfyat
pcek+EybHt5GUWvq4L/B5SfX19FSKXM3Oc1Tk0+PP5NRQgD6TUOYqIQCSgrenlLj
b7yJm4P9jXjElx4z13wgR28vMLM0E9UV7okRq7mPgVELbNW2P3VER7ZrbOMw65rW
XO+B4QoBKUNJ6rP8U+0aW5MsaecckI980Zpr7uaobztt8JVmg/jCCH2vXgyLG42y
`pragma protect end_protected
