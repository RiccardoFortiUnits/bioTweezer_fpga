`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bmhZTfPbkY8myk1EYfyPFo3VSTmnNpE+nO/p+INSlEvuE/o6GDJXyb23jHqVyF9H
NvAfHV3aGU4qc0CzURPZ+RDARw6lfCi3vX+RESdRxscQOqjrpieTxclwDJKoaBQd
IsbYk/c2rMXw7QVQ4pyYs/brnqWK4xKqhLSt1mlstcI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19936)
melGAcpoWpyKTZUOdGkLOKHHZoYSZ4KHLGzzNLG7VPBOo9A2qIZAMLY1v73oyo4w
YNF+rbT2Qy3iTodPu02Uo7vGGQ42ngSHx5Z3KuwgGpuUNPNDCWNTYdRW/pEAw9xU
DRHqgu/VvDtNdq4jr/vrL0QcpGdvmpPorFjLo5BdWFwBkHPXIgAz3Iu7rp64SC34
x5YIlsLC9fS+J41KPWGOiULJU91hQBg1Js0AyQ6ycTxn+9VtN85Hv6uifmD00tSV
Z3Z6LRDOQn5Enf+U4kVsrtC38qzYiJ8KxrRBkjAoNMuAsnzwX+CmLek9Qf4HoCE6
Jst3aI+rPmDdB07h8i0dHy92rqhIkmpYAt0Xe+q41CVSJkU77wSH5JHR4Dw3wRKW
M04Sq7Z1JEEH0J/WR269fpGSCYszwy4bGMp3aUX87EEfxLDb1cM1klY5DhdJrjFD
8sM0MIYFAMdg80uTKz5GZSwuSFkSME5sCoiMF0m+tgjCheI+3o81lYfwk8MBNkkT
KfW4bXxZMOY+o4m8HDS9Qd4mKsZMM9RffV4Nfb7jFuqNdwcbSbrcYEjvuYcF5ffK
d8P4UsRUerq94Vso2seWmpjTHqDPh0NQ8SbBmcYn0J1oo9yIAnmtBZDhkiLKdvtx
Bedj3a8BMxLGpfmwElFE3wrOC3YhqrdgbSp7+fMwu3kTjrIpUieGgQG8oi5r7kIo
jedcFApKyLv1+FJ/lLKd0945IvtOG3zh0jnzJNPXMydgUqCWmUJ181lIxgkxJUB2
Hf+Y+DsXYfpyfhUYmZut+dvbgqesrJgYonxWfiNRs5FQh5z7MAIQZpH0hi4qOdup
dz3J1+TvEPcEy5QlTVBnLLuWidH0Kj+XIWE+3lMqk0+5lL/BLN11oHTQd3Crt4QK
S1Vy+EGbjqkVuC0SvDe1bGF4SQSYYsKTcrs3mWRGGXgkuC6yRhCf65wEu5JGFxUo
xVGWiLWSERswtLwzUei1IsFNCw2D7m3Tp1pzzHPQQxca1k8L7+V8AXzgdOu2rRFz
dE1q56dx5zPHNN5gpUC0MvbjYFDoP5bPrMRvCV49kuu7irsWkd77kJeaONYl5EwL
pzr2HakUm581ar3ECMxxIhQPlXtChEas7jJR8VvBBIt9AmZebxT1H3uwTWGbqn74
uzyycuEQcAnctoouso7JqS8ppmv6KuO1nOmtJzH/xDoZgubNBe1WMC7Q+Lzud/fN
6tjSJiPpA/PSmTDqYDvNs3YycZAPcOxlDKn4vKOlZ9dRECSxoAo8TsAC+LMczFn4
+Ki1UwsInWNclIpb6Qpi9WVwMn8HLCDVklSOlXic7twLcNX5jmKrMFP1TAR6czi6
7IZQd3EvP4q3bfsfixtk6CHTXSpC2m+96aWJu5Dtiafe1gbW+khn6BvPBr+dAH9h
bDYj+nhJyCEcZHKZL6cKtegMYHefB+SmpbwGuBHkEl+iw+beu3wRhe3lcIyTgAR7
yckf5HDoaFHW/B9ydeZXYfLFhrrbUO7JJp9th2JTX8AVkCmltFL4TEGl7HKsUiZ+
CgM6Oz/rqg/EdRP7j6hKuYmnNzGMF5AviASsnEdkY07jS311Nki2nlPBw+3Cqg79
dIaEeOfIcDymZDL2rG2cL/s2UGNj4OwdcnjTRmi9uhMPpNYpiv46riAQe/8xVCgU
CFNVYb/V/ttGr4nSLd9hFIprssVjXDWNbIMi8dT3AEV35YNwHyuZYQappGjfKLWb
bcX/cRoWiERfPbsyyngzNjGGYVT2YJx7nVo8bGE0j87DVXdbWUF3drfd+5upvTAa
jcyKXKzvqmAnLX0HytjF40xAuopwKqd2KZlenY9ETHxeYYVRIUNybUY5Nye76pRV
Ox6jo6LQutSXUF7r+YffP1lROrutuycE75qLgYjShB9PWjXioZTP+SyeLzBdcjM3
qVY6ryQ5wH1h0KgznF3nBxzM+fhMfvjijnJHIVYoD8WTlSde03mlhTM0CnllGqe2
IyufAt4k/hUVgpSAm2m4dcE4hg+fSFFBEFGv1dJsBPlrtK6De2TivmiBo+uDMpqk
k9b8fPs+6rsRyPN5A3zlL3G1J5bbLKqn7pTTWmrn9RW4Q78V74+EYgOFhemm0I0c
80f792DaFpr13aRvu9uKBmEpUvfF1jvwYan8fYwVPVpuTCXEW2bQyrrCIXqLqiDF
wuZN0I/rv4HLixBNa2iTcyQg3bl7MB9m+s30y+8vG4pXp2hjkaTF5w7CnQ73g3JN
5zTrlpEGsqp5v3aw0BkEqg1fEDDpM+FcmVvqmQP30O6jAqqbkipMgNESo43FKfQg
5g+jMK1Z7B6oQExztCxvYdSyRXITBfIw6oy/uyWtV91JHAc2mmb1ucL5XzE3ny8K
iF+J6AW8oP6X6SzbeFNdHLOWZxwVqwwiRqrxv5iBjyDV/KgZhBGXviVRPzwGSUcT
gGn1kbh+xbzoq8pcSQ1Bea2h+Jwe6g6u6oKWCKmGVTcOd4/s+ZXbO2ze8BCupbT7
Y2F6NYfWKr1doBcxGRxu5EnP3j76YdKWu3aXlxIyCUg2og+H6sgALuvaEEpwvabB
5Zb88WqGjoG4TqEIm1fxwZWj3zAqxqFLwtXNp74bSz9M0kM9SN5sgaBK0ppBVy7v
9WYjLvi91r1t3SypEDmeMIoNkY5GbNvcw82V+PxP2r8OPEcdj2V9OYxjYhbyqaeE
wFX7XWxXXjRcKa98t/AoM+UHgr2zmfd2uFiWP17zxsBcTqJZ44TXuUmbuU9YAlSi
/LEZoeDKriSS6ZaM2McNb+sESTbPVGmP8uB674TtUKW6oZintJoG4/baTXFT+EL3
5YmTF6DOLI35HTkcg03KHbzc89Ga3mYNztAZ/BmF7M/JNrYXebeIGUkXovbKK5mn
/vLle3TLRdgmOGZkzI05U+sd09fAIMIy5d02UnI/LZHT2XdW9ZS0rgyHGGO8G+Nt
VYw7L6mJQFUNP9ZND1vSyhfc276WoY8sMvf3LLm2ZSIuh4ZyvyXvKV6LAZcKNUH0
ABfrWNmqvy3+7UL/IjtvTw64OfrTJLSBNQatb7Gm+vcaBVq0cD+lVfSrVOokrkRo
xD5isd8PtKYfaKCXby8c/bE00DvdwGfFu8Q96d/tuS1OxM80+PTQw0ox+VMEYgwi
64aDSezbCduNA9wwhKJZ3Pd43D9ZgUZJTR5xV60DMq4QwKblM67GgzV0H/5IYszV
6Q6GbhfLzxaCvhCu2yWrh+VmE7Z4dirkpS/kxt+H20Mg5F/e7CodTEnWQRFel+dq
Kz8veQ66MMlteLRQVyxMLf42cVxxdmsBd/iNVyqhmCbxKL/ROZhLP0hUe1cIICDs
R4fhWJsneXsV4cZc2pl2644RnnJhk2JfCaVJ9YTxO0ArxnK01cKlAHs/Qo+R6s6k
0EOr+P2eNYQbEIz/F/oDfCJWDszNwAklD9Ql2CBQtxjptPvz21J0DeAb5fp5uqBO
jhn+C0x4QXV6cO3th7XKpICZgDBYasfdEEwUBC9bw4csNsansQR7G267c2SJK0cR
99BnJBPBgkv0rElWIjk9N91xPbx1+GQ2P4oBahkcg64PLa5DsqK2MEdvN4xKkUEm
wiN/g+EAzn71lcRHyS+LRe3x9piN0vZjUkXzCyxoE5X8Bt7Ribar+qoR8z+U27FM
83l9I6lNL9zm5hfT36Vuw9kCeDEsFblPyj6kRG6O3HLlz8UaFq9PbTYdN6QPSIsl
UZw+kJmiLGnnHfqciZ7sDHhOLPXECIGXmGNXk3tmxI8HCbkj25D1nUY1W07x4vss
xfk1q67+58vqzrsyn7uJtLZHay8lunj1ttqBGwB7Kan+HTtXP+XMpLEcNerAy1SR
/xueqslw2oMGMev+PtATVr1CWRldLWQE1SKOL1Nj2YUGvk+YGH7F4c1QCK4Fl64k
vcpdxqkW/udf+EzOT8vODMCg02/eMrQHM6vyK/LS4JUYV9jay5/wZjM7AsxqBvdR
DjYwHwkYeiPZGb9uN9ax+9LLXuJTXqy1lSdg/tKC5EMAwgKUNURmd8cNIGWzbLL5
Vlb27Iva4gFs76yn/e0HYnTEs/W2w/gvW/LZCkQJRJveZsrPtbgjeiNjyXUwISTv
XOQXO/PpqMKyCc2SKn10mZQqZaCzGItWdMIFhmT/82d4j2x2A9OgWp1omzpGxdLg
cN66cxsIOdNcxJIJELEFHWVfmG8q4fbju+nZ2ncQpXiF5EClDubTz5TTRL9bumEz
4VdQ1C3xqtV4mrp4xjG4Nwcp4R9O+jD1zMbGvwOmrPZa0cmeR+TM2Jiec4LerbUZ
xfOZUjXbE7PC4fnqSLapNI491jx9XVkORYqtswULo8n6jUoZxlTmBAcHjxnvfIgY
9wud+e3g2p2JbDbP16/HC8M5uI6wRxunqbNfZneJBdwFn8YwnFiSX50m/1ylCUTy
DrZAIZepJiL67LpAux0iCyTqBTOoIGX6RAGbvJGmA9lcwCsufHjMRlttfJxfY8Gr
87O69yxBlmAiZWXBtBE0UvQo+3l+gQ8niDF9F0S+xq2U94EOsK+DYoNGYSD/Zydr
6Ouqm1chwmGjVSPFyoBfDEpFv8dbbuoOv3v96Ul78HBRMz3PXmnQJTs0sgi6U2rI
7gS4aAgmqM9m8A77rjsUovoO0GgLtU9RRkSIGSXjD1MgGCSgABQDnbekvtT+c2rG
tVG78zmfwAwIHVOqx09QHYkrt54z/Hf1VY/OUv8uiJAXKxHSDb6zpT86wMr06fw5
6q8dn7cpK8kxVfS955cyN1luhniY+5RxYxtgGv+sBD/K312qFlPHGAJSYHP9zW1M
yU2uXn81hGf5nTIiBJxkWQjjLIVCEAw/nzJZekwUX4YjE6KI96Wzh6AaP8k9/5aR
l/tAAY6zdEZpS4ZW9mBLoR1UrPpAz7R/cRMYpORJicT46SlTpUffVFryU6Uvteb3
LO1aXgsagyl6BtyYqt0PIO6+Ny6+eJWuTKZ8+EHXbedsG+r3uTWuuyxtHw7ZQR+n
ZFyK1ZZmh6kJOX2UeQ7lAHYtxT5Fq3DpJFIidN+E7um+rnbQzTgCJqA6necNT85A
VTlY74qODk9TKWIRMrTxvM0Peerwfn3LJWB/aKpHnY8u1mjo3xplO9xHr/mwmVkZ
QAAAOcMshqdPZQN6CHQTxL33E457YCeG1mbtiOai4mSdqdld0yv7FLBKHds/5btI
Uqtm5NYqgxvgQqQyFI4qlRxpf24PDNTypiG/j8Q37o+cYHNx7jhVt77jMowvf3M9
0iPdeAQv2v69+jO9VUjBqBztTERxgjIbhbS6aKIJMUYqxoU1huW6gmwN/gC0SxQ/
wlR0mZQGNuoRQw9ZAE/Xte9TzA3SrKDiXT+ZbfjC3cAoNF3Qi+GkNUxExorr/Zrc
G4/tKKXDqWL0CFa8qZyu+6gOaKqnt9sGJsfBcwMo/LzaZsC3OlzA014V4HeYgQtv
U1AOEzsX3qSbi/2mpMj2Oae6Z+4rqE5KByS39aeGuBmH1yQMiwsNj4nmCehr5O5J
NeGGaGhK+SxWL6ZhtZdJRHhqOOP+CNkL+K0jsGqkG4whL8/fMiFM1f//u6dGlAeq
gjjBW0HbwkG4NKaSIeTZsRnFYifIRPGlXe0HJ2sgxyQY0hvRQpxugCPYCSMHEzSW
zKejb6plGDBPofEf/VUOEN4wOWjS8ZXLiD3wKfJdtjLceCkTwLvskQlSbL2C3DqC
N+2zBgh6EV1yJoDkQoEwTR+Ji+n7sLe4BoUPh7N0ptaDMYwCHsopRm3egycaFlYT
xU6836uHa4AFrdVZgs/AaqehWV49nH/xDutPQRTwRFjJza1wReckhd33MM/Vk3MO
paDMQX6m22FfKrQGyXMBKVeRH9wTmgJ1CiijFZjL/jB/fqmLk+Nnxplz+Pv7GlEx
XpdQOpMvF6WmmBsnYtkE0z+DMXYDSs5dkoI3WZTYLd7XiysAF8bXYLigogk7SwVi
wiwKxWZ84QJZYgs+oIxBf0rut52fenrZcg9wevejWqiHQj1orhUiHJ4+QXSlEs7y
GU+c3LknhpA1FdpcDEcijaNEHvP80EuiLhoCbGGk7MLoncPHyuwCzFU7QPQ+Iem7
olhNQl9l6mlzDIW90BypHwCVcKArR16W2K0HE2xaWEe7vG6pIwuRvWkpgzXgWxSo
uSTEwfMm8tqD0HZF9bCvV0ubrGO8Ef/mI87nS73w5EduEjoPeTpbelPThAGu+5WG
cZpxYJwiLZtmKVqapTGVPUI9dmu/SlpmlFmHk85PMGp1R6EkF92Szd78aFvLQeI2
lR1yeoppDjdf2NzK9WArp1gZPrCtE+foSzGTs2ZWVCurmWgAA/RqKGppn2ImUPhX
R4SE/NYyMVv3Ee/vUedWzuIauD2OlfInGDlRl1LPRJsfXqJ0uU3FOhdlmEOssIdu
7oVMiyjrJ/HnxFpHtkrdMiscuwvegfydPOOjJevZOvYIQ5PV0lNgcLGA4Z59UqBi
RGwe3tpc8669z2Ptxl/rqC71Y3HthmDtlx/GpCpxEXtPiFLrwKCuf9QrR1ns3xyR
LvBbhp7ikQbxOXP2Faur8OdBxaE5InysGD4bxcxMwle6YbjJG/Mv6uxvjO6fUbcd
JrKRqOOaSCZr7lvJx0yeNpDYoUz92jKI0Hh3vI/thmLMV5LIpNI5sxDyfMWZNxsQ
OZVdmlwDVY/oq/RVv5uJYHxxRjRUiV2v7P1+BKjEsaT6O9i6Oy6qpJedKnNXDmGG
OL3Wk44BZ16PpKlpKH17w36Tvb8zWmSR2JfvrG0yVzkdnXAq6JS9g4IBSrlun2Af
p/RS2scLUevwoWzqhg/6/AAjcQj8/yZIjRWquALdgUoTbOWSO/UaDdqJ6sZgiNnY
kYcFUZyFlaqmZNqQnOxXGmtT8hKmdD3XLoephfEnFJQGhltgIpkIFaggcWR5p9j0
lVUHv2JuBA7u40qZbI7p8x8ZfvSiDZR+npjWyFfjZZSl/3ldXBkkzBDl1qwBvFOM
UgPWqAzo0rSiotSXACgJjcAPML03diA9ebbCenMZHD/G2iBI48dEeo+mNfzu09rI
fN4wIC6wdlvCvNNIS4L21e3q86fY8xWDAAvL4qR89WESQgk1SfaSiwFcra8xT4+V
LFPyWJVNJwLpDlghxzaRWPXjh9svEU/x7qN/ay+3p9L4EyBdZ4UmQPpuVuUFvigB
0QbWY1RvMWKfN8Yi31OEujLwzjoM3kEh2dIxVBotauxpUm176izYnrTnCuQmgMVZ
kSPCIVtP3cHeyCFQkh2FqeJCsvmFgxnSfBHohiIoPIqYcgFSIdo8QAGmaLo8nl5V
Vo7N7uLENji2nfJqQGs2+DErQbB/iQhiQca5TxSRMBHic0pgJImkiwN7UWd86Obr
kCn0239RAULneZoMoVIkz4Uhp96kF7yUMGhVdanEDSwUHzXOOkXA6kmH8uAjvul8
FVLaxi3sVvPTOhfCN1dghlFMYSPOjsWvx/6JRfN3F4sqiKmDvS8d3EY6+KYzA3+Y
t2+unt3/e6mVmZSmGXt+qah0xfIMPo5KgniUj2fa469plpSL47rCueZjgwd7s3Eq
3BNXukb8FgOcxpc/lo75SXHOVAX6GDITmA3bBfsWKmjKG1zImhYVZkcYVNFYihpL
Snhl3A/sJn9e+N52sn+tXNnU0unLK836GkYzKKto0RGrnDty74Nco2X0PpFPBw8/
E0wTlOQnbDpCdAEpDJUglW6K5r7JvLWpaWeDIqG1qbhZDU440V9NDVcx55jtZ7T7
jI+4OeSj+tTeiI9ORyOaGoMFpkYTya6prRUQ3h0TLw+6IlWDfGKgGOA8iG9ZvFsK
yV3y6aggTjT7obCyqcouhR3im/6QOU/5swZ3zDJZv7+qFQesIEvMzVxeQAqa5gvR
/aKcPpbGN0BAuL5QSNcbTkDHyWZ4Dmzs2SZ2b16Y/aEdJZysc9rJak9Qr5BN5hOi
YHaP4ScC5BmNenkIC3UTCBZnie57Kbdu89PmE5kubzSARttLvMIslopbImeOvM5p
NEd85+ikDZqblHon6vso2gSdukUwnVh8RpQ4OgLkNn80PnQFOZ8K8DQ2RyuQTv5i
eR0bMGw7ZsZPOLTd2BemSe9R7PHUnnmFrgukzMzknKqJoUaXLNERanxmwpPEo1VE
9HtyAp8b1hkU1c0PnGVZM6/ncKOLMzpVa6+XDVaWoAeX6S2aN7Qn2qt2eQ8Ul9S2
ylzNHSawyv7epudpjDKEW25DwjHVf5xJlHfTDCSRUfN1lNg02Mwhpcn7CjfD088b
HpHRg1jltMZUrPqllVT/M8wsbbwsuQ1XVWUp4M7JFm+lEwNz8u4Azh6lPnUn6/HP
gilwNvMyAdJmShsiZ+N8q+nXnhh18Gfp8vFhBt30eVckYbFVUo3r3gj2+121UO5D
IuyaUbQS599htLGTabF2OqrsHI9ZS4RLjGHtukOqXoBDpkgsGcdmHyUGvPQhiH4Z
U3HhMbbTBMV3cNWPKwvTfL4nx7nIkPecUDEx3q/+We5TpvgXRRMaITKb7zaaWEyU
znETqW4WzdOrIQtgV+BY/ryuMHXgSSLdgPfP8vb5m0fn7x+sXRSUCLqHCMmkad0L
gXF17Tq78xDHcRfMXso6lvRQ75XHOToY/TALNEmcfK9VCxxlXfonqBPhSW2IdD5L
g9Q2j8l4OGN2aponJ8wzQPp1U/mEawdzCeYknY4n99tEqtv66xwsIcNWZ2v6DQQP
oHAtOwZrcX6hCZSOcN2eGElYd4OFnto5TrC47g8cdyQd1/0WgkpwnudH6e2BoWhi
IHz5nw+92RCdcFd2+YlKtWoewvBFXBgZyH5qOGwAaFXPo1Vdk/A14K7ss1do8/Ks
yHLp339w4FGrAIoc/Z/V44WeuGhoQJICkPQtTgfJvIbovht8c1X6hrvG8qHwmzb8
rMSuWdcYj+VwilCLydihBR54mmW1ZwGZl0VR+T8pgMnnTWID4fFarhWSU0PWC5F/
5tPq/+/KUbskEjVs4Vuo8x7aUCaei3ece6wPBr7LpgnkIt3bN/r3Zyj2FLYnbI1a
YVbxEsn74bjVz6+BME8vuNxyc14bM42Kobzl3QaN7ITQx61B7LyPgYUL2nSW3fy/
q/9WdN0RxBH7vzBJpHMxduGS0BsdyUrj5uCxKMJkGDgLfRentN9MeuQwQ4fMsZAw
Nzqa+lIcwlQhba7/KsRJqSBNiRqkp4J+bnhkviWsipftxnTOZI081QTPhiBpYLN9
fSsm5Wc1RBALUyLwe4WVYvOSiQZgT3nJjhV39gKQeU1oi0XsWFVWyHkRMc7vnLSr
fgEUeebWv3P97pD9HHof1HXqm8bhvK2IyDNnDLemNMpZwVBFry+P/nYWDzKO9KxP
bA89ystSCUVQhRCBXYs1XPaZqB8l5jlqXU+2fqwhZswkWSV2AwBLJU6sIxKoTV26
+VkYoZ3Lj3j1lXj5ijWseu6loI9dYkEb61kpN4P+4sU0CO1YtiM8KaKfWr44V1A0
1AcE7KqfTIPva12eIuF9a9r/f8xG6n4NXtnhTccJrqSEdzBg3qnITtxAvWfwYCMA
+8pSFpdK6ZfOl1JPXeuWGxrkER74MhV4QBdlFGqNxjtIOt25Fx6jqweMOVdDkA3e
AjYDXrm0LniUK2YNEvOjA+YIyNPemN5zJdRqEc8YkJCk15ObvNR8YKrF80UJq5Kf
DeCMRxGYDH/A1X1bevPWMRew3w7/ZjhbS383huHXvNGxNi0tpgt6opWshFXEUKLq
4d9zmc4NHIBr7kRuHzIE87OHwJOWWF1/aOssQ/fVIRCDunVGNu5AOYsXe5UEg3H8
V+ZTXqDxVgPsysQElS4EriQbukxvZAqtzBH0ZetEyuzDcYJ/FUWqA6Cs/kgsRzWy
2wD4rrPxNVVq2C1MW/9a7mp+30wZemC+39ACYJq7Wmi7mbk5JjUMwcFbmzxYQ7bo
HLKHHbGSIs/PDV+mmI1DbH78SmP+KbTO1Qt8AkVqLXkSXtmJ6XBJzfaQDnt/w9WZ
mKmpwFjqtatQt5SliCvtj+l2Fi0GSGzXJzUKPNZPOSP4wbPVd1Zw8ifXMlAjizsl
5pkIzd4o35Ym0uaRo8myDq6KNCd+j68mC24y9kEOBvghnP00sNHldZUpjZkuWMj6
qJsEYS/IDBT3XSXZCC2NNiVvX/NM/xZjCg4bKHzhxQXYV2GwRLEZJhTNJQGfRREk
RV9vMFEAaF2Qc/ewx/oP2C/nQwMY/f7mXp4AXZz0pm5fnmuD/+Sg061RlUOpDQtX
+97Tu7Z7CEE+zOFnmk4fileHZRZuLxXbgw4jxQeWFohBKVmFEL5IGPY2TKSICxWG
r9aa2CVIFuceojTZktZJKiX4fJh8tU4E6P9tKgfYDzohvZVDlCnkzMTK68AHgx7W
N+uKJ8NhULbUEpeuBXVQdGjp/5V7snsviX0cOganmtBoHRJ1zlTAK8W3mQ3HWm+w
KIPXriWQrCyc4/z5rEbWgHV++vSG92ZJYkkXz2g5aj0ouryJo6O6haO6J5fIlhA0
1l4nwx7e8qEds53dpmaeZFDezIl2Cgsem4xB+df6Ye+C6A5DyDVsS+LEVJinRLql
gHz2HFJUEwcq7sTxy/FpLGUndP7eQxq/RE6c0r8Yak7HsI72fjgl7plIlNR5ohVn
JZEAtNVBjqYAg///7+g0fC0QLmvCWSENJsAGHIw9wXVC9xZHvxgibaE4izT4kNSo
bp6b8OXrAWgqVrWUbqTjrBRM9qgcWtkDAwZIRHwbBSZt65WqQtcWi7aDdnDYzsoK
fYheZsazMQEg51xYih8AwDDiQU5ovcPQOBWfnZMPC5zEZKw9Z/7VyqdwwUh6roYa
Wk59cDfuUaEnMR1bUhtVxvLkmcS4oWwrOIy3iWnqeC4oPsFoXaeQxM8UfYY3rqh4
kgq/ukeca/MvuzM+f63kszCBPw/rch9jEOAtNbnLgecvZlUAvCr7b16gPI0Jy5xl
eYx+S91e0LkwrHEQM67F4SAX7ykE1TCj2GO+8P6xvIYY/3N5Yy0+8IdScvZ7t21Q
HvEYTnEaKwdvPKJGyPp9V8RFd7CZX0YnOWdBjv01Nc2kTstlUEcWUWwUmCux0ijG
AvAW/wetVLij2Z/9O5Y1k8MtJlpxlcjsgeWTcakIztht0pHGhlgzx4U47Zbit8Sd
ZaXV3idHRDAD7X3vj/+AKlxE5nl9/twPKA5wO/l4zwDifecEq7i1MUg1dUzYdR5s
EYfrNVnCRkCDByyoIdn3Rrk1IlveZwcKQKmjqI/Ho8oEPg+TfVgmwEfqjRcQ3f22
sukTaPJXkYmnOnai9j42rnNG4FFCt2nmH5CeITOQWqLGr4rRKH2cEF2PDjDV7P3Y
WfYM6GXCpuC4TUpt25C2Rp7ZY6q2kVgY3KKze4AYNRpImaO+rUjuDRapUNgZlig9
AkFYcUWkq7RbVUHQhNjULzgDpwa6fjbXrgGUkLnu41mcvcqX6/U6GIZuTe9AwCje
XRxd6SrdTdSHB3PbeXBoWeVXiux8C/aD0lwG3qRYAlh4+gbFOBdrVmJMy0jNV4JG
fU4+Sn4rdm4pLPi8GBihakG8EQbSuuCAV7VbbRnQifwh17Wds+qe0xw1wusYO/q3
OH+yxL9/72/lB9a0f293EwFgociR12mqnnG0IP8kNVvjJEod/Lq4C6dIi6ihcwnm
k9VakvKC0gmR25aG4gH9dcOXSLzyBciv7j7GQEo4ygDFGrRB4x2/f7G31PP/6pCi
LsAD+Hq3gjr+NlgfQHY5907cZcJpB3aTRqF2iBtUfGypZqevEuZlhy5LrCto8ELY
uEBb2VZn6eQmF21xGjoos0QHHLkP8YIAW05liA11QzEuM0QkLTSKF0yHhIJppW3f
1iFuZWvankyTKW5TALXjJ3g/H50RZmZyKwb97EIeS47K9xHSpSd9hcZQ84BbGc3B
LNKdISNAOmk9PSg5rlTNs1SZZX9RcIDDLBAaYJhBb2boMx5VdkNcwlH+22Ess6TU
Z/QJPpI044z61dAPkO2+/ldpbRGM5e20YsacWzT67LsmIGLKkRgVirO3T3GRsUJt
MpXCsFeMOnetWD9yLnfYwiaJZd/iZ3hIuzx6Fgy+yl+4NeEjOx5PlRyQuN6emwvP
qktE3Ds/pUB3VECXU85qP1lVk4l3eORQbEjmjq+lJ6my0+mI294aI/HhrI2Hke6Z
01YA9Qmkdeb2Z8IiV5xbADHhJygR17pdc+/BdFxYQu1oYU7j3BIX6QambESuRRKk
kAsIFZE8IBxM94utDE7orV4I7aizP3YFA/74dXoNLoT5mx6ozxAScm1B0VM6ImpM
u3D8GeJc0Z6fhdTllhfwEjhX6KL9y3S2JI1zJ2mbxWqIUGt5uCI5Ow9edwb3PcXU
935w2gbQLA9bB0za/PLgnOYTmdBEduU6i5UBmhv0vvM1ikR5OItDWkU6cdXUW/C0
gHlLqqI9o892v/nvDEOprWzA2hQ/5dZ6uorKqJQ4fAlZgfc5ql7Be5shKwDRawqI
UsM5fgITjTwIHqwGdH7P1pcd+QWKoPPvNyCskWHcNiC9SumHwfWy2LUCefMRfS+W
V8N2kfX9OLLzsgZvkffgUYk9z1ifK7xgiZEJHOFZDymCjmPa4atlweBIdNSpQAqI
gWyEyID/OGPbG19b0l6dYlGYEORyj+1KIUj5q4qKUclsW4qGH3tuRjAZ1Gtpqz4T
EgUWSqOPIdyLb2qt0gqX3ebdVALY0iQ17VfJQO8ryI26xwHRXSIJmlKcd2tH/kxa
xi8qFL8HllzQJxFOgF/wlZPd8iQr1BMdNQV/t5K2PFTLhBeMe7RQ+jCuA8kKrYUl
F1jyZTZ0PoqHrC09L1mFq4O2voMTnOaUQLb5Gu7Y1r6SOP5ur6DOgJ2URzOiV9TD
73Krf1AgWhWSecCkIT4qDixXIHYfQooV9n7MbDvmSVx0flR1zme+H8l/f1mYQ43p
MIUVhIPJOK6ZM0WTIQ4aCKP1eo4FKubySNFSw2nUbrA6NqtFvne/KBV0jqvnWy5z
WfEw93ZbbyBVopOzJb3yUrnetF2SxZaO+TX+RwsxKxuquRAUIAF1LRnOFBZeFSJ4
1JPqyjgBNk/Ir0RsfmPrVoSAzMXOzXfVjHxecAGZYKciLGTfFd2/NogehjT3mLj9
We0kmYlaQtHOE5u6/tvkzz2Bb++QLZmb9ZmLMkmQCxm7mp5EP2mkADYpST3WMZC3
2jDhLTi31FlF8FaeeX6IYCPakgeRugLq2mUqzW2ryeedSbZOjgBiXS1NNSA/NVk7
NE1nmUlH5T3aBipvAUJOKcP5DklMfzx27Zlcc6izVmt9nv14wFZ0KFjYTyfhbwTC
otdtrvXa5Edkx18UUf0hvODyaRvSVKPq1xSvbl+bMI2gZ8friuE2c6K3BYjyjhnz
qdwCUw8IQ/qVoSNBwvvwUVdOw0fjY7ds4c7SZOYOr0Qtbb8jvzrX0wWg/sgfgiLm
Etr1igapY/0k+jQZx1g+74jC6PSSQaOgmKS7OB92fgUCFft46wYCAOQ5tIuUGLHb
tPRCeLACmZd3hgEAVYGY+3TKfvPAgQMVEHxMddgxyGGtRgKKUwHacraAfOlyeyLC
o6mGi5bO1kRwKekJfj5QBVnbXTWp0tI0lnGQBrw9YieDlE3cXLoRkVsLfFFLf2Ry
vHCSOCPHBPw4+j0pwRvsjRMSKJOdrcFpWp43s6zWGZ1pNzKV5OFGbmhsnBUydcZ3
xh+8JhWMo6Im7ulbUUScVcNaHaM+PtJUn/XnUQ+Vse+V+3l9EeWBpFmXz7s0Gxxa
3tlY7UnYhvm6l7rae+H+C6SQtYtgZAXYuc7xG2EZ7uWNAq/2cVr+3EZwcPYXDGKr
KlKokA7IO9Kxpmz6wvYw6lrLjJc3wHX3qQ/UO8M6JIbHMqco7x96kSJu8e/3RYLt
OT3cKRIoMjXaP1EeUV3o4+Xxn8fJVuhnmezVfxqWIgY7Go5+cMs7O8vamFQV1sta
T3q34ay9EZ8excP+APGB3fyOkriH1ilL8FosCDs667CvqfzqInqcp+3Pn7kbMzap
iK18nJYIpd2ILgX9U6pNmWKXczrBhpblUCMsxfw79s5NeDtsCJZnK1wErybS5EVE
4mQt+UoR4YCOFLIXLbz/SeaOqxVavGJP218k2lHaA5FdNXsaUcKmq5hsKz8GPpB1
32U2MTeJyIBgX0WSp4/DzIEKaFPsx/AJomsZ1MSmu8HujlqKRw4c2i9sdS8DgEjW
CU0M9T0UGli//rg4yU03v/QWrijMg5IyK5hu1BKdaCRC/H4Yi+eICH/33oHUyDrQ
r2NnPPm2fn0Q35cVlvIP7V1ax9aqo3NGy5hMKdIE/j5HsS1Y+8F90fsm/x1R7Cg+
a7J62cltRImJTe9n8cj6qJIkPqrhH3dQX7LZGZwW+XpW9dwUImlbeoWyl1tetuDg
E8Bq1dvfx1xYGCM5n6YDOiwsXJSZ79/BhwU4KUbayUugIe5zhJH66e57N0GCsVa6
QZaR/CTBaok8PbWqO8vfJpzZLc7i4E9tktLDO792y5tr8hNk7mw8pAs67ppSsI3T
B5yask4M5oXyAqU6kO8XnCA0cnp0A6pS8SzCEEpHQPXPJHS8QuWi+lbH7Xe/PTCC
C/DDNnXZgkOsz9JTihnHxQmY7su4fIhngsjZgnJ2Pt7CpCjrjmE2u12YZ+FSuHfC
HNLYJdf+BlTTjgi31mhfNh/HnaXjQeGnR3LGDWeg0qc4cbxH8b8FtFwgKMO9bGIm
h4AoFwdb7LYMD8wjpB3p8q2086hH7PuRNtPsZyH0Iro0olTj8E4h6rtQjaX1l1J2
ie5AIjSql9jCbOTbm6iwspibT4zVuYvOHGpbeNE/ttjEY68b1gsKlp/Qnrj46rdm
3XVR4dzMYfo7QkQodpDso1DSJRCMO8LacnN0MjmaVr3TBWnmKWxiKC0aZPGhmkYy
pxlSqCjmOCZA40RSyCl9jatu1I1Au+MPRawWrnp3kRa2DiqinSSX/bjtozBjfLmr
aeVIuUT1V4GJV5VAte5gmZTHWDF/5UttIKMK0v88i8b2wu7TG1LuayHBB1s1/Cis
+avzcc0Ncu9JuWkOlPChAAWO9xQ5oRpH4cRluHy8DAJ0VDCN0QgO2GlM1AU52tAQ
tPhwWcJV7c7zPZWQyOBcH9xSZknPibONypn+tTf0+4bAGgfmJW4mdb7eb5G460Zd
7BRk1TMtQdemTB5E1P6SYdoA5O4U692IihTPcf0ON5RxaakL22kbedeoXO+n6F4l
/hgEd2ojmTxSVQlpqTmi/h2GKS2YI8aQOzd4aI9m3uLO5cXfUnWaQNwFC1kq4c4g
JhFlMVK9N7axGxRjiqZ+3JA/l8OCtn1jDgBYHLeZb2xdLih5csqOJ6nyYQbfZZ8z
8vCjNMg5OZ9GVVOsGLFX0cGWGxgo+HjUR/WOdeDpdqW3o2t8rp6r75QGqbk4IAXL
GKbh20Q+qOiRl2etiLXW0Mn467RWwbBqwz9wpD3C5pngjalgZnWjEszqi8l50TAu
35b6gdrG5uJB8yT+ZC5tDeM0NB8sBTJjzo7QxL7ZxgC9dL3zttNyBI7K6jgsdGXE
cjEuRWx/6n0F3t8jnLZ+SKj37ow7a9pwZ/sBxbqprPRTZxxaYNZzd+qG+TAEn7SS
hkky3QLIJ1zFC9z7xol6trsMRpYnI5Nqg0epBch8HOrfdPmb5SLzJsCxTGWovb5f
e00TiutaXty7UQXIs3cDDaBeGcN2hAIWiJF5+Qo+6lCkb0CphhTX8iejhgdlzxm+
ghL9pe8XMMKxLMgC4mIkot59jC9XJ9YmrnRI2cNJaMisw/Zm4EG09ZOMNtVa4oV5
hqAVDBYS39/V5B6iU3JD0LEM8DNdcMGnBl8/d1hJFKTbwZY2y1BNEUVBb/l47EFP
GL/Yo+dfgD8qqasHvTYNmX38Kum1YQtDJQ1m6AEGw2RJWa3NR+xqv/x44+q+mofT
4biDiIdDKC7kQDRjuaEjY+pCLqkebTgEijXyKGpZlsjbVpim/qLf7GNDAV2wHPA6
W3oslyh13ZYqGzDVKGq3B11MM0F3NgS0lPeFDTJXJtPh/4DEJtNtJLgvZsqeyrcX
PTfPJGY+/MHDmTZd8Azw2KDORx+hY/pCWQKcpSTemZXxfao+lKfmU6uslM7uhZ3p
AgmJmv0W/xa7BXxzHqcRdJnOyenCZN8GSriDSC5IRgoPpiW7XIMzGX3uEAlS6RSa
x5lC59ohkk4ako2/tqR6XwJ8ho2S1Lzjr7nzXcvMirIG+4PRzPRKH+mQPdhVPXn/
5ntuKA2amUmYq/D7D/AsiFYGYwlAIhyFkvh806hKO7Hrlm+Lph2q7tgRy8c5Dy34
dIBvfmVxjxuCMp5gd5Mc/7hTQB9KOGNTrA3dUJJEusKmKcPTEo3AqyT5sXw9L4hu
ymPfNOmpKJ6VdreHLHe1AKuK/wvu9D02giF0rLroMsurKzFrNDVJtfb3nxFvMVtZ
VV4nzOITd3OdlUKnEuVH5kzWakMbyaNTIw4hPel6vLhj90RfR9+a1DJrBaspeZ5q
Muq5PuPBRbfY0rGIS6K6DAmPIzo5y6EXS6GYTd/Br2uhrKmSwEMqpjPeHv1JNb5W
45IlTbP/npGh2dzdQbVXfGQcG7A8efeMqRwt7ARxjDXAXujB00+7jp32H+wHe9Hf
+VftpqSR2LgJ7SDwTShdjnI8JHVGiwLlGFjCZKQwy8jSliQrDX9GLjFIj+HRJIwq
Bic7wpzDXzNKjBIJLSWhqCt/fxUhJIDg4ddTHDyjbdUg+UtWzYksCaUmJrq2emOt
rhYyImDc1BJ6LzHSQBtWsFyi5r87Hg1R0F++Fbn0M5lMCAAZDxgXVeYJ3I0flgTq
2ZT0Jn9THQ03DWL599AoxzME4FHY+Tplca/nxBarsGhGDAnFrw9ToKueD7ZFKXBC
2trEC1aTcFcNIph06rD+uPfJvXHCTSkCOS78pOWxcELILkZtjdCxQLtoPpXAli5R
iTCStoaosDMzNpyzP44Qn4EKqB4ftY4GAstNg+jNAV9PpjalzLQT4+NSObWIaMpV
97FgtNpJNYas4FBgvIGgzc79AMeYB+ldsqd2RskRfjxMLlalBbnOnGfxfJtqvI6y
YFEanMPiAedonOtIjL5plFds7+SuxInlErtPHBP9/mWS+AxxYClVqmR1u+hVc5Jw
3xNFHisLHCC6QmZvK/4JaJHsxHD8PuxIL6GWutN1VlInyZ44dTIO9jrbmbE3BicZ
JM2a6U2c19n0rqzNEUj8dKA20tyjCFfRjkHbB7SCKL8mQmQlNvknU8JC8IqZ5BPz
lt2Kz7s3skySUBj7Gw6QVL7V6rGwvnKSCXxY2UK24YLyzmZOvcONQz2Wc5Rrxbpl
ejzbFhgoyWXZnFfrRidAAFEYCNM6n++DevhQz26t+nFslPjsA/uPR2p5sqn7KwO0
/mkgZrv8qzg3pRgW8a0dFfMsZphnxyb8jYfFxFjoArHQDzwHNzaNaxPWSH3FwE7N
ldWmouWYVWbEDn3/4vAz4xjPVGHShO9tlx4HiNFZVXTkR9rWfIdZvtgRgz2fzWIb
rw0TXLTsDcurtkVXGCMlQqSMxHy3/XrjE2YBBIRoyqwkQtzqwVq3qcRUiWx6G2MF
Zn+rLXlHInlmL6jV2b4XKlsMLsReRGCP9ZgDxVy8VQ/zID3H0ag8PUiGeeoBkf+I
399f+qFvDulwOYGV00r32NlMlPNhQu7M5JLplvu3VaS+rctKsFPdE3IhXzYKKZun
HcM1OunkEK+AoobgHgE21QEbPdM07R8ao/aeUpzBEiMtuFSSe5gTBKrupq+Qwz+v
fl3kGYSt8oBhHboDdpJ+Bw+L3VDZRAOMnPMm0y23pFM/N8ucS3p2uN+M9tdZdxsa
7LlPeAc3inyNWAAYY08CJlJcuOCbhjULcolHIlVrBNWLwVwMv1EnRbxa2672+G8Y
Gjrlhp4C61DtpbWIRyRRnS8AgRwWmx011h/8rydE0c/stCUqETbw//uXYztV+z4J
l7tPTbR+uXN86EPgIG4jLrzaJ6n3yzvif9SO5Mtb1Tb9nOQsmVyyoVcaGP5NCXLy
r94UEVzVEItBe7DcqfO8HAv8fhMVRKN9PecbYxEq8auVx06VHBjsG9GygSwklErA
DIRyamvWAb7VPiSPluugCbs1TiLuDR46c0f1hmDx+hiXbEokcX2wnQEURALGZigd
aYringQlzX2XLkRjrmleXcyUM02Ej/CVz2vj8HfgDfIw4SvLJNzocFEsb1dCZfXT
oqsLnHtDqmoPdYg65TJ6NlR03BruNlG/WVUhkZo56iE7fKj0CM5ssG4pVto/oXaA
blCk85l6EV6aFJdZMtwgL3wrwkpBusYBnEWpoKiIwlUsizBPEZwzfc5M8xE79YPb
u3Y6MZ0xevzQykDcW9466Vt/m1WWbmJbIM9auAiZHFUGrnCr9umbnIW/WCoD3k+X
oqGFi1y/z1ShoPMjJnvSke7/u3JKk2Qm+iWZHuPtBQIFj9XZHL2NpR0FMmjNNK/q
BvtnuaaRYfT9/ABDeIXXHuLL1Yc3utRgY2kdkVgS500jKc9ihgt/DKFybvOt0oWU
Hv6K8kpt9qHkoQXVYIakjJMFZNsGF4WZnkDa1rf3pNqYfvXnWwXus9w+CPE6xqyJ
8UqSqmFGOwBpQ3PAuvw1Z3bVLR83SCssQXgvhhYnLC7bF2jV8ZXOGy9PhxlqtghE
u9fmVTOrpDaHu8dTPTAOxfRbtRNGtBnShXjJtCC6SG6rTc8sMFIHKZhWIrFmPTvm
XFmBbd+GCDxy0PLC59xRwI6S/SrORShpAM2HDqfY1ddZPoH+ENvMPB6tXUl8uuHe
elRErf8H+Cfobu/envD2QYCTw3LRvq84a/2RQNrp+IjVvmLCOhNzwve0jliqUYHw
R6hr1GvCU5BJCfnI1kXaWLEzpB6Zvbvk738o1d6TsyGPlAvs480JVdxXuHTo+7ga
taB7YXuHb+wuTtZQRzhRy8nPPWPt1t0gvgBGJAAuhEJG9OUzy+cKecYzRN/itule
nbej1l+sxnDpaMg0qaEq63AFDZEc+xwWb6fEyFK+NmAuE8UZyTm1zMpLdVTfkn1V
IqEvDx5/QdM5VW2qcV6svVsCUr7p4OxVdGRHVO5Y9zJ3T48FqzDi7ZQpkSEhmF8W
fuRvmb3Y4Z1RXH/fpg6Zj2EQMAAXveekjmTtz+RY5PNT6qKswQiviHd1lkYsUHQo
GpQdUEMEvolWZfpMXTMSKLeoew1zRtj2M74d1FrK50hTcYI+dS+fE77PxUTrazPo
VIxO/CnhTyQjV/EYXhw9rqIY9DPJZwkY6ZN7jDW5Dug1HIoXiLQgqP9IQOqzva3X
IS++W6nyI/WCLqCBiWnq6ahmF9NbSTcf2g5O4KhWJFLknFZAYs7PBS6a0EwKS/yI
TLzyWGxhIZbY6ffARdwBhpPZ35Qqby0SMGgoYIXdDnqMwAMFP0hwn19SkCBVTfaA
VH7jPQBrjBkaku5jZ054hWUXXx8oytXobNrPucMC6WmDGykAckSN92W+D5GhgRRB
xprOfUKyriZkk6QGG+S5CdctPlbi/81CmgeDov1WBVegMTlleKzXk6VnnZ+53r7c
zIjymXtyJIBXR2egM96o4SjQGU0ky/ZHO5uRh5BBXaUyMszW1UdfQxYgZv9LjQWe
ldMv0Rv/vsw+NlIlXszDtguhTv6LB9E6/qAVSgPR6IY6gZKIjzNgR5v5JWGV2D6d
eZZ2vI3NOAhi/dR/t4NZaPhNJL5ZoFOEQzIouIsBxSRnrYmZoOFfGfXWvzw3WQTv
EPZREMbeUVkNezs3oxegmRtWP72HAyPxvpx9pEHd4/5jK1T0tEWF15IXq2dNt9GO
J5hdThIudbhyWejGP4NaQP/ltsdOc3gSHEbC0iNxncwhqH/0x2Xq3XyCHhYxGj9O
noa0jBh9wwfuOME+NGoE2CalKAPPWbu2DgwaUQTLGUpM3wqfCQCxkKFTiClQbKXo
oD6YNIkAUtzRv85gH8utupc7hz5NbUMDFQxKTAlGdvKQGXE7fc2W3qwkUzzKI8od
ksgEgyjevNir7PiJGobM4iv4wgkhYuIad0fnipAw4CYh2rO/sHjEZzwTeBvN89OK
wUIH9Btjgp2INwizOcmisfahFcREo6o22+2l+Itxmd7I5aUlmEE0yjWh2VIndh+A
iAfGaf/Yp9DEA7GsJmBSyxpyG4WN+wY69aXpmVA0BOZr1nBwa5H40jQsd5zqMfTM
CCNUAid+9L+YVXfqcIRGSW0CPMSAoFlOl00jSeJPyeiGYNQogOHu5vOkVCyHujYO
InIwJbmVq8ku1JgkI8lEWJMWxF87FWd2xRuuTTJGY862fYk42zXutDAPEXcF8F1Y
O2FRrXO6LsaAg3PpZjGqIGikVSQ0B2quBzFiyBul5998WpMnUGpL92gVLD2t/OoH
uWuAQALR61USb+4oEnDE+sOnBRjnN7azdRE4vYXGwlELhAJ44XgmWQUPxYrKru1p
B13pPtx9u3fBIkT85EO5yq2htCcNhAvsgGSc/eUmsDvRN+rJwTFM19BrcSMQ8uRV
ugpc/psQIudCv47pxalqPf3rlRHCWafyuKtzT7omwjIc4MtGNt1OM0vPj42+cx1B
YRrlqLF+BAy9KjHeOqVEJ3j8UXFqzYFcwPH2rSZf5SlBdbXvzwMbvREcmkn9A8Mz
XCkf2a1simwg1QJngplu1DNLLpURuNHj2LstwWkR6jr5cc6MYTmDo1ItSnLRBeR7
P4z5/Y6D8jlEl/WfAoWafEyL5rfvoZAnJfEBxkpGrgLEXdedJfhPj5w9M07dhdA4
XzkCy6VSBKxZQGh0DL7snOSESQs55Dc5noLSO9MS9zzHfpp9g/iGQy4kvuQMtgDC
LeSyKLxACR61L4nwR6oMO1mZbwvhtZ7nY0172K2QTULJ+OKZBv377BkkaYCg+cye
ALlgccwi+qTsJugRECiUWvlm5dh9KcdDUQNav9SAGmMadMQns2V6ym3PKENj/R0D
4oKeD4Qxt04fFuUn8wqAYAw2zZN5BfHf1iBNeOJxLh8/U/9AGc3JoevRCiY15YLf
IDvjbzTgLckvdpDKJELzq7PvWl4ULqGXafTXujDc01m0Acrk1jhqniuF/UcXvvSM
zyX7eRsi6dKuQ7JNonArqIut9jKmcgL5DpkPHYtItO/orWQBmYbLzN7dDjtpbrkQ
r5wLXhZVjCyUSOLFToPPKHYwN/7ebbzKJlbKR7I5kf81JegGmaSzkIEHf7YWcDd1
BeY/tLbpDDsDQaL5321iGf3zQ5blPowDl1kSLKV3YAolTZLuoie2rAV71/Ufadyg
BGZsM7g5k3ybI37UaCEuJbdJgxWGw8sP/b2Ugf5xfgV16Bi5ZjXy1Y2/9s+HeDik
Q+VZ9pcEVTWpkwNvSsm0Uud3l5X+HhIO0cwpAZ64xA9A9pw9Nzji3mVjL9lXL8/S
Nr4M2Z5YIzQ4/nAnBTBNrLWsyCj/w297w9xWwCM3eShoraCeuOSMppjCef5C5OQW
Z2gWWkHHvl9WXcAlxjvEAZaPzielAJwpmDMjRseIDLkQCYm5+81Kpe8/hZjWgpPw
TNP2cJVM+T13G1F4s2LPukiKuNf76hNwTS3W6rzr2bWFX5YivUAPiuatSQZYArU8
bcKFhOS4onibZrJ5HVd80VokZCyqflR67vKwQL27b7j3yxDAYq/1HjTFPzTV69iD
2UHOI3vmZaQYI6vC2iTRkcwMmwk1PF5lP00hkHjlV+g1bPTFS058IYz+j2U0sBxe
OPlwtRUeiqgZatJMMTq2w9Bb8ByOQa6vJqTLFDK9rZ5G0QDCLEeDEP6cIv3AhwkQ
msFyFrgXSSsGyQHU+IAm3KyxBVf4TIQpYu8ucjRk6usyxIMpLbO3Jqa33scAfdZH
gkaaDzckin8WZRGs9lNnFWOJIhXQiOJQSJT6jJ7m+fIGe0QkWuj0NSPWyxP6Y+y+
8/yKR/6eLzAVYxKUpluYW/BG8hJRrjzWnuWPQFuTWUQS82oTtX+5FwI3weaaG2HH
JSscfc7Xa8nBGut3tv6D6J53LQuqWjWd+ZPc7Cl2K2U/vxRoXBFTdVeXxZMCgZC4
CvdQ/q/i/qYKhrTe7vrtvK5sE+AiTfBozVNiRRHPD70DwSu/X3TXXXZNhea1eXDz
piqTgt7iNP1e49Vm4yPy1jN4gp9Zna8nYSAz3bf4pEmS/dX/ZTEb9UAa6XqppzFm
/GSrlQuyQnrIrfqYfnIV5dpyWtKzKx3L1Mcw3AFo/dYDcoYFvJOYqqdvBkFo5V8C
b5Vds50/6+fD/irq62xL4IwWURcFwzpLkr87KLFDP9iYu6vyMYqeG2eeoSM2Ak9T
TmrzFTOXqS/FjjXl7aLA5xImHGUyCP5pAF+FMcH4mPwFrk+72GEwfDV8Fz0e17Cd
uhhZ2SZ0BlBbKlS91D3vNZ0pBzuGBsRhyF7ac9WSy0qqxQ/OUSjD4MXLoqVTI4tg
BiQH+QM+tsJY/u2fhdVtlLTcicgT7aIsCwIWArCoUDrOePbCpmN4dcamiexjM7cK
KeDzvCMFcq2phvI9Al/lnZHotDAOMf8WwqHiiUo2u58LvpeBWI+HSww7n6pwMXXC
Pd4A+BofAXxdmo6HYFJW3//RpOg74TLV2BhW6R7yYApsQyKh302c+TozCFRIHmYO
+QodJRvwgZymOEU0RF/RGDaIW2ULwTpSiY4R8b7hydbsz1btJavkzH5WXAz8yr2h
0gwArLX4QLoU08Y+nXg+UGzxt0YTo2aWP9YH1G8UQODF5hWXCtdlUhLJtogL++Et
DTLtlydjvn5KxGo4fFpnzyGlE255sA6OORo5FP9TnBidZBWjreM9Rugen9YGGG1N
rsJnznEKL8FfOTFvQlAI4L0is8tKztvJ/Q1Sn2U5JzMIO/kySnMucxKAqTb1LKxH
c7R7KjQCMB4kO1PywR+bXCKvdLFrH+pL664+2NsyLdQ1czufoHKGab8Qhsf5YTjK
cvOoa8aK4fdcAwcHia+XvGR54/2sz0DfONGQ6rAW8wevdMfHQWMj/+Eb25gBp0Rg
MJxi5UT4BEk+LmtS1YFqAXRFdWsuC/Gw7xKxOZ+zwV65ZBmo06zD0MJpJJa09gBG
FD8X7DqQNAihWleCiiHOXRZxYG/QTP1DOT3V4PvadJJfMCbjjE+xw8lVgUJZDyFZ
5vYauND3csj749fyywC98p0uxzJsnw39uQbpRGALRlqDGOoIPtcfRu5E5eYqPRB+
8BaCcut+6CLoqa0hNcufQQ7twi2cR78s2qmmqNMiGCGoJ0eLDXDT83uDc/T7CcH4
As8SsWADcq7iEQa9J4RQYZEynqRORpO1r/2B4L/ErA7eWSerxLm9PIMc3R+FzlR1
fSXK2HXsfu/voMgs0AJp9/NKDLIWE12P/qOV8ZRSWRoZrEGpXELHbg+A2lvo3enL
afeAe67+4drD5Qt1iGEbOxnz3mme1BRwX01P6TBLetf6V6iOuQp2rzvFrrdv1vwh
7a2jBJYtNz/nFULJM104KSgNNLpCjWcLMd6zFy8IgxYzDaqdEpzzViBVlE0tCheD
p3K29lhJ3QsBoG3xh1SzEpIdpa+SMfN/32R5EfGB+wwFGRnXZ1rUoZXWW+yY4Rnv
Q84/KQilQQxf5Eq07IobuETo8YwMp9PqKdwn41YTAYEZHrxyWwVI8j/MyrgmQhL2
HGH+9jwi4+6j9maMcSzJv23LEK+b+UZfLLd9yQPmPDyDqXZiXNvqWBy1Q5371/ac
VGMsvgFO14xFBpzUuffn5GDaCuBF0DmzDz65TwzNn4ByhoktiKPswbPYIbXu6QK9
n9X0AJPuP42ZPy4Q86OcrU32IB738IwMmr5sxnMWSXXLs7IHuE5Acxh1RV4uTCbt
RQGzSEmF+MYIzlgEPTGnP54jQROizFTDu7UFJZygB27FTQ7MmZRDxGRfgDaU7VEx
n3KU+nIPaH3H6syGJ4JbUNaoa1E34OqGL1rScunYsCAmVhkWDYaE5IQCfQSfSO1I
fNMpFLE6G0oxt0udP/SW6aWm4ZNnhPRr+WqmbbMLeboTq/uL0I7nFvCLl1SNzOXs
ZlLmTOnTdl6/dP+Wu5C1KI7qbVhQVfDzo9Loz1rJ8UWFnRkvz6JazXsElNyIJVd1
RKpXmfKSqEdAhgxzcW5g1OUozOyTbWYp8sqUCZa8XC25fhb0wChhjdfdSmFfWzsp
AoxSoLQIOR7eelxPkq9OXBwM+8B3wnQkelXj0qNMDGfKdiIrDefK5yhgGVtY4lJo
Z+EvDwprhxZdLOUaltQdNxjVp30UKWyBmodciTQIaNyWug8MTWb1shcIFvG2hCMD
tn9Ao75lyt6Gpfkrvks+4C+HES3M0l8ZJMcEU03dXlvhOG/o7cUogf+mcvOsl6Vi
5Z0NVHxvZ9QP64vM2R6yGtmIuKgxTgilQU6VTw4zSeFx9qoR/Nlydpg/E/C1CaeF
cL35qrr6wPUkar2+vlewvKzzsH4E1mew0Nmu0HFZhcPSKei7O7y0uiIPaQg/8/bT
wqgu925MFmFoJ2kWUFlFGRGJyptG57Hmj4Lqfeh0N/dXpF/s7stAnFFMoplbaygP
kd9lbLCOVdE6TliPi9V1qWHXT2QVhnfWfq5kTOr0n1uD2BBOd2Qt/efQKHa0lvHi
RLc224Xgu1M1LhmKVZr3yR+ycNJyl46PU6aN28XfSNCgyNiDYdiwhHfcL1tvLFUE
2Rhk5Ja4MkVu3sngmCH01rUJqOS3s5cBTLVbEC2kJCJjFIskhMXriMsTey1V5NfN
YWkksDsSyuFRc5MJrHuvzsJECIVPk1qXyYsxPMbTGrEoJHU30wacIgSPIJ4fG2uD
t5bWhXXGd8B7foZ1x7DZ4c000EzfA4O85GyyawOTTR0S2bK19dCahY+v+20ioC9G
0NstRne8l5zF+PPYbMQ5rzX2+kVXdIP2MYSex7kzUZFUZQMfFEgnDMVGDnMIJ/xR
yy6pl8oMc7wYpDI1zZwDMWdtKPRm0BGRImD3Oy4rtZJCI6oro6tsxp0/ltB29RMn
hixtwQh9n1F84yJAessooMIzK/a5oySXKjJpekxEPwjAWcgNkm/Uggmcmxi5IDcZ
xNbQTw+gJlZWzDhlE/aSQ9kBs9VKU6c0yXalSsw3VXfuT2Wh6K1VvKkV5EpYbqSo
jjwshN7946dSMhsMgGudsIP6ZtbxzNamae2VdAT49+td7s1W+IRrAizl0k6M+3jP
jXFkQ8xLelq1Tmq7XonA2TYuDhj0gEjzg8G6G14rruyVyR6IiYroLh9WTK7teqbE
tRnrgy9QApD4fW3O3U1urPxUZUh2BvWXGaxqxBTSguQlbguPDyrhzXv5r9s064B7
RXXbpKyoCNJXbe1nG2E0mNz5olqton4FPyo9SsDDnsyDLTOb8OLbfO5Yd9aNHkXV
irtMaZjM9N6g72MhJHTn+JEaLNDvLjC8Ob0e3NVlZNs6gICIUzvFM774WtAieLZv
Z41hlVYtHOUnjO+O3E90Nx3X/A0ptTeBrTGISAn52IjwbphQmNURrEnxA40SqTNX
dBkn3pcC0YVJT8g54okE1WQkRPhPEuFpd30S80YHicWWYG9pg//3+NbGoTqhj0KV
XGVUhQG9b2iHlcOYhfBWI8ltLRiU/+YgcVrxluSk3MwXYh1J2GPkMWgEYkQBi/Do
R9no1/QxpUAP9tqkTw1wNx49YUhE3AVNRVvLY+pLauY4bBErxurSb/SsGxg7Fa65
e+j/myWdNiY3lLL7b4JvtqQM0jtZldWezY0ZLTjwXeGmJCe6GGeVDWzhwwacuOSq
nWPKF89LTuuR5SZhOudtT/AAq0g+ibmO2gHwwIVqn7+ygALNTUTZXFcQ1z1XFQBJ
Sk/irQ1VaPAerJv0EYb6J+K4w87BcjWrHNABCVY8FhAhhuVqwF/r9Cxis7K5EVx6
LjxLFiSQoV5CcdffIVVKacpGxUaXKZIe9DRQMsiCEHa56FDw/g+OKvBJJbWbx79G
mPPj/uALbcvgknJT2XOACOVDQQVjhuootWlwJJg8PtSrQvu/RuKC6slGCt22j78z
JqYCo+VHDoKPqPAaM24Ea1EvdzLmx9aeR08YwveHsDK53Dq4vZVx27zHcqRa5iM6
K1/TIBLzlBwuppv3mO25Fytnky0XE5GtyxlO5beQoVt7lTdXFYOohQnObIRjlU1Z
Z5HvSHFeHdYqEHgrWtSr0nuKSVExwTJH04H8RM/tpHGdQMJQBiJ4aGxYadKS2WDJ
QGA0GTfpyQO+QYQ1yANebPEWTY+XdiWKUaiRDT0UWvRPZ1h1cUH3BgvqLuimXD/T
ETu4YDrkReYec97xeoLgkdztAJ/emDeFRy/iWOq7+k26HINSrihIV5N0PdqjQaME
zjRQ3FSOcbva6deFQa4DuZkXxrswWy81XJzTL+Gcwy2POmfwjFBBfXsL+heskf+G
7M6R1SmmFnjeUdodByt0EfJA1eCreDWzZ5jBOHUGjglAW2ESn4Jwx4v3EFDstvFm
ZWpgY9Pob+lM3WCfwgOeHdFt5HJVoMu1pQQeUfO2EWspyqAXlb2cp3HdKCyNfKLZ
YwSEUy2KYTWETp9nNlKT7Q==
`pragma protect end_protected
