`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ap1JBJDxBjInXlAb0zPstN+eqxQPJoSoINhJKqmB4kx0vO5/pXwRk1NYm2MwBzYa
/lxFoFS2Dw5l9GsmMbnaDlb3gdSJLCsSgI85BaXy0uBvdPHRwLYvFRzQ6ToOSWFu
8vTLhvR8g8oQKeAWtTMY87WThM8rjp+djiV1G8MUZyM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
NcsTQrsYC4UI59adZ1zUAU1Sjc3IZ1PJJg2n1kiGcj7BTFN0hSiSASHJ+S33wvMz
8KfBUxwYk7QAu2nvSTgFhcrD0p1wdLllL/LLi3Mpc9sNauI+YaiKc+iCcVOKmgdZ
P/Xc+0m6umMuxPQ1LZgdzp4u2KTuZQIqmi2qYYxjAhCgu2GXSXhoVOulA4u4I0Pl
G+3dsp8RUxp+BT5iTS2xIRRMPlhVP0yL7ODAYz6X2Ln5CiTKk9uE89St5Ub679FV
wTds2vFiKQbCmL5mpzYuLQ2lU12AmLB+/hMHi1VeYRAvZn9/6KmvP31AdIjaxw8F
3gBLDilzcdq5qe6sa7ChIlnaB7RhvjJs3MccC+ISnsMRv0DrGKJLbLJGfUTqbCsB
3NhNxMNn/6N+vASD5qVaQVmee+7R3cTo8AEwEJ6t/bxXbd9Tn73nh6Q9GzI6K2pL
K37x2gIUZE6jxpSnTRxCDhR3AvV4N4c+XeYQ4sxP/A893fmYHqMZlHQa/657rySH
a4+f4X+VR+haStXIiHMLUsN3nXqV2k+MqmaTrOlaUGTfYFlW5lPwDm+ln+Bnvl5y
DZQdFOmnN9yoHVDvnm9Uwp7ASL4ZIptvWbQDFpdbg+ZUs7gNn29ug2AGijGDsQQb
XhYoBamZ9DaSAh7Wc2LLLR4NB9ULCPVG9yqicaE7pHGks9F92lGVuPitJ2Ang5K4
3q8YeOLpZKXG5JrCCqsjcaTmfp90+HZIf4sD1dNPO+97QQf6icD//arHQb0hX/fp
JpB/9ZntMkDYEpznrnbWVm3AXZ51L8iVGsj7d5FNE/AU7WH5mDYPy0PLnU20DLgm
injJP0jJZ/9VRLZg3liw79NxaPXExzbm0iGSWw6qZ7zpot50QT/CJAy9r+4t8dbQ
A15JLd3vg9M6nZQbBGIUL71tn04h5IUB28c2XVFJo4Ng9Jh1F7Et0Oly9UWs5vBf
YXknz/dS1Sp/PgAiD4Gefw3FqDIEkQHx4b4OuE17Gl2WnCCYKD+nUbtFI/f2+FAM
VW/EPrIuoTowtUJ9KJDMukLSVMTqJSQkuZZ5qo9Y9jfiBzvNmD+UaefePFW9mEXa
oQtXqDK+VW7+P/2dUp1BdXel1HxyG0isrhQJQABXexFoLvzgv/uf9V09SsaGSKij
nLO8+S1ZgT2XR0aC5eDwTBJXfsOVcKyKD2Tc+h7OFofxYtSchnFvYDEoXQCFx2yZ
UtOnWgiiyiu+/7FtchsgqQi6nQGsghYI81NIigKIJzZ3cfMQc8zmgcUr/NE80Cws
QsOwhfU7SJfvg4teV0KYJO74Pun57eUctRm8Yz7jLmgyjtfNlNkiA0+Tln3Tbcfo
x2OqvB6FiTPM9Yyb0K1QF51WwKxTMtNUOcP1tbTNZgKjg8+TeAmSjE+lNBZSmXca
4m/c6dhPWvHHkxOK49gyGu9drL4xioScdIxH2gokwdHDcCK5KknKMZsEzu/Hyzll
lOyLAeD4hgJjW7eFR/8D0GE1LQFgjMtAbR9d5z34WniM8m8DVzdMdvWcvrliUe+Y
nIY7032aWgF3JgvosPHKjDAOADF/FBJOnl1PP38dZBkqKZ7HD8+dMqDEVbHbEaHw
B7IoT1FDXiDOJBUKmnAqYSXlgGrsEDsHyotd+5N4U6Shj43DcHBJhGU13au+rb9l
cWKGe1ob/sz9H3e9EkIshaKbcivOZOZYvNlOPyQ5tU6r6TETYEhulqljxWUasyVq
1EbFda0G2JFaFN3vaPM+rZl0iuXKk93XNYsfjNuLXWX0+J5Sz2TJgd+CqpLgHm3H
79Q7jqE2+r6wCtHFAHayulrXx9zsrObelvQ/Hf0vjZIa8b6bLSjxiSZ8LTmPjqi2
WBC7BuotaYAFQ/r5b+9BMWIsCIStmOd30i2cX/L/kudCanxXsR6+QRIgkOiCbsY2
KpsrhtmCLyUf1XEqUC91Da1cUswHZy+EtF1Z/8HebMV6u7G4DlQSPLJhQjo26PYC
LHmFjW26bmTbAdXgf0i5yfHyJWim8icgQUxWl6SpQw6aEv8jreskwjOLh/nOz8ar
efjJ3Eo+XyvcUKlrV1O9WLupbSb88QDPiXmLQCFIpZbTEWZFRDoff/3ezC6MF804
xPbgg77J6ea7K1oD1rTmv0jJp8BI4ABv9aMhpV2WxZHwt49Ng1stKNdOsa/zdaI+
rrUgvebEntLJFp15z5etW0dyqAz5YbnTgIcM1VxzazFIwyb2m651nUK+9A1yaFHV
NAUx0S0bdg6nCNGHiE4md8TpN0uocg738opIyDa6v/8JMuHjP0Lwjd/QqJiVdTT4
Tz6Jpzm09wmRhrn3AsxyyHxjC38fVrSrtwxKKiF4piFVSpw76QDE+v4qEAQJBRIo
VaALmirRa+68YOJ8gixz5ctbDRi8/UZgAexhjwidrkeMA7zk7ntACc5ns0O2Au6Z
AIolX9MTrNfiM6Pjmse1Ou50cTbJ4JrJpCMOE8LvpudArf/Rk4xUhoEbeAVwQB/l
EghHzBLeq9BBC8HdN3CE62lYn61boiyUV0n+hdORrcuQpQjm24nuf5XlSMeLGuUf
LvroZw6iT3NjfkBqb8y5VzGQxHiGPsk+lO78lmD55aEPvj55RKPENfabHLx+ZH7Z
+L0UVrRxBSbpaAxWO/VmrZ3OsOU+v4TXwfL4+8Ej0v+amhlHW1nG1s4Tn8iQTvbk
PE9zqFfaM3d970r3fFMTbT2Bx7PxmG7/ziE7nodhstafyEYKribkerOgQGSp3UQt
w+OpibXTfnakk/8k9UPZghXLhIXCzhVmt6cmQ1pFxyuhom8B05wRc+OuJOfXzgAc
ByN90fB9oRCfMnD1d13ZaOHGSToaBu8Dqgb+WbWMsDIG0ynaVufqNhpt+bR0PjZd
xt2f1DVOSxe+ShmwJkCmTaGfm4nRonMbzwFWQZTK/EQvuzMK6hqmByXe7dg7mn4M
F+SkIUAKHkoVNEG2lPjQGp7m6t3CXIkkR8BgRl1TxnuDJszJ8RqITOODKHiwglPq
/JJVNOUp6LU3bZlVzdlB68ixclmSIRkdxiXIx6mFxTJJ9qsfu0Om62IK+dhxxAkh
M4e3WAhCIJxOBXDqm/Bkkks/RJqjg9NTKMrFIxPhKYtt7JfLFkyWTYFXJlyTGMD4
`pragma protect end_protected
