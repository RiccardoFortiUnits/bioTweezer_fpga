-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0zmfkW7W8UokhkNN785K2w956dgGbCcRsvEQsgzOTp8/fDFJzcbmUfwrTQ/Zj0pYxMpQGt+y5jwT
pI7PIzO84qCM/ADdq47nHjSn5c7cIidQVuwOnn/QvmNbpnZdph32isoCSFYv5qcnJ0bCyDkxUMkw
tbOdC1boYOMuClry9ryzqrzfqIDvxAy2JSfKwOb4wq8wO1g0x1OTpwZkxYOawbeqZXz/+AXNgsvD
kzsVEEu2yWG/yexPDsn/QI/xeQr29zksRJNFqKkw2HPE6ekCGmZM27SL00e3TVTkeYnmJ8dSNitl
FBdovWcmoVja3w1iyS9hQhGPzXPtZL0Ul4REew==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3024)
`protect data_block
BkfwUqdgnFxsdFoZi8JoW1Zi2wfFZs01bDNRVoeEGi+dD28pe6ogntH1XZL9dX+qHxqV9QVEhyOB
a6LkcYLU9R8FPafZ53M+WQ/MCuwSU0nVtr7gzHXXl8TbEK97S3yxkpaeFU1kGYCHlJIxPoBxKa1b
302z8/QNaNogMHENQ0OtjEVPbj2VPRW95K71SV3CrkXLXFb73ItG3C6xTPFUZAWL2rIZLHayfkiH
vXkDMYKX/5M82zbP0k3Vv3g7CyoQSfs8Nj1ACOxpsrYliUrRaz5YbVO4/d16KppTJ0NV+pAS4lN6
JBJRpTUARjbNBqxeziBoC6jDcHhYA5hX852/iYq5h/cZ2JMF7a22ISIJ18H+ghA3Dd9mgiwKGkEp
irQVJaRWUgrGUSNzZTCg7OLLs+f5kEv0WA0bMkc5zZlpXUSH2olyDI8n7fltJMRu9JM658sL+x+m
VeNVb19fgp4LIu4tp/tDlHQX9GhHbHLYT8MBQb7msaDlyVjqyWE6Q/KVkVHko16FFwDcx8CkJE6A
6Ce0U2A/UyxNjV4lmehx3IIfxKUPOMwwxYSCM+v5R+gaLYLCFXdqp8qssfClENi1FEoXKhZBZ3ZO
H3R6pGViHq4/8hJC2P3Od/Zc7hxK8OqumywupZd8z+CBFC46AliBA3FRFDBU65ium5b+MPADtoxn
5SB9OuTrrdRtJFYyb4UzvtboZ3NfUYQktUDOq6RFqiqgEGblVHAssKCBqLsLo1NV1bKkY4oCbIZI
qciWNv/RpMi7RqHQdQw0gqt2zLL9AAzLF1wp5f8k8Nt8P/l0qJiOzZakWAIqqm/rqANnKa/tCFkY
5HCrMV4xzmmwxvDaW7g8o86F9p9Ig7xZ969xlYsgGipwkahbtFhIVYNewJMKMz1TaHbqNuHevl69
Qe4BXUJBsmkq65PZf3uPQXf+FQaEviwbCPEzzIgIWoBQQUjFw30DYkwRE6Li88OfhbXK6GZD+bBB
V/G+/V+l5QlFynV/RKZ8mWWhxxMXCSufAm5/8PlfLWC6ojDdnO9W2xrnHLqt2+F6He6KLTxXcMZk
JcaA6sU0zv6HiaP48edBQy9mjxG8sYdJDG5b81k6WrZe27qP7iKQPgG0wi+3xDDnRR6ZMqjvPoE0
cekVHbbou1RItaOhdWNdbFlNbj5qd+YMIwWmtN+gi3rINAxIKAFDF3TiqsADt8grOlAfG0nOPi2u
Y4TApN2tVYqd/tvoj588p2xjAMloyp1cwiy0P++ttQ2hguSArKLQ1xFqiMSkT8Ds/1uViFgAkef8
M4l2CM1Kp1gx36nxMs6A9ERDBiWvXxv60TJ0E/hc9ImpdAWGk6qHltwUuxnZdh+nc3N3GJ6j2eQm
AQxWKAJFQU/sfWDWueRKAkJiJ/91fJ2ODAk7eU3Bvmt2opqsOzo+dRc14MjHC0lv+y3IqmESQ9mL
664ymJ4Rk7uOOgcZvL6eSVDIxAJrYu4UEqCbAZUfzxGpxLwoAiZE6xFa/6FEK6kSIM/KScuxudOq
RDuAXfRlVxnQrWCu98IWNptKf8Tn48kwznVV/3ENWXewbZtSPnfwA5OV2gXLXY6P0bONGnUfqC4D
wNv7zun8IbzqOcSNhuyV3Au38DqKcek9ZdN53BdsBmSn/VPyM1F9b7r4MYB4dnl5efYn0qHqXzeC
tXRoY7/kkPPIBWIVh0WgY+RZDYMimToI4UwTFhYZ34QxsuQV5sKS+R7vZejaijvSFLIpKyLRMd5y
23Ea+rmWs0pIYNe6JcRF8YIs1KAf0GwrcrEjQn5xfiil1KOM+FxUwv2mDi14hnkLp3Jvsf9YKkXp
tPbFBxqqJyGQEDYdz0nRlhxGdsYQ84t6oz6IdHXtMJFrI5BL7Yildd67DnpUK2e6vsrr/NSVw6s5
nmKw1C0oWvscXtKdpEuzGLcftuJqB9TJHrm3aYLjDaLjAHv0U+MVoQATJbphXiEv80mSrME0yt+e
p2AiLxDexFJEwdDLj9Xqi3WPXiSckNqvjnXj7MQjblUq0v7jIuICyo+HWp2CKOkBXN1QK5kC++jz
8RxkOkSipjvBxIdQlG/9ICdAgFFIuDBCHob8JYRW9aBzS2n72p5l52trhqj1agFM0wZ4O+ho82Hf
H8+O6ytMWMDKqpb6XH5GMj/a/QIGVj4qdZ3xHyRSSEb5JerpL5hSQX5GBkZvUl6poeUzHVg1y9W0
Ne6ZLoHciBrnv1dS/ml9nnGf2W8h7BS2K5HnPBiPZ/fGhL6gEwFikRO3vOqBbgfu5rg0nSUCB/Jp
+tPgq+CyNV7qd09INT9MZlejAeXqhSSPgEZha1Z0xUlcnwo+sJi9ZiVD+sqF6nC2StblUmrMZ3ug
+wtZU/XmWNWBJhCYVUQ6+f5SoT95SwgdORmtUts/Fy8govj2QL8zLB595pwzOUJbvBTqf2YlbxLU
B++61NEskwG5vCVePNfXwmDoljB7BzFvHBFbb/8Ra1nkVUsTbF/4n9qouxjD5VxRtvgZVKzWsiNA
yLWPsGMA8fRHTMwWFkoRfdsTPDH5oJroAVogIAVo1JyRrcg+10H5Vj162Adex3kPSU4vmXAWok2r
8orxP/msTU/k/pys2chS40N9DD0K+02cCIzJFF+e59uPTQN6iEOcp+T9mH/7Cv06JcZfZvOmBo0C
nhq5JyNajY9GXDkYNYwU4tQM+WxvH0dTbdWX9qil4xCYLrUOyoHcBqqcmmnAftb4HqHGnEdg0++o
PLMK8aUsFIPOLjbsnSM/lAtwPi57RwJps1JtqkRQTs8IsXjoIrropmgWMVKHUVpxlJvCJMCyFGXA
0Vg5BIlvJO9yuvgtP05o9zX5QGGDsimetdK1gXm2umsYvhG9qXHx6LHYd/vsYY9dBzX4wtV39epH
N46LRIOYrzCYLKadmvdr1S4WqZiKQrlZ0D+kuQDu8IVvXP8JF9B6wv+ElfTA1LaBI+51zcRHxsTE
tUdIMHQvm463Fc8Av57LCi8yORa+5dDbEgZNHE+nh8VIjqWE+K6DnPkayAFjNmOagqwC2Raj1c0c
yyrJ6kY/Qxq7U4eZWoHjEHyAPBx5w2e8sfQ7ANeQFbeYutk5sIgo70WQQrLMWQyzxI2Oeozg5zUr
nGEdADkuQ2l5uGWiZ4Vw0LwHF7jwVUMBIVH3aasKHGEUkk1vlEVar8lDfmF9Yybkjvu2GJnCA0rm
7hjkkv1vf+jyu8E2+A5IhHHGJCGk/UZIueRcNcVvDUHdAMm5+5yN/yylTAu68P/L12/tl2942eeo
83MiM/0Yo4gMYu8PJKvX6NnwhX0UxET6wfTYnTfZvQizi0yuJFMMlJHbMbXb+ooW+XDi7e7/UNG6
OY/67KkxRYOs77mu5SmxfibLsc/qPZxRpmlQK4yPOS1EyZKsV2YMgLM05CIP/c3xBNrk6BoWr9Zk
s/3+4K/0/kjLXiz+3ZsHa/eyBBrzEWvJthiUsXk7f8m0QalsJP5jE3ZeSftnPZDWgNH8SrfuCcf3
X+SPF0EtBTLuGp1De5bP+mR5PR8G9Xn2R42FTjChfJeZagJiul5kmOJzlqlB2GG/9sjlGckP42Ah
AHiYBjTauJpPbvcQkV2xOKDFuAaPjZPcKkBJLuaDsHuWpndPexrzq1TRHX4boyNycvOW9wHb8XSN
FaDaHBFEYBSU87/L6HICvu9RXRVIH7YDiINLzw25h0KElgmK3oHV4GIl+EqQYlKXnXT1JrCcjOTe
dKsZv/GHYFqvW35lfbUJGDsEpcQGe/8sd7SyXyCcCjkriXRNvl0MQQpMoCCjRSTbvefy/19Y6+YW
jV68wyRfg9cTZTuMFpakND+UngcSjvRYCtfpydZy28IXCu4A+i/TGv0+zLve7wPMdAwEt9y+uLQb
5lhmWrMXQ1RsPUO/Mi+2FEszSNK7et9uXZlUKJZzXEBe/q8iEgVsCKUWNLxp01Dbig53dPoxuIyj
2h7nnNgempWr3o0qdYwCMdMYQhdovTkpGnH5dkgdE3QE3Aw4UsUjeIxta27QhlUifquMzigcUx1t
vli0
`protect end_protected
