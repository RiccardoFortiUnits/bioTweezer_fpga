`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o6fFh0sFq7Ha9Qo3Oo61g25FhuTiy28qfUewSVhalQqGHZqGZ0Sza90EctIAk5iA
TQShLdLpC0qQLv0UIDkeXH08SonA2vWYyr5oR8GwPQbQ1Ga4SZu1z7pd2DqyPY8W
BUMMobtOIZKdNxLFGHkXn5IS/vgEK/7OJ3uQ5mtGauM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
IBCepvBS24q3n30z9enIPaGUHZYPbaAOwvLXhjondP30M7IeVIJbJh3+hBPxi1lc
DZBJg9RDQy96wJoA1FPA3WegtnPi5HXQwxMzIvGS8b5b3YjS6OKyFy9Ap1CXdaWR
8c968C4+XnYW6kBx8K6Sh8W93i2clRCKFsVOLRxP2ipXe+wHRaDe7wmeCL0rNjVq
9B+BiJMuwSmWfp7pfbArqTcDiUK09CJVL5bd5gcUJXOmWc4c/rvMLJIwWxXWD1q5
w+/FDnlRmEiDR9nbbaMw7KdfjHujs/vSI3MLIqNrX3XsaqKrIYciuq4LIRLaYGkI
iEx43836kLdxNBjdROlW0//pdLsjyvIRtNI1+4GAQMA0Y4N5GJJAl3KOGZ41PeGB
8tIn0nzHcMF67j2uWFIQQrHQj24AX3jyqaTr35H1FERJcJ81fLr3qGmXbPu8Vrqm
2XnLfjDduv1xSWKprMvMlDcNt45J+z9QNF28jzW7Lxa7G9T1KzOK4Rl/qaHhrfAB
3W3a2VzauVYcep+6fhQMqeNsgyWoILuE7hyudIHU6sOy6AMykir+io0kqvUgRPYc
OcTv95QrWrgNUkXCszW+O/Z1/Rwr9bMXZwdPLRKdsDYLRKTNAFj06ai2dbMVbp1y
WbfzgxMMBmhB9+IrAYqjqRmR6/pg3g0e85xsBv13AmPiKnvtLWDBVm5nAAu4Y0kp
TbtBkrOswppYkz4Eb0V5KFvKkkXRyej5GVgDVa3jZZmjyYh0vpjU7NS5DeXf8usD
OlBzwFvC4c7cH2ubgogORwRJ92x9rwwj8v+3DbeQMEJuH3L+MrVJaF5sMHzfH5xb
SEPKwsl5Yp6ywqchUNMTHLRPE8NOfTspj+l2mFfHdz3dqZnUvRyLGWbuXrqtAiqL
HuMYXy9jJpAAfwpJF2ONWv59brb+9j/dcAePI4Yx7mxncScsaK4usAxpZNcwvnqz
XJaJlBPZYiL1LA4rbdt0ToUfHDdMsTnEJlk9+9nAvfZxVOUqvIEOsIh05/Fg3uKW
tpuvqmEwDb6o0IDMbinCwxZbiBZkPYYIb43pEgbdKShJZ71m1E6s9JIBgWM1nWvH
e/uVs3OVyubrpxOZu6d/78tZ8Ql9/EAcgTVn/exWWxVQCsjcSqUINHsH3sqelHqn
J485mXkmfkl3+1VE8QQ5Mt6QBiH5iT1Bc7nVgBvxiueHBHq4k5IKndkYlW+Z2XJh
5lhMAf9LnEuXNN2QW9D1TL8cmBPjT8xSQZaJ7UDWhdsvfFk+/z3iuh2O9a1wei5j
HiHApDJDaymwdm/LDIw8tTATcYETb2hu8nMmAI+gxdXJqzDK9blwvxRNleU55l/e
e0r/JkxX3dNASfxa/H80eb9bjtaPyr9Q1ZiszadDoWYd9Cu++XyrKfK8IzOVQ2gT
OOmLuJb3tyYTdSLOsLI8gTHWX359qk30Xo5zTt4MHGziUkMqp3F6CQcja6nkK7et
ZBbGVt/2H9rM29a1doSEKnzxcNBqlQIGC2r2A+ySRigwYfWleEtNTHUaqZ1jHsNU
e5MC8r5/gAU1bYzFw2r2WUt447WkSaedx21rRvZ7WI0S0osMjLzifrRN3D97GppP
bdtZlK/OV17TdZicMZ7mL9hHsxSbw1hHuKWrRju1us+eE2RLMlrJ10uKMxcJhcg8
3oGv47pvQyeSqil03lByFhbGGYAiy9xxpZLs+9DAzjHg3cyStKk8WVmrop+JxzPj
dSJO7epr5QT56uE23i4e4BkagU+7dmWExmdQptkKS48K1Um/DlbNqKjrhljgQE9y
p5FseiZ1Eu0sw7BQmY8nxzUycGx1ItQYh2fC8CZEr+bMwruUQIha1AHilTLXr39m
T6dIA/3LEcD6fWkmzPvCN2bc0k5kG2MKHjfdGLRzE6DAn/NOrEoQK4rJLyeycWy8
n3Ks88Kjh+TrFjRnuVh8P6moF13xp9FFQ0ScJz01bOeZ76RsvMHBtRYNdg/vF1mK
aFCrWowCPALF2plJ3FLyERPp6FbaVvK+7n76hES8GcwSSP0cB1NhZICY5pnpJDto
csqYxoE60MM72K7yDLuNb+qirmj0uw9qyYl6XPvABhDInnOuDAXIVl2teT5T7WXM
oiEdKGBi7dPPyAwb8gE6YVxBhozk8NvNJtM4pK4P2zJhxYX5dsCALxn7VueUR0h3
F6lVox+dx9zNnYLkjxcfJA/J68u7rf5XoVJ8lsSZuB1gEdnzegckpKZ/L2JEqmCM
eTUN6ApLJ2EHwMIQFcEWjzaKVyQpZ3PM/Xde/pcUAKfA48HLSwDB+E+ZBtB+xzuc
sEBkeTnHlY8KUJBPDwVj3D1sPmuRWlSyw4NUv566BEdxkveTuqzrqa8ietO8xGKO
ytR0BpbRrnxyCl5M/6Rz4z+RsIzQufM3t0RRSBaY6N5q/b0Yh7cVA68/oijXJCFQ
mV/LJH6iWf1arpNNBFtlkBQi2e4IE8ISX8+9yPbO+kZeEF7w7NEF01qVal6V5E7+
+EJkITVOoGohgoqO+ksbVfDYg4W+wrxY5SESjIhe7K+tSJYmt/i+6/UG6UcVGCfE
QYnYua5znXonH8VxDLvXoEvUfgx69H4IMyFND3uRmeRAYCCOaw5edhSfA3/A/9eF
agKdQcgHnxIboQ82LpA9yqxRifv7J98KxD8Qd9+9GgYKLZjL7flBKjlcUPlT8nsO
NSF0VeT5FG7LxYF186s23acIp0XtnDTdDFWZ04HoLj/UJo/Gs8nrNBnijUwjSM2t
zEIwElz86av9OMlAHtWMS39UXTbY7vFvMcZszEOPX51ld8qMjRCm5OTeURncxABQ
gL+BCzLBYPipDs6T6mGQ1egQIN+S94JyvZJDbpBYERi7e3E/5N8VvOyyPKG8qISy
zwCl+gdjaHn1aZBkI6rOcxpKNxCxDob4UateFuWtjH7kgBzHz1sy2rjFf5eU5QgI
Ps2f7KKT+CRfTFoljDW6tWFtzqxS8ptW2qsPZzeXCY4KZdzMiikep2rj9vI7bIzV
hxytEtwfqmKIeuYPJrkO2mM5y8qC/b4iyBZPEI+w5IX4tAaNob4PLGawM16yXc0r
IGWv7g6PaJiKRDGgRq0X1JCCTAvdVPsAJj0y5l2C1qddU1/H7Y4UgUYygeIJZlP/
KmcTjjgvOJIrL4L25GyrsTKy9T1KVxPxGy+BZ9ffEmqkerwgNGxZXXmSEj9m4aTH
1x1rv9QJajY68IrWv3I52GieNIEYAWM1rB/WFhv5A5ycnyusX5mjDaiTYVRorklN
e6pYjElACmNd/M1nQwZOaNJwHMcoCBy+yMHfTqhuspZo4Nw3cOIa8gZXRyfzaHxu
ZmToTMmrDph3ebABOsJIMRuWpxEZ+ZOATi0lKw2C1EVS1E1MzesJXzVywF9/8Ylu
x/oJE3xJCjKzn8HZLD/Sl+OzCRD2OKFLz13wHu0MPeGrMc91HhmnaTX7Oa4E7hLj
QwULxl/4q861Dro8geu+Uby2bRsfJUAVPWUadfYOVvRZX4PsKoCXLJH9sJgij0h5
MR4dZQwKYKa0XtTMa5LZ+urn2sA/ch6aK7URSGm9DaEoea7+A0C9MHVdnoeCpcV/
r9MUbMwsHPjYFLjRfLdkMg3YK5vZmUB7iB6HV4oWwDfQbiEu2MRfRDVK6E0u4fZe
h5o6k206kuIb/lo6wYNL0FyQ3PugzCzjC8QRQ8M4TlBIUMM9Xc5w2IbbtK2Du7KU
Su4xvymisgDdDa8saRz0MWh02PaPwOTmVLloiT8IZ6sZOXwjTolA4asswGmwY9Oy
tFM5Pcg3woNTz6C1Rc4Z03H9s04a3G+umiW44EfopbgFXb5DJp3mE7ZvoMtjWNEA
O663330MoZ95R+GK12i1AQT0DIi3jun66j6K9eCmeGEmy0Sz/0AR+k5taiw1XQoP
B227HFhtMbjrQDpb15yyqKFipFu5glFuZMquXyyHYXYFaCTbrMCyuuwdR/F9iqT7
98IHd2GGqWEyoW2LlgdQeltp37tbA/tYNmPh4JHvO7J1G+xyEWoy2rZd19YP6dcx
4ZaIQa7iYA4ZykqEU9+t5A==
`pragma protect end_protected
