`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FHarHXIwYXquLgjitvvBFhSG4ptOtxcI7ddRwu2Z/RgEUG+L5v8u7XiWVJhN5BTP
lyajoVVpxOo9gvq4GD1T05oep8lL8pzKx38pp7pShB5bAgdyjcAMEZOnqYEVhg4Z
gJstOpe2Iy2DTMKSOuBgQ1Jldsj7UynoWijmsbwsXuY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13568)
d9I8OZanJOdSIpGhZ5A5KfJzhihnV5TQOcVeiqo/cnmKVqdm62eZAneBEIvF51Hs
dWVYHFnVRCAO8ltn3Wgk3P6yDMi7qOyqIziZrbeFQMoyrW+06nTeL3wqIE0iXKPm
oph/eFXfPmXJ1L0dfgdRPJpaSBiMuz6GLQXQhs0r2oKJxdNp9sjkP/vMFEhq3hQR
8xRCugymDjx7rZ4aSX58/wbVEnYGki3TvZgt26Q1Oab1jid+5y1ko+Gnd4+4P4ns
Owqu5YTZ1YmYgQbK8TxpD5nhV5KJUxHYVQm+vO7NZrnmsCLnyjidMCVg8JAXwWbi
QRSTJ8TcV0RF39EoBUG9TmhAI6reovMdBR0NitIV+XivAS2AbFZM3aoaK9BZ01wF
EL5X2nv1Gdpf7+AibRFZmXFnV8WoPsjY7Ewly3zSuI22FhTiuZ7JqU+48THKhnRv
7kbsc/n0nxad3BfNtHfy1lQiYb76SvMPzl3HjZCZSiKWCvD4LY4xsKMMXjV6vfsW
SgOqAwyYaJliKnT4o0f9/fqD1dizOMF9dLBfqqMjDfCpU8bDipM1EC4BPOCZVoJE
d9h0GwZu77zdO7qekpbVB7eEkeqEkKW+n//8Wtn0dGJEhOe+Ie8nDVl1Gu33ZiEw
K1YEVLulXGgF23B8IbI3lvfF2AwQdtUqyTy0jD7dgVVnGLqlVJ7KkamMrS4c8O/y
PcMB95IaJ+vDfOV7y8+EjdmKb2m3KSsSPSILMVY36LPPGlgSt9EfPRaRbOrPZDy0
myFN/qes1eJ6aIEbCLcqQ4eSwkZuYQRUP1ayQDd1jE9c5tBw2XmcBXUy2PieQs5r
ruVjhVZHq5r9RJAHAJSn4ljmJQ2W30jbttK6OYkRLOW+NcRm2V3mz2fBXqHtklmX
8qArPUhTn8pNXVpYFazc/TP3NchPUKZmPdTYjPiOLS2ryjUNU4XRbf7q+g0yXBtF
80Yyu0rlEtpwbRaHPmYbXDE23vd6k594Dr6BSyu1/hdd18UYUg4DUQ2LYXWjhfC8
+WP7EtOn6IpvZlYAh/ONHJWd6RcWQcxM4048iDn68RtK//akyiMXqrmD0azRoCYn
DYuaqRsacAkEvlBYDdxjLZ4wsWzfruTsNTNbH+64sg2KtG2DxmFMKTHIU2WRerP1
Bmuu97utrt7F3sxwSkFiDOeBc2nJALfBRAPkFFBwK/hiY0ge5w/qehdF9Xp9/koe
mGXzkJBcDYJQPuokZT5IYqLNEz8pana+wGtDCdT8nHseOKV4xdpbjMZfdFXFXGzs
0pHGUTi6RQAMo2qn8Ilkb2ZwYHcienyl2p8ZnrIHFthLavrUMuTyOiPMsRbEfrth
unt+RUz9NmbM/7fiRqIWoxTyCEzT2jZ3es/1MBQnVDJlr9fAygy7d8pHT1GSkVVB
8Gk5DTqf+Fn630SMuX6wWyc8kBEkp+ddLRWy8kq0tfVgpOsR1YdEwUyCvEb19Z0W
C7B7YlgeYb4M1+Hnu/IEaAWxZ+4oVYvx7iiBOaeCpbdzRx9oFKT1d4+ow+6vD0W/
rwfJEmlzyb/DhV3MblgLsksI4SroFk7NEndEkIO60A7wDOkQO1r4Gz3uWxtQ7dEC
LoFqzNrrZR+KSbFWweYEA/DcDFpLQg3tPN7UaTuDk8JjxxXOPdSkOitNUWchQ1iG
+Vj8lxuqpyBEhCfKD8yl2NGmjTUgXf2vCOsCMUmwetsxh9fvN4puIhmZ1iTUUPMk
J2vy/qJXtkRJutmPh6pEcCCxGM+F8Sd6Nxs21PSD+4RYNoPgDOReOX4EZ9QEAlhp
bjPG6PidQwhucH9aoJcWG60kg7+q8dJ/Ci++jKFYfW8Yr8yxRH0Ihat7ZoVqqcxy
DtJGVD1hKq3xkLjWCecfTiTZ+BH8fE7F6A3GgsYmUZH+ssL8a3SV8/ueGPb05iXN
89f3nbzsZEBb9umaN7Rf+Fj7bZlFV0H3N32Nee50GprDdDU9mwDOTBBizr3JJ3ex
ZYAgoAl4+8mEpP7drmiUtw2n++/Ijmqi/ZOvmGf9U7tdXfkKeQM8yDEZU29W4UN0
qJpS0ZYARnl6zDBmFpMI0HqJPYdRJYMDAoz6jGXjwnaj5YrEGhCjfSOokV0wHYHI
a11OYS9SASXM/GwHJnX2k96Fh/R9+GUwiHjz5XsJnz7jpw+kkLu5meyn0WZjSe/W
cH5/p6jocRqA72YhqHXM32BRWptuDEmJHaQtPSp/dmmyBfIsalBThsCf6gyXtXhA
NRkKv/oXImVF0sqbyNTNBE9PqW1UoKFy2YrqYbiaCjZX0kA64tWT1eqGc+Ao9Fw5
0iT0MZqfDmwLzKV7+6x/puEb+ghtwk+CIzLzRKHpWH6hpPgjU+l8vouxaCr5SH0i
tBuGLS/tM4Z+WIZcdTQYu0u1SwsRfTOhFxWKMbIWQeJVhU//q4qqQBHZEm2h230n
ZwOM4pFyUkmpPobOOPDPS55DSWMhqxPo28kij+9GAfppi9Hz6/MhG6tm2w/NU38H
IIOdV2IvhrJ+1tKBzaBRQYtUpXLNAnM4viCoOM2AZogHuPEULoOD79pbQYORJs1C
xd5373FarTqcczanVRBQ7reOprvX1Cer1jLhwyqUtKLKsRJYn6d197OYa/9m3Csp
g2Oh3hooflV/UFlUnIJsrL+k138yY3MG5RnCx/xHvkxpXY0FUH6Kil6qnx1st/ny
lUvC/+SWuv+TKTdTIv/ek4D/zmvBAnBFlYFHxMr2MbfJG4+grs6oakoVtqLawP+4
zirysphjv7gytuwFA7KRq+nuf4aHZYYgGUgB224qcQjifGoXxDkVsh7m6OIq+zAb
ycHU+3nIN4T8Loezd+K6KCzSaU9jJ8V/JOL/o2UMSNHw+wiFUG1QspX5P0Op2RIp
2c2cegQmfkvj6WNSQIiU3WVyBL3vhaiXa2sYJ+f7ErMOdXOR1QFLUJYmLnEPLbT4
RAv5hh6wen4fyTAhFQukHB79DrWOc5tzUjUyVn66gk/sioUqGnVPHL7n1Ug/u4yp
+7O8eqSAly0jGspPhP5cbwk6eX5awe247Ob3Q1DvDJxrHGTp+M9pYy4OnQXfWFG4
rPzixcr2ksXBOAu5ZN11RtMFE05nK68Ih+mphjjveATKJa0Fe0f1LJ8iOrogb/Us
dCdeL7krp9JvY47ITyDI11m3SYKh3XGD+RXaR/7O9lGJRgpl2Ot1AqHvREO44eMa
vazi7FhbAY3tL0OadZ8tNiMzb4/FQxHUPInk9W0iK4cAH/a0OCg3rU8V6/824C+o
Kr82i229PdJmd0MxK0qUf0uDOla/FoBjBI6JDNwnVzA0d+ltBKaVEl2U0zulCFG0
YKodaxnRf9MCUfHfevPuISNEA8hCZ+hF9IU70i0AX3vwLH7pNepTmexobpBV1m0W
zIiJu3OUkQJWjBzlNGfrEnNwuA3lL/Rg3NJr0ZJEq/nj3zShrISzoKtKw7ve4rMT
1dd5CylxudOQQybrsYLI7kz4lDyjuh0CCn+wrIqGWOsXCYK7Cpyb1Onu+ep2PPzm
mzAZa/7VQY3tUe6MGoW6R6bI90DbVak3q0KouthrvlLy7sQb+0o7bJYrHXHgGnX1
ZpoUQDj3EBfHi0MAcxwZx7Y4a34VYDaPVHExx7xcirsNM3BgaEnhjZJsh3ZYageO
5G3I9e/ka00d3kVgKAUIZjB/+Tn3kF6xq6LQeqv/oT3/vAFI5VblRSs6JHEmazUf
FvmVtxh1RiMWv/c7pbBjvmTZ4WQ/ED9AYguLXntdEdXl1KdcQg3Jf+MrsX4H2DsJ
8dR3BGfk/eMz6VGjyfur5MMs0li5bi9KOCdDm1ZbSMOXBvW01y0N8/P/omOHobyE
ScAXvt3NzkfHksOxQoTyJioKX3vwZ0CtOO4jBSiXDUOP0fk0gZr7FSIDi6MHsmKT
IPXDjVG1wuNU0B7B3gQ+kj90ZT94AyEv6+OdeWKJpdkG//vjNRmGI+SAdo6r3IPU
JBvpYCHTjuCxYNReOmcFtU3cgnpZO4SUvKAMXV0iFxdtniTHgFYkzyLqsV+DQiSc
TsRpLqJVziceRMnKm3SpKdMAqIC1Edz6Zo4LB/KqHQYOIRCB3oD8mlh33BodqIbW
HYiTnWmTnRf/hgzMT4FUUvuVkAsNtNj5W7X66gDSOVD663d+1uYVi8LNEh/qqgbm
Pn7GZ4jJ0tPSvTQ9i/ddqwVW6bD8YC2pRCcNQs9HBFRpff8zsEZspoZcUtQ9/Ja5
YFfiQQP/1DXtM1tu0OfnZi+DxQdd5BsaOHjVzlalH9u+zoKxMsM8/OMPBCaZX+W3
ShyXiYCdiflG9DkJd8m3TcDgohOC95BKO62xeArKgAkEvukd9H7zBwIq8WJmJR+d
1sN8aeXPIiiDVb8dSdYT4SxqT0tHOmsr2+Va4SlOBguXd+PGWrCheNVBaSD0suzm
91F+uB3qRQDsbpqYF/9OTfiG2KKEr/EiuYDzdpCyfvswPe9dQCTniLKURY3OoOed
9wLn+83FSEMusRk4Jpz1dbc4zkOcLoG75MSJ3+9OUuKEXNVS/QICR4q9r5T5eerq
PEKFrZ7NtAHJ0jdFKaRFriVQ8++KOAz0FYfHQyxQrwgxdLB/vqkDvj3ByIKduQ4f
mDRUSpAWZIWC299oRPHgyb+TBHjhG8Q07TurjN33cBGamojDIOsbzWLZLiqsOOla
skNLNHofekZsr3L6/rFvClMDsiahJyJIDkm/tPNQUcthfgCvHG19vmHd0CEY5mqL
5MK8e8VbBwOcaTM51mMlGeC6AY4J0yBe6LpKDIj3OAA7sUPMb6mzF6982g93ReaT
VPXIv1e7LQyNuXQxzNhFnwPGDF6trIAiA1+n+aH80uyL/HIDhRzaJ9+Bc/UNeZza
0DJv2R/QBlWvxXj/IywHrzPSCijayKaDNbVYF/EkgrQKB3R9qyMRukCgQftmIyLR
ZkZwDb+6SHSZQZg8iBYFBhGA8BXmrTefcJbwVrUgcDZZavn9wfCv/swr9WaRnkXT
zDg2Dy6ZHILjFzewhDmFPvybm8V0Cjwd6vo+8C7PSj15LP6IMGwmpbsOi0kyfXNm
bscf7TO6NW0w2NieGxeDvnNTIGVho49g8XDDnXuazwzKVcZiZeNGKJT2UQCnRjPl
9VhWMeV6RUIDSltp1vttbUsZ5gv5gSQJeWMMuePDp5NrQ7AMuA+HCmn754L4wRWg
A0CdleqHAjEymLQ7XQ5naHLBevM4JxWKSFB35RHflWggCfkR2qW37dv+GPUkh+kJ
GJkfVZz6IC3+aR6L635q0lLbsHPzYGA5Wa3eg+6c1+/8tEa9zn73wpKqw7qwI67+
e6/3cbTamoEaR9uJu1tNUR0tgXaUSHqH2oPqWkuAzzv/wbqwcx7ZrI6Vj56U+4ae
4n6hFV76VIsLOFWPGxSXWZaY1scbLp4LoaN3igK2jOmlIfPXU3JszbbqLN+otNbe
UWJ0O6+YLtXFB5woIkn0ppqug0Rb391M9lfDOeLguCDSDjitZ5YWS4L7hZowAGeq
YigyzruXGEHuTUuSIxtO0EmXVKigm2pCq37iCaRJDtKjJ71LJmlH6Ln6CGrnIeJ3
C/a2AWRrtYy8oe0vQ9zjdIeGtnc1tH89R6RaMycwYsNJjosYKSfqqoS8bqKhr2sP
q0Vf7wORaWitmto/fzq+kgPgOSM5sE17EItBsLgmGvsreYAooYvAGGgVe9eE8/Q1
jOEXqtX1Gy5zeFRmFpyKH9r5Z5TktdmxC+yO0ASGd8dv4QEunWOkmUwvnBitCdEI
JX+AkN+z0hy2g1GRlRwQAyfIhUGjx1K+S6M6SZRs1b95cSSFfebE3jrDaMz32NGB
6uqLzT9oKYK0AkiYRZ2pq+TuG6MFJeskmaJo3OXli90eihob/VRDb2ge7cYFfRHV
Lx8bmtwGLIbALmi/Ejh1yf/mrc4jMIIXsnTZX1imw5W/WUk9ip7ww//tEYb/KJv+
ThFo/UdeJdRJ/72YlaojB57uTgSMOLpm2QsO8vOpenwe9SOd9HxbRE0fSu5m/FU9
oxC3Ka/2HhbLS3jDOxBvC76eab8NyqhamXWTD2qWozErNuvXLKsUVN+IJkSHqsMR
lpbIuz3BlNRvldIJq0uakh4Nc+OOkgoAPdmWDgxIuJiQwLJuTcW2D9RWDpJPaGPx
QqQZazVnpdvH2yon24OMhaDQVRQs9j6SC+715EtdZw+u2LDFaFyPnANZy7iKWbIU
hqOHdEatpAUwIoUHyXwmuupW3sdOJXv3otir4T1HmjFCfOLoftfLJ6iKIQcEcC4u
pwKkuDHRnwPGSeNyy1zSBuMBG3VM3YEaHbesSoshOJsR0ULbJ2ctNLvVppzcABWp
OTnlCD3fgkqXCZQC6RFzYzecmSPwVfYp+wM+53Rp5Oq8Tyry6z172J+ybLTd4Zq8
Q19kYThlGHoKscei+a31smtyV2HY1cG0zSNA0ts4ErTQRa6vq1EmMAuROSuC8Rjr
lxBiGSRgHfSjCrWJ/O8tajYTYaIBJhqJsJZnzSysOLnFBLCgLwxd0TvcoFkZqFda
a5LVFmDxIKwMXZJsK+gVo2H74BxoVTiBTZ3Jw6CsfIvyncP7gzm2yb28FtDwkxuC
IibP3eph/sUl9//v4BVxBfBFWbjcjw/wZcpHWvaj+v8KOadDaWLpw8u/p6/ZA8WK
7THIeXUe6FWwal32YsbQ7+2eyPd06BQb9oqR6cC4xcHTgldLxCpkDtxfahWu465S
8XzBt5ySTiMmUjLTd5Kaau7eKDGPvntpZFPyAg5zlbif7m2nv1WgMK2oz5QmYnOr
yxFkz21IX8oV42N6MJI+o32J4395q1tHZtfvVKGgAM0OcD4NQV7TKagD38Tecank
emugMzjxSlTWBWXAYiOiQs/srmDlZUZNWkF+/f/hQJvJy3ygb3bWq9PILf1rS5+s
kI8YNA52mmd8AUplfUL36FhQHzrOyXdiXZGhOmCRgvAy4gQR1XQNodG6RWJ/BdXO
X+ifczYfFSk4AcDxroslYoGkGSRy0r2ZFt8FAqao2ixhLbnz9hMlk5nrUlsRdbFq
F4uIYQq+l+uA/52TMT0w4aAP8qHGvsXfiVxeQTgZvzIhCubhXd6YS5tawnRT7+0y
g9Y4vWrIpa71mgYrW4ICLrk9JVzhieirmM1shMK2hZV/15wA3kz6OejKkb4E5Z94
WXh2qO4MaGRSGFTzqFCj2DBa5bWTCDfB44w9U8le2rSLxv/OdNJtlnoaDvRbP8wa
ePxOhPhrpp/KBkwz2VWAObHFcfsmOrUAS0UzRHlBRkfkra8CU7a7768131nzGSud
1GOUPRymljwVCOV/biNG1tOxB0vv2bfjQ41iHCejXzo8x+Pukw1yrchvLdQuEc5N
OBSUddKUVCSnnUvprogcKFm2NSnXomJN+DvvG1NmV6A4cCb7LmXJeceiATAenRUa
owFk/RFnfeYTJyTn4mr1AuXev+1jL/IQczenTa1bxDEwSbdVzkKWKPIyeyu3JUMx
ROlAxFBHiaeAE6OFnk1F0Q6bDkhRiD3SXflUlF1fXTeAxXDQ02evTJfUoPWeDWgv
O1uleXb1d6/K9HnRsMl88RR62ruyUJ7qCXUBerQ2ulB7PuO8WLvGfDxz0GfcqOPc
r0eu7gkfBx+UZp4huANHd3PuFI2GMqDLWRPmEZWAE/CTw/IXNG8GR0CVpyYc4cNU
ZFqQBs9UJge4DH8BelAdpw6ER5y079aIogq2yvcdLgtMq9RpqRcDGZWS/RY8evyO
rD97S90cLEQ45MqCyHOvojMc+sZpilF19NbaZTUM0GBo+KVRrM3GlOVpF5jZC/1r
7scrhwvHF4UVRBnAq4EqrVX9mEpoNRKQ2a2m4rhuW/v4N1ulumnULgdjgMkKwBlS
NFSrA0JUhv+WdGF1G86qj5rcT975Yg5TPmQ9EOH5izIj+VoC244RiCbBt/e33TAo
AcbnAKDL7YeYVkcLcb74cJgYtIPKt5dHHxsZVT2UFPfjClYzR7hvTQkuosmTFxS6
qE6Ab8I+JseyEITvbmstUEMPFsayAVVF8qmLdgDp9/ydu/PYUmQe/+9xvtYf0/5w
Kc0KdrFEsU9iP5+Q8nL0dGiCrf6W4jJfxUmqc1OGRMHD32bEQziS7Iy65ZFua1on
ATcFGTpb6uZM7NuxE1Cohj5mZQxXOB5j9u6sMIzhIorVaUVPSY/hrIPC8kwxwXW/
nV9Hv+S3x8KO4HQ1+Qy0YUqlRsDvGxyrJfN6FjIRO5hpjQJ0s8ZtXX7ydiahYQm5
3kyZeVys7D26EY22Uc+bByFRurggeNCyjGxRpskMZkVr3Q3xmuv1840Zz5rQJJUv
IEHrWfE9DklLYYmnNbv30Qy1+0fZ1OR5jjiEQTGu3COwxNrDRdGl0dvtn8Z5VWKs
YWsCMbirt4wJO0uxgDPdLIn//J2pGJiAsslwslH1r7KOQvWSJ7XMcq1Ur1m2N/2O
lq7swLfA4pjkV2lfSphi0YjWShHoY/VKhsg62jbB9MPLJLju2FRryz+5IpOBqohx
B95JC12HrmAjqi/89C9kBGTaTDF13S/QrBQQJXXfO16qlbQdtLvVnZcqBjzeaRcS
uPIk6HmUc1Iu/7fmQM0QTZ3JfpuA9jwOFchEvBfqJ9YWqmKs1fgUqC4Ls/bS2hng
QO50S+KaqgHwsSkglRTNXcFsn6WDT6NYL23L7rGtGUXPkx4ojV6ZOkxLoSRSR6Sf
d1oBjqYxpEbYz2GbsMdVaRTL8DNwjXUWl/2w4Mfc0XH+sL1EDZqlCLhkeAKHxQdN
mZrOQT+AYNpMn+f0vKbDp7tAbDjl+JbH3QhMeRWFRyYvBHC4WHssIYfV7wtzZbKf
tbpAB2hXGwWcbVCLJS18o9sRwOPPPI4ejwxJGtbCrGQZSjmOD6lkSLbY6pALFiJF
+2dnJofmohPz0DMqA9KpcflbmOW3Pw4hhS1ojc52tnPkpu1cOR+n5KX1iFamX/iN
ZImEXoLy9UzhZWUu/DDxfjqSWpkjmbS5eDdWKy5FYMwcT3TLjR+px9UTco3l3jeP
DI60sZtsh+YeP6eszIYZpJptZF2wbH2WXVm5OOqO4UhoIffrb4xDAXjVguBnM1xf
xgzBiEIcq5CnRPkpynlVrvZT6E8/BS4nj7GwQY4KlcfiKTfe08PAG5cjeFBurfuD
74qRnExU1yE4uoGComm5L3xRfChZ/coP+ZT+ls9LBEPwEvH+CfvMo6dELy7F3nKX
vMKL1V2M7w3KIjT4jDr33Dz9nGUcdK/qTBwpYZQ9DYsxOTV6psusSOR3ALRUOVic
FGCVRHXvC7mbyLcCToTCBYDbVAro2P3xdxAcC8Ln8jxd32CvOqXM5p7HMOcsx/+i
pKCTXDML0Eq5Xjb+90Nq7VEb6Ag7kXnWmSLz9AAltD2Gg9Ij2PoqYFJyg2/mrqPV
9kucjlX3nwKFujnuqZE8BkUGWZzvmnvPB8Pv1nnwW8YuPJZDFUkx2JNZH7dpFBVY
cbpqf6yfjBxP4mJk8ssppMgWYL+Q5JWKBxQlwHgFgMJNOo35FTh80HkOXGFqBp56
j6p4f9Ywx/gW9E0rIoSpmlLiJcB9kcUaYudn/a+A//oLnibctCgY+0DiOaLQzYKC
vv3yKvSg9GVatajFQEr+KpLCHuVfuMo1Kh8w9Zx3oQSv+w9jAOLxhjwlHU0P9lfp
tLntX6CScea0G2V+OT0RIsmFtzRXql6OmkNRwrCZWVDBUZUQkzD8pDOHrsDGL0hE
4OdrXhfmZS/PD3WRLSRB0vle7nb9oQmlN2xfMIEve+CBpzaD4rEwhwa3oKPqNZeG
+Kwo5Pahzcsm2y8e9yjYYEEGcqWG/zOYt1Smdmyfncvxz/fh6WEiqoqq/FgWgR2Y
+ctRI52r1wW3TN7cSccT5WMEGGGZ8C98itaCbPzLqwa2+fZ0tzOn8bmZrXKFDWP1
0+NBd0YrbuTPerJ6bsJTbM7MyjjjEaWvNqOvutsIy+k0IW8esZWVLY0VQLHjxJ6H
U9FaRftq7bwXlpeUmZWZaeXWB/d7UEn0Eg11BEEHbT+ZhuJvZZjMtf26sQQtZhg9
sqFvpKG6gCsti6IMkzc65qif0aKPM5Kfe/82nBymxgjPebkPdX54qjQXVfi71H/X
vQH1e6x8GrJET0U3pVovg7klj/5PsI2CwHZCiMg/W1AzRT0fmlZlzNVghdmNu8rD
4c7iqmlIBxMIXE3E4rSkH4SJSVmUNoO1rPjsWwKUXXp5pcBH9B8keqZ4awUCxYLK
gff2LXm0wUMz2cC9lKlVCNfp+6lRmo09hJLweVNBxEP0ambgfD2hRYl6cHq4KSdx
aMbFYbvD49U8lK1p7F3IdE/Adl/cwMmeqpphs8NyiSOobRf6T9kcw9/EVsuWLN6a
jvgu4hgZFmMN7Mp8GrJaWjFngIayLJB1bKZ0H6UeMvgQp5/xVjsruAkGt15as31H
BKnaDV3FyaGd/tO1GT2v94EP9waZiG9Sz8AEWLryfxXBQ+0S4Iq+EqlaoL99I8LJ
RT3aMMjRj7MaTqj77kI1wecrCCfV8Hi6mBSwDKM4uOn5Ugp1m2DnAvTmeGGrURxN
1C0lsCPP1niaBL8Hpgb5V9DFhvEBxwq3qCD0kyybjyzAcjte+MqQnNH6Hz+NeEF1
qPUeaIwXOUzJMtTmgJNigbF6Vj0mAOiZHqlfvPMu4g3Vd6W479sYe5QH+tWfP6aW
Osp5Om3jbYSe7kkKw3Z16AzrdDdHb8PMvWbYqe3xWmyDGrFhLz/sx/XOtbHv5W4L
9WGl08kaImTRWOOpJYFnLXNi+kVy/+GP99QS/XabHD69gfE4iaH6JjTVilf5SEBK
SfuKEV9W9fTAw9Tvv0j5UZHbAY/Pzy8FGe2K3+XgLhuITp50S1vhhoyvtZY8YwJ0
sFZJiIKsJpRiwBxKGKmKasgvBY2xCagRgOMC8OM11qOyrgytrC/JI7LFaG27SH3d
8sS8Ss8cioK4dzQkhgxn5pU8Qy1PRDVtoNFo5rXEpEn+NjWSoNPjojcQimLr1AfD
rsqgARNGSDXV5QfnJqJB8xyDpvx/2aYbEWMIJ02Iij5U6GFqyuGDHwgibwtLX063
r66TNgLNJRkDVtA/3y5SQ64LAzt30R4Z/ks3iHOnf2/XnNAKFeH3vTXWbHeo80P2
yb8ynnDDubkAqBB/Hi09H737h+poormAn66ZMTNyHIDJWim/FmKBMBDJylI3bgV+
ycCiPYPZf9xQXUeZ3YirSWPA9Z+OLY29jMgx2jDt1QVjzMNK3I6lAKXBa+udvZIk
snZN8sFiYBCMpZ+c0ttIepCP516BPZSnfpXzv8N9kqTJEGLJ9p45SEG44J8Gmi87
6huKJyNX768wOo3790Krk4A7bEObxunXHruLE+iTvkYNIFsKSSIeaqsdT78+s7GQ
tF+sUTGdgyTRmFPDmAlG1DkKfsGSeW0202rsxuaVPHw82bAtM4+JLAdisjokl21v
NwYdd5F+tH3rG72loAdD0f+JN2JrnhRdndiwfWJMxXyU7eNSMHMYQCIDXlisRCHp
SfK8ia7liAvrHnWl+qhMIONER6+UggQ4Ty40u5atjOhEDOnxo2kF9VA2v0pqrhhd
1QxBYmEXttI7y9Jh+z6l5v7D7GoT76VTVBLwTnxqApDuBAU0rAZtKGkXn+i5yfjQ
ieNGJIWNvTt3575T5UgEhBsioeu451IDNu/47u8SbTgZ57WpfLxZ0jtVgyvHCcfR
arvOGg+lhRcEIEa/E61qq18SDwBvedwVCZ7au3X9bNXhiZttF0d/gHABo85HxAmq
3s/Gf2wU+puZF4AvCAoj0cxTbx3WfQmMnHjio0ctb46x9rJmO82kEchs1mWhzqlt
jwCSbq4vAxlkeaJHEgnk7bHVjAz3CXNJtGzXxee1COjm43wiDKTHDiBHOplDwGWZ
kSbKpel9as6URXqE3aKcgdLeON1gqCCr1LeF8VxjbNtCkZKTFdAWDcV/0Jf9Q5je
04mH/xAvy6l7USrDm7myeqPtMkA5xTJX4DVAJ/sHMBq4PEVT/wSL+Nb2nln/k9jy
ASSN+5VSdEZ1AvKlJ+yRMRNPWXfdWt0kz8s6FOqZRJMpis94I/cgfRenv4+NFMvX
TN4qy7eyPCvRj7wCC12r2P7+Mx+SIzXMSb+OxxiaIq8GipxtaZCW4f453KFCXRUt
SI0DiVEGze4td/ROv6Q+6g41OrAbGgN8ztBW5YdCNXIVQ3xl0v69lIvGfkTJJ1y3
qq+K7Ih5WXVBUc/Q+XG60QotPmEA5VgWLvF24W/c4mxVMBCYDnkw6zcfmcEQpKEd
T61576iz/Ed0Uk/F8UkfwJXBUVx5HvoP34dRQH/EybCD7eliBcncdmCjCAemzf5V
j/g8cwCrJpop8FJUbJYo1U5RKHMi001QISIYytbEMl3HlX+j0GkdqVIdcIO1/PQC
wwnB66fv5BMCCDUey07g8IdBe7sQ+jILktOWpmPPSpJKPBoPIzqDHHUbACI2CRBW
VEEFhkKyiAkcM7oIZOYwtCvsfteEGWoFhde71CVdrBUZce141oD7zutwmT1GiWgK
FCQIXb9TRaVYeVqANqkRKYKEXgthhpqCgWPxKYXJ8Q1sVtap62rzIk6XGN/9D7zE
OOa/n9A8PbyHTgDc2ZwY0lf0vAQ08Gc3GF2bdcIlT0eCjsVMwK+QrWmICThFHYcu
8XRHjJnBRWwDOkw1qFKr2vuqShFlHYxd22uWfbQjIAnAKiChBSP8doGvJbhw1HGH
YwjELPvRdcPuibWHTMrBIuouZ5PU0VPiBaCYCY8MhwFQ8Ob5E+eDn1UTTAHUyUVg
So/JbiwHknI3wXFRKcM2QUoZcBJx0ll2aQcpBsY9jpkayK8tMM57soOGGPw0hq2P
9HtOVdL5Mv0wJwm7VdmVwO8W57GMjct+UyY1ggQYj8sfLGmFNlR7rARXwahpI4OA
NSFl0d73dgwh3PN1mVzB7Afvv+gbE0YlgNC/FNubO7pCBFylKNsSNndNm39DNyep
A3ZEDXrHgCvii7nJVcqzm2qsyLN8C02EU+VpSQb3lVIozkA/kTud08eumbhWcsoS
PyIaftT6lQ4X7ndMG8IDBzg5lh/5Ju6qKMI2GGSBjDYJHEsOjG8nXJOxJL1/DbFc
v1l8lRL+SmVcVAwKMbOePN8UWYmkzXaVNHgym2v+bf0h61di7NqHfxZGk1sjmvTU
icSnhVWYtUshIA6nOnkzbqm43KUrAgl4T9DZWP/pkyB8nHn9pbbyT/zhHmMLs3sc
uMJTWR7e95ABgVGuekMu0EbR28ZiO4MYhaPtK/RbbHBkfq+3IiNCSxpp3ckMOcHc
U4vUAgAHGZVZlMGHTR2ftk6w05F8hLUcJ/YJnNhxGuYU6R6Ub7yqfzZoEyf5skD3
a8p0fzzsMV3l+gSFC9WlHQjjbONZwG7JtGEQzmP1tV5nr5LiYuXO6Qwx8NJiwj7e
BEB5uMYnJlzLfH1IKCDZYdZ7xK/puMiFozZwePaAYg/+ndA+ssc0a0F3vgo4pS7v
8WlFtzNatpi0zCbTAx+5zkm9eDCg5TgFE1GWA2HcUhECkKumarqQxINUUY+TqNpp
SbDl0ZmCMUn8FICGEKHjvChlNEDA/ebAobOGZUDgnYZkkj3ubE2AI0YjNm5dy72u
oDMnPTWrykmYFKKdpK6hYHYvcoTswMQzeLY3BM8jkE5GLq9UyR9uoqY35OyRMM9V
3epP4286ThRMXGlJdMKJ79zuG7m6woHKEJ5ZpoFisBD55fNkm9ZfZyNSQnhnDrHZ
I4E122SyN0CZlg/1uN5SWltvSOIwiPjFKYCii3eDqo1n3vkqGIUTW2LfSqTo6X5H
ySwH+7LQyPFc3XksNg8zGkUIGyONfJalfXP7ekg8ZtAhWB/gBLWajNdTgl8g6Bp5
KToyBouLTN5e5yRP5YltHLNhcO8YB2ATfH8rKlta+M4GzNoH+7PwzC89crMBpTc5
raHG+kuXhdwYvo1vrMbE9Py0eK2jzFba55RpxPs6sGJulS0fx9AvV/IeMcF7PRia
Muo3Ej2pkDZNcKhMsK/1dMwQ6BczaxQAK3fGffJyNPxNAs8pihJGHVQtwfmL+G0G
lUa7qxXiJ/ulDU+hkTEhwq3JrpvCv7BmExyBw9gu5ZtMtcPlSVW3eti06k+fCwXk
pEmGtDggR2Fh/xfYG3RKJS2gSEXrDF/3i6k4bcFEeRoIai8s+kehgTreuq3/EhLY
VecD4S9V5AdbpJBBKGFMt4b70luzxJwsrhDFS9KaAF92/5X//suJ85ovWUJV/rio
2cpak0gL47hB0sauA1zQ4Ja+YFeU0rvzkFdXcr9bOWUEWIYgpfAnKmC877u7xxmS
SE+SPSNWS4LuzQnmuouDOTA1mO5POGRPzOjw8c01DjlCkkGjJUx4sxoVkT548Q+0
XrT99lnWHFSWOgyM+0Lfkrqfrr0AymwDMqPESHJ6/FT3+skiFH+B7I1Cid8J86uw
Us6Bu6MhjHckP8vbA6z2USNRmkmorvzFabJ2v6pYDTFCJ9HVsVKG0/QLoY48XrWY
isXHzlvAQ2EXgFVkOGYR3xJWfxdbBoxMpduS1MvZMZho0bwgc4kpWcq8yEMQYZhD
Q//twQT4Km984geJVbbGVCqA8WplBCq8h60J9ofaGZQii+qFDKL4pe4UkOiZPh9l
vPZ7IrnmhgwLjg28Yq+GyDdWJ3YDMFgFdozJdfT/0U0BhQKkKPgAWFbHueULQwbn
SpylLMoOD4Esb3oyMJS5TaZc5R1YPLQlRb/YSZsq9Y0dKANUYtwyjCFm7oLg6aZK
8oskB6ZZyg5aSiMkPQLnGj6w9I4VMbHoH38KD6ahxblLBncxw6ZXZVtC681ncXNC
OmYjtbNQCkAeMFH61x4knkZMoVHPdjU82VRhOpbxaOD3Cm9w6RvVrB/8fH48bQp9
T2OekqJ+U+6MfyCu6QHrWKwqZNbepGkHaqd5fj6GUhIFn3BURlIrmuM6UztAzK2W
Hnphl0vrALzfSl0PXau4/GQh6UngOlXw+Lu0nceSCsdfSyhwCeoTc+nJ5g3M5/iO
lowcGl52yxfXpx8TdfdSZ5y3Zux46bIIy4sG/eccOy7AeHxmLaCXSfBpXQEkbSy5
muGvwG75ZKkSV/Re9FYVZGcXoMIFQixaNccRajNhSmNljr537Fj8LK99jdbN3Dc8
kk9nOwhAaTH8VwyrbLLZrdPICjq9VegaP7i6r/xO234WXjGDo4AuLuBPorBFtaPr
o80Q1zxIgrXZUpJIdaHh7SUCloBaFGDtRCgY90oH+RQ+Tq4syDqO+8Rv8YQ/iL2T
sD+PVYHQDOaaBcEuXwUd4wwWdizKnKQHJIehRag6eByS2j8nQiOFRte2Emr4h+MF
sZrjPYXWGZHUFPRA4jSV59TaAWE0Oo4pgn4FRIB4HS+JPLJKFMeEbk2xJ0Rd6dnt
m215LqizGmT2GTpITLAIKBZjEONrtp+ePJVonJkzdblPJmyO9s09K2Ei9hppqBNe
YtORP+2iBojMR5MjbgVaO3mukOwD2Axp5pwqGpHMV5xCSzP2XdAQvb8ZmYAgDiUg
/W/DRDPmtzypL/RF9egdAmKJpNByoKZjOsp2i/xY8AQVVnnG/HDzvjII484VNaye
sANq2fhA3Mic8NpN+lF0aRpYIWhWur6B/i58LdJ4gWAvRRfYcASxqe8Z1cvCy+wA
D3hVI7EnHDjJx9M4DL/qJ/1Fz940oyLMw8Fj6Fbv4u505oXfb97hNCvMoDddCa/Z
A3gFNmHAOAe4chIL4SozsVDRrcQXbLH5AlnR4ytZgmUTU74wUi5H6uhgzNIRVGq/
43anLXhEXlBPBaLsqd3wBmpt7FphuwntHQF7oiubulDQjl6a7miBF4Lq7tHmRkMl
RAQ2u8yO4ta5NBlcXQ2Ahn6HSdhr03ffLS0Salp60ARh5p8K38lsT9kc2I1we/WA
rTb1NjBNB2auZleE9NmCoPZdvMZsCA0MOIG7fwIIyiYGBM6B+WE9blWIeGR5WyAi
as5e4TLBypCbICfnWQGEw0M40iYQIhpSKOWZZNwLIuvtTaQrGD6vJTYEjv98JtoQ
zef4zGn3Rsv+3L63ekk+u+SceKxicZCqongUgqzRX1T1MAw3IPpOKdkNmEJPl9UP
eNjtsUW7cGyM7RHJETxzqltRCU8sTXWUlL9li0fznX1SMo3vRLqP+h1jgGWT8HwZ
uPP/KYH0OOXC66GEdvIsvR5Tl30drb7irnpITcEkJGtBde9SmWJOm9zQgmTWeXOm
aNmJd2GbxlBuu7fluD9AxmkmtkVYn9j4Gf7gRw+sw7zO7S2v4DOXgfXdEyUC23fk
fYaR2bE/39q/OimPpwn46bgXFcQVtgXj3AuTgfYrYUQRVSp9AEGMP5qDuohAt1aH
hvj5TmxCW4aD9nemaNbdllz+b/acgMJnCB3BhwNAyxTSEE6oKBYg4QGp2UK+CObQ
MCz5qRCK+0mhY1gEVKbTuaxSClzFGcH/1OaIht3emzUyKYyRjGmcUFOwPwSxtQTd
U0hsr8JVYq52MaP+eXCNeb3HgsD5+W/+04uuFuXTNOHJsBxlu5JNho/E6RUcSo5B
D4OOdRrtWCr4a5Gt2zh87AxyVKO+Hre6zE7UAso4UWAOeUnW400yZz9LKkekKl0M
+n5iM4uexz6JKFzEWY8mTm5MZYSqOFfgALTtlnic6GR7N3xxRHhHtlUIUC3DSJ0O
2WWy3J3g6NvPjzMmdP1mQ+aEt84iVJY/MtiAB/J6n9WsNcTzgwdGfNvAqv+FwF5M
tz64cSaQuvlN0O7qRAYHMNAQL+7kTbthACCjdMmeN6kfVu34Ryuud0EyZxfJrbCQ
V8X/SMHzlJjTTiEMOycVmz9YVwNd9E3pcNTNu6a+pmxrpY1pSyL60zLe4jl5h3pH
CBRRCjP+vL5N3jvl0aY9DghA7CaLSTDrRjkgNVocmfd44BvR2bB2RQi+UIikpnAY
eJGBFgwHFC2RSFMSt72bSCucUYjuPhAf7NAJyumQt0ed9XL1qZN4uaPk9iZG4CzA
+ALrtaRhIlljxA62snrexlcba4PhtxyPTUdq5YK/7WXTmuIQMIbQMUQmL5l/hgfq
RJ9B4Y1CILdsBUpoJoy5eMo9w4nJdl20ntHhn/2f3kne0q6qGE8dkg9g+DfoOTWI
gCn3rmctfS0mW79IqFXn04rVhg1vE2ZpXHic/nQsCVA031Q3Yt3OeKkPoKpuaVZ6
6LaxLvHTsDFq83vfTS7B6LFxqPmj+rcMn2i+06fn/Ohrl1mXvqkuEhUu58NrG2ku
vp2vehuusj2WS0aVlw0kVYpmRejOTaG++/0pH1FivIjZn4XInvwBVn3JIzmv9Hlj
aqwKVQXZt1895RUsBph9QIQwqi1FleAudos8fRhrP7aBblIsEyBzCuv+O8EDcB2G
m8CSJcrp2sQMp+YjXCIW3mKbtfcrDO7IvDVw89YMTT/Ss6N9LYaO6QrsZLUXWKXt
q/91romiUY7J+b5x41N3RAi3k1znbw+ogVVSWrHweT3zzJpB9/92bSCuKxI6ArjA
SSa2N8g6Vb/ILOEMNh+AVFC1AdQ/ALufLEuYML4mFMycGn2AchCRUG8ppk554hsz
7LtExbMM8TbUTs0Usysyt+jRYtu7Vb3hIke4u3hbGJDHZKn2iqImwp+Hu3mVowi6
sUWCdPXofegTdQogcOGA7jMKprhNR9um9lYM5lZ+jZbAjcmUatc8Skf3PqDz6T9S
MR2FvVy3eJD73xva6nWg5kIWQqAK8tEEot92Q30Tkl62m12xGdLjsn0HSQItvMle
ufho9EOGyfFkG6NkAqg2rabmU9RC3aBAgY2RziJwxLaOyaPNjaWldub2w1dMxkci
zKBh+8hf/LgnlVJj8k3aRftCpCrYwPSpGMt0D9SiwGFOT6JLV/w4J/AhlDYrNZ+r
azlymGn9ohvkK2Jd2ImkwzloI0QngDUdKCpjda4o87BCrmRNGgqjJ2V1tLZ8/rKE
orF+ls8UpBFeaBRKn8k5jM7f22Z/u4EeF0lGP+mEDHCTXW+4HsQXljfBVmP2FO7E
S7PxQGt6umBNeSe98x7mwtnOKDh2aUsOxkxJjVPYm1c=
`pragma protect end_protected
