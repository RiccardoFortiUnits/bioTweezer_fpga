`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y6m6HBa5hsZzgtA3RGb7ukRysZGgmphq9j37iZS46kmY4dthdKDSWGnWP2J9JCE+
FInC1kLlLOEZo6UTXbjMRcAYLTsHWxzqoN5L5gVcuxSc6p/QinkL8rqDVIS8GK32
4rk9uNQH9V2dz5abbJJJUh51AhNy/T2g+sfzH9d0IsE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4848)
eLZEmanITZdV3GuvGGQpceOgDffhqqHoW0PHVmStri2v1ecsdshrnT3ajtMdoia8
mYwNare3+154WfoB2eBdWhoM2FlFPuPS/H+2l8oj/DExrZ5o8mz55rDE3Qq1m/Ss
YW7mVw2b2Arpp65x/4Ajm/+tvHALZrKM+3sny+7CZUD+izftVQngMQhof8Olnotv
Gjx1qhwvw2W1mEu4GdXyzBeeMpCQESbvDCHHMF3rg7pB0jYGtCT3JcTbbVPml5kY
ntvz9XFDJuPibT3XjKMVeB1OLrXd/EHc2n8FCNhLiO4IQ0i1roQ9n8ZQXDo1szEp
y+21lIkdNKDCpFP2wPRLMivY4UrlKciQk1zz28k1wVyV5MHWep5cFvlbqgR/KQND
LiOz3gM/sqcvnuU7IBiITOaVMc8krjLTqHu+/8JOGf8J/RUn6wJFwEsPOyI1yAll
Ge2i3nZ+5WjOvwEtVSLnie+Uoie0AW5eSvzxq7N5AolDRb2+gUoi7H68zOCpthf+
MGnSUufM/TEFrnq01Jiv9Y9eJk/UV7C3oQ0N5eeoP7NG86RbHNNGfJ/Lt4frEwLM
3k4gPQ0EfvTfP+wikkJFoMbavfmeZo/pUQM+9qP2b2YpsMUxBhGN7snOrdbVe869
SVTBq+ZsBKlIsszitkdDgnYnNvS0z7kH77jt0DdVoSZyD+oL58z/jswJwQnsHzkU
03sNaldnfCzJykfvf17J+gqsSH1+h1Qxti9fOR4xR+W3Y4WQyQsHmJ/ehYNOOcpn
GyTeLDgGl1URgMc8QPqySvKeLq0ra+4+7ddBkKI3Cxxg3KEIU4aEI2FjyyrQo8rj
9/f7YnCF8t18RL0YAyMoczvkZCdOCSv/B1bEmoATbe4eVpHfEys0GcZ303GCL8Jw
ozfq/8jSO70RQJE4Z+YGygsAohtXZ7fusxzZPEIqwf0Xxf84EL1QWrKfOaZpqGC6
IxM1L4FafBAqQxsNNgsaMdnLf7/dcztt7jzV5/TwRVELPJ6eZbXmRWmQyRur8lu3
e+s+ivrgteGQ7WOQqVo44sQzd55FspM1fyr46/rRCy/A9wp9koG4pqq0jE5Jtqqf
hIH7q5l2BvuyDu86exq8Lg7n/RAxNbwIfwzb533TfRDcthW2qx0gXvoc2IGcqELQ
TJbd58UKelE66CrOsIdOecG+nmrTur1WkuxZ5GE5eG3w0cSEVKj128bEs3I5aJcL
BYbxKsT5qmCzqlWtZDup0abQErLRJIQZypbzVtA5/BbKLXnt3lq+QSpwtDCiGe6N
sqevaoZr0SjVgwjMruDMWZ+FJSZYWejQeOfyHWW1XWaE6szvdzMw+/e36pwBlz46
gpNzCu3Lw1WNZ2djzKifbL79nckI2RpDXul3lChX04APtdE5NyoZXHN15MhIwzo/
55u2LJhPIbKnGl3YVP0CFCe82Tsrg1LY+7WgXtIyEESxEpVFeoLtL695UJHgBwu1
bOIKcwDRCDxfPHgW/6tyLV55Wz+919Z2YGc6BMw6G2lZpdNLT/2plkCXWAmrAuNg
yEoncLOxMkarAR0a0u59H9y79qHJ/JKKPLDJUJ9su3RmV4RZc6GwQtESF7T35zZC
MenQn5e1BmE8ylY/l/0eLf/J3yz+hJqWXDbbA3ogkJd6MFhOdQ63VkJ4/M1D6HHl
4FPs6SbzJa3TibBLVrp+GR9rhxR20f5LEbUwyopU+T4cYssQAMqVa/w2A5gzl8BE
ZYEeQIFUiUt3qSou3/PuhUYn8CV19LdLZRKB77tkzJnzBsk2Q2wSW6Ok788blL7J
HA35P5JL67h1dmCp9/3XAnUmovbHi6rdD9Mhw+lSgeeZiIBvdUt8pNTZaoyAv3tv
W0MVDOqDuZaOkokPYsW1AOhGBTusZWrBH6PszG7A/PAN25Nss8j1nU4JJ6IMF0F4
kg9kZNteDJ46jBUmXNBbrQZ11XKX3fkEGqDUUzevfuRg3hZvLmefB5RDUmdcjgiZ
Qv29cHoz6BN9lS8h3byhUwkxJ1N7Fae41m3FR64Y2T8btoGINISgDIkw7CdU1C6M
0fAWzvqjLLzv5M8gSCf45slkLFIKXGE1VDrNWSWCFZKGjdM1BC+xxGSpSGqlngQK
5JtA1w+oG6Pn3BAZwbfLgf7WSH4XtZIjf0umhcLod4U7o57lfHGCH4WNtucelP8U
NmNfy/YI56ipBzgna+e1vVugrgML9X0BXAqh4e/x4mTmMQx111D3eD+u0jTn3Nm8
D6xE78AZAr0FqjXDAPyZ4dMjA776FkiXUSFB/f4VD60wBomd4S0qWwwy50F641Er
Yxya9Varo+I4XyMVtNiMrvs8vk5zS+wzwWboIVzndZo2uzgqHPIkt7Hd7VctFrZs
5yAa0RHpzs//f2ZGs/WAVHDvJVz4hO3qXo3Ujdh0Z9xmlUabLwP4aI3vg7iGp94F
WtUz4+oKGxAV3RfONU15mCzXI1BFbyIaYcoSfEp3lk4H/ju1f15OQc8jjhLWkLw9
6N5bd0NIkxdDXHNQDNCYuyebUfsxZ6s8N7SwZji4z12MlrA/hoS5DDgP9OkfsIBd
NCRX302hJB81JCgjWnM+vJ1r5YMr4mIYA4pgH0tXmFei1CgcSdWY1XU3+U3pcMca
FinRSmXx9wvIpxeyJ5PcKnnBVuBWVolMEzWAIc4uCyZ0iB4e0X9q90RI+gqDHxVk
VqblRUwbOUBtZfNCLEQnOBmNtExRCNUM+MLflEsDVp3mWVMpE4z3RKEGXXhKe+55
A/B+BqOo5dGgiX+1abYp9W9M/KQIu99+6JNpXxVRt9COZmAqVhbiqr7FG/Fu+N4Z
rr+hO97EkeHmTVt5p0RH5w4D53Iu2fsEsomoeHn1j4wlDmI6qLdaCLKT//uTZduk
uxtArAf41vZj6YfbnU/YvWWKJoo5jCohi0yHVOad/GPqNQeQZNc1qvDe/rE20gNq
KgzWqQo54np+tgpFUlZ5iu5U+5m8VN7FL5T8W49gng6N5fKpZmaYhmPcHDBJQ6eT
LfmtjpKdcWwhjXDja4Ln+nTcNTFLFjqN7Xs0pGwfdR7hVaarX8znuyOcYRFP5aC6
GJzC5ViJ7gD+0I+j2LSEOrJJvtUuLWCzQLsAH6/s90ma2matoiAp9XHOBE4HAm3y
PcLc8RAJLdKVxghBwuFBWfcTbDZUrxJuqi0l1EuDVeJ3RyG+352VgMgi7bB8Sp/z
9r2jxZkHEjSg7UYK63qDZYYqHcnI9E5UMdcAlR/TtkfOfRwkxAtE7SOksj1yqfr9
UUyCjWNBOhyUIOIygKxn0QD+OobY2f1celbYo10alwS7aLSH6NsVm6bt9ecy9PeU
BRzgMFLPez/OVVF+X7A+xJw4KbLHkOIDR+5j0m9rTsNJ1V7SBPYE6YF8AqLHN43Z
wdeyO79m/ECv/78m5GOUqFTpW7rWG03hG1MSAzmbdRFFw9jRIhB4Bq7LhQRkILYc
iqDrYPeYYuDPGMoz5Rps7MWLJX6YAT5kbs4odI7swbsK1WFzri52jrj4DRWhdKnP
ASwmiFzhRCgYqSsuoRTv/nmGDDtNfewAbOX3FiNe+e8p3IK7rCujMRKMBITfKRiB
k7XKEr5xy8T4erQNbhbmOn/JoeAbG4dZwXuvAT/h0lZWEFG54VN/gHiv+KHMsgEf
dJtoZy8g5mUqCWzeT5dFDgmLrKQ+TVuhimse/1BzaSaeQwo6DXDzKUA6JUb6pttP
kZlnh5DsXs2g2sJnF/n5iHhS2vRWasGS2u8Ec224pfKB6wicLEDDne7QMPmhjSRd
6rBi3Mc6zucXCXEXT7jThiz3Esc+BM+jwi/91dFI02r1iahCH4N12rzZ7lLGFwlC
2OT+3Z3BMSDNR4ShAYJkI90Bk0u0HfUkWFwy+hiLA/EP/KL8Dz4vZtGYtvdq4eH/
JYK39bSLlg4jnvI7yCOgp4ddeRKLbgyVNoItyYZWqmYkag0gtst+tOqrQg1f47nj
5jL6HrrUFM14rQW55SGRUYzPzqtWn8r9qrUUYTwzqEd8VyOtbElQGdNwFhVQhew1
K2P4/du5MQAIqA5pturP4rank/wwcA3izB+ZsbJrj7A+AeN1l04JpuPnCntcrGSz
+OPJiTXm5Ha2tq9V+F4v4ymHhCSbhrzoDrBga/UraaHTh32GCqlx8jDB4RdE2jUE
H4P0TeDmJ+5RrUxYrdfs4oavumMMO7tHJBXgVJFIWNuLXZfymXflq9RY4IVrsyyR
XstqWAHdkWIjAVUx6efDsxRB2N9wNUPXuj4HPUCPppSMxNNyLgsw9HJHF4ruWCom
KSrjrM1oMKX3dpVnMNQTFEb4aahd5Cci04wz30zWbbsYVfbAke5d/j5AFKcM4xSe
aaoK8p2e3PgTq9pccegHrwEmHhxldeekvcdq9P1uW991S4o9PFfcPOrSPIDtJuvi
41xhQ2Sn/Q0I/Qng+qPiTwult+kkkv1TNTVBOvvnhwLmTcwzni8Co5uHniULfRy9
yISbbif2s94jxBkfCctTOtMY7N640lqEhTK83sEHqVUQksjEnNN2duogzqGzUulX
IFYDyPVQT9REQrv8zNCzCyL3osPfU0QvEqxaJkOqvVK5tXyF8ExmyG6nrw+wKGle
k1Chx0IOkfP90q/ZXAUKHPEYpN1U68gh1RyvgNDvNQdMD7qGJ8D7ThfBmNJR4uK8
rkPZ7Na+0l5HI7Wu6KYrPKX9pwN0szzJCO9FgbgsIp2AIX8QZzM5dg6jl8bwcSgY
T3FXLSVtn23eFeVKSuEODnkX60BzU0rkJ7y00csAjlrGisqccBw0UtQ5w8eUp1jc
psXLM5xppe4Y++/Z0wQ8JhJkyN5fPK+WSqUDXkF3vyi0+uv/IK2aSDlYiPrexfrc
AxfbYNdFrK7hyUeyn1OXVeRs4hv9zTtdfcjIJt9tkwKBmTEun1rubPrm1fjewRYF
BulAM3hFq4FvRXX7OXlOv+vB5OD08au0+60FQEoxIYRR0N+StShkw73QykA6JP1S
9/ysR4aw2A103d7pN8FNdask3TQhZcqzjpvnU6JjtIyDj8bQgNPfSfU8Hscga204
y6XO0dkqBuuOdQSVWN9a/La39H0Y7Rzkrp89WVDtD0PE/LS2hsuwJknkGU826KIJ
SSgaoubVsXKEC6JTkJfbGJHHAf1omK1yPxUSlSL6yLreAwhd79j00btpwb8+9thi
cFrguyO2jBvLYVAFYkCK7UJwJub3DcHomcrWkBnPi2fpRbKjoveXnvw/ryCMHqs9
or+SjDDA+io+QeZtwplP86hHvToBRm//O0edHmbaqsg6GADUX9KlHiP9uaX367OE
u8DpW6oFMzN81v+NIueiAvHf0VSOx3j9GO+L4PjrNBQt5t33A6OBukAn4mmM9n1X
wuwCpeMf03TaFq077pONX8Sgpmv51fzyfWNpICTxuImtao3d/4zBs4WrgLAjQLUX
1relXFt+dkoyv1Q+o8sRkgD1FQCZXX8QOUw3swTz/xl9ummCRgHKbvplcTmWKfQK
AKlfFvDeVfNtA8mWqXffqCs0rzTleZsmmI5QC2tmBLVgzl1SQXWT87l/76G2hWuS
y4JtGEsSmBQrPDAv2JYmtKSft8As28T/0mBI4A46OyI6s1nnMS4scJVWt25kMBdk
5BWaNg9T2N5JGlJvJ+7c5DtJYNtmHHIzJNilXoO6sYTfpoJJWdbt5PstH71pNotb
roBVdu4aiaAvEpt/rBYclnBnIZVyYz3TzvgdlPtEqc5gjvVDGFFwLHAB+HERd/nW
TLAB4/UfXoTgT7hLnHW26UqrFWYH8iDZisv+VRMeWF7HkOsBBSqJz2NSod/MiWwV
bm0T4JpQvBTaB6I0NDphE68p+B+RF5/baLeYGDXgVUEnGRfgq4YqVx/Nni5l5czq
BJ+eJB+brLYZUBsDQ1SaMvFM9THOuuC2Mn5XvAlqPdqCj1LwJqIHa2SvwnddMWLC
3sH8psxI6pQ7GITwiWHosX5K/BcKWTrA07i01/ye+eOGe0uQ+Fb1/sLM21AYbITq
Gl97Cd0CuXYxcOfB+ubBgqDDUsdXDuPIpcE2QQ+OwCcJNxtEh/RJFZA12Quz8OqE
onz5xGpIrYyw+7ys1Islj1RT5dA7iGH+ftKZA1tSeZzUhnmKrmwvw+1XLS18Op7g
57CkiZLsxsnlkK5FYdn81epsGX2vXo87KAU5ELSMyfnVZDQkIIoiBVrORv7/LY2p
Lyj4qhccm2Uw9pM4zdUibCFDEDOJAM9dvQ8Vx6YGn4dN7orO0KD/BWBvLihvgSyu
YLFSH2txmC1yzKE0pJ0q53uoqAAjZXLNauJ7eTszUnmTBKfSKKG6I69ZrdV1YaHt
9m8gjRN14KsY4Zp3T7OUGOHBw0SYfdx9dlIsKrk08Rh5uKZJfhcE237spi3oVBiD
vxN5RjRF+vlaS/NgbI/yLE4XVjU6r+vGXzO43XeVzk9xiSaDVCxL/EX1XPm5UcNk
`pragma protect end_protected
