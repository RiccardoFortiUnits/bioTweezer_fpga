��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��x���9eS� ]�_g�Xh3��1��63�A�1{Վ�eb��9��d8_��g�G�oWs$㩕�䫀�*Q���7е?-�@�Z��.޷�0�Ȭ�*
XL�1���-ec��D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2���f�[�ˊd�i$j�sƮ"*�ne�����Z�e�os���Q$��4�=;7#䒤�T�E�bW���ֶ��eʢz�x��58񜖷>"�1Q��u|t����l�;�V9kʚ�1A�5V�y@q~^# 'W�b���\��)h�7B�Or�"��mq���
��L�2�Juo��]$����EwVp!�, ^3��P�DPh/�6[YYC����L�pO]i��X}3վq�m�y-e%���x�HA~ovo(�Ig����3�*��'~O�w�,Gm��j�3*�F!1�y:�[]i��L� Z
�i]�s٦&��R]C�&*�'�-^���?O�>���]̿���Ң���m0
4m��,���e�D	�"��~9 s�<
�Eڄ��96��+�Q�&*Q�ˣ������Q\��QJ-7u�s?<3��"R�`��[�8��#�NB�Є��&*�����DX��W#�?���i� ��T )OW�x��gx����Ќ�z�Y`R�"$N���S�@�|i���*T�JQ@�(�&1'k�k�Hx�c�;�|��y��Eݵ����^.�Z����Lg��ު�멡�4-�(��i�/�%>��cS�%"Y?��>jB �d1���%�v1���>+��'�q������;�Tm�ɝv��_��w���9�^rRb� >F���rJ��P���*DL-�bۉ��AD������lX��{���)8�a�t���I8%#7�va�c=�KԻ���5���y�Q�@P_�o���ݓ�Hᢐ3��?ɳ)l�L��Xݡ��,�#$W$2� ���t	��<`���[�smc��Dk�ׅ.X��W�.G��}�A�!�@׾��O���x�4� )=��2��(������W��q�QI�,<�E�pl�$S�8Kg_�o���	��	0⻑�f�?�\:�����xM�\6��R/k� �[S\B��awWġ�v˽g�*��w|>s����`�Cn�?C���?�*�Ӯ�U��-Xb���ޢO~�:�A��͞ū]WF@�{f�|�
g+�ꋙ��:fð�_�1c������6��f{:�_\�Od����h��3�__��3T��rqdK��oS��_�#�,Lu�6�}��1���K��B[�?�a��4��xѾ*��u-J��Q:�'���Y4%�\0�m��d����ivq9�0��d �7�%]�"cy]:pL.��mj�[eZ�TN��C�d��T�-1
��!�Yޝ���g22����������2�9�_�I��k�+����
0`V�!į�:����ںL~(���R�yA�E�.��V����(P�G�t��1�|�h�@2r�Q���8���.V��8|CK�Y\mU�}s8�,P	b.1IE��p���,G���|�.��V�p��6pDDW{��t��4���E�Z�<|�\&�(��2��3�ɰ�1ѬT�U���д�(̨�Y̤Ű`
����sY�|�D�|gz�	�i7�ɩ�^!�~=��<zҢ�sO�g�7�ir��P��P�}����`h��H�vM�h7
�����k$�B4�_����xv�ܚ��X�-+F�F��:����k�g��~+A�~�+����֖�kD�� B�s��J�~z г:r������N�K@X�B�[3�S���^S�d�Z�O ��2�7h��]{,Yk
��M�(���T;&�G4���(��4�sN�d��� ���f�$�%��a�^�,0� !n�Z�#E	UșQ���4ߠ�.g
 ��U��0���ɿ|t� 3l�b�i-|7F�$�O�q��k��jQ���{��c�e63�u��u�W�hU:��E*�b�P�-�"��g _M"�����r-�O�MP;�����@5�����+6�
G�������%e����5'`�����Ap�:g�S�ꭌ�wP{�EU����K�(�M)K�������8�r�c����uq��m, ��B�ϭ|5|��j�:��R�B��J��4����,�>d�R*�2a��$����/�.F�F�3b�8�m�_y�D�}���]�0��8sQ�y�_윺BV�ͱ׍K�BvX�^k�����x(�jp��H��h���.ѭXF�MH��L�F�3㚛�29�c_��~�<�^_�aꁪ���5١#�at{i�q>���{��;�-��в-Y��(�qs) ^z@=�Ǫ�sQ�n���OvMg%ճo�i,ZE��xex�ޞ���nL�R#n�X�
�'��;�W<�]���f5z��0���R�,����"��-F�q��#�Y�6��zJ�S�����~%�(cNj�B*�C"�A�O��Ҟ3�?;�Q��D./�3�B���[��'����;�p�!����~����`k�X?޷���G^̀v}Mݖ*�.9��5�旲֌�����qe#W�ti��Kb��Z����ذ[���J�-5v;E�A�x�I.U�-Ў``]2�|����h�L�)�Rн���x�D�����ٟ'E&���$��\Ũ��.��R�]GsgAk�^��m	��1�>������v _�R��HyW�/
 0��R��y�XJ��i�%zHF.}"�>�J�B��H[�z$��1c��N8�d���zL�
����ݞY�ȳ9M_�T��a)v6�͌�&j$���WN�\t�"��",9�tu��1���ԏe�)�7�^����S{Y������f���tVT(����=�J�ƕCD5y����z�ݕ��,�Q����r,��O�S��z��G�m��M�<��E���F6Q�Q���]�N��#y;��_ҥ|r���Ǿw������*&sC�G�**xg�R�DV�
ˌ)��'�&G����bѺ��؊h;Hiȉ���J��އ԰,ʄ��=�g���Tޯ�� !s��ˈ�t��n�F��J������ٹ���A������گ@2���곍R Ph���8}i8gC$�*
lHo/�2��
����'��A�b$�pw1�����?�͹�M��}�t�B2Lj��}:/��}E����J �]σ��툇缇��CǺ���Yt)�*������ �E�/A�d��4o2[��Mu��rǟjзC�j���Άr��3�+�[t�g���Ēe�z�&���P���V;���Y#���Bp��$:�t�h��E� 8��&S�K1�\4����ru�*��Fy##���;�� ܢ�Jk�����>S��+6\���`�$�j7d�X� s��v~��Mݡ���^e[e/������RH�#�dWT���֚iCe�ü͝���&o	Ү����#������lM�2!>jza�[����c<8ӣU��AV�3��'�t�Ir�=w�ŕ��4<-�
����Y��
���uz-1~�����Jn��O�3���BB�~�٦��Q9\<XZ��u�b�����O���P��5���mN�&X��go� ku�Ė ��e��I�͙���u�df]��TPm���-���61U���J����[��2�\���d2C��HV�F�$��_ݤ�fff�T�X:6O��ҭ�_����]��z6��j	
�y�Tw��g�����j���������Q@�I؆��U��ʘc��=c�a̖��ܔeQ�e�|�w?�ohhe�M�'��>W�E�8B	pa$S��$���->���R���+���l�^��7�/�r�+�jJB�]
���['Fm��`)mea��d$c-D�Bj�����W^G!�/h����5+���@R_�e�h��ܠ����w���r�m#�EnQB���������$I�LF�g�Ki�"D�V��C�Ik0�(P��(�����2AD>Cx�z�=��m��}�]��G�S�݅H��/�jGK�L�S_*f�\AR��-F���)Cie�:}��QdC@ٵ����`d�S`Y�C�u]~�j���>̘�%[�3;��x��up��Y�x��Nj��'<��O�.�R@,v�[��"���kuF�r���mkיּES���xZ�v����T�ȿ�p�v!Z�>���jb�y��E�*��o��Ǘ�:��B�^��Q q.0J�X��[c#���+�8v~�Cj%{���3�&��=)Hk�Fn�
�@���=�z�bʢ��x�Iޮ�%`���XE6x?A̜�Ds܃�*�*6R�1g�z>��C�J��>�'k�6���R