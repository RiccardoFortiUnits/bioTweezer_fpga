`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VHWDk1lfodachVgKKSNPAG0HE76ZZdGv0c5QrpZKam7jGprWRiIGq181Vcokrdb4
Quz2fkImtqOqzxqZk+te6YPJSBpHJMbdKm/X4tECyMS/OzZHQn4JCOSkMTIOlNE/
W3UgUp65+OdmQuQL65F/91GRcPpJx7+GEcDCG5kaO5Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10960)
92o48DOGK/cWaPXoRWsu3LTfv8Ix1zl5CeMr6h63WN0pKExHNNWB5NShJVAl2D6N
8fivMLjneBGtbjkr8WquHMj0e0XF+kiXSnPEe/lDYBnHXiH+tFHTeUMeyfFSC0Tt
hMhkfZXQaudKLkSdofAf21aDh8TszQSQZBK/CRnxjE7/T9Xp7QCgh9tPz9O+xglR
3RzrrOcBLTNb5EJJjLgWSBW2sAeccFLa+tx1TWcSm9TV6E6h99s13b257vK/qk72
XZi5wsoFbBiFEiJ2C9HdRibdvS91G7fywdhhWFig9eD+Mysj7YWiamPazqVKp1DX
M0eZMRZvwwYWg8+ODgF3I6Ljs1OBI1in8mOt7B0dRxvVBwpBAIDji1SRvwh/UVMN
TPkogq8yxzRKWNRNYOoVYybhXdYbr33bD/cZhr5PurElUe38F07zlQb8HFRRhDPd
x5GMeqJeNsZBngCsPzZeqcqiphHndyo8u18CEqS0iJS9tjs57mxiqsPt61z268vc
wCtcJJVjZH1PXJN+YPBNhP4IyZMNwKF2jsMnLm6Gsv3u0dMgRcrB6WfeQn1H/pWn
HRHzi2EeG+StaHlMgCSZFLxIx/NG+PDNmhWaDP4yQI00klKdyGU7E1+PCc16TSKZ
uxOBOwxKQG/ZGDd3AoU+04EU9C5QyItGLMhb4dNU/FNZJjggqJ1LABX8iKrrgcPw
2xZM2eD0pyytsHwMQQMWhRNPvxJm4WwzFnxD9AoxtXb7zg6r0knFyQbk1CdQcl1q
LJA5AQ1e/XoFy2a1BFOIvzUD3v4QKlgRMu9DKjN7NQ9lLiFO38AlWGYyYRw3YjaA
CYc9msvBgdxZLQl7MTv/kyzWrjhQiYV1IIYO9FTnrKmdFklGhfS9wJzM/Lejrb0w
L5kQHDFe5TgpNeODvvfK9ZZgxK/7SoAs6NjLD+1/l6YA7SrjGW58jg5J+P/Pu2B3
xMwWmB8quth0wllFNjwzLoVfPQ7YapCEi3yWZrfR0H6u5YjEPXFnf0Do7MPB556o
gYvv9doMju7uvEOLNbsk9njmULH1DgkLKmcqFFzbJQBY3Wit5bqmvGbj23MBmwJw
W95dFbuwkB6deNVvVYro/zx/M58qfWMCr2BHUGlhJ0Rs+H2rtj5aGfvxvEcS6q45
G4K92IwYM0sJY5qPQe+iMvMeEKH1aggoYFkvMzoVwlijYZxFh+0LepYrRXzBJf/W
Dz9EWEd8QdC7Fz5jcxGt8ab+oQPUJwAHXpyV+zn1vpsiM2mnDTMAwMMekrd0sW6n
ve/ciWp9vXDgtZVIe3Q7HGxpES5tA5GlrpKPJ+71KVoFUiOmUTuhIqLnhXfzIBL5
8lS2fvvb4pubEkRZnDItMhKSA+oUYExR/itmkuAoeoNmj9KFwzHvzk9Gz0g34JsF
v7sWlIfDXyHgxXc7nyEMNHye3gcqb80c8fDYnQV53JaYBxKxI9anoxVJkl2m3M+n
BvsokU38xTBjT5/UILckRRmiy4eIG6L51N6XFSjCmj7uyG8zSoWrFg90N8S9cFFj
jjoGMRMjDKEd+5x8zBU9tl97X1apGsS3fRq2hF/p0qQ0sg0buQaXUoKgVL2960OZ
AF2CUJ2TPnm1pKDuehmvzwAkCXvLwu7n2jWMhEk6ZgAVg2bqpKvi22w7OKIBNKIB
+vz3C/tUj0uUE59cvZ2bxymcx0hxGJdEQawDiNmF+G1m/BgxJNCoefdgXEnIDPkp
xxzywP0VFrLE8N2TCTwpOmp8ubYLiE6giudCGf9qomOTkoC3q70YDBS9PJlH9rwG
Kamb/0cKgJ/39MGRYV8N/aBz5/JgAaF1d5dFGnP2s0mB1BxP8X7V3IqrjM1G1SVW
vEUmxsMkoFTijwmq9Vh6fBqVOztOuDfDAFeAUxutjvcZFZ4cxzw3+9Tbc3GoeBsm
I2cW/00UeqIzInJ2T4FmSPhSq0oLnmrhKeHtXVgz0bnJY7MHfb7NjRdAIImvhMUx
E/XHE6o7PlLnArn4jxqm7BsQPPdP/j75GS7J3nSeKe00EQb6KYvE63P+MZ3n8Op1
u3RUHJ1m69AiqIb6QNuHm92twltVImpwbvApQ3WA6aeLCz9eLsBBkxXapXS9BF77
xOZlE8FawHNjSlZwzJVWLSQUMXdQ6sQNPGgZDw8rd7DRXxssgP37L/4AKvxPSu0t
2HPCgVacp2hb+n67Ql72ImeMdRbhNEAa8AxiXuTAfCDOZcfEYorpH1BPlFti0RNf
eHNqZaSLxeRS+BG4KRkdrfeayU5n/PerQ3b+RZ/PoyQnK03jkW3ufLTdNrfWDxyv
Rc8gf4Aha9iV1lY3Vmphk69pKZpMQCAhRguC8/k532eUB0wtEqtcdx8JEZ9Jk7pJ
ms9vuBcuL/veH5tld9ifzM7lsy8pQeTPv8XZl+unBWm2P6/t2YW6SwkLFzqn76j+
cAmY/UW8UtX+9cfyNRfstJ6yxtplokqe9x83jqw2aVnAFdEM+BN61yze8VV5KwCm
J1a0051SLh2BYj5/Mx41L5MP1TqXRCeCqrdLaDPrrVinUPHtIqKt9eZ6IFZUQQJM
lw+OEWVs9mc02t/ZMp/EOZA4HZpbxpGkrv+0pF2t4sBH+hlxfnNApuU/8cE5X7RA
dsdLlPa/MeJqSFxLuSAAvqcN4vlUNauEKv4jQNxRqhtM+2QWZ+tni55dVN8WfOY9
L/NzsZpnfUw9u0eP5dRdnaOTg1k3Gd5HYZnJnAdVGNEWJ+TsZIr9ESUknY9deOAk
6PRCbYHnLrmR87NWL7r+ibp84HeAs1t7ISE/gaii+31q8OzvCRepmRTfgc1gunqM
TmMkOWBrupz2TsgZddsdvVBrb5gDM/xfUdbIB3bTu7Q2PL51D1Kyzub7o8KztCb/
mPHlwldQ0+dZz5/nxJt+nNKhWH7Q0Z8eLj6YTMeILyjxvLFH4068v8jc+OgowiP1
7bb9thCetb9gKIKgKiXsgNAER2JnTnyXpj2z70uAPo6OMZN80rm8x2EIYxJl2yBS
nLPiE1hcez5n4mj+t2Y2BRW+EFG5Y+7QCP8DtgOmHfWGneVe1BdKGf1MSCbPScSr
S7154X3i0gO6irUHSWvF1MZz3ngbJyWQx4X4QJgELu++Kgo13OE/3quDpUBIl2tw
TT5AYFtQImCkwd5Oi7Cccl8U/b05qDEUcBqw/rCtyGOvZvTd7QOwgjipUL0yDuKz
sBAjc9RHZqjiYK+1B8KC3jVmxLVQIoqzoOqDiWIwEdYVe8RuEvtdZwHcF1Bm3vZN
X6LEICPrJX2JNghr5+kZDo7vSDMip3VSkk7TP5NbaUoEAv9sXHxp74EHJtIxkL0Q
Q6LT9x8xLj0E3yxvpmcbF26mi2NPoWnYtToFnHU1uA2lox3NKyGu4kLlQSkHZt1Q
GiiYqr4+6YKrvFZ38X/LUWZhZU0TPHp144yAvGjbm5GrQSqt/pB8Z0mnWeytVavO
L5Oz/XYTByen9YOpEkHsyhbWjBL0xTNYh0tZo3y0yTmwZVYUSgacj2AB7YDAQbOd
YX5mnWg6asDAwpdcoUP7MlNAQUrZTxDoYzv4gHOOntOHvSFttZAWg+9Y0udWRyDg
iGy+hye3NsQ17q0jXbVeZGzivN559Y4qEwz3Hg7EQpgw3R9JI0vjKusj6Why1qNt
1DY3RLNSOU22+PhIUyIXSVm9KfaTUqH9lXyml0nBT309/tXubyBoWIeOuxW9lMOE
KGDwd+DOjBjl+yfWwL2qyBX22Qe4JoRB3PSr1AnZGhHP//jVrBcNZ7ZMjXK8f57O
tedKs5SvGrHBplXcJrLaZVZn813hqVscHqXYGWRhqUC1AywX14PfUutYXQ/EU7pK
jfeWZVGeNnvMpEcouwjyWc0bC108z9PRZtaKBE+M9KOSLcHgTdc8ouv/mxO/YnZK
pCIbXLQg1IVn7P8D77lpjIZ8pBmagQmAHwgYBlCYBwZgbSWwbThz4uaMZom84ShD
U9VOZ7AEM3DfYuIHIuOsA6yPSV6/ma3PG+IbsSNNqgVVTete5Y3SYz8+8qC/8pM1
RUYb4agGEZg9gFNur8uhVPnPelTi8PPN37M1Q9pOyizABS7pA4iF7LsrGjQckoms
uu+u7KoJMzX2FftyqNCy3lcibWc2z7vVNTFkpMdxUj8SPb3kffAjLUWGZA0H7YGi
ocsPWL6CTQd0QAmTHobpg+WYTffCUPMbs72+a1Oqn3xsGSXHaI+bTHy0kCT6pL23
OiLlre5AoLswuW3ERhQTu591uwsPBwtqlUmUxnpZcpWf5eG6048lmFNMiJh9qBFV
h4G1IUXwS3bWWwccgckyJOg4CZnZQOj801ESPGLq2otZ9aB5wrpc9MeeHC0dfduP
PMCe19Mx8csqWqU8UvD7fVhvfKT8oD9GRKYcH5+bLXbdU6AWudai99kLJBFI8Z4p
apwTZFIrcieg/QNql4B2Y3DPZxw89QEDopaLb5QCzN+bYltWz5siDhxfJ6cTHVV1
FZrZzwyeOMDBLEeJsRMbhIE3rOZr90pD5gWRyfkkPNJM5SUEsUpqvF9y4ShSx+Vt
zY3OsSYJTVzZiBof0NkAuw4OuirUV0lVFOUubyApPqmGEJyL3JWQVJTtzHIDLcCj
Xo0f2zRB3xFgp0/JivciwwbSa51jnJGbGlpgzybix9fKrXjz/7ABMeKT8vVjj4xW
eI/7diMeihhCkDYq28gOOa/qn4CKfJMsK3D8h1b8q2JN6al5nJ0xYJp6dZizY8sq
6XrSJmcu2W5PkaZoqR+bAG6KXnl3NH6GyrhPZmONvuKJTIBMRnHsDGA2jE+vbBsF
fWeLJVkZKo4S2L/QSLqoHyJtBeCZ4a1ZkUT3wgRev4Lw/vLU4aWsxuds9dwvEzcg
uNshK4Hx7F4QHMIK5PAaEKBuYZAT5NipyCy8Wug+uO8Vjzx3J3Ks9h6dpKUGSiTd
VQKz3AX7/LW5XxyYOh5QTBR8+9hkkjzq5YodLnoUkdXVylno+5PnfraYsNoQACxQ
lE5M9gk2LP8JQ62Lgm/ug9leR5BLC7VRAHZQwM7U/vcAC7ok8ya7XZR29Dx1/ODu
HWKaVbiyprPkpsuoCVPem9VgPzbJM0ZvVStD0QWdonIi78xPI9iEYz/zcJkWgubG
sjK0JSKcpanbnSc28Lu1Ix/MMB47SVY3lqHuQHWaiahxdQWuSokpyBZUmuAfJywP
JJ30z9JK/4LDIrEe1RVs7tJx/N0ggT4T0C2FeeAo88aa+P1/v7p0qp689FvRtY3G
A5c3fuz9y0edsNhaS7+mp4wV0Q6EddtjE575KM6+kXqLTKrW6EChF/CewX1tcMCP
JBoVaZL7bhfPHjiN1815ZrjM0uSxvG44DiknOcp35bPMCVdmYK/8nKjDIZFFHivr
D3bFoNrq0vEQg1Or8MBQkTh4pZdDC4J3ok9K6T0gNvCHGR3/wU3H4yq39eXzwIYQ
sz6/hv+j6sZ9goNo84towavAP12g7qCRtNCS/llJUBHVu15JoiQzN2EQ0EvGwXIw
JDinSjtewpF8iyVAKemcojT/+ChLwtWDUYjum1pFPaV5ElS13JSeLUY4XvpaldrD
I7Iaa+jBuPdNrLqfo9pCMTy0CwvW2y5V4442VOzzL2Joan6PtjCq5on5c9Bw2/eX
gm4snuPwjjK8uOEOOMd0kOOdxvIEIpPWYa8lU4KYNkf2Lr19JXal4DXyUkDn2Rt5
GDk+8qpEntmiNJnt3BNlqfJYN1J4L99SjP/nla8aToZeIKXAuf8o1LIHr6p2F+nj
73Gh8btniSSH4HShsrElbU/7dsofA/ob9GyQBJkfiOuFYEqtfyGT0Y7RaBobv83R
NjWO3VV0jjGUBqWGSTAvmViy7i3GJ8kimB1r6scG4LOlUkKUlSJEglBS3YYBQXwU
rWeOIpv/E9LpGHEI/dsTBnNVMWouj8fmc2AIZ4KuKNe5zVJbmtvWs4yTDCANkrud
hPGivJlNZf8knPBFV1k4qx0wzZ2b1ySNYCm0GHPCjNMWX87xLHGrNNEP91AD4IFM
sLhZbLhs8oGHEmIk4nqqWMSdTpAm9IVg9/o95+jb7w1UNNJ2gcsnWwPhGB0SsrAp
pHfVRsm8v/7f7A8S2RY4Vmy2wmRh37/i82QYKeEvaTCUtnmaNU0I8CI73QnwYEIj
XfttP3iIvhP4UGZI7DVW9mAT72ClaKS9s5obTHTB/tqOTQTk9CaWzyYHl0aCGqGn
MD6DoWjDnNreZaOGJ4biyM0JobqCnd63eh3TLf2VGZFDRdcEJ34leNSIkDVvsElV
92hGV5wlmHtppM4yPNsEmalmvfb9m3L8bBOPIUE58KAkGkLSs3q3/Rge8Tt08nrV
J2bk66FJlqWUZyFl+B2H1DPncptwUWSmaniXTLnuRznaBBAtNKu3hkGHtfCxfRux
A6Y/vpE5WWGZ/9bzSRxXCfoG/qfoYdaSxDJl4wpeTfD96PTzilp2dkDtVJrL+xI8
+qIlfniIbRm/4bVhjdzujf01Mw+S98Sg3WJU0o7okJbOIfTEdt6gqADkAxHZWalv
ZYCrZWkf8liOg1KGaUGA3qkh4XUG6ZV7d4642zbI+bvBWtrNQM/JIg1l4h3Spf57
q/QhYC36OsmdHLeQByeN8VIyy/J2v0tcSfkyTjCgamgJGe6TgY4uzXMpELr/v8W2
WMIUzVfaBN0QZvlFY/JsY/wrsR48aD0MSng+cGjjzTfR48Aatcoiy5LIMRLILsew
6VpIHrGN1IqnOKn+Ej2sqmzZny4SR4tAEqlhBaQWQ6OYrcCSUMLs99zlKU/dKJTT
fhJbOIcN9DDfTrszZvBUU8w8tdS/RQ+FSy6gxy0r38XpznO4EKY/3ODjKeDaDP0d
MGxnXuGUZ6LJL03m/qxH0jyKIcn1oCATOc0SsYe5tHqH/Nza/4MII+fAKlVAtdA1
ApHCEAgBMTtcpIdpEvCZvbIWzK/tRTnAs2Fe7jslaMfWzbeGWigtUZ0U8vM8zDOG
oZHeuW4B6xnOOAcmPS9OWMxT91P4uwY6FJIQqtiCzMDAqcWoe1E5/nVcOxiFQZhv
8INFWNehS7aHKtc8mzbnp+ASHXOmQCxiqOM1vjUBy1pLS+JJgGn/t1YoYNworHDM
MkAnHXsppfOwX/zAQl+PTVIGuXCdueF+tZMyJ7NndX2gyDfJO289x5vilwKhzNsL
B+o3KXltWYZM4xjsGjtvflupAQstyoTZaN2mVFNh0QyG357onSneBXtxk/50tVrt
rH9r4xcZhvU4/+LEflzq9bfUpJZOholwKViesdf3n98wwEPfoPi85RItzJk5w6rB
JEqDEkKvQBibv1hIaI1nzm7FfnW0oBCBkKm3ohpoxwkl6qBb6QwoP5Oo6QrqZFTg
Hl7NBJTcVlTdyIakIuLki4B05kV8Z4NrECT/Ror38xsZedHoU0Rg0LUD4ayzZUdq
ctzYpSZPzSQclI4qKIMToZ7SqEpQGATnbBTIrqrY7EcurABP7V5Lr4C2/ZI4sWwI
GZv+TmJwvamlkoIwDXL0/lyq4SdS5TKB+Z9Q0EOX3SNRJpXYQVWT3ttwvv1A4quZ
zaOMvcXzDD8CXLZbz9XflnP2X2VDNLipUrGZ/K0Oo9WN9bchyWHRJ2OKTBhGets+
IHIqqSBzqeT5Ei/KRpC9lpFGdQpcq15r3DskuIdWxDrdPIwKjG/LrfeVJMxouSdW
KJYZrrU4BcQruPAsyYNNdp8+pPhmsnVmOE46w3f03s2bUH/yc39PNFkRWGAQDcs6
bzj/Lw1XJFUdDiJSQ10Ir3HrYlaz+ecbyhbCMZD0Kfkr2+Yn+ixudi2VRrZz2ssc
T9I4BNrwE52OEpfQ9Z1l5LGP3zKc1anISd/e7jcIuIVhG9U/O7ZPzjyH66+46aUv
izDc3qmbPMv1W18+qhIjLvfQcldqWNeQXh/sdl17wTVfGQuFKT3o8glWVwrY5hwy
U5L2CUjgFU1+vc1i9IKXwJHnlAWUb24pX/7RD5QnWZG20RsiZJByrNsPIE0+3FsJ
rtRWunb7UJLLT00vjqoXE7ion47jLsi+BAf6O3dZqyC7J60BmZl80fF7jcyFr6RM
4J76CD2xKDsfKB4viqfk6gdZ/e64dNCcJCjHGmWW7ElMVXBcAB9qdyDSAjK5uJUu
aNW8laJ+Ndf9qlCArsJqGjWVzzvnyea+V5LGUF+UkQrkBeLkSjL8rGXzfB5RtiRv
zff6KF2y90wYJJcE3c2BzNKBmq9KwpVc3bjVFpCuThYxIF60SBdsUePDyMIH8k3G
hdaJZzvYGmYCHJ5G7pujA73o1b6pMUyTAwTu5sw1vYS5raa+/iumSQ8RzS0oXgH0
73DjyfizcvENE2ObGMqwByH5gYdZV3ANKIf9Z2dCmxuLvQ6eXm/ztw6ObaTTx6L9
sQuT73V7mGsYxq6FGJ+7yHB4VRY/FzbQEHdhtsywyos1TWC6ouKQn92KSp9zx9gu
3xnI0ODm+FGVvJpR0bgnzjgSsoGp8228Ax6lkfwncFlc3hIf3dgNIpARqTUUFWxQ
aYfBsHVIy17vwBZfuvmxgi38lytAYWArv6VE04gZ1rvB01gNkfGzHWn2akb7UCO+
mjNUl+0HHHIHIhf636TlCZnVtrThCZUqt2oHsFpVSrjEwGnHwJ1E4dwwjl7VIbEx
Z4Ui8s3YToa4UzYO4jeCn2dfy5Td6RS2LSAErKY20lBoRYOGCJ8fOxPaVEvq4l/P
dKq4iPBMFSPtKvw7cWmXUxEVYtsdq7qS06sgEY6Gp3lf7C+vXF2bLSjhv9Ueah+h
6ouUa+iBhR696V0s26Nbj79YkwGIDcGKDq/nU1XjFzZrK+usPJ2mFsNxXd5BAS/i
d39ypODkCVn9HmiuJxnKFaURUkdDiQrWSLYNpzgeeYtQ+76s/DWNBfS2wbcicHfE
erTrvFAGQx980mbB/cFmHFK1oCZ7th+a4sEL96p5ZkK3JAAunXTBng5TlV81lu88
WQu3EN4Jt9MvUdtFUqzqvC5VP/Fj88YqcdLbiV2H09eUZZXHyZOD4+rqF0h1n5bS
O5DhDsfXgQp6evFHcRxd2et9nMWcrUkdir/o0qGm7NHPTktzy1m7CwOLh6IIDc41
3iktZ66I91/PYExlA+RxuaXEjMQUQrVyed0IXSkcGwHu+PpQol7utFFvEW2O11Sb
iKx2zGv2s678bWyFICEqjdw0NLU0nwVc/L+6h85rWNAgwdmJ3Ah9OPb77h1x9+a0
F7Db7S6+n1joAdIbSGIfXldSnSuNOOMutc2AKupyHMXfgqg/3VPXiE2i4OGfhqbl
ziUTdSB/Heh1cTBuYbY4EOTFQgbiwibE4EqalI/T2cXDjpKSuuHnVFTdedrN6t7I
OaTWEUPuX6j284IYzOpo7ddEzSgbUKD2yLwL5ehOlJFrcuHiH0msjpe+j3VS1nb3
MEjP4LscN7XNjuSpsuL9I3gnSFfoRBKU3po0zYb9mKRZih87x9DK3dR+d614gfwU
aWNzCxugcZSYiccengHnozLfuIJcLVgIKWLFDjzibdPoQRjlS3lyXynv8kBJnlGE
NYgIV2jivrNNazrZzi9P+Tp8mZZqoaRfvwtp+XxWY+YxHnxmGtDouSH9yMXuZIAe
uGKTz+cAuuZeTy60Gi1V7wUhX9Un8nZGIG9++q0YuhPiEgWwD3S6TClLNjYdtUIa
T3V5373yi+FtPJF3uXHs/S6PwQtvt4ERXYYsjP0RDTdmkTPtuyR3SscpNZ3tkkaj
I2E9GYAOGwCitALoUrbcLEMZR+plYB5XIbIq1Oa2J2ACkMp+uUUz4LE3eF/THx8N
1pqsCVAQezSmKtX+OwEo68LmYXIMDIIQ4aWzNNdR0SK0fJGZqBrH3ySqZMb/XLyZ
++uDf1VtJwOo/KhLgYxakbgVUArYjdzRg5PRvze2NmtLiHl7N1AXYbVOtpfVdN+1
+/yZe4TFI5kwTCfyjBCz6VOsLxwf5sHwUfPzo9dnSTcx2szmLaMb2sGweOUflrbx
PGD6sWbV0tj9mcT5kAghdXEiZf1yXuGhaNGjJGVaXURJZsp6kC6MbT6wPCdyjc1d
+IJHwEe+TdHkt5sH1wD4WwIOD5aKtBxveH4WMaBV5thxSmXnjAR4fJuaKjmJDlTq
T8TuueT9Azn9ckYDrWWzh9YvLXd4vviK4Lr8eUmmW6IDxVZt39/BwAJguaetltjP
wQZDgr4FsPooue5IbKJf9xAxpn6CdGGppCvNsaTmZH9+SgKXoOBafTskeuqULZcg
DI4mBjTwfebNXIl4+mLKC597/nOetjlcD2rA4QBUKVddgMv0upSmuwdOl36QlStx
Rxevd+ynrjcjXldB8XJgFLJV2kSPvvnuSzTjHy0jBHaHfR/unqLjvVTH29GL3p4R
7fzowDMxI+GqWTTrx7RNZYF+ft++b5dgDefeU/eSWOYHLKvfF6vkaOdW/2GGle64
wjFFV/Tezq1NjxBkQCi7SHZO96ee7f+FP8AXlX7f69kPPD9cna7qB4RRNJdEeWT2
/p3222ugL8PMwoRMLDMXYN6mhNpcFOtQUsdC8kspixX1UccDWX1+KozHJRhHy02X
LkkgDl47J86MxV0zKYCjvLTZKfCbcMi8d3aTwAx1i8csOLznXXuY+y6RG0ygaDPB
QIpzCIGrwJ68UCNOjjlFJDr0RrDWjk/yS4fO2xqjjXzJ7y2fh4zWQg3ahLh0FWAo
Fk1G5OZ2APtXsB4gQN0rUkMi/KTkRRrFRxQwS45UxGok/Je0BKuXv7vXIeqNWFce
njd/yUgqKbvUCuAYoUM5o1EnAghuVQB82CYJcxwQQiiK8avTOVvsA5s5cc8840rX
J/249tPKE6G5jW5MrSMshymAowNtBT73MWT1ZnF58ajAApe48Gj6n3eH2gk6cIWS
VCtT8ByBDsbd3MFlWKyZsP4aKsYJdEMFjd0fJny2lfRWM+4YW0bqX2JP2TT1JDuL
oXCH1qDLEOmCklJLujbLhOT6zCt+pcna9YeKxyRxUxPAKUEmfxe8Vfse2YYiA4SZ
4XeZ2qNkgWuaYT17NvaUkwJ+67Xc0DPuQwssFXPnIC+ODjBTDFi2GpU+D30BRtdz
xtZT2H4Cdwg8Wuzllo5jEWXviutk4T4f61BYc045xKiCPtchflGFFxrKnmwBUeR3
z1SUQ4597NiSvFfvIUOkKCorD7sjvFGFie0TJ2H04WeFUK5M7Dkkps5bC/lVzXru
pi2zZF6UU9jbHOe7wfQNnNWIich+cmK7MAL+c90LLv8z+HcP1VTgHxAOTQnxnYYK
Yiopz+6SBW6YdBQnZXF0mWmeTQO1E6yYgfxDF/5niS5yt+EZbcabYPI7j5owUAWb
yRlmKZM9oZ6VJIUUqBvAm8PKMIs68bpnbgxgV+10cttZjr4iyFSRxrOZ90n1ekUf
sH0cEi8V3WE4vMZnncJn2ymrf0Vg2e2e1JNBk9EQbq2IUChTf5TaIujLHG0OlfeH
bcYX73ZssXLHZ5ii59mKbVAKxszi9YNAyvAbB5TtSNbB68Rrl5enb7kaQEdrzBPy
shjLPySiTToQw7eSfuJ/0TBuatOXnOGT7Jgkpx6UZdmiWsPFyIF6tnQZSXWxuOe1
2m/BTzfqpfNudoEZeUywdZSp/oDF+p2xH5qJsWXKly/uOzJQWuQ5djq558ByR49P
0b4IczJiS9o2+Deydzhh2411xaZ75yyobt+z9M1d+K1bPcuNX8DVrLWi2JkYe+Vp
Rz2HwV0MY7b4GNMeAqsEavOpCYM6WR1d7ItlJVGyo2vYDg9G9GuKDKWIXFDC498r
ZMoSIxhGpcwTsUFIcOyZNbkhRFYgjQDPGL6Eulv3r0d1UlAif9m4u6yERP/nECsW
h4QJKaTT+8+zJTdzQlu7541CsNiOIq5NGez//NdLIQ3tejnPpQbyBYJvccfOfFGd
0EArtj8X/wKrFWgsoP3rH6M+03ovwZSeqAtKonEd3OeBMNtxXqgGJN6LjetVpOrq
2dy1BWsbpx1LUM9ntI7QZwsDCuu4KiD9PvCnhjoy/HA7aO7Ej65zbyupPsIWuxmT
ROx7CA+abLlFdfdkKpsQZk2fdl0t27m5FYdxKPbyYGjd2cuWqaCm/Cfh+gGH6a0O
+0JZ7tCaopr47/aWO1aXqI3j2ii3++Vj/TSxAECUrM3uVBjGN0xGuUCQEO7PFYMD
xjl4yO5HCvOyqz7SUy39eHXm2Ix80LZYFheuauz/X8WGWAHd9LfWiZN0LvHtvLi2
dsQkBhcQoe3s65FnOvJeN1SV2U1RzTvaloCD6LVymK1Z2+Kkn9kl9VUPi0rkQScV
VwIYxDBSK4oqF+XP/ULBHuTF/tI+138AbVl7i5148w85qB7Zbg+Uer4D9uJmJWqw
uVrJdQ9FIBiu3OdRAXl9Y2dng/l1YHEcWn6UoMgNqwaJYJw6UhHD/Ec0Qj6rGGwz
FuQ6jwy65Wi2ebwgSP4kQ+2Ha0ew+RCHlOVRn0/vh+OxDVEaC+hUUUVsDFbcS3H6
ivujco3PapXUAXGDSwiLLrdFZRB5SJKj+CCAF+Y7VVMEe19P04gBnhrI3B7dSaoe
Smh8aSRJObnsP0ZVnT30Hd1r+4cJcDEQBFLV6iP7LUh2fao1qQZ9TDq8uWm/SNMe
A80Kmewpo+95vDiXiESm66efCOJXavzcu4oSJwysOCPosBRx8zVvZbqVNO99/T9A
G7368EDXsPrwBaNGJWMrf3Dt6Sx2njfp/cnpBf4TGtU+3ZjWvFZ1fhYun1/TSAeg
ARfkzSWKcVBvQnaqETjQk+xhhTCQZqRZcz7qqsuRsloRRpm0FU0c0KwTCwB51AdK
MRy04kAVynkSrwkLTpz7eoRGcIZyKSY6s9TcihvZJLKNOZVFmFFGP9dFSeXj575e
+n2biALV2o/PPxZdplZY2uxds+FK5NfPpWhil+/xLS0wvpMqq2wj8SORy2CcqZd9
puo1jKkqOpI69C0+9YZ45Gqhgw2UpRp/4kjjKZpLrUCuC8F6OOCVPVVE+93Ew3p+
nb0ZW0dRiOGIgn8SWdmakn3QKu1tJ5ApU822FZS6tGribcQn9eoupgajZastlb+f
YAGbpDX+/Ddgck6ljIH96K8IshBmhi/R6RCwQhGMbZJpbo/ihls2YZfh8nMPVIat
gnuwQDaRgbbEfoqvEycI3vBn9ZnfjEKZTpGAW+6sL91yUUjlabFGkbebqTMkeaCa
8+Rs+AOIqAI+saozJdCWZ939z4AF+PsXkcWWwZmlJZ+rrINiGobLUzXEg3mSE3qX
qqGfVlcA8KOiP22Yf5D5lTAgnbzUOPp5MIOLJqlTsB33CVL1Tyyy7oZz+TdlonJq
UwxVguBOX3hnY2iE8W/0mcpgjx0iTzYAPl/9QjqTi9n2Y6TjRV6AeVL8LtgwPAPH
Xu795qGlb7gmcnK73FcRcpaMMxapII+TzhyYXw2MbemYmffttey8RNYUsNXUiges
xQpfODoSGeDXyux7bybb9tyPM9dv8X8yL7+djJ8lYyhh3Dgw9oeTPDMHl6THfcvs
5Io53YYg4RE5Cpl/6uSnHxb7hgeutWp5yhvrxJ01Ab3Dbi566KBS2kMynIMltwNn
QOc6xl6PnBHnkJrqg7GOqrU/+tJF0bWHlPCyFrikWzL/xLJr8x4VzMTzLg9j4cG/
dnFaZW02XD7K2hX/bDU3MqDhCKRyDUUe3jbM0LeJRXtDpMygM/aKsWNTnoFkZR5C
0kwOE3H23O8FGx1nstv4/4gc4xrb50E0eufov9r0UW3HyfQy6e9HnzW1ylsPnpz/
c6fpDDQrENvb8UXcnWGn0WYK8khcUE1lAklRxzZAK2qL/CU0iX3ZAy027sVa8CLS
RMBzDeNbhS3lbYnNW1+F/l8nRbDy/ubLDvDFZG0TB0+tEJO8SujsgbOo25CW5ilV
AAe6D9RcS0oh51WJ8LU7oyvX8zKlPNIANCMZz080qzXMs21gmYItT8OfnJj0z1Yg
pEdLKsxNfjkQkw7a61xvDwbVPz6bVv/qrouKCep4ezeCzXe7yiL6E0FWzADUoeOU
En+cXj06ABRDQILldYdp1xhWyRagcSdXIqyZuEYPOLvW7mcnlP0qDFXOIvhHgCtN
nM7H3i/OCg8k8DMwdK9VWBJ7fvYJXmZ+MIWIjDxqcfyJr7puOikCkHnXF8/TEXii
KR7jVzN2nP+ElsTtZyGZerdGWs65G6TbwvePgshhgTQbYusqCkQ7e8MGfh46TtpC
OF14E9NRqiALgzIjOBx3p1MbTOQsgsJ6mggOsYqgSOnFmbJJ4IET874IGOha5x/a
VUD37Tbn29+rv5UMRfe15VUe989UilHOothRyNI09xKGcD5num7Kf6ZDPIXds1dh
MO4V5kJvLvj+yZPM8StvLVOCaxI79mpsb17YNV++5QIEMwCrv3ByM5JtkEE7A+ve
drZO9P3eprc2CL4+nsW9nR/Y4/CcYKuqLYHUVarODxMO1FZ7J8nKjZCrKvvNe5px
J6aluLt7/5wjTucA0ZhmqOumZZtGWg0uk+KqHbPMckClmnax59woYA7ZZNV1I4dm
kMliYOWkSl/uJJmzrObEBvYZwauboeObuxkk1VAOD07NdIu2nFDuw7i7q97tNo5F
ofeLeUftrUCQBZT+c/2cTQ==
`pragma protect end_protected
