`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eJ8XWHouVCBz3FhTDH9npTtjl6KRYjm4M88utUUsk6HqaBMlnUjug9CCYQ35hZtM
QfNFS/3XfJSq8LdFaXAYNVU3b2yAG/huAYJ8ob3pTEE0HGO8ecISMc/UrsDXJjQs
Ri72YROgp/ohigg9aJXbR/TV99bEMTKO6SrL9E7aQ0E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30832)
4JSXy4qPQgW9sE3uy6R1bqAL6RR15xb5m61F1djT+OMSZ6vKl8lCKmF301Setf4L
lv2RcUO6j4npc7mctRbvTQi/cIqedTGqUwaXhksK2QH+r3Bbz0dKU68iwjtcKX3w
6gjRDwD0O6sOXLcMpoVLUxjtRY+VHN4LowZIdj4jX/+amALRWodhsC41u+LtZnRn
4kixGFae+Zm6/rQ0pjWmZvN3n7H2gsKnooF60IjnhF5RXSIYHqppHaRB3HLLbFsj
2fCpf1oBc8RcP5Xyhst71XLeam7nOyv1dNHoW3PsNrou4p5nir/YYR6P5Dz2siMk
MuHlWhv735zdxD0MgFlN+ySKxEQRz9/6Dj441pqA0qVuLM59b6FPp2/uEB+RQnn1
oJR4YP+1DCXNT82pLO8nCgbJHiv03Lijrme5xxyicNm2WqYR+mxUx42seqX6R/Pi
l56JYp7PdPnTzBDz7kZCwxgm6ICmYzctuUAopqCh2PPG0ykH2N5t3HQ7vOkw+SZs
9F8AvevbvSIxoI3mwJ4sp30f61LMt5YqKJsrignT+RmXsQtOwBZM7tIx4/dGZ/Qm
aYbnj/tGwRho9yIdCEHaCmuiam5J5U7yyAfuXZUcB7y4K959FMAsDzZ4rvFoxPTa
64+GwmmR9JezXpelMJFNomK1jjZe3vAd0XxPDPN5tss8PF43vQ3gnvlftyi/U7b9
YzGj3/dBOs++J5qlzWnkmHEAe3/gTvdBpAOXNwmJHRNMT2uUJYArGF14d+pxeo0u
LQjJHWf2OCw8eIZBBuVsaGxSTwRpaqAmcN+pD9yIUbHsk/B+zsLfY+ExmUEp6ltP
ofT6xXgQXzaiaLQObVRho+Sc/P5IjHYZhDlm29JYNzC/VYm86oBy5nTkXYZPngVs
htt3iG2NnUZ6C4CfMO8GokDUogz5304r1TIxRoM6VJ1H869q2T8Ui6XDK6dQQq+f
B/hzZwdbEkHkXz2CIeQcnLru1uScPY91bQayvulU4nzf6FYxVCtkpOrxuxG+LL7E
zlp3KvU0do2ktSpmL35xSlPqA1PtwFAJwG4GwEETqbx86KikDmyiE9pEh5EA+Uzo
JZfzlglYMzzCI4VM9SoqoJqbdm9GZyDCsi1QYAMGNaHrEHwyWD87qzTT8wRTa9xs
8JM4eDu0evMZrW2CrDC5ZOwPthlwXwwCgV2vPhTLpIdTHnIk+QWrk9QG8lRd2MEg
5Uy8NhmPWVmqlqCP/E3kVqwf2kK+twL2O1qO+vvPrQhn02Ip0AkK7U2e/xaTaWtm
Dm3ax93ZsrPYSUzTXDoXQi8TSp97+JLIto2GyDheX+dQst/XCYvyVTkn6BVD5hbT
yGy0tFsCe/lmxk0UXuYLDza6LKW3BEc87PORPSP2RWp6ZrCWrif64zVwvcdaAaBU
QW6tNFToqri0JrNLOSa7WossMrlG5dra8wtantLqmWEwLc9DfPhgP/lujxrFgz2u
RS6feRUWnfGgvsXR18hyp/NiF/fPETrbpY+Q2hRi8Dh0p3H4Mbl608F/J59hmG1b
kSwm83klR0nLJhThgAGbJ+mbxwNlJLSCqNJvp1y6G4zyge6f+bzNDA23WtdYSnhd
1EqzgoZEXm4nCCY/DObQmCW3cXCIkU9nlFJZXIwa5t4JaZ95T8RG8TkiPPjsqQVr
xP6lg040tfhnLHPr3EHBUNCsOBmtoGE5Np00RVfrJKKNVxixufxYuSEkR5KFL75g
oECi5H8xhQHO7zqf/Eo5SsPqZGdPB78C15D5f02TqCIe8DxBi8ULEErQWCbLjtfA
+EYQlM6I25Ss7nF7hQDuF0LuLwnxx296WYCUtzURr6gV7VDcWaSSjZB7c36UareE
u+Btij7YSuodeAp1YG9ekD6XuRMaTsFyYHsAWYMMBInPqD5K69rOXeD7ARIbjMiC
ueF1Tx4unGF4pkr1NS+MRkEa3R5m8Ptyq5NpjZ8p1ts9DvVIpkFINpAgrRXQLcbV
I1LbRatAg/a2MRQIE8KXCmDa6/v3zpQPRzzSfBPt3mAXMgj22Fk8EKDas7JZyEPL
IZcB6GMW+B6ngbgyegbq6dUhJqHyXA86gV8w8X8l9pLeNxQGhenLyIdNxiqpcRt8
fYW5fDHz8RgSjADf9KVZYMQqXlgtey6c1BI4xih62+g0WHxrlTnZR+ccfUr4BMFZ
9bL/zU9vW1pLWIQkjs85Fxdx5ZTl0w1KNqq/7mwCxmsFG4HWy5ChM58NWoc1hZDs
/txtDuxCjYSNUxoTpXRT5rC1d/wLWVOSp4s649A9w0ZAq+xzKeFt980NkcCYHs0z
ijDOoU0pEOGtLccQ6pga9+zFhbeMBh7T7rv9Gi0JZc9cowzIF053wSRJ4ItxQgTd
K8ho8y8uUmZGd+sdYM68sU0W/xaxEklZZatEaN/Bq0x9YJgjyDzuGwB3oYn5firv
widHBqFEIrDzQzmMlqPGqDmJ/EntwTnNS4crhEsIV7RKP/pVCj78NDthkRt3rpZz
GRMA/7b6Gi5+t0bgyJRyCb8tf0khNa0moT2wgoZqYGbUrOY5/ZclM/IN4MvXDrHB
B6I0iybB5d+uWB3VOapggJW8hchfxAPsFiCpr9IuLqrs37RkkvkqRW+L4Xmx2D5V
Bzt941BBSEN11/HMfRO4LFbKzgCn876AXh1GZ43kdoTHPa8ODoAnOmRdpHuuqr9M
MgrSctH8/Zh+mOr5aNfR5dzNZGQUizvWgmShpKT1TiAdgvUDxpfghdMuu2jJSlly
nn2K6mVAfwftgx9aBuIrBpvhbxnCa9swSWBQk1Mf19XN+458PDn8nydnfQTRXAiw
LDQKCICfH6GrChFPee9GtM+tyHh7sHRbqlogk5lEG5O0MhCGauXdrWcK5FbDytmY
qYJz79F1U6uYWOQunJre0JsiP4O9JanULaaeqiPnuXXorjGcC6XnTD1Y7fzkxX/C
GB/hxGxsu/atIjRWIGHcdZPgSHhBwrhq7EVU4ZgMVvW3HKkPIPOGGze9xDp8Su/J
/exB5so/AUxUBEZ96U8eOstTXfmDsbK+93PAuxd2FuHXf37DqovYxvfcmFPhDOG2
oi6hNLNJsQkh1tc7CpX3t+ksof1LMwv2S2lGrOHR1qhM32mWkOp94G09LNnCCaov
XjdC0ueXprVxbwut6/mYFA/WxBLtQZRRkidBfyMzXU4AcJxsiNqplADC1I9/d2p6
tTNrbe9cXt0vsSBqGuuz6uwTsHkyROaxQaB7CYbB/DD5ihIoKh1qYnvnr3mb+9y9
lsXErCLqtYykXPpPrpfQ8PAcMPaw5c7c+T39G66oXrCqFsdCvNSZuMv7tNY6fOum
5wnMmny315ZygY7xTcZPDFudojjtbZAs9j5pzXs3rIuIY/1Eubfq+NkqHCgesIax
XBa1H0EgLFdH81v9GpV61lo11E0eH655fh/dYTkQZN3pVApVMePz/n9hXfV+NTP8
ygbuR2xruHgFndyTKXzvdXUhci4bJD6anfJx2drGJCaS3CHkUjy25eE8xeg5jd8u
vYL9kB43a4Ew0RATzfu9qI+d/OGNq1JVxyaZPVDh7B0TtCxjQxGSUv8XOZKqGdC7
82jMzuvvI2KcP0n0WR5GP3YjtP6LykTgg1sC1ITdMfs4+osN0Mo3Gh8T/oCLHoQ2
XqpWXXm6oqEE8f/k8hPxFl1MKc7tnt2gHm3F8Zr0mBWLxuJZVUWasSPVj4lDCl1z
fuGcWQzn4mZj4MWSClSFveZcZBTY+H0Nejeo7FJYZuzFUz1kaeE/5GOIfwS2NLJW
SAIGqoi9dGtVLHJC0Xdv4JxJQ5Wc5nrWVC2icUhfZSBX09suCmG8PzQcBsUUZI4B
l7TNeOhuxmKoVTw94SOT/DlzWNtbuKmENI94b5zO14OlW/EhkosQ1WN02/Ls2wan
4z2Oi9DyKiXg6Xomn2GNKTY8MtR3xUuxkpylgGy0DwHwSewz8u7CoBcHSfw4N+7o
2n2LvofqyZ2vIoCg3gZOfCLqOMmhowGrl5VGhYdN7kJ5PyCOpcLdR3iVz5+nJw9R
ck34jYAmTMRVUI3JxiuzDS449q8+rYmG504pJc9DNH+WBZFjGPhBFIXyAqBHtHOt
OnC+kpm3dm7Ps3Jv5/2UGu3iy+WxKIi/sZHzZ5PHqSQNHIHmK5Ed6JfmbKR3GkP0
J2AjEjYB6Op9CAbb62gG7mi3gpNJLElxSB60ogVHEQusbU/xPxBFRCc0NnQaldfL
4CF4N/K8WBwoXBXS1jS/96lWzU61I8DEURgCRTuhQx/sNjDYWnFiz2QD9ilurclj
ADNwyE+vasw7PpvOhZi21nofpyqPiCVJrEOXwA+Z25BvKEGK4+GApXgTPv/95LQ/
V0W+sNPVsstbKmqLe2PO891aAzHpCZn2O4pp1W9BbkqpyM3s8b7BB6no91fW330g
f18+r3ULv59eyqc48WjX/BCiStIcT7oKwPswXo0+uUWj1xR8a/dVQEEJt9D0oZkF
T4TZQUFvRAQ99BD9JH8frPc0TWAeWjdCvUgrUkxqekKHcO6Yw9VgzN4x/disp2yC
omOopOn2e00OHE8JKU2AEBprak8xPvQQTH7O66iwTVuAhPtw5h5j2s5J/wbv1izC
VLPTwAOTjTaAbxJSSmenyZxphDaTlHUqs3qwexWQDNM+0NZLoiVzu5jQnucbGAlo
xFyeIWQPVmMcLws3XDUua0lNxc8czUbCGxbj/rv5rCMPP47ScO17dP9LKgEHSw0J
cEvcojzLF2ZyWAsmVad0k8TL6CwQ3QluPrOlCeE0d8tKuLNjBiM5jkyc2GtIeoow
OfjYvUX0W88mqxExdj477c454XF7cxaAG8F+0ChMDt/eQgs9akonROMPU+gZJrXR
mKriladu/nPdxTp0BGq0G7/FZjvXrFzY5+xWK/1jFz35DKc3+8ch2fuMmyx7C+u+
NuFEy2RDlGFm6mXsrGcY562LIUx1hsoB5ikU8ddeIc4OeFPIpM0kq4QvjqnaJw8K
ToOPNkM+bLg34A+Ztq8o+9/5uGJw+iz1L40ALOi+LWMXdsVfiUEhX1J2DVgtlPAx
UGB0ve7ZitU6GHECCGhKFaXZvgal0AuDbsNGvtA5VUMJdh2WUsPKCsmeeVPUxEJH
QnYxzUAZrYyCiWQa8gDlHl6TOnWWaK+Oq9goPp9u4E1LDCY1Mf3f+f+W/vudblKP
VJs9JLMymOXB1/WMQHkKdwWjWbrp7y1IKMvhQ2DrZ2N3/ozESVFKJPlPPvG2oZ7A
+gku3YwXFH5Cdlbx/Qz4umxFWwlEb7tbSJJW5CtCl4rTq79enfs9yeRAbOExSJ1R
Zo6FbpdPJQ1DvNNwTxFslxJDYIzUX3qSKqgijVu4no3Kw4z4oOrxZXAMVkRc07KZ
yLx+LE6TBEDr36Z2OGF1Nc88FPBX/DZMJ3xb8lQcEqhufTN233uXKD7dTFyyNf7R
K0O4gg4nvcanAUBPbmokJTtYWvusLVmxannh6h0alM+Ky32yzqokgDjI6kozigTS
F0+r1sIpQ3qhcJzJoi/BLOPDuSB+w7Ag6RjiVdraTe0k/4biNEGFaGDVkv0P3YpF
8lBPBAh8vsQ+Fmkx2uCd0junsA9gDQxEe0M/b8AISaVALKk29FLe4h1cIhCf0adi
GGx0hxHe4sLM7gxZyboxkjKGeuhS+eSR1tec4zgN8+ZX+DJyhe+YVLechUsOh5uR
baYUTQ0UYOAVR7H/Akp6MxGQ8GtYV0Vgkk7pElCX+yEQPWxWTukW5qtWIjB03tIt
70ZQrck5sLTMDC7GdfjAf9kQOtU+nKPr2x5fZ0ji/jfJ7RzRE9obZ2E0Upw6yi6j
rP0ImLEv/l/g1jVLJmexL93iKGEEf5hqAGDtTvQb1vCgCNnUdgOiSzL+E97HsiGm
w4qb2vZzk17M4SW4ajTgilT9Sw0Pgm0kEN0N32y+cSuyPXzTStgw+Cce7e5AZ6JF
Ps/m1blvCal+ign/0tdN4WfblbRRh90ylPQhHNa6uBUCQ6fXBMO1H2WidwsRHwMW
PTFLmL+J0/C96nPapioDc3vCpEg979/ZqOd9M+6HJ7xfWJfNvH053ZKwQnPFifS9
+dFP8MlmRHbBWFs1DCx8gP/bgejIk4jx3i5KYDc/wuenEIBx1ZHNmy5mzgjLYnpj
IPj56+wLygZB/Kk/UZ/ouZOOd8OClgaLBf3O7ijRN4PZOydaIL97KOPeGXgYPzL1
WHwaj51pkPlE9J19n0FyDF/zZo+oOAjZKPkT9OlSZXppyACTHuhVIGsAYwpzm0xT
ozl33lMClEmPMakR1flXgj0lQaV9ac2+3cCbojRKZJpXWZg0uy9gwe9/s79lPAZd
c6UnlSUDY9mj91k5WoVzceTAEhVfnpfsqxJ+YNW7Keci6Y7O6208oeAJ2JS8dpqS
WObhro9Cqghv3I0C1r0NMHp5bTtFRaXQNZzU1Pxs2ZagPqoD2gH89jjK569XJVHy
eEDYoHyd0/8I2WGi6WoEt6ZoBKQRHwReO5MsH3x44iU5u7sEvw7u+xgKjBx/MEj6
zqpXq2YBO877DT/eFKmi4XjBufofDCbJWFEVpH67m7fPBHyF5pHxUGEgX1BZKd/c
Si5FcEfZUDc9n+0ysF5g6usOMl4eMEPoKZPftvXuEgfGnmGxdwC36Ysv7JRjE0AN
uJgnFXcMhTTUVGfbUjtESsMiOk3wE+MeV9/tlsnrT6h44JRdh7o0bVRLgywAC3uI
FH93nkqa3WHMyR3ZsKOQT1KN5wt6qo/0oNfAmlT9KOZWl//OZ9hSSR9vHEY0JcIy
iBqGHGmNMj0xybt5wPjLiwtipt8zmIpe6hLopOwm2U5uWQbfLmPiePQpzKRG4nWD
qTSfP0aKTZ08fozCI9Z3FsufAHThpspXjuHNA/xAUebTWlYKwQEX1qe+pnNyxcLH
qFTcYrtlrb2ZmJL4jWKiFWJDZPxUKMFEZOsV7IkbrxowLgAFhA1HCbVsu0bdKj2A
YRhyOHYnYONYafHDzVi6/9LQ+fARUNlfes9Ge6LJMc/4OoVGf/P78qZAL95HW6cS
ieO7IuPkbjUeILAdDt8d5u+ZW/zWbw3ILlmu9wZCT6lZ0NJPKhHc/j9IqaNh/Ea+
3uyrr9grmstpb1XlUOVlGbjHFsW1rCqHS+52gG51Y6lwhJt3irc5csYcbiTWMXsy
mSEeOHxEZ+NXd8P/ZcXtbE1w2m5DyVIhQOUoeLYi+xWwVwONXU63Vm9vDmlWRiJ3
6FZiAQw8wLaa9IIDgD7LeiFoksxXsQD+qIX9K/UYS2pEEu3qaoPiCcI9q38oW3R5
5UO4NJyVAoIR982THOVqsBytebpFOde0LMpx0PPbP4Y5k/g4fBbDfLnNJj8LpNsL
wBUq0dNftl75MBYRo6M92LYlA/C9PdLFO9/pfiB6Tj1H375fDaInGG0ft2A5LN5h
SE6AvhRGezMKZNAi8SQft030S/eXO6jU56CYa5YDpjin6zuh2eck2IR2F9eY6Ur2
dX+mqNJtRXtPf/HRkzo0zVdx/rr9uYcLSFjuE8OA+xaqFyoYdq69Y8pavpYzV5kL
1nzxZg5LzJ8fEvpgxk3ihk7QGSTbiN6ZtWQGH+iDelUqm7NC/SQc2ncg67oTThzZ
cJcbbCgM897CqpXKC0zR5LsEu5kgvVFkOcuzEmA/QrzDsazlkXm06yTLIwGZaW5j
neBIwLW5LMsao9Fi3/UYCU/BxI52okciuJWf+fjgEEnYPAshi2GgV1igkWUHne5T
ta3G7dPuMNNZIAybu0fCWySF+gi7+ONtmp3vUh0wAvVzFOnm/k0G8zWiEB/vwfZv
GfM/kOjRqlRpUNExfWe337NfskLZULrUdL/Cc2nZ0gJAZpgtxpoUey0SWHg0AAH2
0ZrE7Q6csRSU9BJdFgNrKmpSnVK1w8subQjiyy4GK6tvQT7i/F/gxfP+iRG4KYna
6I6rVs/b5+ruE/7a1Ce0OrtY4Sfn4KUkFkuAsr+i5R73jMI/EqpXZlXbZ7EC0H+Q
50w22+XqX4DmNxb1ReckID+7Fv80aMmqslsGe2r5Jp1DTbvFZ1IE9HFcpJ8dDzau
kJyghsX4Y1Rvvx9XeMwD68/OH1Fx73KvS3Y2Ly+9Ev4wKrfxx2ZA9iwFW9GnJx7v
Ss5HzNQZ/KAKGnaWHGl3wuWEAVRUPoPocv5YBGRowSoAyiU26epZf8jD+b2kaPKw
kJw25mbg9LCkaQb9JoAQmUMOLyk7u8rpNS7C/QINyOyvv6G0Cw1JjXz0URGur0wC
5awt3ZXUlhGxZktqPY0nMGuUxPiXkuqgJC7UShwLrQNDmHEbpppIZGYZ3TV2iOlS
ZsdOHDd4Ng7JotSGDV7jal6ICj8HdPey4m3F8i9LTQ4bEeEHZJ+yqS1QdupCBNId
lliPViWKusdWalTyOfitgyq8z+PwHCagzdu62opd8EGpJiPcQU/PIyUd2SEj6ubJ
t+1bQGce0ab7jIKeCsiEq/OMDE1zAL19TV3d3KWEOEsLLza6KKY6YpkttxLhi9PL
8A4SCzEWuPe3WCCQFP+yhKoRhzoghsvShF6w+aJ/BGtrleNgvuI3VlJK8r+6xC9a
LSi8bEYbVxKTsckPZ/NsTT6CWF7omB6otNtCccejmJ7q/bQ+YgfjEwHxWK9gKfcR
g9Gyk3a1rQkNwgVmmYB8GJpWND6M0ZTMShYQbJXUQD7VbAAei52T2jDuXKX4A9GR
HTds/BVF6znqaagPZ2wxVroQ13g/o7OGigVSZPPAAopJVk6tZamffC6fmtMXvZ89
NtyksVSEb4qLllYi3O/xWmNLimIEvNdnF+PM1xwUbfylFhN2G+/lukBnhcEyuJJR
T+AS3pBgk0fsszVk0qC6tvF3jL2Mdg2QORRKm4dhA2iCG1TbFL5mQvy1pPLVE6Lw
SnQk/CC6aQrJJZZXqr/3sKhCb6PUoJ69nFSNdOoUrZaGaxitFyTNen+d7hgSbpEw
MDqCp0mof7dtuAS6KbJjSm6vYUek77rmY0Zp97b8Fuc+VXRfvaLrSlxg4dpc2lO+
ydNKV6uraZLl5gkVVVOIeSm4qY3Cb1Y1fjbeZDX4m2Rpr9ke2cgJ2m9Dvqu/YMp3
eXI3JGR3p53/6rQmM0pE5G/u4mPkxpd0o8aF8txsk2i1A97Ji8zaxC5gPyUBJnep
Kt/ie6jXdaDR/6zgjOfzS/H46SlkfAFWaM1OPpq2Wea3UBSYnUBwr4mFfcUqNs1U
E/TR0t0K0UzJPaUolNxylZPwihXDELW1zcqam5jbmnYimY8YLNIybMyCNKlZUduN
Sm0LptBya4NosFRzVW/ib04HEPlsuE/ITyFTTn1Mwykraaty10i3fq/xZZWYbpIL
F3t6I5gOB7ESspADOHf76sgg6sjBELLwYQlFXIbKwyqm8I7m+DTYd970a2DWBbF4
WtJ5vld0kEiKEoXoJkI2bXP1hLAoPdDyqwl0ShjYYQZWtpqwFY4lANPGlkOX1+/q
eFu36FoAuQ6ohKPGfcmRQzvZpGPfRVSqVFA/ZU5j6UnNUKtTr1xCMqN4KiYGk1l0
xTEgle76dO5gsHG0DiPdVDPW8wQS6Xsa/bqYcyyjb2vGJDit13fBj6jHJL9bpGLm
QB1r3Uuk7T7JFSzo3KkzEOmMDclajq+ctEqu9S3E4EeYCTPzL3lZE+DdPNEzCNN6
X8lD4tJj+FsoykDJBGppLmjFyeDGhmBMZQglWhwFNjVGEnAIWbu4kAVsMznbEvNp
+q5nudwY4w6ptcKJJQUZYEgM31BaEb1JF86MCd3eDOSNRMIxQfNuGcHN8tUrIZj3
dQcqQMeSc/YfgCznYgCLd7r0PliM7TFmRpWyuaQ/zrDs5agPP++VtHstSbWrZcGA
OLh6t95XPApX9+7ao3ro5+VlfW/URysARvfRf15gtC+7yNejU40iTYHK/JAHIXcV
ttSMnkT4X5i9JdjPEjk74JbESgqqPVTg+pE8ZzGMCHw4d2UfKGkORTPKvz2hIS5R
U0MyqsLpXiO4TAawdGwDDKtSjVm0TxmlnE/gLJQEfF4VuPzx95AvWpOjBlPcF2Oc
8FfTKmKBWJ7Jg50SQgL1YLr2ZzjRPzFHAcq8CJW+bwWjI8t14fMy/HH65sijQXja
KNi1OWtUWAiK1DAwvwtbN9sl4QvxdfMuOl07OH1GbRgOHIH3iJ3cZEeFTeNTLFN2
hGto69dRqydfbWkJYS3Ub9Kbntu3Az4H4kT98Wj0gQJSKZXTLX8GmGMlJXOrJHcI
2Xb6XDBM9SHxm1NM/NWcct8rDNO/+F5r/sF1YKuHMZJ0oA5JeLx5up3ihkh11Z3/
5aaVnrT6SK1hMrbu6cl9PtkxQNy0320+rnssCaD/3sf5LiaDeiC5U0qz+840wkAq
790lmhbTlOWy1nyAORz+9GN8yMf+fTIPsvfjgRlz3qePWtxpPdIxXtAcjTBEQfxI
B7qwpJWLcQX/vV0+b3z6xvgAz0/HeS6sjrnai2+iW2ylE6hTMbptWKmWc7GkmOEQ
ywC5R6BHT28zA8zf6WOa5TEI7C9zIQVnw3L4AhUPaeYvF2ZpwOJHRt6U9zfmbhFc
nzngzN7udVGtdSg4v4xWorFPrbvBKVx+pAhM6K8C5hmqxu8r5pdoc3kfiFhO5lyE
INVwpwmh8Goz5+s4nFCIQVQGoXtr6lmq7QygI4IDXeE1HV4H4UuQu248HBkL4dS2
x9DrSwpTw240OD2wL2JjNJVlNx+JwwvWFkIbHBDyX8UxNkiUfr64meFVwZ2rFPTl
FZot+BP5S6EFLLDpMZh7LnbZeJVvKXXLIOqeJsDsjMXaqx314lADUEt7nJpsDqkE
QM7FIfIlyx/ITI3iP1zGpVe0JZSJRveOARniLmhbJYjhLwuG1nSehJK8ZDMH68Cf
VGC2AXy7fuhH8f8oR1hOa8WM4DjteGR/VvGXxqu4RzwIegf+gffehLXKJ02ZlR5Y
fVhQStioFybb4rjVEttcUMS4E2K09IlLlsVimmGlfAoq2Ik9qRQcRH5PlUzS0WGJ
43rB7jgyRfh16hKx0ehQetNYlTjO++irTn3me744BMDLW9Bmh0wyxt7VgT1F1FOV
rnhoPBX80lDn0P3rHbqgwdVAy4aYT8UtduyKBqMzMw0nxXCgbYyFjsgE2eksA0eY
zdzXkIyck6g8eE5SQ9np2wVii4lWwWpJe//HkXS9VBlOxYiMfjuj3iaMW3Saej0R
vabG3Cqc8eeT7Z54Xbl6EPA0Q+lAyVVrLEpQjCLD8sItc524gHelFGGrcKIfD7H/
W/qgDvBV7KmKDkWXRgBHivlKD+I4VgqUNkd5O/eN6VyN9mvw/Ydsa8RNJpjGdRT+
MYsWvyebsFC8rq+4jnVQsBiWVwuR/J/DwMQvILBZpmY8eQN+IRdpbB25oZZuHKW2
XlcAHulGxRcrU/9jZk1To18BJEsFE6W7O6CWQ61fChYb7XzLpUvcoPqXDPInnS0/
YnCKGgOYerEi3c5Le+9QhOKOVu3Wgei774qBQ9TgcAKuR7/P0+ZPikXXg2Ya0R4v
PrIKgDdDvyRN0gKzdbjIpnfPREv5yk8pGQyXhsbo8tUsEJ/e8kpq8QRtSZXuPzMq
uvs7gvH9CHukbR00IFaLkoC5a3gb6oKokHaLv4kHs77t+3NyTZv5tKmumtPGNOyL
Gig8RKOPZoa7VD0X99lf/zNDVmKMOE3vE47CjoNhFqIHAf8j+oirpOaOh7iPj7Np
S8YDMg3j+hc4F9/0P1eRO8f/dd2QOD6qpbPwP3Le9ENlRfY12+OvGoJT44q3p9g8
e6QaM6pgnoUC6bxE8cxRtoxw+qesPR30/CMLxAtqaiYmna84/TUDPYHRNiQnQ54t
K6VFPMh+dCvnTqI397Rg+jCfBt+ab3t/X8erNlbR6UInEHkOySqCL2blO7X34U2/
hVlQP1AJuTF/7KAAmaaa/N7fusm3h69kYRy334j4B6GHRemzdYydLknBw/UiaPNk
4S7UStVSMezb0bm4VjA91/2K4PgZ8qWK+KsBJUWsy47F3b1s2peQY7o/b0b5mpFn
BODIBN7CsHs8MGRyuofSCOJs2dIWJBL+i7K7ioBHHg7rYvrsI9xaHvvF7gDMOI7s
/psJDA976Iu8MIKHhssrV7DoBdeSKF/xnz6MId0r647UfRvyxLMgbGFJKvMqXOrr
pKnI/pJMvISTYysTMsWc/f204Dj4cKN6KfTkoq4nxJHL6ypIhiO7bDU85AxvOEih
hRwtvICD3a9MRv8HPliPL7zS25cQsY52M8J1C3E62BlwoNFjVR+mcIRizaYHzCun
NKdrWMtMCo3h+yE77QLraCURBXE7+l3lw30ijJqOJxtMQ5oanKVefireza3fZSEC
dAM3lOZj7hhtZ/Xr+PAEcHAk9gUzaC+qCA7PBGcBzP9K7vKZIULWykxUwu6ilmbZ
KXK8uvCAk83jU/kLgAv30XVqm2D01kp/IRRT/n+zchcPnxmapxPqiiviVnd5ZGXD
D8lap5+C3ijlp9D6E0ALZjboV88ZucAnhobD+BBXnZp+7NpCL8Z1ZDhpIVh/4kpv
wNdhkuGf0dJ4AURav865G5XgDMwINhn4CAvNCa06PByfbJaEiWaxFykfxuDPQybA
8ofk1qe3Ag5z4irmlyyJQ8CBpSLscPlZ2y3fu0M0JOgncKGh5sJaErwI7VRGETNx
mNLT24xkHTHxaOgwWUt2WkbXENPSN3kJ7BHH8gB2DqWmkFlTPEavdWChbiuVHOfj
YENePZHkZlKNwBNuc0r6vUn1QiaQvHZCkOaEsMmRkyzGj80sCjDac+qUePcsMFi7
h80CYBbdeowggQilRqUEtxLoPI/SUjAz83aRe+dA0X0xk9jSBKlYp/P7YcEaqukz
zDF/nRQT0J6lSgY0xSfpPZ0hDfwwkcmitfqQge3TAx2S4cH5oxiGpRCrjJfvB0hd
6sIZYEShzXm6FwXzXhZVXLn6paP5TZIoSidW94DVZHi+4hq4n3ULfnGR/vHywT3R
2VcuF7cAVZ5cc+wDN2t2GFJpYqoZJE6L33Y/QXI9T8h50CL7Hb6AlLZGvSXXH15k
hINTV6WDi14XsgI41D2Q8cDaH38vp0qiHcSotwk8qZCntw1yIUsOJ7lmV3wCDv9z
ZJDo/+pp1DF7pmRxFV598RCALuMR2JoMxZnmghFam5qye278mvlpRAaBjgbtWfz+
ou6Seq11An6nXBiVDW91uMu9KSlg0UCOG4sohrdWpaBda5D54vkrLB6C4ysRZWnv
MzVpE79gfyaNI/IU93z5YUjVnvkSOJufkXD9SYuP5quCBbmPXlKkp+sS74Hsy6DK
1ZI5izzMfap5sC2c3FtDeorD4L+Uzhiusg5SkfkRD4IfhhlTEgTQm5bYeW23Tw15
uchxcc30fzTiB/UdMr8M2vGMaIWpRVL4CuCmT8cJcASgyst411pYhGl8PZ2YmkEo
YzJgPq3FsLTJkLmup8mIB2RxRySubkXnjVPquNoaQEmDXYT17Is/iupftfcQTf/A
oAFtu7t+ifyrQfNkC/pLrkmM9bsE2Fw9yp2C1UkKEUUZlFvVT2E31/6bdnczg1qu
aG8ZKoFTFDU9/0VQhoemjZPPMPFBIpfPwTsgwXSduBudvGpY/LNLSme0uf518lDb
4cSsF+ZRLa1h9x9b+d7Q9Uyeda8v30W3R0qc2L8d/fOvuBwEdfMdkVdbqrh1yTR8
Z78KTqldQtmsJfqgIXmtmQgUMvBjxIvfORALNDPR5D3A79OIFlzJLBluovvRWOsf
yj9tiKxGozfp0Us52cW2CHxsCN5ZO7lUPAsW9368Jn7rTAiER/hKL5MfQpJd5vTY
cdfROPuA6oL2ldHX8FIv9rlx3Ccu4mEE0trruZcRtkY5zkZ22tuXy8lvDiEglytp
xAkZty1hV7cVCHZdfTYRakXDAOfsiHuk5blYm7Yy9k8Yw6ZSflWHUg13gNvUr4cy
202gvmUTQFe8kls/ZbkdeKW0UcPxoOsT1M0r6FPPEEAhoXxBy9Fp6nNfopu3agQT
gj3OkLEL47/G3cBn306K6aNMYouK8cq0nO+rXoLk6l64FIm/BgNiomcxVm0k0scA
3aDMCEopg/Lo3Hiu6CA/ZYp8pDGCn/eEQOL1NWjEvHpQFXualCBaxJO/eWLGG1NL
u/ozbvHmESMiLjVpQ5Yi8z8gevvVPxD917SBzkM0YpJqpxWf9oW1SewjcCJCBU71
+lczy+aza9XopjnG7Gt7DGeHgJkZtFTG6B0ebQ/NyFiAuYR/aPDXSSz7her3jidB
QUuBMFJTAQpCcQopWIl3VMGfXdr3tPMnuQ5VpVDwLO3fd7gGFi5vrXKcAw3RfkFr
PXj+S4haVy5+p2dnWGEPZOkICylnNY6ZJiTwplEJMl0QXTHlncdUj3oAuAzriQTx
Iqp3D3JkbUUFl7OjSy8D5CpXpP4MVZr4SJuHWmbxhRBEcn/FWIpat4wzlfcipgFF
FlTP4C3SYQkY22y7sFwZYClWLtN+kTA0iUz23YaSy4kLs6mBOy7Ff+PjmnhIxGEQ
E2TzmsD92w6mRce3G1q1+y3d6VCY21Mlv6dDOTClrSur9YvdwsuTz/OTKvVJpWIJ
A/ppPbpaQ2k4O4IYUF1IzVcP2iGYGsXuqA7DHGKnJN9hzKRf2D0VuGEOKPxFPyFf
e19G078VvFDWwgKBN6KK+o3wpX+sq/LxatY3dBloIi1xq4bVFAyl0i0s8BwzIryG
72o/j+bTOs/pO4CBsj9kOSMCq3g4f4dv+pDhGRuBDnrb4Iz4yOmwXs8EvkZ8uf9W
1fiCVSVNr1Mbj/k9bNxdSK7WkT9hBv4mdjV5JCCZio2jDSpIHzLU7lel3HoJvB47
HMF40xa7pqSEdhbHD7Qps2Y83QFKEQtUVOFw6ZMi+2tJ1yaBaA7lrMYI/sFbp14J
f/rMUumzkmQOWHefmWpLV1w3ciucHlsQIHRHeFLxYcFyo34cGFWffrE2g9mxkVhQ
0/lwT0eU3p8PujobYavEAmNTwpNS7Agvas6H28SglSTXYT2RWeWwhvQxfRvsNZSP
f8txYmGnu2GKT5FTFi4jAdd4kEetDGprPK3U86+HVD9byEE5vdMJJ9mhRd3Y89uT
D0tGxjpy2PtmVErAizmEAGk5QGT+uNGfEKmV+NYNX7jD/JfOjG1L/6NpsvDezIoz
vi2FQz46Bh5F+TNbyOmMJ67KXjID/JpkG+1K4lUFeWGJnVh4InBdQ9fW/WYP3Ox7
WMnYy+FWllYnM4umJiB3dZX01tbzSkfOk728oQq0ouIm6FDXZun/Ot0HF34O18/z
e0rtF4UY70irYkyJ9bINybVtlRTq+8ITcAuckJ2GIQ7cEIbW+pzFHEeZUftdaHQd
Pevev3uXhohSQX2fc6vpjih3YmtuZMHo4TkAPJcVL8LDUAtGMX5biYm3FUMZBY3W
kTuo4KCeVtylpyoVqJhmoB/3AhjG1OKniMak454Xy6ddd8PocM3hTej7GZH4tloy
VgL8zza7e7sd/LO7giQ7BlvHvl3/q1oWk/LqxAXGphbQwvGSIEHO00e027Ib+Hxb
WrUnpB0Aws1kDU6v4RaqNLStArNjpkL88MtIV66D/fpUXPulmzp5kdCVMljxYPr4
c6lT28UH0pgbTMP9Q/qHdyTwd/z3pM+Wwxe1xErv/OCitkxuKJWTBTD2X6NW9wH2
SE8ZlmFeZ7TtQOs9GYY5oZMuhVxFbJfBAmclF+H4GK3sIgmRMsmLy30Z5a8TRO4A
rZxr29JH3Dc58Ox8Z+RvgabUQXLrnc7h/7En64j+FYtXt1IvsrTg0qeDtyYcVjxW
Zty8Rvj36zSHDWK3KXTY2uG3qTdsRSo4z927AsPCwQJs+Cnr+ugZVxnshWPv9lnG
uYnRPefkjhUR0EUnGSwh3SPnV4Lf1BW2D8yhpUfYF13mPGPvI66Hx8AVSBplUlFo
RPLt1dzMjjf+PhX/kzu6Ge8jZS2zCtgKA5ptR07MbfCD/C2AixUBkTuJeb11sa7k
WCMcLiO0r7UNPGFeR43Ix28omyTqwcobAD9DbO7mgArp2NrsslyUgHtRoTcydcUY
ZoHGlLI+z1PpUDt1o2PbXGpKptCX88WoqI4ghziLDUzIIZAH2ntfn9zqSJIRL6gj
oecgGOnjCenOArgY/xm0B+9SqBvQfXjk3ykmu4ic+1jug0TVHYLMLyr4TVIlxzXd
zxKM/FQU+8L2kW40kZ3y7HmLhmOJ916o+QckxmWIpEtGi7SPrvbGcyVmfalnPxqh
ok4FpBrOM8qBiFTgMeN47HeLslnVHT+UWg1HKPVhio/xc++rV3nttGCsP0haipXQ
WHO9rLMZZYIR7i7p3lZKKiG3THhNTt+fs/5GPdEYPJ6N5OSyemylFPI2FVuwYI8c
1rsRQVtGlWIRWQ2nzDBnEtvT7I25oCpLRYieL8cTFcIZkV4EUaf0PtUUrJfPl9mO
rvQcYPrD9mm5yab8QNvcDNqEsPV6m6bViTwrOQpbxOW2AFhro202Z7prEUgxqaav
PvSWZrR/G/zFbBGbhcrZJQdSe+apQqePB6RifiIvA9suZXZgClcVicCU78nzJRBH
dEHABNaPGD4mvf3gY71PfLqIjbE5XkxQcG6oXRgph0bi2/ymI/BGIA+oole5+PrF
HhCfrrnWHbb2Iz8rXyaDjuJoJiLdXzGC3irYKl6aorccgynDYsUS4Bl6Y3y/l7o1
bMz9RqKNFTWhBdVjDyWpPYfI0StZj9q4CNufHVWzPxy8I7JDkz2+FNDSLHIr8LXr
nzbOibMZdMjq6+WYQ3CKamM6KPMtgI0mewKVeJQNihr7XZ2MZKH7nTLUMxId5VM3
NGFfFJWplmw3a3VTjtHRWKyxPEuS8wswGaTtDahIQqExG+inxaMWJYhpNNyst5wr
1nLysaeT+LK50NrLj1EjocWwBMARtzLojwj+v2czH0gf7ZJZrjhjMuuwtp3y0Mv4
HQvP4TD08akwTNhmzpPtr0KTKE0ASAV2qjV5rtcmykrnFcguBJrwSXmh0APXpkHj
OJQvmpIwng0ITzxLyMF0S+RYeTixtbXt9uu/wjy7zRLXgEmVYY8AZbwcLHAb28/t
kCCpByjJHDgWAReY55vzs9wamJsrTWQz5O/v55DL4u68N9PyG6/i8lKOdL+GA1U7
ly3cyYVmSptQl9wgdNCa04pPujhjaFn2/e4hLua2D6nm5gOmWxF/FfkPAXamGlsK
8FRLmVHfAPvCsQ8vxLVWpcRLzFViTXbOKGN1TyoJz+ApiwV8GozkSJIJLT6SdXue
TgRRL6wj+c54ODjdqOqdK8y3p7L6PMhELgLzpKIg9VM/n3tyuUcq0r+EqjNV8jKY
bSEh1oGs3/IGK67Fw2pGerPTLItx5bHa0HG6mq/BdMK+KH3+8eIX/ZWJnVgF01w7
iKClD8VHI6pcI1clhr4vnPs8rB5ePxK1HkJxocHBiT2PCQ0PWMnPWMHB3VOgkGSw
QNPntiK4WZC8Co3TfWvfBsVw06X07BLy4MufaRLZttqxE6/hSyJ34+A4rCnb2+0O
LgE9hiKtKj8rAflTC0aq+JG/qubKuzFC10ln6xtIq1XkBtKq1At8uD+AQETjPtf4
J0IAOtc0+ibbYuLX+3rvvLH49kRnQLGnwv80w4iq021FSqeoSD9I0dAYZtZEkSIT
k/UmHvq2JgR5CVsjUSGFsuNIuBC1p72rSRPxHTgPbCTsjXtMhY9zMu1SfbPLHK72
xz69DLUdYteua4n6d1glMGkvLcdVR9UsjXQHFMpovItvIXlo4/0yr7bPw3HC69fD
bqW8iLzUrytzlPm/5qIpppL5L5uJEWvxa80UcLlVA2oHeKANnDD2Usz3wAlvM+Ev
Ui1Oqec1WajxnQLD3nF8q4YDae6jwe8AHQK8Mb86g1YB+ulJ6ooX7jBWgZRlJOuY
5UmBykneJx1lrLsxcOK1FM0ik6o+QodpKhHyWspUEFMOnB2lCJZEF6rryloVWlxx
9StXs/6bYGzPq31oFmhraCAlpK9k9vVnhQOLOSvFyiehrZtb/7UeOLV8j5JnZBg4
bejruxoeh5L26tH6JzTobF92kXyc/ujC8tqDIwTeFnHBrH7PSoIyJG4msoxLHZMJ
CjW3TiyJHQTs+QyziNUL3E71CkIqvwGbt6ZkEvSdPywFmqFzNlH0wcg8I0Q1Yz/x
XLg6mAlcv4o8NTGEOodaNGiYpvFIoK6reERgsFXxr1iHU8Z80hx2wOjEiUvsI838
3XQg7ANGTXkrVCpjZ8UnAmDjvZG06xRayNhdnBCgGxAYftnv00VesipAkOYaStuu
NofDN9LriDbX/imOLShekEe73wEo3R5ovhum9ALT7FDpCcz2L+deDx2wVv2bNUez
M+01INOeWxMVgrR0Lz9GhP82m5rjGJH3/20cTSHaJxktJWxCJbxG4ndRAqSpOJMa
DuPxOFt2nrqiR+HNKUEIGAgqovv+w8fWdF99529db+4vUp3RR3L28LqiPUxUL2Rg
YPwvy+NZEXDpAT+1kDH2GwPneSBr9Cp4TolAGhiWefD6UaXiR8h19mXsSFtPGGBH
JyGU4xCxcJBwF12KWqC5p2rjP4MW3wmF2Xp0jf3sH4FIbXv1za/D9OqKhZCSH9xE
kfREfsVVG4pA397F9JoiT9PhNqRUaY29o5rrqTl5KxsqjAcRiGWLzervVErLqRQY
KvO3269uHweJqn2ZOHNtGJEF6WaVK8vpjz/naIIdKh1bsyb2fWdETcFvRrZao+Lp
4L5UWAxN86VphmE0lA1WVPE/BhgAFZYpWEbD3V7z3H5RuAQ0ZaF61UPnwi5kwTsL
tUY39bKt0fC6zxb/DaW7keAiiOHCkbZRitA11DjdTKqHPy+j5SJvXAflnLbZxUbP
4v5JKWD4koO+aQJLOJYTYY/l9Mwgz11ZXM1oOOzh1VhE1cAVJnsdH8AJBmW3Wf52
K2tLqi/CKrqccsVOf1ESpHRSQhlEmilK+NdqOLm4La5CXodLWmBst+ybWW0mt57t
NsABWXB24BojW45WFwJzVbMMw25zujGaHwIvgAYck9vf+e0/Qcx/krvNn1kYRu9Z
DSrsU8spgxyUWP2qPwIjduHJsZxlg0LQtJcxkfLMYsjjQFw8Pi9YTcsm+p3fG+V9
fpp2MiQ+bxKMqKe2wvqlarTcJNQtYYIKPzhJUOyhbTPC+tdOLpNWJRsybS1YaIOk
24nRq2CWx+b6VPG7AML16zhLThR7ExZ+HD9zUO9qkYdK1zqlZUl2tHQzx4tsyQIG
7WL/M4W9YhJbltPxpil3OTflLHDfnieADPQuN8+zPO1ufdK1nth/ycoWDHeWKc2+
ICoGy8ksO9HdoXNXarvljYVybycHwrIiGiFhFfuPmsPv/nEFe4IZgs7thAH9vRGC
3NhrGzIjXzY0rMnxjqkcAR6EBLWNgQUL23kXuzUj/jQ/XfdU1RElp3VtWZECiESg
B/bkPS3LPBstoIvshX2qVsYC6/mp2S/gsV1AWBOr3lOT8zvrEHgCQJ7pBmSZHEY6
+oA9RjobjCalLGWEM4x0vjExDcaARbA82XanyemmFnOJfsYpDvFyoERZZbuEJR9W
x1rY1k4G/trKlV2IeEbRVf2qas3A+2a7gnBQQUwO4/6lm6xiw3nXrGfpyDZ3Kj6z
BOHUE7A+BseNmYyqMzyciSUhAWtfJWInfxuryHWVDmtbBnobxMmFbiWhqPzVjelH
AABx3k+UYWpe61r4ri5ApZEE+zoxMNcIIlKij7CVV/3nzmYH2Xr6aF2dtUzXQtXX
otYmc4KX64//8abUaN8Z1WY4Z4LMgTsclwRcdiHtxnIqL+udsIYZ6RILnm5H6+Vw
tyOl4F/iZei9+z6VS5zsAbtjkBKHRJOmfpjU7YcxgrfiV/h5DUnrvoKWOqHjf3pO
I8o0SxKYGJWD8KIAZtW+1VLAQVYvGuz8nwMmjuRMdDR15SItlbaiui2PyAGY697B
0P2cK9PcSH0qCIOoPnbEfgmcfDtiIPum+qeF9hCKzAY6xrmLn27NjYSvaKBXoeKB
6sUtCs/FWTzcwG4jdXbY0aX+LOuTSM2JxwmAf+LV0yRWUvOpTA3kDW4AdCKGRG3D
fRiJK5IEHzGzs8r/9/72zwFccc36H6my+rMASG4nD+2/JrkbhMoFWZF8+BEOzSc+
2YjAAckLgtycqaRCB8JIYlm8bFk03ToqK0YLAE9EgsnfhA2d20lzGYNZW44zv8+k
JbTBFEJx3mZ7OMnXpqt7HaJAHTFBrIddKwW/zJFo/ilE/oOs2LhsDzYnOxxhOGDL
85FlaQe9Ktek49lKakBZ2O8JMyWEWy9YKVH294GLQnYL6Lf4PV3aP5qjbGTHb8eC
bavsCBuC3GtPitwXvrwwd8ZpVUEryuCQcizovgQeyTi0tqekoncBMgZEeMhTw5E6
ewHdGe5UZNlV1Z5CxUrJM0QE1m0yvaIMnISqyeo6bCgx0KVzuAyH9BV7wOyHgBew
SHgxMpcvbzf367K40sgUbsH6lb8F8fuIQzbMrn4eHRVUrpFdrEXUArGmnzhi9nM6
9G/YXXqBzTgxjT5H09FCcoSsPSkIu5FMSrI+HJgG/gQGkUIPUFm8omepGfiSOEXk
3Ky5btJIPVaIAPod8Aph/ry1gLc1lE/qE6DyOcOcLE8rJkHQahXLLmXt6Q5UMv9s
P5vfYVNbGM0t5WBJdvxOt0OKp6noqQgDzKZbJynM3+G6ADlbVz0l+p9PTiUJc9ub
g2Z6qp2j0LacdTihhD5AdxwwUHUVBmueeRbXWR4Fzeudtg2DrXj3OtvNj1OejkSa
myZQXWceY4wqiuhEeD/VRxBUK++yTkbKBbXetR5o6/GbjDULY3rOK6W041mNQIVf
7LqZceQKrRAlLs63izUfAMZZzNKxA7lp8ABQN3lJDMuIkimR+mncnbzSCz1PKUYS
igASj+wQOtji1co/UHWNa9R5pGAYZDLKHbNk8b+fn7K2hHbnbbuITjltpSxZn9Y+
app6q/rDeVXTtd58/9uVygAdYul7r+1Ru+Z7DYO/nTZOBOra7tt82aUc+4hOVPWV
sSmPnVMmmjJ/V9UtV35ZvWSrHeuJIdn9umTPubiuZ1s/QClt5qYZExFIkb4HYcnJ
9hpPjkg7CYiBKIe0tesbiWaa62bA//4mTx9KRp4SpDI+3Y33J1f1fD9BsZPIy656
08ztIGhj2Rn6LgppPkXEQenq+IsPD2pNpSt2MjlC0zxosDrGnXhML52q0vX2dxZC
k7gdhzrSPvyDS2gn2y26hLRDngpZfb6kT45MMJhkdDxgJe9OyXjdBjE7zr02UyQt
owaGuQOnnchkZz0WkmjaZAg1xKKIzOT8L4Zr9+vvrKVDlnDBN+3irj4Md1vrB5Ty
QTpTPA9spDWZYKzsH8skm7pfFdzOE61qMatDiIGAjfiAZY85INIWcl76P1GoLYfK
KYGs41stEP7R1r/ZRotFmQ+uoEA5exVN+eUZ6M2qbUtzQbaZRtp4E1annspO1GDe
QKXSM5x5u+Evc+rr4YjITtiu06WVTJJg25LQn8L/Key1cgXukolrebcdXxIZ9aAh
hDT+VQkEzHJL3sDxkVOzKXgrLKsSzfM1r8eDmAPTK+97ENwAf7VGkXV3qrt9eOnK
eDb9JDM1XhWYpHY3vzwWNgZr8TpGjBGinGMLgZZ+T1C0LhSK/We3N6rMWcfJaEwf
HvlmJ/eDo8I/Ab7rsX3GLYAmtXXwbCNYWkULkcTzRmIc+OQz8U3TVJqTQkI4VHJm
aghAVf3eeapiuRko+nWjeAOofEYlbA0/rwQb3CC/65v1nlIp3ZCstePVjKV7dwmc
3Jp7so99/jsjIe7vZy+XVpFX4j38XrkWHxk/293RGe6ylWjuiAzsQ49CQXDloaig
j2YKkBERihhR/vUb56bmssjpWdnwuV2UGhD9xf2GctSQZiXXbasNw1867wlMF4GE
SbduFaArsfzboiqfZA3rg0Qb9Y4WgDPfl+2Ld7uZ604RyMkchD6poTbtmuvhAEyS
xbGoyfYw6bStme+0aARkNw2LIR6YSvH3BteTpw62SaZ2F7cQsG/RfYesLsl1Fm1m
0Dm/RsDCpfSYUiSopccYGmn7TYPLuWfP22WhI42H06I2A1kOOJOzG70UIjq4GOq3
B//FX6WIFCVoAWuPeiMc6HGYBW0uVuUEpvWm/WhmE9AvJyimX4+RkKSw0WQiZitk
m8y6o6saYJ0RqkPRXPkLQ3R0MYWzujL8d96y0YFAJbfRjMLOJ4qW0xPROpz7kg13
2yRLyWDmV2uLLNSMn/iTASwnvTMLsqMqrBZHocEhKA4ob5Ie9GMXOz2nEQeaIUYa
oLpLzcZuhCelg3UrBwGFiuGyjCFuOv+vbxvJdB/4KGQUigXtoY83vrQ7jh69phh3
CDuVfsKwWeUZ+wdXm22lAs0otlVVhiwMmJiU9fNQb+LZKyCUqf9eNg+Cp0WPVnPd
6tWhrRSTSw4wnFoD5+nwPcXtzDpBCyvo/0iePp+yt8zTnuuov2pZCShzGfHM85U1
uAcHKrq+nlSqyRUK/AWav9OmUepx04D2GhJDXvPnlt3maArQGEHfvEwEhM8ZaYXs
wI4A7sehWoNo86tBAMVRPhuNrK++teSYaXMP4tupwCKF7M1xxYOLijG4D87Xxu+k
LXGzB4FBj64uyBJNM4uwwXGGJ7Z8E4zcAY8pWuD0yQCJLbepA+KEP5M9S0g/o7aP
wgM//MxNNaf4RE2gtlo9DHofjD3J8OGAJOipAiICll1PiJzsv27N1JC14KWiUnVC
q/5TaUgrFrLnxaQBh6vYFjdAbjnTX7xu/tgB2ZEI+yIPdHxX9PflJRWB2DgnRvOv
1Cv3bBcTq9ni83B1z8fGJ5v+ZgRSbbdJtyCdPnD1ku5ozk501sNYKT+oHHJeSQYB
7lPDaAhSmhIuW30D1YS//O8ZdzjfUN+akAukWW4aupmbVsqIXSvTzkasILotFO/1
8LGS9I1njQ1HLqoLh6Wig5Qk49TWnELIRlUS7YjbvK796jFtiWNrY+aetdWXGC0g
o9FVIeYUT4BtSRy560i+VcwjHS3NZC5JyDg3TYsBiALa0VH6bEAMBHiR6iTrsN8f
ecDrE7sW1Gd9YiUnC0aBhZKFaNbUs5nLW3vaTRS4TefozOItIhKw6Im4gSUZ2K+G
1+jEWF38YjoBkLibRE73iXbOrqlzW0802nSRqR0VZ0uJCkoYlyrb6o6nzawHxp+x
WdBBO7ej9IoHHPAl1uXQUMB72McLYS9hD5/Hl2RWlpyEEVeCalmQnhA46AZoULiE
0bf0GW5QlXdKiyyBZ6LCGq14sN6FcXLiSIMzsNfnV589TDW2Ou7Ojevn16mI5DlV
o2FiHilQDN3lujJLiDyR1vGYQinwMN6awYHtJfx/CfdmYmrnyeTqqqJvQihhuc73
ZVekCzAGEQEtjB6BJIhg8pQ0dh4tdtDWoP091/FGePot3o+GE/CCgIWJ2MsiKFUd
jtp+6uafovITkJ0Xigoi3zTSUjEEJW2D5rJxM9qtqDP9NGJmqUx2nQJ4AtJqa8Tl
4wIGoDbS3OLgXZtv7P/zkf9enYQv6EAMZ89OSovgbP3YMhNSmFx17z9B5UlssnWs
tlzTPNpj8dnxjz3AVLyaiYTi/J8OrjYY+JEDax2VKNJ0UBW0v4FB3/9ZrqKGvTDV
FtBme1weEgpE6txWhDTKN+lSmF8AsdAH9NqSRRpFelyQtsxV3dfPiloEWudFV3iB
TXiuRTskDa6TaiS8AAv9C6/hlDy1/R3twlfOoGjuM52qcT1PzfMf5dVkaCsoaaan
+2n+CVmGksidXx0q5imY50k2X0HdsJpscIvfI2oH1ETAVm9Zy9rv822Gxc8nE/uh
aZTHEAOKrvvicCeXFXybz3/3yFznEwlVQtFOkl9OsBedBojLfW4jtL9FN67YCsvS
CXgXEc7w0bqxQIfIHA7tGD/KK0ZdqoNGmnH2Nh4Gl1fBRb/mnbHntfUI7fnXe3Eu
bGgxVKEffUId96X7CXMuNO90CrLNbOIg7A3RZJrKKkUe6hZikPC7NSZo8cLXTEpK
Gghq8QkphtazUO1ZHnbVo+xhCvcOugYNdkZW6RkSwpiV4tA1Tm07c7bUw1pUeZd5
JIzCGTKeyCzAw+JDE4qFTC57ZRvT+RHq/bRpg5/AwqlsrsYH7a2b8NrtogJ87Zza
lxHOG0Cudf+Q3A9B3Nvg5lXLquPER4yWhIKOOw1WNPK0MGquS69BoxH1mZfqa+OG
e3Ry7hWelHsdQXTeKcwXX9loaLxUbQcwptk9Ff7PUyjYv4jJ7hsr/Oylrgw2G4dt
vmSXt5sOCGaI0BzDNyYXpc1HRSzE9mxk9hhFhlvLgUtvcsg7hypuMK6WQ9zCHywU
ouKxyuq7rQ/nX5PI5qa53tzuZkjIch6eMinjM+Uj0ilSx3GlZYrOIsHcDGTU0JKM
OAhh7Nx+Hkrz+6VpbRx7FCRrqJ6kUTxYPN2PD8ahkpUinkTy67Q2C6KjdqKO62G8
KFls1dZXIGc6HwAO8scxv4UJ+QdY5QDEQmQEhZ9VkWgNY29Gk2HsvTWbxA4a6C7+
7Hx7Mv7Ryp7ZV+Xh8/e2ofzhXRCNk0MrGFgyjIiFloDfprbcfwlGTKPy/WOU/Wps
6Pv32T/eHtkN5aGuO5qrR/UgtvsSloAjNoJd4g9WjftQ6t3dU4MIpRT4gjbUSRB9
f0RTEktFtdfINt9iyd52jJn84OU2iImXSYKXjPeQhxG9w7nBjI8vtgfhSMfzC/sM
sTPW/1L5796PHUL+77AGzPPaj+FEJKou0To2z4NGh/+gRUZg/H/j4mFEc3eZRyxX
tuYSzFR7DhC6u8LjGx/uOnXHbq7I4P55LuW9KbCrGNqWeQXbz8hJTLi6n8ktDUTQ
rP6MYmUsDtTsd95wx05UMqnJ+7HR4f4hl7c+yWzOG95+YQbj782tjiJ2n7LRzc4Q
zoqZ9uHWYOZEpBxQOb5D+C/uYFKlFHiiEdXYc51USzpbYPDcZGH/s3YBymcl0Sdk
Tv5hkIalUlNSrf+Dp7pVrnvnlyQRrSBMjDj9YlPZCVg7XSQrY+TBJ+03L04pPGd/
b7xmccJR3SjrRwnyRGHMt13+hZT4LJUPDWWNPGfGbjJkoMGoJw0LxOTrJMX+SM6+
OCP3SoQINskKKnIW4lVwr66Bn7FsSJUkAYapTHP747r0vqbguCQyEbA2fuVsKmit
91r3zsh2MagQlGOzRpBziQfC60oW/hki5m617Z01INPYVwKretET4es8OGghUfgu
6U24uiK3KFrnrW5wTQK+Lp1ptXHgAV3lzGgTAkpiQgsqcTypxUdi4vjhd8dfPsDJ
OHBQLj4F97ofv1T8bEMwcHst3q282R360biGyB/hhT9Y/DMn7oACtNsesJIMAfeM
uU2oN+ID5mXm2i0Qw13n1WqOHtGlNiKWZKgOteT3hhLp8WUSE+fgWX+Ohf9WRAq0
+NnN89/gjTlawaiOrY3AdUbsgXOQJr7R5eqDr2DnuOqV+kFGXz0hsrufuBzAjC/q
WMzlsxCGwbEMeFDIrdoPDjTR8+0NSQ8xg92vz/Wv29ZTPAb/so9EzweNJ3957uok
lWubsawf7vdhyOi9HJvuuo8i3G1Ik83EFVVg+el6d2j5oM0pETQuXY20YtrDqqwL
d0HTaUiv+A+W/2LqhX+ChMR+5Spkb8u+G1TRAIOiROOro6RnCa2Tpdm2PUkWaMWD
aV+YGn5YedUlbUp2Ez+06gWDGj9/pkFzvRqrdjJiKHzjz29MEdLLrhPKDQP2WeLY
SqN+bWnRkEOnrZ5Qtl/1krdx42ZRJ846wVXlmYlE1p/B7TjMKFn66ZW5gYH8U8/B
pQD2C2zm21Twrr5jv54RF9l8ZhWDyGEXbQASC96OlrjwdPYP2/SO0swn0vvhFWwP
sVgAszEmebb/jpyizNXVbiOjefxSVEFiS+0t1Uh5VIdsRYncpmz/J6GeNSt6CPxV
VvZRO6RATAQizyeuM3/HqMK/M1upYgr9OML6ESNM++4ld4oJQIzjt2ygqJsucdko
kvSr1Wnyc5NDIynYF92qFxXYnsAtLTM3OmIRV4GEPTfx8k/wt73Lrivze1LIrdR7
ZZ5AsNXTX+OyQ1QMqUdrncCOZm3wuMAn4WT2wBYMol1XxRrfCb3Uu+Nlk94kK6Mo
js+HuiG/y2QocZ8Y6l6vq4p7cShsQZOoMD3X3v03bxZ87Zq4TAbSoIBNgG/vvUVz
Y7QvhAA5GisTm6ZIwfPu4G8ZjQQG8QWpxxWnFN8DKQNCuECT0vE+irt+cLy/Ui3C
Ag+Z3n7sDZMCtEwwVHlv5PBuzF+9UsHOL8Em/7T2fpdToxlAF2P5mR7mbwc5jpU5
lo1MeN4Dob2QkkSOF1eSeIqQGwjWVbi6W44QYdqdTV14OYWdLHHAzMADMqZY9Umv
BSl4OrWHD0hCzINaXeIinypMFIEK/+drAWedIZKUd3A2WQIWLgm6AKea764vDdL5
17rfzoJ0fjghfBrgb/58jgluTek3Lx3p/gsLXddsoTkl1AYIjxbioVATvjF03oc5
bXajHb3vE+zbhsluFKMkYX/FyFJo+bnMcITeE40cbUUT6a1REjF79Tn7+C9Ik//6
18EhuX+X80LP7sZj0RqjyV7GV3ayTre50blQ/f4Fgl2JCPTajeSI1s+w/2edqzkU
nGJB+mwo5VDdPNMU29uUX43sXsCj2DTGSU4vML3sM9y600a7IGwGEsFzV6ioHx4O
xbCMuZRL9qhejEvjkfTw7r1+xyMNb2nXh9uJKH+KJ7vieON5AQxqPzqvDkBjD7jz
Kia/DYUBlBd9op4RWxAGNuET00pPcgpb6QUqItK8oll9h5D4aAVpdvqJf5td80ml
8PSaaZpWmi9IJPW3fZTUuqOgtXieCWettM9NUIbZXgOVTiFyGFW5QZbkUsuz0zKi
VfpvVPfoc9BvTy76Uupz6iUnoh7WFr6h/ssSp+O58UetLtkeYDZa4kHYbYoeEN0e
FVE9d25D9AP6+LcMMzmFHDbbYVJhVaPNc6rVYAe7sG7YggkhtYY9fXwhqI9hoaEm
Gl19ZLDojM/nlMVaIdU82uPJIRAnQAcOzJ78up904R/1vLhMDmqECZfS9zz00EPs
+E0h5lS2xGyo4YzHYXhriU4ySjWpb62aZfyTSt9KIzWOG3UinTJoBuAZTwm3Wer1
WxZ58hN5f7XTjoV87YxGrlc65ES+aSW12bcJHMSWS8DZhj4Z+1UD/Zk5QJANofcO
yZ47RPKEs+VGWwUx5xOMl/lelRWFHJLoQ3V46jJ6b5pTNGtFvIa0ll022jzWp8cF
dIlIkSSQOu6716HQx85ffihbHzRKdVgvB/BM0weoEvEEk+Mz7YqBd7fAlkkXr5/z
yV9NVVdGJ5zovW+Hr9lBYQYsmeHQAqDy0JtfEEFeFMNhKeV/WWLMvAJr4TTgqM91
IxnVX2HwgapRXjpR8KSJ+i63Z7ORGIiPuEniHU+0zXlO2ifzi1pgbag25SnllhyQ
swYTPtGLFvHte/DnesPcjHW7E6ViTLeBZPwdB6nsdDdINjHNqntKVs0kZjbRuVbP
JSsu7sJzlFZ08q2ByEsHPJ/UZ/4z0MGMEH2nM/LDNi9ESwBPe5vx36MYISDA7IKh
YxMQC3dACSektaXKAVpDF3/feZPeozGChIPktB0zcE4t8zphuQ+SgI594TI1Dx2L
4QdK1RWV7dzSmvPm1v8kz+FXz3qEOPPncPyXE0sit2om40fIGz08spw4Bto/L2zD
LsL10Axlu3UGT5atmD1l7cf+8DTGhtSlKpoE+a7Cx+eo6OUYF/XzUW8BIeY9yrqs
FOXSFej4ZjdbdH7vECuhA8+Xnle4S7hELLVbgYY40baSdz3coIEBqlVi1MF5aWLE
8L2ZWywseDnbuT5T9mzRAnHGrcDgB2gYJo919zeg4Zi1v7Pew2NGeOUQqEUOx1da
1UAq2dsgLGLMCgzwJe3UzWsVuzuG8XBh2nE84j4ZVixxiFZC2UicOJDvhcYtkNLw
lw325a7bnz4TC5YqZIwkx08lsxwFVF+wJNF+k/aqr4ABSZOrHrXZco9zWT4nZLOA
fZAE9fO3xoXpSMfXuAyOY33QV6rAkLDjI0u8UVkyNTxNRSx3+K7sKaEhKwJfCI9d
7xx0JMN2F2yuk3f7d4kn5FXF9amjc7olvqvrgf9NyedLXZOFm3YFgnLBLb5UPLvR
7vq+zoNB5PHPLKspksg+J09W+kFe3MVdqCEUkr9xYthFXAGt6MKhH8bu5Zk+UP2/
2nL1ymeB2AfY6hUvY9np/1o5MJoyq+xblrFMPP8QBNYFr8IdC57w8XdXzLA21jLt
MvyL1fvphy+64e1f1AjUAV9ywtJKAnF16iM3r47I0sHwiE/qbou0qf2lewpKDhJg
jOBED58EpmJ+9tTHzss3NR4ILduwRW8783p/shEnFeyuGHiuNh4SM77SwhaO+rvS
gVmwoamrChXPcRot4EblrgJYUvPDCRIuIMCsPRLGMIrk/ZcueOiE0ViC9Ewsu79v
Wq+XkUlsXPPQFF99VqXkqr4oDJzSLcc4e5dycldwS4lio4YncUn65cWpiJL92JP0
uLxwVFUFfpxWoI1cpkvTAa3B7i7r5jA0kvyYNjxWSm15NYevOF5bLdwpXUupavAV
O6D/cMhLIxxdESufhixpjtTTPUxM0lHSBDWCUU2kAR5KGakV+7CtYHuIODxGUo50
7W40kmZGntwNIsAuYZFikUPfSHYsYPH74KYnEdKybpFLslUmEpRZQzT1WeIfnSnB
KVz3kAtub6QK7A9CLmeASbpSjQnju9pUhrtYCELFcH4sUjKQdoIjSbny2L2M8u0O
hfidX/V4rtQ3HQbQ7xo+J9YbqogMKW++OFFuINmDOHuGjSsfS5pNYTDN223XsHpA
61wgtRxpmg2UO82Abs8DzODb820QzxEoAM/5Yb992z8MmKff+ZtMd+2hBUf7VFxX
XfW4vuI4Nt1SlAp1vT0ms8jt3TYppbGg2evzxauyOsI0ZT2J50CyUZ8FZxoB2CFY
jKgblg1lmGX4EQopgWDbvuW3t/tgEhMCTiaHu18PI4SWWOMhvQ4XFyW66mvZR6oM
AbCPwHzvpG29OjB8YvdB1j/t4lGM2qq+mHqzD8uD8oWwQIG6Zb6OL0fxn46vGLzq
N2lQbMe4afBqNLiN0P8ZEAwrldC2s+FWWrrfC+rD9BvjCp4rqHuZYfKSorkWaZ10
IYi+v0LFWGW4169RGMINsf3YL0TDNdhmK6gwzbOUfj7lfJDgfoWoItJUr+lAPlcN
chWEKNJ6Ybm7K5ZU6hs69Ww6XrQKOsOWYnEzUEV1P5IDjWBw9vLRdEdOUq2lGl7J
Iwgd6vqMK2HbKKd/hzt0zV72oTxgUQFbquINohfQP4WQBwAH15P9nXt0pHBfwalf
28cVUjWaxhpPTAMhuEmmO8C8adkRrTCYBXVhV8jk/70lp9WC6thQoOOyak6KqehR
m8CjV421TXU7yzRifNYHfKzetYkdcRhNgocJgT7pB1M37sWKVY/TtE9j0PIO2auQ
8ngypSv2R9NiGuvn1GwcfoOYfgYpQQS3BOU2xcsCbXToTAiHQJ71kPtDkas7Jxft
nx06OBwSRJsP0OeIKXJrJCsNxBpcPVs71ZnL5hAVi71HNpddWdF+0zWli1AFhcFl
SA12bXzD4MuxGx1pyyvBeq2abUttt4rgoKKM0YEOUwzXoskJxZRZCpVuRDDe90C+
jedAxK6/9B/KMIDgQHWFyJxlZsOagCO7czcpDC7/RNi2nuT+86nkIH6qSTntBW5H
4k3v8EDjoHtf/RVaak8hXghy/1Zxl8jGWOpMsEqCJkuzQH39CMgRPpyDKN2THKGV
2C1ckV7+Gr1IlsqwQzOIJ7O/DsdF5BmOZkqzE50gW2c1wbpxhGjP8NlRUQkO0g8r
+QJ47RjUrmSY0Gf2eq3eTYCt0ck8k8zsR7sS9s0yFt79meCFBh8muVwQFScPcRoQ
Y32YCEm3NhtFao1qoehD+Dr9V451nHVIrgi+HTnmd3n3bd7loW1Pd/M2mizN64wB
rpOK2qkpuIvx0cZ+LfbM64keoJDB8NkowfOzoCqXK8PwipNNtDti9V05M2tV2FPE
JG278qALJHQS07TfSPzm7HkwQHOQSC/TVmVHiW5K9LTilzwVf2aHXqCWj/GVgnJ4
bMVg4eHrury7JUYw1al1DzSla/psoqY5yyfSyVVMJRnSxyzx+Am42D238f+p+9tO
oqcj0ljvfd06SG67q0HwaBp00nurt5p0zuWHRTpZ4C8czBIJ3EhGDITbbPp6maNf
JOZuipVe8Myek8SePCXptvz5TyUadlcaKVlkC0q1vob8ws+aTRmzEDJtBLng4x9d
DcKfO4E9EdTWSTPJl7+3dD+1dT1H4C9ZTlBV99Z6oAc/pMlhm/3wk2A6N3Qp/4y2
n6H4oHDhPijLOjTgy02q9Jfp8Fh5YXWoAsNnmEWl395HQ27/tgNcdPt7PIyaKzYT
QeAvidXCVT3l0bBTKA70NkcI+U4OpSSSk8ThXib4stTu7lNqZW8pV2/VW4fEjyt8
a1tiPnSxP9iw5YCn4SfCyWYJwtWB1pImABwvAemFMDkHCaoO9BlABhVu63qqhFL8
D4l6f23GcM0RDUD3TQN69SedMPDcirhT73Lw5v9lPWVWgT/C/bxyCymqm0WBsU5G
Tt/Faa1vBjHR1I9Gynpi7uQjCF/7YS5Q8UjkuGYbxZ2ph0XG/eUFB2y1jLDtDxZZ
LZVmEpglalNN4Zjb7PtAekVi/W8D7tGA2tMD27869qnKtfF1xw07MC4gw/WHIpR4
gOAzvHU1QN1UsOyri12dDsh0PqY64eMrxzevT5bKN+PWZDkoULDuyzsCxHESAz0d
ddAQPV+YMn12WproMI6BGqvcHgeYOmx6PBsKhmXiXjIIlIzLw6BpyeQGeR/zRxRW
qOKw7zFdr+59EiVspxBA5jOlHx3mdB1oqs9bYaCJ2InLHEZx43qFBiG2MF6n5PJC
QyHvTfoBC1BhlGmpgqTdUytgEF80hnqoEAQ2yAWIG3idBWscSBBPHcODuGwnEjFp
7qXtHa5Y7zgCdMCDt2uHeXf8Q3f6otJU9ldlMYAkolvkjYv7KAM+6XxmLtSAz9tD
+FtCf8ABrUATji0QNnJnjkKaWvz7a16aASEVz87G2QSlN/cKQdkVhx90CMNNBWMu
rhSXxMN9g7SegoBhN5sh1mBLEP5/HfLCzuWZhYvQZl1jQLMhPBySAaYPPYC2A8xK
pZ2BSz8ztqPkRfSI7WauoctWqafaS+seOxvdIgc3CSjkxLCopPGT8AJijy2qlhIO
Ml6tkwQgtiR/PibDfIL0I6tBwNnw8PXOesK+s3/bltwBIjkyt30iVqC+2V3y+kNZ
PBIm4CO85o/u7PHLOQxmAHM70dLe6AbpZjB8Z+6cJqRqAR3gF+ZoScGLOCYnLljo
bXwS1ptgAx8St6gMtdDArdjzGoo46B28ezgt6/sFs7n/h0MNRdOULpynYFrPgHm7
9p7ic86aGXLcSFbVlpo4+fD3BG0MtjWTj0qS/IbUny8s6gG/WnWlRw+IGeremFKp
QKt3s/v+ACQVbSDEldfPXYf2FzgjwuDybdl+UX7sSKJ1ocpmANitYI3WSvDrmJhe
O1H8WUN/74hOF6DHre8uMTSS0D7tAO1u5+7aIxf/aVGczEJY9/wGXmBXPi+Fjp+U
jq+/F2saBwalBAdNxWrbrSW07ORTbCdw5gHSgUj/f86tPEPtMfL9KYhvuDwXPAY0
QY+xP8T4jlq9658xF5mdxnt1FbuNl9au5dCqTBM0ScXV9e4qpHwmbl7D5Te4CGYR
oW9YaorTUzAUuWVyd970mY1dJGfv/AXmXT6Xd/WHTHa57Ajb+AMIm97d9WT8cExv
ljDnH6O8tReKCJbDI21lDfje2iOSt7VCvdgaqboarTEsC9TKQMGMtpYnkkJjyD42
Zba9lYkOExAbIkOoYX/AHmlfSkdNpkn7jgcS+MNqGRTAv5vNnOaa9QBDNDpauHxP
ohgIiyQ2LopCImYfehNxEG5kimyYB8nyp16r87oA/wz02rrK9V1skp2Bg6aYqrxo
CA1CdbSmj5T0QXDRGhYvM+dWXUXMYHhEWBdsPgHF2nHLBDo3OVGYeuSIUhVu0x2H
0WREdllyZdjnJWFvXVD2DOFDHmwcPTcEeagxIZAm2lRkagd/HAV5VFitNPExOfFD
NvalFcRjokx6Sv3Pq/wD2EnVckVrN0lAzVjWVXetCphi1kxC+P4HeLsfrZsecnl3
Ck5FBVwk4ihbxtv81E6uhOkWh1rJkKwrAUqoB+Pz+C5W92V+l9S9uO5ijwm7fdJL
jEoysoEoUtEB5sf6vL09XBvMWH/roydcclMG0LhD2EPLYwzbjAeaxYbExh1M5jnt
Z4SPi99cDOlIRZG0oZ0mRbD00NUD6s2pFlGEKOIa7J4WRIhyNGJDsoheeTv57BCZ
u8H+y0WbuN0II/rL41AVmAXRZqHCeLXDwTLMERrhMNL79GdACqhS9TgXmKTxMxKx
+ewftcPPUx2uunqdpMSVs3NesV+z5SNGQv+5AWYA70QWYfcvECKmRYXvZwU+fP9m
ORvELxFDyAJk+yPAj+k9sZokCpHtkaoyIFu804u5SJm6KGH0F1RBrLL/HYF6hQZW
RZIQLz4I+ECUaJ2rk2mD094zFIMn3aVt7ScCa7dyDry6s12HzplpVR0zaSw6teT2
tD9ksa10dsuCMnPp/mnrFsah+I23gRPdZDzaBqdMrz8JN2wWq7W09ZxwDtLbaTaG
GovmOddhDUbvtPGUMXJ9l65TBrjU5KwUqv6i9G8S1jEc3ZiW2vaxcQWNDFeg8gxH
wa4MTpcvWutrywpB47Ep/OtiZGDLnEVTQxgRtWqHczeLsfy1UoB72lule7EIexfP
JwAPFGZr8d2EkTuYtMTlB5Ka4DYAc5U6xSV/DmqY+maaVAY0Q+1yHTAaTJjPsbek
RWEZMEYlvt1PVkCnz5nBmqkbx5WqQ0V2hBuX3lmJ1fmAKgbqIzsE5rukvCOf9esS
Mh4kBgB44gpRG5k8a30t5YGzmT4hYd60XtNftCDL6/kyNQdScLhJ6tOp8bMJnjxp
/pYlTvAHr1kfaGK46o8rXNJDCp/kTqCD1HEju4MzQO59JhoaZSw2jlHogzm4hmAN
rJAJkmDF5NZCBhYDe0mNEptdWWLhnn8ctQ2B1opXeOpMW/6JupneTurrT7Y9FZdc
2lSvy0Rsdxq6A3HfA5QOSCSz0LhleDsdJCf6fSFs8FLj9f7vDnC4TcgNXenTphnu
MWBZOh97PcjadgazY6Jf9MqzV95JJK3WpLKXrGXMGzjoWdUZNxCJFPTLiNXpQ1aR
23Hw81lFehdsK2YAmH3Fe9RZdjcAyQW0CL6kNYSNdDfFqItVd5+3WnublcJmtsr5
sdrp9O9/wpbi2uJzzbwtaEMsIi+YeG5YbKb32o9lSg3PSg9JUayX6FW63LNk1lOF
gv9vUuQsOKg4mQcmArLkvFi9X1zQcLEgIBtThDDaOLFjnfEoN0m32mr2MX1NMphX
qrFbFvjJCQbRb3zRmeyW1rAJ7D7re+vGcmdxWhx29GanToXLLHxNNlGagjkAPcFO
L0GBAg+vYFtN1n83qqyoxbYCYEzEE+v3ef1a4kpOgXVJpfrf0kj7w6DE8rkcVE0x
3VO09aBJHHw2G9hYc9QGMPmjfvvt8bMvrlRjWnzJHq2wOo8ucAfaCGIX7FxNFGE0
Jgs8yucH2RSk7yy8sxnd+eejmtGa8BnZocpw/NnmaTIzAoc7eqbMJ4hQ5H0TALQ7
YWx3PeqHVt4jfV8SxSGnCUfywvHv7Xsnl4jzjmDhtbmUE3yeR5dlnzTedXJKfT1i
BOU6kbrcd/O3DkzuN4aPq8Z3X4VfUKAPkqOzYbuDf7pcCIUY1nvdWQJATyQ4jvX3
U4cAV0ULJM2138xVPjpcbCHxaVC7KBFnSqHGxJdsL2ggfnPijBKi6UEP1NwYhECn
xQcEAVbW+uESjOF3wAn/3aARc8ANlYCHmdtzReSPZ5gb1fgfduWF16A8WSwV+zDF
+KCxU9GFvfWAssrr7ANqDkGiz4KRExriB4mQ4fPseIO52V6nSkahHyNPxQ+5PQ2k
rQQ57GO9K1owt6bvetaEdOtoEFN5yZA5antPUG/cmplO1p58sgIxmAO2Ay8s2xz/
gJ66i9TgDOPmEiNR+fh4uXEdYILKhOr4LYZGJUKDPoIwdyPo+Aiego6ap1HDDT9g
Ryh42z5AAh0VlM4df2eaqtXBgHvrGan62/7yfI2fNnxQDqVfr3QxNK54s9OKILhm
p0dnXgZ3wevDk5TGVb1qd8g38eOXMgJdYlkQ+tXyqF4YJs72Nc55WwhZ0gFMfgat
HzXGgztTxjGOCod5vLf5/Fbo9aLG8U9tEW05pjlEbq0Kl4z5l6rJAWhZKezp3vx+
7gBYfy0qtgYyWcZtFQ5/6uFt/yYWSdKbzkSY9UUsf3fylpl21RNn1gniUKvxzELA
dvU+TyaKee6+0JwTRPPttg0uZmgOOB5R6Npc1uKyal5sRpViI0hbAH3mEUjAp+Pv
YP48W7KESABULR6s2Tk48CJmiAFxbkWKg97wyx9acAWG6zi2LU1+eOtz5RU/A1h1
zay/vcn5tHv84Jl/4+bwS60nNjXJmbseRMPPM+3V5okrMYoz0GJTzulSZrEPfvgs
iQ1nRH40pBViDwQG8Xu/FyBGYatnUwz+yQUKwl6ZmZWuvn48avL6Sz7kVX4icePK
45i419MEihhN6EuT4LZk4M77gbCgSt5nyuZR505zy5cijmDn0vq1fmtDF2S6IiQM
+bklziX7PyvZQ+ka/uZuypoKDrCMz2tHeyAR9kCO3V35nVQbCdlM2vVtBYHx1GD6
QdMvuO3tTaDZgdKkYtpcHqi/1BQ/7tranKzM6L0VbDRxRKZk7ysxF8ugjkvLwmxA
atRNj6uZuqVoPN0zbyhcxkvz2tqXWrrzM9zAYd9MZswgQFqJH9GBczs0JOLOk9Ln
+1TZGBABKAGd0cykpAUz4p40QZdRk9lR31W6FU5ZvRYG+idvWzsskrb/FLq9wZUH
DTYIARMxdsry7bHke4/SqncuPQUcMApWrcgLiQkE8c1DtJF1ZBlsJhpzdUKfNFAJ
9zGp0hJO36JEnKQgpmtwtYe4R8g3BtYn6iCSganMZdeXScKfB+wT8R964mlg6jCI
u510rStP8ViSKToxn8UUolXItAaGdo+Tlx5fCppoPDjxwLAOhE4LcTdgEDgM44oj
ZGxoEWYAhsXucCL1yKg71yzta8rB6u9k8zG+TbwoV27E1T6laMIOJOInwcW1w8JD
WOdEwgHY9sy1vKKNKzTLp3DLK4RWxdi90KZZIedXVcHBr+fQzMgWM3F17Wmbcizk
nYrXW5ZCI1fHb9uU7otWwXAuZqjYSvwwzHFQW4fv8i8tOtHRTCd86wIka80bAQ0p
gOEMWCZb4V4boo3R0NMufhq4NTKbYS0JY2NyLia9gv//jwJXb6Ze4QWxwbya981Y
LZumt9L6ofkxW99PCB0VBMh74XcLJuzrfzw14W+0lZAZQmYI5w5WANFZyzeCVb32
c9K1U2We/EPFHlh5Bb2POX/cUAdNj8ihtqM84+6jdTqcO37sFwaEH0IvXZtx7EVa
QzzO42rBMIiVtYj1oFN6UjA7PNPrPE0xIbeLBIyyypKhMXwZ5zBINJt0T0aVEXQr
BIxJIPaeyEwiCQ5lJq9DRcSDj/qlt/3Yqhpe7QTszU5GmOrOPqpzQHqrkNUeseX0
zkY+P/IFtK1goR774clr0i+aRWknk0zCbm3lmTpRIpv0mLmbGiflUGcuQD/722L+
CjeqbQC/v9YjQi7qyJI8+mHs2YDksTVXL0E+uM+Nvl2BtXNpET8z26GGozBx9KHh
rHFxlsHgOowbD9tn7TwCRFoREY98GjZry/uBe0ky4wpoFbs4SrlzsG9ScBtD28DD
fxGnekCWoBbWgpq18meE76lVfvMHhkezBNWNQadQO1Slkt5L/CZxf3E8hMwdkupM
2nH719qKJC/5Fb/uWWkM/aPNZc2mRiA0KmAP/PhxlJwxElOiHWazvICWIXVlfjVY
rUX7vru3JYYBGtFwpgYk46M6L9vAGpy9FAWGa8x8ZQBnwFy/sntvNd12gVQDDkD+
lDDi6TDJnMwsKS21+9kvreZpB+rGzjXIXwKq4ZBfRCpmcZ94CnS8aL78agCKnlSC
4D7mATb/xMKsygKC/6b9HTxoKnOMmR1jmBBW4Gx4llbjWG8oUSndXeHtSXdEb/Sp
GbbUA5gbTOf8pd0YcYnB7eq9aqTARD4IQpqqw+vRsxMOOYfrjsIPZ44t8nApNbrP
AFnEPp2RpjDSE4E+tYb+3twq3ke6q6meeKshj1UiAFdd+G7xENr6ikC/FS3wakaD
kcy9TONB8IggR7X3KW7WHMEymF066YnYi3aajCA5gxiEqXpZCM7VzsR/whAPGpLN
ZRQDKVSsxeDzXTFWjMzrTq4Nd05qTHMc7xwg+wBpz8yOJWTwLu6TbvY5jSRFsyNz
ZX0z/2cCu3GZFLZS2BAvz4kRF5Pq+9+4HVgizbiNgH6g+H05FQfLjyk5hDT1nbGD
citQSa9J/DAFCEJeDAvKdmt29wHKnKH9LMiKC2j/hwqoODyu3nzv7p0/ywEiulWl
MklNxh87zRcpA9y9OdHCI9vkpJmWTh6gFM0Iyh5Bk/+Q10dZu0WBN2VBqEkA6FcX
sdLhZmoESkZaauUjpHrnweEHYcJTLhs+bepncqG+GicfiTRWcVnGnonQ6CnvD9P8
e8hjkaosHyf67ys97vVO1kAqsPbuYdNCkO3nWrMAO/AlQTM3gxrTUTvU48Qd5GGK
t1zjzULXifC1nhNVUgf2wCeGCv7xqLRb+cCQyewq2XfNu/zUHScfTJ82CHhVgvU6
3JGvw4+eHbJ8kwwAtSqeA2FktiMYF3v/Qi9HXk/2FEmVCM5hW3rqKppsl7s7MvjR
klC25dX91pNU5hOgb8nR5XtQx0e1IfIwSBgtRJJvdEthkGeCCsrdjV+OJebR/4F4
lojK3AyFyPglQI+R1/hspXYAB88Q3robJuKSWWlnX7JGSH3jJGwixntp8DTuHE+x
W5aZgQujn7fTrvUwJmbm0SHmnMr2AXFjRVtJVHi3ckFj+9VMkTCvgi/2gX0T0+83
XEVqtOepFtJ1wC0ilxftGW3NatbMyvijqNE8OXo9srFSCMxAKTAIMM7vrXq4+JtG
C6JSbC373BT0E4y1Hl5pQOCMj7Rxr3Y8108Js22z1YjnIhttTfZA+EQB/kNSLsOv
Xk43h1PCpiLWEMGTODKksveFWtsssLE0tOzWi6/jGviAvN/+0x4hjBFziiG0+S5o
0VJ5NXXkNNJY/dSc2zKazMkeFXJjvG8mL1SVWtltkQR75kiadAIj9vavVu7Z1qUT
lES+L377gAcx+IJ6uzOl6vJoLCgIxZK7iQlRn7bdpFsq7gOCgpwJeRBwzF3pc7HZ
Kb7PYIO5rFauXvCPDhtJOPO+wIQ12X8SG4hZDziHQW8wuCAkIX4qFRxdQkZE4sHh
iT1eexN2YtcJ0v1GzHdiApXaosByv6n45cikgFPW2CDCYaFLA4jhHtMD1cshNAFs
80RpzQOTjVZv1wp69VPOezDWqVJ4zL+IkMCZv1dyX94ruKNWz5UWQ7LXChg/eqo6
Bi01/Kc29Nagm0gHuSJz5N9LsWdMf1Y6IQcUwFPn3T7x3gpuaf6GVwctgCZ4Tckl
OEQtQrBw1L34XuLzU5JTXsJcgsjmDKrZ4R79ZYPaWRTKKzG7RsnZ8tBPe9TeUOoh
qLywUaEtvujZuYd+ToPCZ5ovbOUBXPWuBKDirX1vFopYsTl1iMBeNJLWuOA400Ni
mfwuuRGGBksCilRyw1MzI47XSgAFAN0iUqDDutqzerupSyJe+k4nX3fJ8Wx2XuLv
vbkgYBP+jbj99AUJ46vHq9nyiwzDcFxiQxYglkVmH2x773xB0pklwrCRsX3OXef8
IJ8rwkPWPG5rF875WcGRsMGNedCYz8OKieSUEAFz8tdFg5jg6HFdN142NLPIU1+d
Hsh0nUrOBhOnomlDF7fh9DI/0Chzd5xRigCuvcda+Va22GMJrEpr0TAtw7CHC6Dm
0KYQSa02blKl1wuSYwf0cqVSj5EndStQ1rXpWw7/l7VLk3EdY8URblqz9zpQqEk2
tDr2MVvRu45f6VFegO5Z+XAns4wtPlG+K7ktufwDFmMMTAaWcZIIDML8lkZGnBjq
F/A00RfH85Lnp85/DMrJXMFp48yr5m254UvK2KHDz73QGKZnCjDrYfLrXiD6jflG
cExylVy7HqBe22BWywmyIegxFvGU1m38SccC1k0rbtROGua1R3lq60FvbYY7/rXM
lXPjvmCM16Y8Ly0Erkdwt/p2TYWfG4qZxeo1V8Cq+a8kvGutCdwMTj8Vw2TmkVIH
WtAtQhSTcrmzG6X2bq1GFf+NDma/5gyqgSUC9iz6KQnHfSKt8rqDfMByCT4bj4M+
2ZnHHN806W9LBDrnVu9K3C4Lbs3rqUXHii4RoRhm6EQUzPLdMQzQQzR47utdsvPg
QPDXxsZrnBnX1Ch+ofIRdgbWLOkZXn6IKU2rISg1D2VUBF1AxbenQ1L/W4SJuyA6
TzTHZUUb+cXjNboAjIr4Ht0aDG6b2qAEOBVv3WGWD55EZOYOd1WQU/jNKyN4/c6n
H41IjKOkhbGK2OoCCCwlX5ce1lHKN9eE4iJAYvE1QFhudyuRPAF9aOeurZz3xHtF
zBk4YYWc2XSHd35xfUyp5o+aSMuGarSyDqYfVxYIA5L9MVc3zYTK/k09lpGuAALc
WzPwP9bacJE5IH7Estb0Tvd2igYzjoprcxySxrckaJf2NwPs4oix+bMZz2RKvh9q
+vKHgnnyc8YMe28aXCnxFEGDUqtcw3Cv7rdkZaqkpV0dv2GDuMXf5iw/W+K3mPIY
3weNFob+8HLLJ6/vydjWw/EqC24YHFlqjWlGkWkzgzFHHz2T4bSd77GDVQB0zkMu
79gIo8NCR0me9h9xNTeQudceXz391JlRe4QaszSZhcuamHNZ1VKmUI9DwbyvxIAL
vCKJd9UXledOPDhdOq9iCoIqJD86hI6dFD/aD98ABoqHHqRW8PTu2hNo4CI1mc5/
PwLg9HkwHdv/ETM05DdEgH21Q8FUk2PK31RRhscF3yzisSds+rmNFDI3b9WFUmeu
RSPjtsxO118J6p3xcXprwWTEwaoV4Qp42D/3sQKIjT773Tb4R2LjTMadv6tNlLMN
VhUj9g7rf6EhUcgGARm3JRGK17Enus7se/iSryGaIiAqRx9iEgpqe0e+EPp5l8Kp
7+aKDIXDdI+uPD1hKlzpoPfkrbPqQJS+CsdPnO+5M3u8iJbS/wCbTn6NO3BZfH+d
fytoYkxZIbLKw0w1AcfLaDVjKPOAG5nd4rEXRiBa5fN6Ax4MdczM72VtNEzWSUCw
J8Dji6KAG8+RLWWi+AyD24NlUZ94wArONctywF+10UXswc+3Lvg7CQ+EB9/npUZG
UaPH+DR0NFUPbElqYsVhHGfJh61IC2UwosbcSDbaePKSOKXzszdslVuqgbZNrpo6
tlg6gMmB6Vzf6JFtmg8p2VYsTYNrwvtsEBzVb5Y0kdXFlTYmt9gn2fkFTMuT8mr5
+x7qTmBazYTmJc8Z+Wk7Fb3M1P2+NfFP5GZojcbdc5eOXthJk/u5/DMeBMTIbGwG
GIH8rQqPOG69OgIDXM9pzCqF0Aok1TC6Jby/d5B28kRnEspvySfgeLAh4kTnJbwA
69qXoTyH9tJF2/gPwm4U9WlGmop7QBsJ1kjcv1AUfj0FraFvQrLOmYN3/97XHPH7
iUE8wkVpKLW/fRJdb7H1yxGT/cn344zeUNVtmC9y+qpu03m7YAKhcKz1Cig3lUK0
Bjs5Gg3hT2CrY/T+WJqQ+qXD1wgN4wDIBWRFsiPU3MmILDEIC4+iw+jYzpCtCAhS
rmusOhgImr0A0UabkbHRyLvOQbFyTUyyPTfnVMbHZSvSXR31jorY/RAhnkDZzWBS
Twh0+ZW0PfEUU9c2GGcDONbDAJjJ9lSpgpRbD/11qdDdSBu/KlWkcWDXD4tIpnmt
p5IBLHVnGkfZKg7WjLh+DvRFPKGyKhCFjyUke+m22GFb29e7dGe38lkGcVYKYG4B
s78cSboPsAGsIr8Ntzu6hdvgPMrOdbc6Dop14GNCAy9/y8G3r/5EhV2+0a1NZCnD
FkmRL43G8aYtD7w2nVwpRVUlYWGlIvXN+uJEwAJeAKxpmeRNqosGvQcCS2ZTJopI
pbWESDYjIUB5/1kagC9ZEQAYs4OJAVUVC6ijI3DqHHed/2hZ3tG/2zqir+TIwXAx
PHIznCdasq740JdFIWMEhWmYGinDirn7l8RDzLqEE3Uks/PG4Aavz2CUqplcg5XE
tx6A6UZQ5xdgdptCXtIFY2TqcZCBxQH8BXhBdbysymccJHxUQ/XQmQ7tgJq9Q0+u
GWRy7XxRkjmE9O3D3zVQIstsoUsnECNepFSpBks7/r9nEKYT+hJVvsFMbiOGF+Nt
IyF8SeVgdZhgW8vWbMv548H7BMkJ7Dwbd7G96dV7uY78CpJByGEwCd8ThoBXiqJ2
77eB9Kp+fgieMCHg3BS0QnJPyj370TVgMgxcT+4vJ1QYorLxqUtmPRrsLyr3n7rm
dH1H3A7ZF/ZCgyQpIcgdhw4C4sRtjtiKD/rxVcInIb8Iaf6kAzsXn5R14l2O130B
2MM6Xzl72bj0ydtb8zov7saDBu4mCpPoq+bxnknJS0PzeqdVW+b6Bp3J82v2tWE8
Jk8sn4MkKy/PHhdD31IsaSQ/9R5GwJ8vryoP5Q7uoPBb0nce3kbZrVse8aqJWJdw
2lcvtNPe5a5jerkwrr+O8bJAPL7yG95G8RgzdoWg/9Y2kSYq8AOux8lXhX2CQKxh
6tIaGf3q0unBsWvR3mqskr6cotDx9ogko4YQlIT3K36fFjAC9BG4kL68D64ZvMIF
aALDWGsEKSIfCFsL4Uq3dQ==
`pragma protect end_protected
