`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fOrMSpTUpyd4KwaXX5GMY+oJThdm9jWLa2BFYeeNBDL6B3Cg57eK8KVMSNfC4icX
hbrRfCkV8Of2kCTDg8AbBVw5PpcNAc2W3eqAYmknjh4zLy0X4TEwZrlvkH0RpCVU
AkR3XZN6bPA5I3CBoOEP05T4l/0kwwdg+ci/jRdVaDM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11632)
gQqqnu78vdEgG9ZNrl8B96CwI/mgnYrOjUzu5rXHiPAfrn6RdSQ8TmPLiCgoltNI
y3jnSAp+rQZN2jq44/clAdzQiBXTm8ENj2moKFfhHO5zC14d/4z0tZd0tvxoU0tG
oRdlzQcsMsO4a01pRAkv/ju88hXFNQ9AeLCbxu5XN5aKpRmmnjZ+nGTo9ztBKjvN
03UbnV84mVOIHleIm1Vyaio27kCOouo8LmXDhEQ0iBd5ew3DZmGsiMmYYfDOkvSR
aI8iD33LN1x3OQ8HuptTfVfb25LSWRg18rbPQ7sLcFDGS7s/3He80zpC0TKBYHtp
N0st45oH01sd2hzgbQlqr2PnwOKsOWDkwDHVq6AEkqvMP1+gH9rMYH/Rg5zaWhdP
aVWKMmEG12EbfRsK7hHjSVzOLeNYNUWoBi039inDc7EgVp3+jmsdoL3wdUhxfBd7
uRfOj3CtUgpPIGndAYqffA50HSwHVUQm+WnZj84lToG87l3EHkCwVj5oKzBHi8N7
vUU7iK8JGIg5z7FwZO/IUEKihsOZEFj8++MaQyf//tOMKBPwxjAE55SIh7geyzEa
6g3Drg/T/XiBVp+5r40SpB/OCqHeyMkbZ5mPG7i2sDi5mKu8w/mVZYHCF0Gzm0w6
n2C+Wkf2eMHVulLKrxjqFTBpX4k49aBZg9TITRGWiz9KPReKN2F4ntkIjJe3SEBi
ljBbR/fd5+EWPVi1JPDt9GlRX04GOnXVKeFS5udyTVZi5qUb/jidbxTug70x2Vjm
+xwzKwgmdjTf+EajLewC4sg30ZzI6i7VLu21amippaaXt+u09QNFkl6jZLSSMOsi
RUmEHkcdP3oppji46HeHSSYLDd2JsKbxIuUXTQ9scdhzT1OyXCSvTT2Qp+zLxOfB
6/7wHMSY9ftAmsTH7KUxWXSolXh2QmArTQ1gX6ixFcw9nXDeDDYOHEkBfK37KtTn
VeFHsVEHLxT7NDB74kULC8sJQxWRLr9XT8Kt0/KSeRWDbnVNWfQ2ZxIy9RvvMRrG
k1sPbClcOh8HWa4LDizu/mRv7v6B3PZfe781Tr6743tzpOtqNLXD2+PN98Au/JJq
gkB3W2rVSZclDpYYNoUaBcF2Wi1kueNAf7PavnlrbJXN2APhm6l6rpIVqzh2FpoI
CH4rA8xAnVgpIs8qtDfXKV+WZ1/El/m8x+KrZt/wpUiviyP2wTS+Kq+KJLkxQL0j
uWY0g0ZP5u6WsOIwetydzfSpAgCJeZJpXSJGM6VaNyu3K1+2c5bgXYiJTdTFGUaC
i/R3pC1prADMwRVlU1bxEuetuQxTOlcTjpdrl6Y27Sgu9CduZcvhBcdeTRe2E5Pl
8zbovBimfCtHBLoeaQumegRak/9v7/FBDzt4ZNNbyPqIAHd5V1MBFNnt4hHMSs4x
7y5vl1Ys8OybStrM47CrWRp4aNiCDKqzeTEaptmx4I1AqarCoGj9ja+ZUB85cv7B
/1DKbbRN6uHi6PHPcoNQwoNTHizriPKj+2ueAWm182Oh0QYajMjxuHDQ/xBU/tL3
6eQHQnSLk6UtS0a/L3h0G1M963kIgapl6Lh6OQ9ZQVfDERmVP4ItMp6/YlIIcL+M
+hKvrjNT/CNZddCjSAFFTCdDOiog+ZYJnBIRfbqDOW3uYTaUZn2LOfoxQ56yzttD
pSPJmgzooSkultdvv6nDOzZc/5kiJ8ancetPHvEPcW80ZephPR17Y+sabCb7Aclf
BzqI1sf8nHCoyu0E62gqcyPt7TAVEqmzCFjcD41b6+qFMUtecZjcXmHHoMZsWafx
GVSNDdMQMZY7gI2Sgckvla2ifCPL9nkm5ixNptPNZwjXL0Wm8vxH18BMYUkKj2Bm
GzvKo/Frw8qwa3GuXrrWv1jHKU+CjbONroYv+eSxJcIGvQ1uUENPbvEw5hncXPiH
obRFBliiMPKhFr0NWRvnC9/gClzZvPr+7SgckSv6He5fcic9PNFzmTI+e833YkSW
tvRRKKXRJo0OtgunxIyoXg91G8DLvL+OyhthVDEpLYEfqWQynkpLT+rbfS1zn/hH
T0t4pxl2Iiw+f7+RfyP4l9E089A/wPs7wPsAZ31y6OeTrV8OVbrvq5Gt/6sp7bn2
I0GSZIW7VFGIUl6XzKqrtlCwX9yis/pkQRqU5OvKvgTHHdyEZZMJw9Ky+edClvEE
XszE0gci6Dtth3NnhkLDaQ0nlURyCobVz1WhuBfDXY6+v8gK0AVnSJHCmmI1KYyW
5EVnyUygocE4vSi//65VT9FITGAK/LMRmQQ2jv6PpQpR63Ydxc0+rGGPbDukPoLR
zTWxyi3PrXOOIj2M6gDpv3WwQhaDOjuqMSM2gpahTsyP61FlBwzPKmklRVjeg0tE
5KL3U6XlrwiGB+ENYtmHIzWWzr/tzhaTgrW5zMKQkC0B0NNhlPcmvw6UNAPtl13J
STnr/tGx6xc8gqks7O3JCU58t/YRjjgaEanmi/4k4XyzJ75fyaoLcA6TQTIlFMSY
5C6e9+wd9laNlviMmYo44sRBZE4FLy+SJpqgPgPvdnqcV9vGAJAhCnF6segwwBmV
ZOBfuynwNMJD4BMET36gOVoYAZoZmPkuc9wXkFlP+9mmOyydby/WB8fE3WC4w7cf
nwAHjzoTemAfZXxPmJfV2AQZa4lPKGEHtv3IUO5l5EYb3tSf1zjaPpgf+Yu6yIoT
gIBeE3jvDf+X6fXzbhjObpqHvdX80vCjsz2P6x8LAEEDG7/EuLOGMTGjv/x69AQz
vs/jl0tuZQhtV6uKccz8RNpKi0xnBfVkQlltxeTh60cM1n20e5/y8PJbcnaXuy1l
H5eEyJIhIwg6NMbXJAgGE1j8JvAOOwoE+fMKhOjSCvGPOzdu2nXs4OE6Qcoeem4E
UIr/obfgMx7Bfzj3RBj7LYN/rlcaqPNRMGQtOcSnD8vb8/Kujm3Pc5TAqpxQl6os
3mZPKLf+wiNR/Hwy+5MBg1GmYDD++Jy4MZbBUDfgv2N+2nYrRP/3tkGQ5WeD7gvC
u42oqYdDzNtHyn1GRhS7pdF8KjfircfUygXEjgvjGXYtmBDlVEQXKURy3FBQOh5y
k/0MgRRpq6pIh3klgAEfY7BSAQbLmOVwbovc4wD1MifeI7o5WWn8aftYFzbLId2R
yCdTJ+OUN6lGNAfqHs+Cl37Eai0u3PuklKmxQ+0C8hKYXoqjQPq6knVWKbmkUTBm
5LBVLYLgQ85FMpe6LAcb0Nbb2I6zW2z4Mz24bHRtOY+gz0G4IHmK9IB1dOtkPGKy
+9JN+g7KscAGtO1gL2lyh/Fr7b55JwT7AJw4Ncxk1wglHcUMB7kdwyXAg4do26H9
8ieBlDwGMwnzrZYsUfM5OKYsmTtQi4m1ry9S4bq/HzglimdUNMPEiCyTrq4jFGCi
g+mLo4898kNjumskhE+8csm+wLvNY9ro17Yifp5iGWaDwp0S8GItglCdfEwn8hnl
vafBal5JtP65W24Dek4Wez5CFZ1vjppvHZRRvm38SJhTHSf+jAHY0HeBuSWVYvAL
HT+nKFDjEDoTsOtU+9Qz1VjQbLFRC3qyi9jKwXpnLQ8pQrSLQSiVOzxxotjwyixe
Q5NggRnMp8LTuhtlZ3g7lCEXZmteNPqU1C4fgNrSb/v2sM6aPgKPP/7szTAKr+Ij
InQLypkAnsaMFDKCIgt4gTKWhleXtemYBJM4qv+YchXdrqme5bjeB1h8zSQbDLor
Ij1nyocjlO32vhO9P8EkmozwrnSnaFMK7xmsIobldMiFsGHnxGhwoKIgoZSnVi/z
7V9wkGTmbtH3fvLCUCpbuHjAzHVFHVy8gUBxhLgmpEI3dHJXHvf/n+/ywc8G0wNq
b0P5xeGCl1c/M9lsQvnyJ6AxdROjOrclqvvQpsN5y8Gw6lV4pAeyiw5CjT9/LcYD
Q9e4dlcqHy65OD/QCF3bpAES5DgUyaN7C46huCpt3d9b27nDpOuI8TZa91zVA6GE
/2Bvyjo45wU+OKxMWMUoVmZeSpjmTwfjvFr1IewWbD4pVQOBIgSHBauk4UFdFJFJ
cLlkErmMWeQ0+uyeJ90+fyvW6rdjnEHEfjilHutzyiUicVKcq1GcGFrOawP9kDak
8GZACB4uz0SNTRN8lfB25qlPVVCZZe0tcG5I5WI8aYiD6levWR+YpMBYB3mmR1DT
weu/W601z6qn98v25VUBqFiYbbx6inCTOtGitHKpOLRDjPGchfqPI3fF7zIFW+Tr
Cr14RavMny3SpEFtYhBsrPjMan5rxltEREuV1GfY9gbr+w+rP1TAjbuaRZTibad9
5P8UeoylKhyN99aiBVkia+NWMD+uEUZkAKOpTCi2pho+32JXkv/oMr3BFz8FTpKR
CrXDHgrcKp354nTtWW0bBMeB7jWKIyja5bMlpgydtgsQDybG/akFE/NT4bDxvJw3
KEfci2pi5BMCMWwCNdoplfEtINTEthf73AHRAluXHe3vW8JCP/IODriuOxBCte7b
2aIKepx2l6ke9K8SMoLeAjnHl4krNa8skgwtIrWVnbjnEt1yy7OrZWyRvftAXNc5
POA6x93TK/ZNMti7ub5VMIViP8oleGeK4pGdmQXenTh4L4rpRewRaqbXpciEcsRX
R2j1BhZ/Fn50kYCjdJlwGN/xzodUvIBiDhlBw0q+PCtac4OJe4/BJqpJ6EfqMGBS
AwNWp3Ll2O37lkgr/UwmWyJI55J/MdArUxJKFyUp02zLFlGmuOf2StCS/MZrrve4
ra0162mKScCj6YI7s8qWIlOrUjFqd1tdm5hImmu9kSTG6/pWRLfbMo+TLKbxZeD7
ISc3eo2Vpbw0S3Qe5tL4jRuhgt5lcqEdP+p0CFDECWUoUfdbp90pB9Qk9SMp0kIo
uSIK507Dh4Sn/tFtn1yYp1p5EZw8r3P1yNGvpkyQaVS0jZOJbuPPuNN8V2wHtTls
HAkBa/QT1eAEEiwxfidU7BsuQ4od2kwrkyoFPK1zGc9j8CA1lY8la8Hz2GGjznFU
ZUjcq37DeLwyjyjKnZaVUCW2wn/dYYlDmKMPOo64QNS+kH7js8aszRQHIwM7kb8f
HW6Yz+WIqDwh5VNydm5YUSozZBTU+q1TmIlhL1gOBT3Ct0rOMStoIrs4sNl31uUB
x7VyU+IwjURJZ+28ZQcbJrv/mMu192Ux/Ke79pkKfc6l0t49W8hg6KWThUlehxjB
3IUXA39bAaPi2HYephuaC7AGTstJgyUoxfMjvU7RY8L7c4zpMW9hjgk+TWTxEE55
F3V79PZoaw2s9hqQFZfW3o5NpvyTeG5zc0swHyt9MOIGxI5d6G7ps1osXcUultOe
Qvbb/ggkJ80JJGNNJg5oni/kb74k2lQFT7vfJE/hysitc+5t/VqRK5AL9AnsFuo7
3Vbz0ucxeEJYKpn1C7bZa2YZeyl9dkNSS+Z4/YeAJW3DTc8BRkrjQ8XSEXi4Spgp
x7zt2XfqBPxhVildjF4ESKECzvvAK5lafPSrLQqAgHY2lFRwKfOMA7iNp0MsVtcy
irrcBYdfttVu/iQn6IM4dZdm6isbyXSaOF+l04ZP6sKOp/HsuXCnnTHj8WJRHiph
9V91GNKsVcl5JlDfkobctM5m7WZC7wJGQvVAZqge6HAE+MuNOEFnHug9hdbPF6F6
WUH8lr0Tmg/G5ZRvwxu7Y2Od9rCo9D1XCKCVuPgYBEtNES6vBidTpbGUyLzy7Pdx
6vMWIJteDLpqdi5VnPfb0XxQAfi2dkyXiVh2tjOMlTrQdUt2NUBgD+eqRV4Nzlig
4EsOqI5qSiJm/stUe6zX5/FaktVrOYl37cvYPTxKzxNXK1Z4cDx+fT3xfASNZ/Wx
IKJbJYcVDXSbT02z2NgcFaqQS0WEer8/urEiyaCDN2523TanZ7Hx6PYpKpGS8gL/
NyFWBn8relpVZgslk+XM0h55jRomir5wBABE+rGho4ZcRll01kWqtoc8+aWvLAKk
iDrg1lwm6U/A/XTWD/YtJbsm95rNQPvWIYAvCh8J6LNMq3IVHZSUu1j/AAuQ9aP+
QTlNe8qd+IpSqozYINGk8Ceb/Uqgez1J8xhmRSfZWX82o4fbSLY8vEWd9xpv9R05
srJvEABABjYH5uMrMQEEXPwwjAXrW5kUPqGo+g72Hd/vT+z3oyFR5cOSrx4IivC4
KKBvu59uVub/68cEyL7IOAWHN4t62+3Smt6veum9WUDtvSIUwE5Fjjsls/N8DTee
g7yEl2klIWNnPVa4ox5cCCMzNl3o264e3IVAXsHMF+Ld/1ve2dDAOB1GzNcnSFUJ
PqzFf7ErsWMNs4jeiVFRglgP/fS+fywZxiG9qOu1+2LkEQEFyecfSFEG07fzqZPe
QCopJfiLiFu1ii0gFxVlWyo8KkzLbDJcf2+w+wR3z1ujeWHc6OKood9BZ00Di4UI
kLXVGTlDTsUj4tHlac6IDa7CBUS6MSZwgldN+LiwhGlOPBq4kkARTPpBSiLDnPaX
+lf/BPL6wVYPYTcIfvf/AZxwgcFswdFUPUuKWfRU3iPnIlLkMSrlUy746Us+8a5q
6bt1AEzPifOd6O59GnJSpz14TlMyJawJ7s/1lY4RSLRNHvmSOYQ6wwOgmX2x8Y5W
kgXjDOtgCIDfNIqXoe2mUOBYUugAwruyliGvw4JY/YIa+lLHqF8XHgTxun/kpqOP
Tym4ZtUz/zmiYzByxWbozStv022sEQgJtqJLFzmVliISScoNCCdN0Ft1l7p2cs/a
//XcnaSMU0fAZJwJT1f6k48VwMv1lggxvGcWBsuoAnFmAdlzE4ubIX21EQbtEjSU
QvzE9Cv2oKutQeMdqrhokAa3q5Koglc5dzZYHmDxIFPaFd5xwIKd8C99r+pR7mHu
ZPqRPno67bU84CkSjscooxTcAARqvDHu+5uNbDt9l96uTQX5Jowzr7wN4KEcTcHR
ffc70cZ09Hw4rsXkMAFMk9hSmAMHWEfeSaJ71OZ+Ae6n0OI0xIDZQHTFJ2r0XIyN
dOF2Gz/+odknvwzIBvwTp1Z3YK0bWmVcY+tDgDsFaoIrHTP/Q5YSl0qC4pD/o/zs
tLebsesLA/YTajZ8aWvmhZF4vG+sbLh1xZaoOuTFIPwnsHbQBOPYIGU+PJo+Ep6B
K5xgRQm4HqrJrlBY9rAwqxKxD+6jLD7JpGzmGKxG+p/cg+QU2cWUCkS6iGdgUMKs
FXNwriXh0Gu/cCXpOV4Gb+O9vWohMRzPxUB3YaMf0jq1wwB4PTA8WsEx0ghr+Nk4
3B8YZ2WcqSmIEZkgb/LgjjZU+FUle3eiro0tvk4/Tax5AbV0pWS9ScoN3kZ19VTb
EemYBkssXzhu5IUeobx4iFyHrIzBcc/xaVVC49C9iF8S4B+3xyEDl3HnLp7MmObx
gqRE8X4qGC/PoZZOqcSi7LIeOJRwI0bLebrdmUIHJ1dG7IzwBXsR9Ge6YolFEAlV
wLwXj9x6bI9JC1feUtDL5UgZqF1qy7nkNB2znfHxTBRdrIxB8jVGPPJOzFX2sGKW
BF5ZqtPhEgNDaaG84JmfMISLdkTjt47kce/ncFx9UXzqHsf31qkPOgWfPQpbHjn4
9uyL/KxzJzi1qGz4Dmb6Exq53GTTiyzt1JJAQbK1cUXtPqvpkpI1fzzCEfVUONfp
vgEiLQxvhmN4YJ5N5I10VPAmxCW6FpOn8ddBnw455V23krJFuDTPhnqQ6McU+i60
vIfEP5FgPQNk0m4W6cR+gsjeYv9ZtTTT9h2dDwfLtaaXhDZVmLnCnEIPHKeepc1l
4BGhD42egC+jt4wyJBkttPTVF0bBqyx2cA72SBT6CTflWGcQmm2D7CX1gLzAxugE
1hgA4RlCEwKLwfJGNBvoREAE517vAFAemhhJS5oqCyFSQ6JsVdIU/D8DVWMblcMm
jPjZBrUOkdBaTsqVpNfuFWls7l8jR+5IhafubICfafu4ChsTthq0vjHugb8MkJIw
2U43bmaTmyflBuB8/uyCXgB8UWhTZ8J6+EfOKLxNsUlw+Oc6dx41pxyAE1GYHsJ2
nxJsNBSQwXpKRGOn53ki21wro+lsK6ohE41/InWfays+K2r60hpz3UOyWJeLcwC1
5b1XPU8BvPXF0lBpL8f/SApT4OSYDxafIRwUbhWHWriKaVp06W0VXoOxaPzCcRFK
Ld/jYYEmeSIVEeh0mGPf7zbUFjwzbz6ZcG3JMPcycawHG80oeNTic6I6KDIuVAUw
83BXlfe1Tw3UgexuuV6ReqVRLC6kqOWgHXOTQGOel8AyJUaHkDj3262FD8JvFaIR
TXQWEqougGG4kswYrbTJc5yokBNLsD+m7WGt9vPMt2q5JebV4tIgXcwHQd1c20XQ
joQccLNgehtDVi1GMVp6Tkrbjila7Qd8TiwtTn14bwA2d14ySofLaPHyeXYr9pqj
O/Rp98s1MP9UHRnedanfbqpT4YZ8rJUkrPJtBjB96F4E83cHGOD9kdqDzEgsRf6x
BJFoNBnI+ZFvUNCUX23TC+B06CP93BrJywXOJXRbnZ9sDNc/17p6h5fKRcNqPP4q
FcZM+8WgBEsXkJ8yxg44WZd6ElF1eXhm0exB+3nTl8wVPOmGXiF0Nr4d55jqoioX
VyDEPj8JeEzxajKVNCJGSnJ9CqejScI0bmz31Y2plZE7TlJ4zo55Nwgr0MkUwyCQ
4Lfvvi6FPLJVVLiwTPPbc7eWSzjDwMa9lZZXFL9cy2RtlQRhcdtRLkYnfJ6vovpv
SpgZiO13OkZvuuU9BhM/96FsYBAGs7kBNDADD5hlzTDs6A4kGfwM21nhEece5R4A
25luj9ZfJI5cG6i9VFJbgbpCw9gvbRa/94TMgTijXPyXot+wmlV1LObHHT7Pvdcw
fe+XNADEpeS4ZlfW/XG78SIFh9+jw7Z1kiqnmFPMBNU2Kd8pYljjivX+gC1AFoC9
JBC7i8GKj+07NVlzbhx+179S1wIxAkmT+YPcQCXX9AaAc9BXx4S1AJ5IHY+pqHRT
KdPcPW8qN/FOz45MMv2NKg+5+rRHmhtfnODb9RaQ8ZnWHH3Z2ANVPqbY163nsEll
PHIoE13o02tekr+NqH9jkoiDAE5h3sPPo8KlqOnSinwS7xihqygxRIGYpYpXJEO1
n/pVF0wKDWYZiGXzxH22XZdSVH5RU3NRzU8xWuCIGumRApSKjY9hn4NCUOov3gaB
WSDjsEh7oZpxsUOhanNP81kG+ZKsgVfeyE/7pQkxyRIlJdt9dSCcRUJdHzH8aQKa
hBDH7Hc5JNbS/OWqh9RYo0ab12Jtk6Uos9NZuvoGjrJCO8vWvCCUVeCi05TF0tRT
9zPVFYoqsSVAGQov39jQ8NVDrMiSk5uxZcGYHDNptnxqexlnAFWYP50BPq1loMwu
4U3Wszd8J7c/+qHXrFNACxNnZ9+dzbrNeiCjLs4LUgUQZ2YKJWee54ncfpIgXV1R
t0H+DP9N/f+ysXiKMIZ68hd9y00OsjnL5Oi0e/LhZTrtbn7e8c3vy/oNvo9gxVwx
1e1sqZavc8CHcb2k9HWgTZ9VSSz1JgQYIcTDwxvZo90ttXATzeeg7HTOCSgOUCqu
KqCOGbeTlyXelrLeIQpQGpFnPyyxsvDjcGHw992SsCilvs+l09U1MjV0Y31WrTzl
8EDEDvBC6EpuOq9tzK2IirJGWOTQ4VU6V5gYq1I3FP27jW4vTHvlXpZbGtSS3ylo
GpwSO3U3MuiV5Wjyw4clKqb9OIfwApGT/oLIMzn/7pcNrtNvcvcwouAItwnCVa8N
IxQH+dhrHyoZuT4zu0XRmOb7sdczkq6nlDvZKhAPUKMIOvqzwHtaWQdq0Iv3t0bB
0NbViCo6/AFFWay9XzGD5ba0xiXHgv/7jdusHRiBvtPliUTRHvujqiTSkNbWN1Zu
EKIogkCCa2IUmL9mo1SIYnhu879CW4BVexFnd8zdsVQjLSBaMM7yD7HJzACALfgs
zRD9BQCRvG2jiAQqvbLEm8ad9rcunTS1BjS49m2GsBagddPA/MP+MAg9uJFLrmb7
WAyfb1CvpTGql3z/MyEu8tqtqy6BzHu3iqrizlohMzI9RrFrzt+c75xMT92X4Zci
PsObN9IRW6KcCXTIBi6C0jXuA/J+tGzCW8O1W8RodOZmhxbXaJA36+XHqNYDVQFC
U2iIFVmtfcfRx7E3creWNsW2n9jsnzZ93i8bXlFOnLuAg74butvrSeKHadAIo+pI
w1pzCpUzbp3JOrsc6Me8YxIov0dQYdrzdPiolsFv2BGxG2AIfYa7TldQ93zhN/Jb
2Dl6AYAv9Bp8EwPhnLstQ4AV/Ef+TwisrzFd/FsQqKK1qT5LHc/MUiLTfsWP/u1r
A2uSBo8tLHjJFg+OLRReyKKbYrclWxPmy1pVW9x6jq/PHGdjxd9JS1QoKNfccqyh
JeXfxlHQkmg8sMgifI+FECia+EkcsYoR9L6XvxUaA/d0tQpgKSjFp0UmtnV4q/yk
TB/jd0W/vqnuLloqrR2bSiHDtKMo5qoaVKWJoiEs09Ym0jorzXoi/FFFLiwxh3qA
jGmxLp1jZpKb0sXyDndrUZdEVAGwoiDeGHJVy1LBeHte7fK4bu8keXn3RIBkGVAC
4BWP84fUgK5SPWpyf4FQukP+3+US46RdRHwfTPiHOPpZ1Ynd3rsC+oYgbUAaBgmp
afUov3lT+xQBdPaPRl0ruxnP+wP4givjpj6V87DKpMSTo+j+hh0pAU+BXCXgiUGi
DutdjuGA2/u9i4s0DgY27VzTjDbu1wQA9lOzF0vI4pRd2l5qJCfWJZIILnxKf7df
tu19e+zDeup//DTsog3sgmyMrmkfr8h9boa6BjFGe18/JiVDBK/WnPJ/POYAje+E
PogkQyuO1k+wcl5VfOjDA5Prkn4lVF/ft8MIKawH8nQgrPBXDghMwLfzVVe+Xq+G
nfBVAw4rLy0WGp1E7QYKbRmIfd/kEgcaYoo8tKd89byEky2G6Txv+lDsZXHKQjeC
1p2nwXq1U63bhgnk4oW6hYymoJ6kgo1+mH4ZlenI8MZMX+8WLgVxtweozKSYpt8M
+ol4jp5JhdkSFWirQ/zkrMZC+7qcrCMkW/Cwx+TOIgLu9zrpSd1QAdWBTnFthKd2
9dm90J7UWQ0XRiOrkri2gkeHcF9dkwfjjEIgwOagoz9WppRmKXkrQbfCLTk8uQH1
3ry0fBZUO88W1U5PdfCIkHWZN3K5KXmZTrx8LmpiiedLDPkw0YELJR46zyAe2koy
dVIUvF0KQ0ZcixxEq7cmoAJS2O507Gn4z759n8IrjlL1q4RwIDHeWV9uLG0Or8D2
r1oyrypwjj0u237A56s1KqrA0QdOpn/ANeqMoVmoOIiOLJyE6T4PHw6oZ7dV5QGA
YC66kM3VkMZ0MDMUDv1zCLUwSR6vMyRZMeanEQGSCGfgcO2+Ot1ckuH0bPkCFNFu
yv0gntHbjP+4kmMKpqk4c27Os4+Utme91om9nns1EatIltxNuWrkB5FqS65hL6rT
GPeBwwnKhnXN0U/oC8/ymbcDl8pdmuP8w9wf+13gVFu5V8o+DuX1vLXTLUW9iHsj
HuqwJVIsKMvE9op0ZOXDxMIPVBV2qNd9Y3ztYoYn9hZbbvDZJ2kjtqpbqSdTMBks
r+OOKzKjlF4LuniRbNXA1+D/TFi85oJroElFwwfd33DjNakYroielIBLLNoC8MVK
z1g7BdsQURcSs45KGWZ8SAcUmgKGjTO4yqWWQ2fAU3anajINFuWNlPT97jgremtk
EVSKH0BObdtq0jg7H/3cg8GInGCqLXsJn6b1OkohStm1B+JPaDEj+FV5UXamT/sz
sujyk2PlnK5h86ZXTaIrNHgdiA19rRLM/VnsCIbqupJACculRkam6o2HP/XeZuZn
kpIjDXWvgdUqSDoP4ZK3n5U+H+JWp3NenqnCSE+s1bqk6j477j54BDPyO2GWQAfu
h72bNk5AhGJUiUd9LR7ZsBnceNVgcsmeD/JuMyfrfIhAid/OjmM3wsl97Gurzl4Z
yRAdqsD5DMafVTulnMD9LyxO6YZDCZG4SmpY7IcwiDlNyyXkKrhjX28c4e/ZDn3c
qewoei7duWjhdMjvKMDZxk+A77pfvRygvB74QPaOG1x+2ydlQMWtwKvbwML3IlAP
9f842+ZZ09VGhio4ZLgfRxHqkD1oOX+cezyXgtS4CUyyH/Dss9QOr1znO9rOFdEq
hXQO4m4ESJvmZwrkXiVl//DzNEqVv5zX8rW+1WpUbtg2UYqyQvoKjCxBkzsHGe2y
GXbUPGD5b4N1dC0zDwOXLPxQOAdJqnq6gNvIFHgdiLPj+YY2ZPJXqTv50p2wfLHV
1JsmUaFffgml6jL6svJbHqF9YDXl+PjH6VUmbkDzFCfyg+1pWGzCDgs7HMjjZ9BZ
0Ix1x7+XO4OhohWxgievPYcMD01gaocEJfNSwmUC9STxfJzFesOeKi0XfD8dNHkJ
1DRlylXbgZXv30/QR/Ns3OzypheZitYhKkxxSh2UVwKXXIiEuUYtN872pDlbA2Xq
GrvyY5ZzmJycwf7fvTcNiulkcT5E6An62Wa8e/JzMmdFBAOGQMPNU6b8M/PVz8sF
qwBJZp5Qt6GSb8/xdjWUyPmJ52bm9DtocXF7pVvOJo1dICcwf1HFrKQfnGXeyNei
END92+iFYTalS3zBfr2KYeKy8ai0Z8Rvkabu3EH+P2RfWyJq61rcVR5DV9XyqBTY
geyz7kmEZFOCgXe9h/Ff8XL4SrKHiaC5JVCX+9MUNRd5HGoXMlKgPrDdIvRSN7Tv
6FcCqPh9vYHQTZMs35FVKuWNMDfyTjM7HuMolHAeJiEPH4YOB525C1+8DHH6sKrp
2dblfe1J9uSDfUoDXA1qa+SlNkyeIE87F3ACuQq+KQOC1z4u6ZQqoJItqQoc7V6X
Mu3Cg2UMPmoI3HPBGd2mXdvO/FBl1Nx/KPSUvIBaTTJqgIfSNmXs5q8EBSGKcrKv
guQ6M5+A+YfS+R5p95CQdW27lG7jEMsmShtguvuHD3/UNHCj5GjpqeZtcBjpeo2Z
tU82oAGs6590mKIcIGxP3Uh5bwPlw4tNrZmn86/jSQ/BOtCohyOQQRssn/IY4XkB
CMxRQ6ExiVOseXZwarA9nC8uX+veyXZsJy+H970a67PbpW5qT2m3aQheGHsdK2hW
8JVAa/Gu6W6OiDKOmXkyS7CyKLDCu7P6AcXTzXph3gHP/M7/vY385SrsStGCmHHG
DGqQnL/JvndEBvQ/uhRpbLd+GxYhrQAcA2rqVp5WdDJNzYAWVQazsHU/S+hog1Zy
A+eU+Mkyz+XmLOpD8/DO9/7N4f+UJpc1SxbBJvqdjO1fzUsgvpqp7fxqkxStCNG8
xYt8+3vlmkKwGt/emDK2/Id+mnY/Wd/Nf1qDpcUVaOwLOCmWzWAGTzFZ8gh0V+WZ
kQDIRY6oyQArKYH5ygaDzmtBCJqLQUD6HsEhUol9wA1sD/RHprqF8oI0ECkkXseS
qk6H5EVKCgo47ulwGDbFHMMXdejttD3HocQ5Em+RJEQgpEoW4cKxDjkHhmVqkWmM
oRwlDqTTWTaGCphjJXflhZaP5zS6D4+jlyCZFmzkhc81zFjKgpPja/ktVuWDwk6H
mfoNKRK3g4NbvFWoqczXirc6ltItXw0GO1DGb0uWhMnaJ0I5O7/3Sm7ED7UaOLpL
9j1gRitnepTciIMFlAtQghmvQ1ewV/iKOViC5HfvLTq6a8LWnQfs7nHfbB17/NEO
L84KyS05MCig4OeWxxrwVvcqe5sguEhV0q72pSE7YyBht33rmGvvlsBw9f0G4XSz
+B6RwVzC+NpTt1/roE0hDh83vZkg/nyI6TF6Qf1+qTPa6Nz97g8q8K7tqLUKKYmE
gg5Ou5++LYWjf1OpiuGHBXrJqoF5qBK99JNr1X5vAWNKzhXhEXTo8jpUAQYSo17m
fYigBRcd6UI0LNdv2lP2HxZwm+uQAZRzbwhWwTOIvhdIM/3FO7bQkQOFOR8PXNf6
ZgpB6JYyFfP+KttlVSJpOvS0mMKkujpc0AVbSfyV+uYUkBo2bphYuERVQmdNTqsE
3ouUFFWhCZmna/iz6VNy9i4wBP8VMJ7nAg4NBwxQZxvyRZ04fsYTdCUiGQ4fjHwq
8z78Nptbpymz3ai10FelNXWKHAd+BL9sMBQU/VIUN8FEN70waV3424FH7ioSKuHU
Py3J8V1slt7pcMAdKrEL5UiCINDCdZFbxlBuNEx1ORYrjAVxzzH1MTBKpZqbUvmI
unDvNVbuGH8uD624C1zWrpjwFpkV5kf11hpQVh/jedjqlVcqM+ljM5VnbDRbeiO/
AluBVm8Calbf3vSqGIeqcawd/JNJL7Dqq4XeDbUfG51porMY+Uahf3k5+Mud+66v
vbmROiMGW4h2fkokEFzE2uBvn6jEcC4wCCbhvO/ejev9SqUpevX0K9ce5zNgTO6e
FuyHpPFWLmoJGl5BUKRqVByFjXT7JIwsa89x9pSm7uBJEuDoMx9xUny2wYuz/T1K
dcA5Hz6Z2xN7uiWG/mekHZ7m71MnhNLYqOQDIg5SN+iPeN0NVvwhTqYSA7nlJ9Ct
BmhwO+Su1IKTrKFxDYL1nVmUvPLs7wy850x+Z9i2pKbTdojslOCnc40E+V9//HgV
CEkNI5w4h5W58xMuUBRvWscYJU7q0o+ML7YC4IIT04t7FEfbkPio6irCqa9e//6M
y7FPztihhq1m7dkmvVW39o9W3ANVarTRxkCAfcV/TNdMTicrg51Nmlef9KEoktEi
Eh9X6b7s/4S5y+JYg/4ouujMfh7vmZdWF+7CVl1mvYhe6jqQy1dzpplOMU3ZMEnV
uPgpooVSnZOvi3cVwI45PkBQMLqHZJ+Bqp41v85FFcDPFVS5MmiYIiP6bYV1wJlA
O/wXv3cWgC7keNEMQX44oaFAaolnrDdwgES4WQrELYePrvlMF5jE3UGTUb8+Pdt8
fPUkxPbRdfEV8bk2A/sHGVHyjUbfvRSCmHUuMEoiIjV62zWXXtHhjQVXeBwTK1jd
XeayLY7+1ODum20S3azD3c7oXKtQy6dBCCiwx2YxHUIUt63lMX0yHhmYpJ5fhtNl
Zh+9p2eQBU0dC6/wSI3KrFLx16GNeNYQ0ANEG3BZtAOe2BN/YAofMVUviwgvz4pv
HVBVwlVunOPxcqJ0d6OgtsZMF6LZzrOJN3FLYjrIE8lUUAmnWAUQqyUcaeKxeVZR
A46mSNm6MbzzN3MiHCUvolh6UP4LbwbK//8MLd9e1bTmC1rlY/0X/Q/bg/19FNX2
8CP0K6aYzGKphMCRpp78VKPY2tUypire/mI8GiSi3K0onRfyfDJfQOxG1dLsxAjJ
d+IHClF1d6iodSgQG+kpiZAS5QkQGx/rekEJrn+4PHRR8hjiXGWu/+hIjmtOoeLf
mfrYNTn1TJG7a9r/16+tOf1e9+Ne8ZpS9/3iby5LBoIoYTe2w/lgCwTppMiUAqfi
X9btExSIdRTqBqE3yK/PNS2+Gi7JkDXxMA3P68OVSTguIqa7UAC2IimJLKMnC445
ouF0BIRV5+h0+pr8XMns7Q==
`pragma protect end_protected
