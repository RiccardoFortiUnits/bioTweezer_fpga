`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Gj/qc2FiT6detPSFTejs7+buI8dq3twZ+6wul3qbUFLRkCttYsqBQDHtewZupyhF
0QZ5we/gAFgMb+oOLJF98h9a/z5LRD6/z05/mOjhj8IwHsaJRLcS/JH/Ry8Gj6ue
QhD+bZ/B+1/SfVo5hS2aQumyzhSBNXDLu3mdkjaF4mM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7696)
NQ4qP+/PdeS561bczMKU3soe3MamEmdhPJv7+HxiadrS5sEY76mORWCKvEjjKqnH
KbUGNWn1NMeeAmp5KD8ZEKfCBdE0h54ihBbFoHFKl1p/c1EdrMjWzT5lw8z83aPH
7OrLy79lnkQoV+mdfps+0b9XGJGswJl1g6LnxOGgSTGVmt53PtrsglJzyQ5cE8/+
FgRuipf9W7az36lS1k0N8zivamxAKqGbJ0pskTmwWozWRISdYe5+FCmVK6AKO72K
a3Mzwi/gMt35rwxbAorblgDzFyTrKsZYSEyMPKk7YRaklb7gHNvWGO6ai51O5J/B
xYIQu0qp5oI4mHuv76p172n+4ij7Ck4lrgzIRGQCKCWRHH4oRcM5ON0GgtEeGXyp
UvkQeJjDxH1mLeu2U3vt9WFFWxOARXXZCfssch/bsQ5f1SU0tiEPsqOz6otzD5bG
XD4tsqsqlcy2VBhfTC9V9idmC6siUC8Wp8T5e8M3FHN6+prE9UUhJU+KSj2KbDrO
gxZKvapnJBMROMWXwo9cef7e9xz8C8bBxFkX9FH1fCCLVq0RMgYum0H7fqH+JK2M
U0x6jNEl6yGhMY88A2yDYfu7OCucPsp5e6aks7b7BJO/sXnWqASAnSeoKQpZ8uY/
wqbVgNMNAASMnkiEZYKcyarFVs8PywK/tB8w2vhrG8ZFZKQshDh4UVTlFQfnfyL9
aZkpqXaAySrL/zsAFxfTW5/Bxsw93bVHMpBE7nZeVkVhDZNGFjtRRwV9P73OqHQy
EZ3Lr2g44yMBQLkjYowensc3jfAw1o14JpCZ6Mg/cGy2Nb6ox3+gYTrIYbbtwome
aaLKMdqsos2SigY+q05sbvr8mvriIOzoz0qnfuRvW4sxzXjFBbUyoKPeDyw3AwhO
BreY3fau8NdMiZh/Qe6rhfdAV4OnS3pgWClCwLY05mTfsINS+zhHkM5Ijlbt1MEU
Ca4fa4HNKeUeWuNZoviOhx6swJS+S3T7XCF/nvpKCWbylnw4HHSArBs98sZv4CEd
5Vg2Fev1yU7yzDaxsYEM7aXProqzmAHniqkOLfhzqsz8O+O5kXoWnCaH1jceNjki
basg7jTbYeTGlafoP4p8lhN6K/RVNYmvrSCoVaszGSLdxhwEicoHFg97e7gNsrW9
MY9yib3Wq0VbLgx/rqG+H4gF10993cmqD9+4PmABFPQsXFMb2goTJeYSnm0yoYoC
Z1LOwUHv1TfyFNet598DZzK4WFlPZ0ECXABrb6g6qP+oFOLc3iwrfeXA0VKNK13s
muAjUieFnXWIhit4rB1EDcoCjVWg/Bm7o7SMfM2QyTDQr1zKIhT2QV34mzXfLhhl
MTJcuBnuj55B57nG2AGTcoungOwxDBJqMYFsaFRqxhhnU9reVIlKgpZ80vjlK3WF
0u9qkBlxeHftTJivvLxmso0hrPke9DcFVrWZe1WEp7O3+CKis3fE+KNs9is2Vio3
7kfMOPn7HUbyezQ/F0gLAu7Kux+SrNmrYoLjzuVQN1izUi0VEAW2FTTA0mYyoND2
JKyZSZZYxx4+xTsQ0zw5sSyo8x41FRZH7e6yZjIETrQwhNZW1kyombCoig3Wglwa
bIyHB7K3wVyTpiEgD2bS5s5yg5Qe0ADfegNP5aJWDk7ZAe4Hagn5gYAC5YtnAOxr
QaijB0kIBEvV2TTf/DeDD/LrBOy/B0CIipBRd6vldTBfof5K9PScPXVDOOF+XEeq
d44WWMiR3F070pYAdFECbL13gNR18pmIu6knSdM28otLxyz784Ane4U9tGlLZ58q
qxjsxx0+ySKJQ+bHifPLWoK1VQaqmrW0M/TTuzbOVgga6e7tEpvbvDYp0m4l3GXL
y4HHdkkjDB5zvlmR73BUJ7uYNftq5G3uBDMve90EzdOHgeg5iSQqlR51o8GN28hI
A8WUEdkRBf7yUa+q5eoaIul0K2VUe/4u8KV6bhyPrEWUTNUT9TYkttyWlM1dAFRR
Zd+DlcqF6xekoTVbEOhu42Fp2s4QNe4/JdtWCEt0jL6KdFXUzGN6BXghzv6bCxpV
oHj0WAfNkn03u2jgQaYxdLvrqQWZsxOl2Qq0GHIDwUGL+ijGrLtHZi4uxcix9RZT
Ad0okTfpnm/lFD7AxRFXDHPTVFMq0iI/tzmyECQE52g8wVy+L6tQjY/xvE9lOXsj
qB1C2ZWVxgPE4DiohtoiPpTw1o8Cpcg9D4gKZt5jiwfdeQazOtRR5p55/fFsg8ZH
lSJFWz6Tc7EeoSZzur/w/FK7hEdeOnJPuVyu3wwsCzurksWgoxJEu87E1zBfKsEw
VWtQ0eKnxc1LcDVEPZQXGdoYyUeMSV8wgbL8DhoDzxWIs9Cuse0QK/6nzhzxWuQB
y4eYBQzukQ45lJIBtT4Bp5Bi2Pm4Md/B4M2ge+lDnb3qfcJfL0PyjXqTx5BO6dUp
x1/94j9sN+DdI+7wBUm0tZInkRKU380ppLbWax6Xw5h2Afq2XJFv9mhrdyIkof81
HGTeKVmRAdCukdeBzi115xGJ/aWU0ZAQUeEtzQmnMLY8R8OIH6CbbZN1uyMsVg4H
2T9l+fASFBBtZoezsQwexsKiydSfwW6QkpZKSvhv6b2fwbnUjt2YBFM/7NpVso3c
NsbgTuJaMqqAMfn+N+XvT4+so4V/h1+RtZ4IFP9oToXnKhEzyPfbOdRDvDe/ApAT
em0fJtPQHrPB4GOUisvPk1CE9tosU0PV6HyzRN4wjcxB/+nZvzuBS+jYVhIc4Evn
tO20z2UkHFNTp/RhMgETi+SYnyyOxKQy2YkYZUDbnKDSoiGpV/8JN2fOGixmlJn2
udHlnYFYr8v+gooNdcIgSbtytcNQksoHtXm60j+nSbAK8AsXxDI/ka6fRIPWibaU
nI+7xF6j+xhErtn2OTwgzWzgTGq6odLtoOiPSXXZypuCigTHJXD/Zej0M3dC2quw
yvLN+poQ+X0ORE7SYllkbR5v0V4gaIqTnc+DJQvWXpsIcENL1MqzCMwkq9RqB0qF
NlxJIRZV3UJP2FrlZPWJ/qA1l9GYKHBpveK7au4+a67X156VbhssKG4nvKPab9Wc
F0eMcT07QRPFPAMn8c7G2WHmDRX79AWQFQwz4xu4a0LT8aAxe7xJKLIDtLq6wXwc
00v8BhmvCpLVaD6YS4QzjhJUqt6jKaOsHzl3XQ6dNzeYUCB4ZFc5V2l4V+2HXfmS
awmw11WC83hCxYQorg1uDgrA5LuqFYNBfrVJKZsvHgf6W1srEywoZ959uj+1ix/Y
E9zZjNFnSIulpfAMn0+he0tAUShM2b79SUzdKy0TYFuKM/vVuxlNmFmS4d8YvAlz
nqSooD+Fs0gLaYTTsBZG6QLa9nT57KpJfHJ+GQRDrAgyFtGh7TQeeyLWS5fgZKr0
GimpQKFuq8A7e2AXQImp+kNi0IC3AG6nwTHAnf9rbiv2SWEB1WM2sn3+qYmDQbWb
DnSpHPuu9mjjPlzDiGYsVFVhE6syIOUwky9706NkBjlCtK1VrAKKIRuflwsMmo2w
KaAOQqhh1LPLH7ttuP1vGbZgHUASs1Ris7bh0K2DK6ldg4vbHHjJ+G3cTeJ5QBCq
IYc9uaXK4CrBdaS23PoQf/+YeEvMYjBCBq3tnhexu+UDpH+NvK8Tey/BeIHYzuy4
PqnyTSq4vQh6loDWlS1ECSTm0hnBiW1YEo3o3++03wqU2VYkzDseyQmsCF8D3hJK
y7VBIrVffppKGqrEruZMhAb+DnuDylFCtgmfoXHmS6kQ9t7oTLDNIszcfd+OWjUt
CJMWUUSM4xXWvLHmt9hB9CadEuqqYjFYOcgZM9Z/JTdgDrKyWKE8gmYJiDiDSf5z
9VNRFsn5Wtsdf6xDtNUmh+nQ7egdizDiG9GY4re2crZ0wDmKB7mMrfWyDJ6Kio71
TaTvNCLolGTuFJ9MSm4VNsRhWfaf5/6OVdSVK0XRfC5ApoVXOQJoncVVJ1urGxj1
CN5rQvi3vfUBuTClha7P2CweLWC3Rq80SJQolWaYLutgIcmdrFTY09fsu7UgABGv
Vuz9ApWhaF8kBywuvz04WCSDxOCz2S6cxVflRkEYBNHY/jp3P4BfXb4FbcZVHrfF
mhv9kfWkrT1RVg9g47rARUjGCSpFYWWIwiArzi94rvHClO9FKHbxfDN95zvAco1o
i6ugX8pz27jYQHX/YsrrjaJ/jaYzFOh4tHu9kVNallv52EAaQVDaVTLxzl/2ID7l
malqUNFJhqk7jz68opkSJh4b0UfFKD/b7MiL3LNPgoDkYMURs30NWhtrFW25xYhx
UDumA96mDMazGZuE9Yk5kwlUELZGwGC0hZvnOBvEMPmNfNCzVPAbPjWD8rJTPHeK
fadwL86JGp6yGgJyKlxOj2cnvPh0pCfn+XVmnHtWs7iOszTtPExkbYaINxr6ztrU
2Dy4wPibOfU2DOd1gFaUoVLO9xvU77oMm3GzzvMFupCUD0Hn44kJoSPwcwAlFWOU
7xWMZWk0p15Ut0eF64tM9yhn1E8J6yVma8HPlEOsoYD3cagMl/+4I6v+X1GsR+C8
Vaxk5gRLmukUVIBW/V2bWx6vGf5ifafgTgCQ+95uCql05T90a43b7pH/i1r1pb2z
LPSFadoJQhH6NclgyRYNcEaX0UMPztyznI2oDFMZ2MKqpOaCSl3CUyXJcYvTUoo2
68zOrrqHT5VStmZLeDru90Uhoa+MgiaOjv6uK9guV0ZCF23N2ccIx2rkdeP7YTTh
em9f7famOU/20vVJYz62BZCBvO8/nIoekimjEoU+ufAmpyOFzunaspAymxFQzG2i
keEnpnHUgnpRFVxVFVE9G8+O4C+3ezSusDgmvRozmR789jxZWHTrVFZMgf2sYH2S
paRq0iKGvt8DTKyBqnUzJommrZrAZ8qk54quqCQHoP2dMb4+o0hnZQL9z34em4Yo
5j2GNqZyDm+8q+TJV/UTC+lpO8tW5hGNpM52PZDx/ccM9II2kSrT/o9YFJNQVVSr
wpwBr6e++iXVdXF8nWluGqjemc3o/4ZfCyhCUODllw826j+FWICedgf0eSWcR0xU
unWNxgBewaXnJa5HbUs8GYpeetZP3iYPcHidvB+8rSbOUAfZrUxyBm8qD9W1VwvI
XR0KsEPiNyeCnkLqcf+NyGSHG1xqReemBE3pDPbKvePjQYKAG16QQzvv66S2zppy
HIqGhb91y4425l/D0fjsC6cfIx/1HO1Lp11dM9b/Kt/wdMFPerSDb3rO1jw1Wk0B
O1/YW1sq1xjGOzRobcyuLK9ssElZDjmAtSYJr3OI34RO6iU+IoVnw0iX9Bhar2lb
y/WWvJbXfoTtkiuvtXtIa1xSYOnLwzL9za+9Np+YyOuQjE9z3LXQGMJbT6LYKobU
IKZEFEzBIpKLx5lnXXabvkd7TpNdXi/vIMSTVbsLSfqXN5wKfxWni1xmTqWYXQxV
PBBF+3pgDJpz0fGypmVwNiq1jqKH26aPKMQnBGkeXXiTw6CFnozSQkGpu4WLfyNV
C2P+QGLH1ZLx/f/o19gbMXdAX27CIWRerh9pUpBLYIeykSihMrznE8FTZ4JlGrbi
ad8eUSHyVyFj2v36/B7415bjW80t0Jv16A5ptgHJBsUOGF4e+wEPH++h+aLiFH7k
IKYUOVzu+9M7kH4FkFdhuYSe7Y6HybPvxZeDN73bWSRf+zlXcqlJo3QxqPAJUww/
yYucrUfM/wxrZlRV0TjfRppcdjIqSjeyV1rzX7ry3BEveG5oznwSyZgWqUdssmyO
yqhs9CEVWklyS0lNSJShc5kHRsKfoaZMO22eY15/MDB/SzHQMGd5tuotqQ3nnWjF
mZMQT6H9sieMIiCV9kzqRi5wdtb9Vf+AONpVNxQCFhsPn8xdrMu7JOSUKUQyeXy7
kRWYfw/v2uYK1chzyA9Sq6N6u7VQfXueJy6A1JCcHL+UHXzbGQi+xbAvboebcdZD
tOrpbAQ0IGLlMOCsVYibQnijHP6titSnV5s3UE5hfQqmQuz+ycbV+ftdDl4ctrom
lwFM2jcaVxYiEbeODIbs5Be+Ed5LAVnWjtcyfKLywpSdiNljrxRcc5UqI/5LYkXI
yZzed7rc2BFazmB98rQmhWcMzNbeSyEVsifPRb/q5bik/OXfypT4TtoDyEYWvOqJ
h0d8bh7q//Q6g1gw027iVX2YRWiXqmGdXHByHGvAk4eemQ89rW5tUmN5STx37XKO
fIoZb/FC4LVVsvk8hdwqs0a66HR/y9/V2S4ELxVotd4gWi7A0U6AM1MkojKdjenC
qokq6ndcAA4qRsgKQfmHZuw4JQTEDY6rUpPD5Iz4bUQEaSHnjdXd0ZqgTgPY07XG
s1mDsKc3NC1i9uw1jY3PoZXQnBKRM1AsuI7NYObGevXCQr9zZA4FPCOGpin+Ke85
ya5f8F/FVn4MUXq5ZMUHTd82Bw8AxLMVWe/erBhDrH2r9kRU7BKrcIwlNXW+tW4D
rEGdfYjlL0cxAND7+cRBJVCaYNuqVUx4Lft6EisYNWlUSy1G32GtgrKGlGyVwPYR
ZMgeYqMr4l52GcW1FEuGN+Jo0HhMB4Pe5AHy6H2X8BiePviqv8mDrxvgogplxD/e
fCQ/PRPTfGtKx80pfiuW9nqBZZ0fRn4bk5WCaGHBt1Y8QgVdLfuGBDEndgEwIUFR
zIt6MSJe8YwU1MkIsvNd9BsSm0yWUoW8ZkyWqw7hmnwzHBhy38gOHDQbyt3xBPqp
U0hD0pNQIPdybDZQehQp37Kyj3N1iEvHl8Z2jw5qckg1wYrO9gUlhjmWczD2dhDj
lfvq5L+xO+KOWkgOoxOE0xaB1cUvAAV3DYoIY5a2YiLH6OnzQH9OL97GzTZBdMGr
/r4eI7UXAUEm7Cp07lR01hQNFcQIEDEg6QIv4pvdiVk19tfaDkVabchJ4pfesjaC
ZRMHpU8qq2wM8H6OAzRJCgCSF70gn59f/q3/NUWTX7iuMhYPVzVAv/532ZdeczWe
CgOCnSKB0aRDUlAZgzuaVtIDCG4kfaJTjPVw3A4pveyfWBjvUlG1rSCWcicNuZb9
ICzQ13tSdPvmdN31dyBmFOnD0TziezjbJziTLSWTlvk7tsPAl6umBvKMDk9nvywL
n7vvPvm6c2rpcPZUmA/H8rJF2HEM4dRna+XTt4nJHhr6nt5Lo5TjTvlNy+NAP0dE
aIjSqrA3CD8nNJaPSEcJrZaU0PwlTKOIxvwoFEage8GvUlGaFOW71uzxJVshE0Ds
jDazgN7PjeZaWbJCBpXgnDQbZinTGKqqTovggUrFQ7tC1ZNH4wb1funrzhNHhyGc
B0iIeRCJaKWQ9jwF9YvHg3uPzqLL6VUi1Ckji0npWyWkXvLb34OQqLe5CLzjWmjE
FevuFuntBh3audJaTdl+jwNMH7Nqwyk2wezca7kq8rvIISEdDLPt4+Fpdg4IoV80
pMrcrt2ml/negGUjcShREJpckyhooG6dnr6AnOoV7d3NQ7o7Asu2HxU+zVhu9376
H3rfMJICfuXYJi1EKPxmfV752NZtShf3CqGp6iX3sNMZ+iNylgFqoaBEi+cRc40t
C/jdKWYbOy3K2FUCaEXda2ss2HMM1CV9+639Koj/xk9KcYC12WVaN8jaNGnKlG1g
bax2/az2pAc4SEQb45jLsIZqIeVfOi1xPuCT4ZJtoecpGbctD49w0F/SNcJ1iJGg
axE+VTzfjzJRlKy+WzYXTxcAeHoq19tcRC/PjG8hBVXQ2LiJbe/Vdj6Y4kV+gtHa
qeP4xcRRICdGW8aqx70q03fvMgqdaRhGrDuaDLONzKvy3fQJ7u295oXxVFMjGmw2
x/vrg3ndJS060MjKN+X+FyIY1SXjhxL0q22rzH0LEGb2qrMY1L8iEUDM+2gckZCV
0fY9hMpzIkXueTOXQkmy9Jk9LGF5HvixYIvhjjJ7XVzIqL2p0rJ/gy/Zmm50UG9G
wY/rjncR+01jtvCUTaxnXExFjiVggcZhK6HN4iolrBVrascEe57RGlP/4/FNx1zu
8hSPRBfh+tvqF+CgnNzW+/7QLdG6p7aB0PLhVVqHXEf/sKVfotKb0xQG+D/4TFnr
gIlj5gN6BMheuOMB0px22ENmzLyPewZOlc+vXBI+MGAfA/yy8YSgpru9isFz3eK5
+CE22UiVguJap+7CDlkHd+1xI7imqPLG48ChhtbzWkfJi9nsHp3RJf5jSjNBU7cT
0DujlobQYIYEEj0aFNmiofC9THaVQF+cxPTlrx8ZJLhvoOnzN+GeuKIuiCFeRhPc
KfaMRTcpYdxhB/Ah3LD2L5A6Odl6N6em1WCFbZFVqUe/nI8SknhTQmtKJwwrda2A
bn0OISLKbsSCzvLIaPO+If+sADEKYSmYU/Lu85JKAaPFc1TRbnFCWHTuNz0Lp+k+
gf6D7/osV1mcQQs75+eSOGbfiMSKQZXn6HbQAa5R4mUBkqJpAW1WcOJoAkYEpjWe
AC0pybEHzcXnPL4aQ7XTKRMmnktuUmAPyvqKQScw1NMFXpB+4c5i3QOW3jWHINfp
g6+cjs66QQ0dRf9rU1zDuS21J9gpGIaRdyr9LBH3rSPs/c7oTT0BMEZrMUKNppON
3XbX1EbK2RIsfQelIt3ABm0hjnnwRg19EfCrKl8TLYht/gtQRP/3uYx8YRl/ohbs
REhl+Tb6lbRWKXsE+B7Iynw7caHznL/hvK2kvxd9M0oJEjWfE5BTezMiqnDiYd8e
XSa/TPoDZP4NFt1AhpwwfpWdVu5+4vFuarhPFf6gr20uAZeanIep2cg6IcC1SwDS
lUio92mj7ABe9vqrmuLuC0nN165eGdy87IMo0RWNlfwjPlr9/DGOtZWDX1dt62aK
eGvLvujOrvOQGsGGdEsvU5AGkog5/IvR2arWU6qEgoC2xIZf9teqsuJou8X/8DNN
k2Z5TTJdJB89s1Nt589x5fPRKMs1zopUo5PxqmlltoUU1wUPQLuhw5OA91fWPSkj
CDvvfkQ9NeJomcfNrIaLJSt8d7llrcqbI3DPmLIwAGo13XOMszuy94iHiBAEq/S2
u8+E3t2r30k/ldiaNJ0Ip/CUKtEXI0UwZfqRRpE0kkF6dz/FBtvS+vCaqZ5SSBA4
N1qi8PPKhAzc943mWu9ipfwh+4Y0bUUpJwtsltarKDV6tbSYhHxLPUdrGmsgIo9X
++eXXnnLcIJ6FKhywuMHXnyYis2dlHfUP958XDm3L6l9olJSe5k/U45WO3mAGFu4
i9vtxBBdfFdPB/kWfE01qbcNdAdDUewk7gy+E/+y+FIMNecHY8N2ynzWlcmX8bl2
u+ba85NdQKfy3GrPlCKDoqODcuWNK5GICsmTOB7HukNtmXQLX+utPGhL/hXMyqia
FkYahXPBRuZoCcxkWQoKjC8SO+yRcm02ZdU6k8LOTFN6bFWRopf0JcG5TOs8JpnN
wHeCEy/9cGGE1m1XhMZuiFEAPB/sRlov3sOlWxAF4+JbVyXIMbDTmdS1qT71qdBt
gxOX46ZrmUsF+vXklENwQ1iEXURDgZ4+ozAaf4EzYhJtXBZVKSJa4Z2NMfc+sdQE
qqX9VwXAW0famipyhbj3xclPfqOjrXQ67gH+CCq5r5CSrzlob/5esoDLrj6VCQ8s
0EZisZo5UUXkCQRXLT+w2OOeNx6RVl8k4/X9brRZB7OjDTS7DBhZw8Rdqd9c2oSc
tYgaIxi7bBEUIqPr6k6ZDajx9bejnpzWI113dBcTDL2svto92j5NyOoTLk/0+f6K
t1fi6TIFuOZCY+WsLXaBxwlwBdFebxjYt7XXKaZ9e+30qd2Zbzrh5w7zQMhEjiAw
s4HRv0AF6QvSZEqOSc6YFDSHmT1rfIYctLUvx+fpYK5WU/jsJKbb+8YwKbbaGjJd
X7Cn64Q7MMwUf+delTt3N0+O8uHiIGirTIXlPO5QI8B0qEBT6v12j44pCupq8M9J
BFSD7tfn98G3KCXnsipKzgt62lZyigBHnO2zB+1KwIZfcv7k5ok6vsYqaGRaItEC
UdTWYX5tgcRpduIA9D5/r19rL4TWiaNvt34Lhf4T7FHTnSXfjUV/MlY/kCh51bZy
ysqKxgQk83gLpJ4iot1uSVpSERFzdZ0wYtYE97XMV412GT7F5x4OqCn6KQtFc3f2
MqTOLbYNtndQlPuMOImieip6+LQWiE6WU2oXq/9AwIAcb2k88owAJ9wsygQ6b66Q
jdxaY8oTFZSqhOE+Pywz251NvN8nVWMSIcY+n49BJ3a/DDu1W4kU6pQ4Img1RiV0
vTwoolmHXMkWtkV8kARmJQ==
`pragma protect end_protected
