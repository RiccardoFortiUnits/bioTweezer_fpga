`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BrO0/Fo1ErDQJ7F4h0PELo/2wwKoQe1d5FGxq/vnzdZMWzbRjzzcCf8zoFtjhx8S
V2ROh73YtPy92wbo15hIMbiS9Lfeos7jnjP50GwkwUal0n2TzEedseWdaA/ZGkej
krASXj322zUylujtzLB7RRbEdZ3mlpN0ChlswGpq1Ro=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28160)
7cjfOGssy+XW9/feVaIHEMsiU7G1wgwXV5hk4sEcC8pq+Des2JknJRyOG5+zgsxf
A5OqbQcrfaLvcQStKHwiqszFbY+yvMY2TfmnVVohWG8wKnfYDNHznCURDZv/j/Oi
w3GHZ4OhaMv3QYmFG3/jnIYTd3TNg+V9RioWnIif8o0Y0129QaPqJpK6xm45LPgd
F9p8Xh+47P5JMPZ2pfQnhJbWkIExRC6ObqQrlsn0AduV+/xhan2+9nHF++5+i8WV
rHj2f5GBHUEvk2fRSFQi8xV0grv+TiL+biWgkw4wMLAnF7V45tJPpQ9mU9BoH+Br
KsPZaLZfAYd9N9xS+gbS56NAdfdNjUl3BTe8VuFdV3shbUf8QoLTG29ZnpDurlLv
NLec0HkevpXxdV3QQ/+hTMuJTOOKu8m7/WcSLJNdEADeDHf0IRUBsSs0fdqyfVwb
FF0lcLPwk1r0aA0GcbTkxX/cck6qJc0/NjwBcUmVHYfg1HLXlm7WAgAJoOGZgOFw
X69HFiVyt6qdd0HXs7yPwrFEOXR6CBW3h0SNO+zL2XKMF3eeEMHOIuZuB8mjMKc3
wbeQo7dE2hV7Dqm79a9oYi7Z5PpImFiw29/DeOKSDw5XcoLrdyTM55lj63K7UbE4
Et47m2kjLUAaqIB4JWSRI/04q2gept0dEK4zt80Fg9v22vfR/4A24glrBfzHKmJN
b1nIA7WDcx6FWRDbqQXrEiE9CGi06Ti+Eo+EOeQ+6y00s/tDnSHhCeHxhF9L0mk2
1XfUS87a9LlsefSpTGfuVBHWLf/szEs5E2IeEEipYnE94OxJ0yA/ErgpWfmujto6
5nM12n2irJ36zbJ2y2VTRc5LHvrQrFYrVrpwM3PfxU4xJYut8WJz3GP38dhR82Sz
G+G64q8AjmxCMAD04wTiXPD3LIL2zEnK5ZJtwcsiq8+Z9B1co9T35NuE86ElX/Nv
NpWu6V0xFey4quhCZye4XQ8feqRyicQCdIpOEdh1qLx6YjH1l4W4PZUmdZXFeMAB
xdrKT+uAcWSLArSZoywJsmQh5inGG9V4b3a7Uc1OpFYpwpENRAwRY9Ndftf4EvRk
Qv34UcYU0VlomCpO5F/OM8vOQKK0Kx69VcsagZHxS0hOj3HumkYqWhyjE8CvrS7M
FDsUMkKmYLgOG8Zku+vTWMhGWHlM21bCSHv7xkhhSKD3lzuX9zluCHiRa0k/76Ga
+VUSy52+nriHuk1m0Fh+VDfsSV5Sxk/PAIL09njxxR4ODUm6Y6CDkh/H4VqijsGr
G1rMG3OHm3CJveUvJuqmdM1BKavtvuzV1UKmlx8nk14QRUNaiHAtVz9UxTyNLlAw
/HXsnzriM/LNYbt/2vjeDoQaRFD8maoTAWscr2tS+Lm132NNPQSo+unl47k0a6aO
xc8VaAS8GApNX6l9p7rOoKt53pJ/tli12pCWhUQ8gtt/pIE49Oa35vTlVUETY9cH
R/AElZ7gaXQUhzBD9MF4W4Ff9KoysAnWh2FI9F4nIbsQfAWuu+PkMcQb/nqutsZz
+KrproC/RS09Q9Wz5uxbCud88P/omIxAEjrbYurr2GYDHXkNcJ+jMZ4aCtUTkqTu
Vf3Vbr1Pt1HJQL/ytBY9uTmWeHUFu939Il+tfX8a5QHltbwetbrLSg5o7QfVzUvn
1C+43rhWpfxBiWjlCP/iPtLDeS7J/ubQPxYruDQ0K+yCw/HGvKA5LhPUH54v3SxY
yo5+u59F2qp4KG/iYwxGVTgvY3LU1wcZ33v2tGSJEZ49XXUK8t6HMqvfNGoYgj0i
FPzKWoCKExTNAYbQ2KuC9XqHV3rnAb7MfR9pnfIiT9LXU2do0T3Z6TD66zcpc8wC
yGmbZpQFvXvOyzm2tArxYzFldAvlmeD5bvhXMflGQulO0W9Yug2C4oRIz0Ut5va8
tkf8JqetYsRDOPVOpwrKpLGeweyc6ygoa0xtC0faJW8d2CR158NTuhwMTgS1bR2r
u/peB/fGROk4KubGFaHSIZNyKzSGDQkmCrk2zf/Bh94G64ewSI9C4+xx7vhI2KU8
cgmJQ59KGqosW7SQFPy1q8TMm5CzPKjf5moGb/50A1uSjklGymJim0NhyISYb8XT
gBZQOiWRYXxUHyINXVcwWsZ/K2F/iA/RzQuyjU8uVTN0yYugN8Z+bMg5v/8xBzWJ
Su++pKHIejoCd6EZ2nVtPclBcfAf/ZDJBjP66bnp3pfg2gdk6iJHFmiQBu2y5P8m
lTQGUN/BXukbzqu9UkzX/93VM0n8LtkWAN2f1tciB4hEFHPjX2Ec0FMaCO7EeNzb
2a52zRwp29BLwH1KSMAs7WPQRNAYOJDS3z8CozjVh8/Ufz6RcbZO8cU5hWe29ZzU
7CLVRDL3KAyDzqngR+m3JKTBOIKwb/0y10LlSVreuB6asZwfSjU6vOFuqXc3nn46
EmuJ/jJHhEhSAqnnNYyXeIXjAiHH9ZUQUyTclgZxLYfLMM801libUI7396Ri98U+
1a5eylMvmvMAqLDMgD+eJRgHBV9Alisw/4Pv6LHgOnL6yMeICq/M5wHq0AHXTHn9
tA1qzmt6bWiIhrOnWKJNmZZqFnTW0rgTV5gFPwE+MwEM6/RLUJGe3qs6TiFORNAf
lLmbbSgWHkZ6bJ07jcyCOtP3z5DYdGD7BIYK0ZHMA7LYHCCIvF/CA8UougMORRdf
y9QI7faC3pHKQLqdDWPCZZ72LoR4319sOrsMtT/itygYF59mLBUBlPJDuhqWeIl4
qMsruHI5q/FVwn19VIarMB1h7vNE0xEOVJLvjeMNwoB6XbQCwZLCHPSfL60dmnqH
vGqHF6esjuV5W4jVXuT/8pa3fK2YBqB+zxD2eZ7Zv/VsqDWFj1rlZ2PZP39Hte4d
tFN1ogEKDy8pKJCY0p9PHzbTXVlYyacUOEQ53BmFF1nnEXyTPx4pd4uSg2gwIqQt
aCNfWMfHzjCeq6gLR9MJg/KeFc6gM0UnohXx0aFyNMHgWkqzN5gZb3/m2Lv0UlCO
1XGk1IsNBNnRjBMXsxnHtk08ScMIK1enREn16mBl1Ei/tqIcpYVfyzMie4iNBB/H
ObGBiAxn/vHw0PR6/qX/eZ1ibT7cVkv9ghPXECA3iDLA32RgNcuhhfHPVXUCIKQY
zqZLoWZmmavpwFAGzlJ+PX//6rpkkgShNlkMH6ChQ3eN2iyVJf76cAkPw6fa/wRl
ombzxo4XYttaspTitOyZVvVNztzlD6gHIhkkv1Of1TeQusOJugGeUcHhBRMZt3AK
+clXisIGfs7zL5LpTYhIL1LcH3AX3hrk93HIB09WlqGZc8kTJ63C+6PmCnBz3Sk8
Yr/WS+bNRhDkIXAL28L4B/SawNjKaBq1hhrPsAK7hT//RT39WlCOJIcsVLvMn7Qd
Fuy6SRVawtFeQl9F83FqduTBNukYtn8dYhx/jg128c91OMZYuywk3LwMb/jV/Z0g
JNuSXAw+Cud5TR7dPHYWo4BDy/iKMY4ylAs5Wc7dcZidpNi0lA47wT8Y8lqHwmkj
9VXQ3+RWtEO9ZMi1TmDNG4qwKYePek+c/jPKsj9RE96JsjFRABFKrJAj01JF6Zq4
l6h6hUrh1obAresN7IvJgSE63KBEO0dMBMApEtXcpNdFOPF9LKaHnuW1GPAyIwvl
NrEo84FJEmhHrt1ZrDhyXhs21NoBrEP0uFQztegUUst0GXePs8If9YQM/sFHC14H
VEOXfg0kMxSDRy6p/Jl3u8L8SAva1k9S9XlT3BArJ4vLhdpthGwbkmodOWFJQXuQ
40hUsAhJGdqcsSF1W6L3Wrl5YhVaCjCYcLEZDT7KuXfGfP0ulgNu4ShdHe4eFomb
JyZA3lUdeOw1BmSgpFdhwv20AW0PHajlgCQqAZvvQrKPfFqfgcwtfhQeqfP1yC5+
XMLQK6dG7m1ZdMjBJBErF0CiQVQ876Dty0zVJ1yFzowOT5HIp2U8BNC0sCNWc6qt
x556GuiqBxzQ37nUPgrkmdCYZAW+/LfrUn79svtMTBbc2hIlhtaoIkbhD5Wp4cMp
+qDNy4xpaUII/vRKHIWpm6e1aZbY5dz5gYnoZrZy/qq6aWZ9AaTq+tmj2uT/m7pk
cF8zdl5ShdSZCnmE1HbTszzQDNNNppGxdFHl1CPg6cJUksBojdBjZTyn8nhHz/k5
+7OjSnzlN/PGXXW9oOgYQHWLsSAVck/yXYGbJ+oi/p5RBL22WX3X8o/I3N9zs4gp
3cznPHlofB9OQ7UpmhCZZQknzPHWbK1KqOfdqjW0E20G45P2KNpMCVvITx4uyJGm
M2FcYQbYpCJP7FSBu/pPxyH4nZ7J8WrTh9aHygbwvwTHLrF/66HChH2V83/7a/h+
OdYEWAd1xEKX/XojsIvWWOY4odf3js2Qrw7J0jM6Jp+8xX7g0wXBNxDrJP/wZgVj
7+0LpXPhAy5qk/eTtTzg93F9awjBu3UbahUvvIskOWZdT1Gm1dovYcG0IlYr5myv
GIa12GEh6qCgcOeQU+NNgfNBfkwiOO7RrcPdsgQTASo1kiPC9P5M5o+KwQkI2C5U
I08PPdb9MkSR34V5M7h7sYrsERz5hxj1OGBpZcz7mw4n4OBZz37V2lpzrLBZhrU0
VRUaw95MKjnn/BaFr1bQ85hAAlPS44M+IRLsyZptqvVdxqLgcES7pzn/gzgRnxWD
6ehX2QYHAAT23myiqo9xrEcsX9mUki56poZVipl5rECXyalsx+YHShmh/QFEMGM9
VFZMEtM2nvgWz4Q4dtUT/S9iLHl139bKEfqSqMYjxhEKdDjZedUgTG6WpGTgTkub
LL7uJ2T04s6QbSJx7m0dZ0tbl+cQ7o1K/UZhJzHfMbQ70/ZiLB1h+jfkE35f0aTn
1dAWMaQHsIa07H4PxB4PkHM41SkmwR0Zh5JUIock8NXApO/T3pQbi3JNobgRlvtH
ZUaIPjQecgR8hWI831nQmR0lLWtlqi1pTSeP/tX9iJW/ulDdMDVeafbOLhkFmTf7
ya1wOZgzQGonznfZxv29a/W/Pv5uWYJ3kpYK8pukI42bAthEzF8DVYwY6Lb2wBiv
lW0fVh9IXUmLwVcA9oYFMyRhemkqXNoIzSSeC29FwoVxFBgXC0fWt1zLgILTlvBA
72t4vq5NWoumYTPK3yumv9t0jL+YnnFAHoBwy6EXZic9u9gaTNSf3M01rbwcqZ7p
KuWmyQaNHTEVWc3Os0YAvsjqGjYYbCkhqnqXggzq5H8imRNJGzWX22izUvd6M/Xm
Da+APiawNqbifwEajtyC4FB+viTg4YSwGujoQGSV33++lwN7OImn61VfGHUEqAyq
TP6KUH+TRuOhpjs9nUS9Vy3mtCZ+2stiyZ7kunr+cmqss45f2G1I9btV4/WqAqeg
du9e3tDCxKgz+PlAh5NCIrfsOpDT/ARFHIEWVLVt2t/FCN8OzwHZJB5Oczf6Ioh7
+dCuMJ6z6BW2vtBhNp+efF7nofwo8h6+JihB+bEYHKfcR6HzD5HYrXh6ls60YtLQ
7BhWwkFbQ4wdDU0ynNwIzf8+uN+jJM5YCxFzkyr3oEQ6gLKcNZWyD+0uAZR6vxoN
TIep1C2TCV8UiCrmOVOsWpquRQTj+9UqcXLdXhn5q7EScoFaGfPkGQykBopRa2rm
bmnT9WIeRPXML6fQPWOK2JfWlA1BZ8LpRXxbaX6VleMzV8nDKtO08sEcOFNTZhNI
qy6G2mvkrCRDsc+iGQxMdzm7IdMODKxbq8Jovn9mxus2oKmh9yToEWjS7clPSOjt
RecvVdrY7xhAnksiyAoLjSh76A8NSTWc9W2qDhlEMxWO9ASpJwp6weN3AGwUQw/o
6o+v4HKYsoHMebapx1YIMtQXvayXsUgLcG29itOo6dESby5/6UwH6RX5sBhT66Mp
jz2uH2jILZyUp5wriRwaYI1eTijw3j6lwhbGnIj7pRXdaRWF+0ycZJgHAzhozlDJ
bhGZ33JiXWFDdtsnB2zJ40IYhreMjo39PLDHcIPMw2mcb6SMcP988ifPK3i7l1LR
+Rk5CDCkqiT4La1LXbOkshD9xrTv5nTjA6dca+tczCZ8FsUQomcj7A3uqv7P1oXQ
sbURZvvHuZFPeDyEYTXDvEUYuVLnv6xCXhOhWWm4Ik6IAtMCSoCcjJOXpRYxQ4Rd
jYzEs0fnOMktzSxCS5PdLgl9xyrybV738f8BanVeGe1WXofGQN3YUYLp+hq7rWuJ
oGtd02j4TGZ/jBoDT3P9Ko/6nzVSm9Ovl5EcyZqE0v4kqwpj+gLE8rIqWMb9veui
inaej+bFiDvjZQxu4e5axIngN+x0icp0GrYorhUPoEDw0JKKUMO4IAURuUFx5abw
x97i/OUP6sZrrkS1tTo/zjshLzkUwA0IX6EuaJ3umHbOswwt/0eTkpss/N7DrFBa
qnphM0M4mw3AtM1LORuWKMo9xyJzKiYpxkfoaYBuwQmonUNTHFnHhsXaYmWhxghk
2Zn905AF57NQ7+3opfBij494dMJuAmdqsrB/q9/iXXr7IUc2S4PEE8HWw/dbuhRG
MbCNdMMZJDVfnD5fjUYI+VDPk0DuxPqQi37YiCSqADp/mb+BHl2s09Up5CqRyN+4
NUM5ikXIfpjpma5mPGUS1JwNZzbR+J9256N7gmL0pGqURVnCxsVbqsM6QXA/+fBt
YW+xmX8GoRbFoH2WhjX9s+Zz6TEqHoiUGjnyIU8ZzL1cnJqqK2feBu2MBNEP68Kw
NFxQtI0pM20E6GblyoXl8yKdEXCD/elRQi0C/Oexlh8T7jZB3/sf2QNWGYv9dYok
4jbN1FIwj5TdLhfpQX+FGdnTJ6tOzf395enew7vgZPQ0VVncUWfu8RbT6i3HPLbH
ZqrUp7PNJhSW9evwCjWvQiQHXEZfbF7tg7A16cHRp723NaGuks7t1lqb6xZaRkhT
D0/1owBoRNpCRV2t0419CXj/PSchn7OWi7EECgh/Kh9NDXmocXbf9e2lFbtE61JE
cZOyJ8EYF62Lpsx1LTObn8a/+JIKAJUArJ6CraguZXjamur4knqU9wSEtuRjZ5Rg
LTWCQCwqxSwEFan1DP+T3xMSSRZrPtzdSMwo6eTQPlSi3JFdx3sf7NtaiSVFPGgO
6myz9gResg16VjliHDJ9N5fAsdYIw8ZNa5cCZU2agyhCIk641efhaCqcYOV3uu/Z
A3wfLDlqEoZnn9OF6hCPbQZG02ET7dvMkWXWj058u322+nrSVxCdjSxUDqukBGQa
eTPMzKRDYUzmifiIM4mI+NDsq/JPqLYVGLFXDqGBmO3DYSeSS2q3uZrJAj7LSOGR
H8NH5Spf3e5BMN4rzHosL/fqvK6iiZLDoWo3KCkhkpSiWPvZbpmOpNHI92/NCSSK
R2f7iA+Euh59QSn3Wu3NBU3KEocnNcUJW+VeDfGQl/MLDxtu4PLjDI2Yvdg1aJMy
rvale5CO9Cznvf9bJycGtjT/jHqnLnkaEtc96FsiOMyWCeZF6PslHFU6mpimzL9Z
2EDNKihn4ZPnfGibmzwHIsPZ2IKYugsTXRlIFsLLoa6hcIiC/B0togGKe2afOI94
FtZ3XEX8r7ejcxiQbQZC/63rSm5apY1aXFbYwF1P8ISMj0qYm9shYihGlI4zAt2E
5AMYY6mVRQmrmh/2BbagSeDd6Lyo2q42R9Q+DPBelDU7qfN1e3l+cBxXDo8gNgRH
5pO0fonP0cCXPPJA/xPP/a/xX8L5e8e190V+FbSU0HFLkRk/52l/L301u/KocHvh
2ZqtrgUnK3htU3f0LMMVSkWEuMtZYKhvF5W6/op2PtQf1cDQEiVG+aqsEZB7bfXb
U5GZQjAwh0L6SvELZkZA6W10L3U+G/MAImpsCNVfq6VBxjP4nRrCWzAPdSJ1n0en
L1CpJorXPt1pQikKkwm/3dssqlOKx2h8xO8Pwalh2BDXxQDrDzpMEm9oR5gzZJor
yjGPYAsTQSocLdoVUA7SIODhE7tACjsJ5W2cmQx0yl/oYJ/Tkyx9O+kqkLamZ8+A
wNIrdvn/3zW4Lut+jkOxxx9oga8svEgNYTkoiMELfQBEoMkCJqtVVrW0HW6HTqg6
Ja4WyoXpS8ZPq/xG3NqlqjjpGGVJDFb/9wOoEQY39x2bEtHz0qST+4zCNwjVD6uK
senhGAgvfK8s3HMsFt/qW2NYOtgJXgKI+XiqMom+4BbWQzeFo0+wCmeJKl+jJzo2
824yRQfMAcfDZZB65Z+n/Q/7cOmpfPcW2wrY9mXUZ4FwQ32bTuLAOhLrYfY60Ugo
X+8Watt3n1vvaiLcrk20wokSNBd/3dJJ9UXMIY4M9KuM0E2yY1Yy25u0MiUmo3dD
llTib6n96uN3OYzqkf6vrrYURKidVE4gmTvlbzdneNZjtNWyNZXpGZ2AJZqpriqt
Sxddtt+JZFzJKRlBACVFLOsNgQQzYr5zAQhBJGlXghU15b2NeVP1r8PVV7lcJ1Xx
VmBFQKEPhiXT7UsAyft/8YJafeb5FovxgDi8Ylx0FA+qB9fUJFTWxbFZZhR28XRS
u/s0Lro2G1R05VjlZtSxmOajv/DAumCL2YagfpkK5m8uIS/p/MCTXG3BNTy+vSpq
sIL0+iL1IDd+MOwZet99RB+MFl7Q0jraQ0RvmyjfBxCL/hjUao2YVIAa19S36xSQ
D3OrXupY1Oi18kpgk9Vk4+u2OTBRFFDaMttPsU6ea0HtFvyQV08cqXCL8Vf9rhJa
l0GYaH/1x1oa35QATLMsqjEkjbdcHKQEwDQFxBHbuksj2SOxDijgLp9XWma8q5LK
2kS/bf454wopFwkslWY5J3PhxxRf07f7ZpU2cSmQl6yq6P4xGAJi/tVfnXrPhBbb
1BZ8BImvnvcUoUKLBhRhJzOt99PHqYcqQlHfW6OfvnC2OJmbfADlsqyAU82gGk0G
2GfKuJdElb1bNFhe0GRLUaEnnesX9CjO7DvbHT/i1gUJrbY9xt9Y9qLom7q9Rk6y
YbLZbcFHbtYvfRZRigQkhCrR01WAG4xQGLhPzflCPnIaFsHo0k3WLyQYC+ZFI2/m
Q5PUPZnr589Fx90dcMXzeSNQnE4pkmxxFgyzvC9MUGZbXgnLjFvAPyk8VjOd173P
OuUJrl4hHD1Hx5EQ7OKLpoBI/cttiWoHtJUVPrIQWwF7TDdahFEL1cu4cRCKnbbe
r+Ga5ru5kF2blmGkl9QxJpiwltMmnro0at2RwEwVnnH5epjMJ5H7fovG/ZZN6zoR
TXNvBHPVhXLk99q0gUfzzMQ5J8LzJHmc7BAA1hbkMkOpw05N3QANd1nFOs2IkbaG
9yRe/lR3yF6m7uDnku8bWxzkC6TdkfOu3UGrBjpiNyWYwEWU8WiLxzyGcZcmcPpe
pC+AKp+kQCyX/uX5CItbJLYGQW/wEmoony71Jp8uGxwPN0qwoNfOfYN+cL9mbQRV
FGqw9GJOZ3ChOLu9+xaCUqG9cPMgC91Ur2y5zDgjSuDVM1pAQJvg071cWvFwEPxr
gYhk5+kJYd0wVyAS1nflSw0KjRPlMXqq5LtwLkr9LzaUqf+QSMDLTymihKmGz2/N
q+JgesqS3XPpX0g2rYPC2BejrM+2YD/FW9Z1HSbX1iM2tKrXmnew6Q9cKmfod0aP
ZcWAiEPJ+dtKUIX25SfG3CP3s0q3eGN1CRLj/GQjvKgkYymVKiRoaHy2WvHYTn0J
TnCyvTAMAUKRwuXsQqzEXG69oF4qTLQmCurHODfNTBoyVyZSUt/82jXb38jatge1
1KkkJKv6yD4AWOGeTZdMroY9dTBd/SeXfe0/naYymlVwNQZR+2gBb3sjrejoIo98
HCnKn+EG3AqWO4j0h0DpsNLCKzM9tzCbHEI0zgltu9nxSiZdPe8/NgxEXbAnXZFV
0JcDEMlqYnRdCZOxLGw8zdDmxsOUGwNtkg9HVmcm605iLIhiR4vsfQW9/irjBOIc
g58h96S+rDmSxC5jWRwPrtItxczjT7cXMdsxyj4+aopKG1WI4X1RPSaIjM1hF5H7
10oxRyaTRgShdgiEsTA8PSWdOYCkLvCztmZv6tRKO1YIqWbqMkK1Lbmi/0Z5Fdyc
1fqvcjdBd7g56DuQwMlXrO9g5Ga/mjbcwN+YXniU8X6yyqhTeN1jh7FIa/umRLAY
mfwjrcTe7zR6ycv+lH1TcDTUv+QMCUklPSCMtAuhNFc35Ud0OiKu7eoeOReBHpVM
nMfSDdaY8rlhmcPu29nDEqYDeYvhLRaO3pHBmR+du0j8vTCUKiid8Y8h9fqCkxG5
Bfvbu5ke2d0ZqNKz6Q0S06ybvnRs5+r91xxVtt3wuZFKzPinmXW6JUBdK9j/DmQx
+YfFuHF3kfPVhv37i50bko3hVcB617sASeTwAsilXEYEgT4H3NPUMI28k6x5eFt1
nVgcDMCAo4ytVbWGTZ8GNM5uopTFa3qTAYhPHyBUjHKz/TwO3uJVAxp5jU/8upMo
G+7gUz4E1nS/Vtq+kx9/sRu2tH5aQUH3NbiMQUAy2VuWvAa2Lbng+Jspu5B70Mkf
SIP7v3XiPdWQwRIpn/EmT7Vp8fnh5MwKZjKyyUEe9CI794Mz3pFJ6PS45yvw8aFj
uI3lPOol7EVRU7G/u02lzjbIo8TyFnUcuo+0+rEvZVdq2JVmyBL5DUhj6zp32O1/
JJEF9h92y8vL4gX1CrHyL6d/x3dXym+AQ3CiRyde4fP8eVXj2lRCM3NnZ+g73CqL
1uFdTyo4T57fahsHbjwlO3QC6XnIVh/qEVSF8r9QYpMEKKJ6JoA3IiUcZTYmBSyL
7vjRsriuOZDFFsJia2pSiOfj3Z9yuQgLkKg51gUIvTWURXMVcaDC4PeTIottZDIr
nb01rbBKF+j6wtgo/U49gSTNVaivu9pEB1sWL0Fy0yJGO245DX7wy4V6200pjE4J
IKvHsKORmnIEB4zhYXauMqNb1YY6Y0EQ+CNXYlzI2UCyegk8w3bCw5rr3TDibDyZ
N5JQ3XK86qMOOBkCY8ZjzODdEqc2Kjrs3kCakrNDg1Io7Ub5HjUST8rdrJY2y8yb
+cQVFu23vv6TvvRb8geppOvpYQvu09TmAwNNcXYxu9ZC5HyK8wzvynOBEG21eoNM
rCKwfxa2YpdUCGS5tA9iYu/WWFxHdwV74a5D6Nc8hzQfhHoIu5dIGkVy3+g704P6
6K+YR76C6obwQaAQ3q4law5PjzS5CR2Pm29UFWEPq+s5wq2XSyBEDtU46p6wKOzQ
Kp7oiMliGv5sFlyvYr9uU7PhMGvJsOxOy87qn1XfXxIkwPW04pWpuyRMh4Y4Wkre
HXcyiMg4MV6RNNp9sM1WxcRfcSdIATnQpZeUl5Sm5QgziqQoT+GrdTwFNqmjsn+c
+sxxkflFcbvpE6ht9nuF/rqDoBHx0hoi7B8/qxnSQEEVoO4HiHsFcqiTVhmJPJoC
NX7NxeQAnGh14EChY4P2DHo3PCdw+dcJRWxAdb9F3GE4F5ZDhxrdpQ6wcnACEqva
iyt9Sd5xCQvGPC/iTIjxV/tSwc67wlyI7sm3g27CLNihBx2rMjzRlYKJaULzr1X3
aBphUxKcU40o3RyoxlzXTmcuO0m3ruZsyt6xi3PGigFwq+ZJGmpG3oqb/qfazb4m
zZOxZLtl3eytTH5y7RoSZ9npqK6/QXCKaDZavznHzYTuH2E+QuZWHnRrTvWil2JY
HJEQFHHBH61FKILFMxUt9uO3d45XRhqvIDv0u83T8HW0kxBUokr7UxwdFio3yCkc
lfPAt2EzPRRrA7gTQXEQ5jn0ku7f2pncwCzrMJBiEFNb8wMPEfFoab14d02wZ9KH
/hXEtT5+/YvCQJV99ZmLFXWaycJMmumwuNsjAb3XhWCL9O+oA80SkTMriVh6AD9C
7MO/3GDiBBqtD/w/v9HQUD8XyJVbA0cOf+yQkzzFo898vfEDcMf7dFAd2Pr6y7KF
UgrvsiauzZPLitWBTJJxxZWVoD5FG8cfNpuJyvGxdpQjorkwiOV8CVy3qutEaRfO
FlmldMcWF990IE1NV8u8pPPclqr7Nj5SFG36Ib+6vcbLpZO3yTfWVOm9QY0VvnJ5
1CXo4xwOssxrUiJBF5bbMkyFgotNhuihSxOxMX9Jkww6xbzzIRP09CLbykegq86L
dAdcSg20i6t+aCHFqutB+DUFRMgZmkImEo8+pG0KRKe+rBVAxZYrEtVZoRNs9W+l
bkFv7GILz2A/JY3G3PX/bFt/9OLW9La9Xsx1UwaGeJi/RWQ5Bc34xLwuJbWG8sDn
EsMuFVhNVrDcQzWk9exwyW5UK6dcugWHFrNcP5By7T2QebtpFlN40K83Epr2RGgm
vEjnJCm90808xrumTNckKcBddTAtmzjod5FF9c/iqzh1IUFdyxsF7KBKq/6pS63v
TtIEnLMLWRREZ0XuCyOLZm11xZAv4iI8dUGIDgi+XzZY8t7HcpK0AZevL+LReQFX
2/7W0S8UkN+GuzrvP6CSMU0HiCAMK68iDdWfuoNx2nbLuqMvn3VjFyn+UxZTGZRV
sxYXllU3qR1AU0pN5XhiwuSAm6uOAh855cakEap6aK+So6xG06baONqxJuQ5ZxOA
b0hve6J473YE2+Q+cNZepPlqVfnIBOyUI6+zzD+b0njot/cQbXm2lAoGZK0zZPuj
N8LiwDVYIHnI9cP/MoZg2Do1MdgPSoVrzATajktk0PHCaYNi1pc3XFNG8RyRhR5W
yd0dYTV8rge8tBqJ2bS+9Kntl3hpRN4/D4ufGc4x8WxudBsf3jpoutvxUXMiPJS9
A+Hj8XwtKQbrVCG+xOZcIlOTXkI/XwwBYSRmaZdWFIjtQ74wL3liZWeGEvOYs5t+
pCjDts4Rpnf9jRTmie8rQap/nTZ4NC048bEKVF3Hj8ZmeQY7ORPykA/DtE59SsJL
ZvmajBGBGwlw1ev0DoP1Z9EHjknxNo09Dvg4Ab1T+DwEyZPPgT10BWsM3KLUyIGY
lSv/qA+nlQ3YJ9Kbm5lFk92K5+yxNV6sJbjbSPsoVwH8ZVkEDwCzsi/HluUR6SIq
TgE66D3A1uKnawvp2xijh3CqT+ptG/mcWreuQBOZDFbM3PCKpHPT1laJ7zwPqqKg
T3wXR7bTesIABkSZVSpzamG92l+ELuIO0j9Yo9SPL8xlpAuqCI7ERasrDApBpSSp
5fGGPhk5VqmBMvkEJiqfE9qHh0nAjJCHEO0EVHvMzAZDwQ0cuMJbXDAzdbQyMiJ1
VsRtaozQvczboE0RgtdGzNMmuoVg1HggLRM0piW8Edm7vRbXHJLgwJANp16OD9xh
Ww4UuA1mU3U9+1tqVJSLOFx9mTtsHIaFxntwZ5sBF5WBEp9lw4zS1bz+pS3/RaX4
9Z7qSWnqHpth3UD9Y31p3+8GdBHBAngML2UI51lLAZ54YTtkVs/Bc2/13JujkyOM
e4KWofd9NfH7Fy7hgIGdbtaHlyPTVLCUQ2SZ4Nl/Q6E5g2lPSVTVPr3w9C0+PZOT
TyzODoNe20aEyEh+xwx22LlSQYIv3qfGCRIXfGa1yrUzbOj9BDH28oQ7qpjb2LRJ
96tRjmtAsPw2VzPooLD6nBGxXJCHEhDc7IWwMET25bkYQDAwIafLwBhajhfqRSe4
kYhNsy2WCqeAUdTErBA5ijUATommMAFuSAZKaj+6BAS9DB7QS0h4czCa8x18HQgE
q6PQNnj9qQ0MsojxrP6cI1UBn8Vinhl+CS/FmCMnzM7zf7xUEy8ZMOdW56F69BfH
o82D5tn41jp1YaeQVtxceRzM6jY7XZEcXdHTLUhOuUkfZE1y/m4h/nGJjMA72rgT
5zsDf3oVJMvX2hw02cqg7rfWBWzXzHYbG2IKu3W79SbByXvb2mLXEzKm1pSw/zGs
ytrr0YuWI36BD9vLtt7M8tMTYTYFa5aT8J9lp/WcPOSNjV2AreU6j2eica/GXT9Q
FW1p2ZWFrVyEiZy0ICcaOmGWJpH4JMV9ehPitoOgFhZatmSIyJlU/ep8CAy8kLxW
HjMHRyiOFQiAdYHSjq1HlwzaJNDl3CTzxUB2cwEPyzQBv+Twwy9Odmc6xhHLYhLe
DVu/wHzKNta9eid4tcHC/1IuDvf8J8Xa67mr/CUcD1z3T7+homdNBcrjcAj2euTs
IoT7m+V9BfecmmcpsUtqWd9s/q9HF6YBmMK7uzqcZ/v0kANZvPSylSmbxLVPtI7t
BgtedSOKbeqCwr0vorj04YqjnoorCVSG55NZLyyKq1tVnKrWvoyomZilCqdqWBGP
h66tyDJjKKKeFNGucNBt6rpDoxORQd53pOjkRHPOWdBv6d3yIDis+rXEkl0LLPX8
NYykYVZJ4rk7QUdnGxKr3YVxjKnZmxYlN/UEd4FZvG/O8UMsduB9NvDvlGv32cT4
D5MsAX0R448OD5YaflQ9qRHCO43rcRQh3vaAqzRYKI6OytlghzVNVZtNM0ssWIX+
ge58LeIVYJz3b+dvu8mrYrY0k7FxAUGrznO52DtRc51CIFGLgiUZm2FeBscHSN7m
c6RlfDa0GZO5IXTkiLD0FX3kalbc8xTTKOOLXN1L1Q/QoXF5tZxRfA/aw8mX9uO1
ZDk64Tm0mQ1eI3MkLmFk68QM7KCLjnCbjosQo+xJWRAxgy/+weVd1884tX+BorUs
HwfElL++HKAcpfwXM2uLDBOShyTP40hbzTcmopdpk6kh+NAGNf9Ntf0jnWdPt0uP
2+2U+T3xQ3hpnfE7QZ2PKDiUMpO480cr9LKwxyEk+HGnnmX30IZpS5P/rn7AITTG
MMJGNhYrQjsWRcy+MvK9wuz9uulNkXAKSdgb48BOQAVVAzdVOMqPuyCBuq6MTYNN
KLXSZF6b8ER78njx8qROMLsUU+2LA1mBCeaiju9Y+SatUJMQ49XHvzLZNS9/ZiBy
u82OyG1u3Udv9wcLTQukI9HxD313OOfXTZrkk3B8MD6DVb00B0yMeOh1e+oxeHwY
bVfvP8by24UaqflZrhO78rbZwX7y86GnRfDbkS1RPdCczvy+mCOS0eCgbs0Z17bM
hytHjbZk7/SIbOLYIaX7K5Z+DMiK1U4PboXf7g1FBDUMqvvnLF8tRCraO1MdM9K7
PXp6qfKtDWDLmRQ8VH6cYaKeP6N6LhWYCmhEVXp+lOr1ZocH5XNXIrpVxP55lRpB
3CYiKswgw7MFp55IaxpuN8eTeF0UpFxx5yxLPS//pCy62vQ3byOsZP/ml7ZXJ/IZ
QykmteC8MTiV/b2Zl7GeF0GFGrdWmT9Z7KxQ30hpwdrU339gtV2PSp+Fpf8J4BIy
33BOufizGq0e0hPx+6SG1F6V6U2gq55ljFrJsKCUOhZasAN6dha01FWVwGOV5WGB
kN2iyGJx10tPwQBJe+PsYYKOMnUFbmMQl324TNAmoh8KSfuup6xJbUPKttRqExPo
aqCIDZFLLSkjtxXFT0SUEnKvc0h1yagBI9GnMuu9haPbaTVAU+ydNCq+Z0LDM8tO
3KhIQkUiDje1moeCzT0DxLjqb7GQuOGnNTcjgl8iPPE7hQOspLmulEE9ZFjtxVVC
zwf9M6XfIe2tQqQVdzTZAoKRshF3d2G5oITi2Ez3gG02aRvurSJpivSYdsw1GvyJ
LLEgM1ELH0sgQkxmk8FouYMq85SsyvulIAhzMaDXKgE0yOgbVqzURsxksh8UZ0ZS
fZSEZeLVW/wsNPUADXbus7gwBBn6HX6OWaJS5zE/knh8NC8896kiMmkWOkKJWSqU
3s98p+SyuB/KwrbQwj32/UFmwbD1amXjHXKR7aJLvUyFIWy3a5/o2h0E2jiGpIhm
Mq1PVzWXR/27u2IAvIgeJXxPftpTfOMAzc0Rq81h5i93yXgMPX0mjixe0r7TwLqr
SS2zlMCI+phF144BTjRBHIeBpqfIZ/mmO9ht/+3B/bJQb2C+IqPsb/tnjG1KImeZ
EkLlt1eecqQvKM9Yq/3N1VCU2ORk1LVJfIXagCNklAM1VeG3/TR+71P7l6zAmcBr
Nx/Hx6HplSg1HLaT11GkPk872Ge7+6ea431jXO4HIPIWK3iXIMPJbkVwM1kUI09i
DrKJkygaYYN3v7bQEPyo5qpOyNzbYi1oFTgtvtEKOppR8/Xgh4tfHjotaPEb9Qgi
KQFAnoErp0E36bMU5sjbaB+Ir2rOZwNc3Z3hUmm/RsgIoPbYXgLR/ZC9M6x6m5c2
UvHZng7A7WJJhTeN0UnyjdkRIeApBoNAIyBugJ66znjg5r7/tM0b/D7NAp+bP4l9
knetdUE6cGKP5Gmntq6Z2FblllF8h4+hvwHunZIJzKj0Eh0NPKQyLqHqXcB8Acdf
T50NGTRy3/YVoGyF/Sxe7C9up+9cJcxBC/kGluN/7zeGtgixWuH/OsEKmLGfiZIV
1I1e2qjqJes66UTc/X5CS04XsTLYzjwev2g+KiSgsoVFM0D5upYsuH5VDMintxov
iMH6UUnV3bt0OWWj8ghFqzwCGPVRHw+rc5sMFXZx8C1jIkTpmG30mC6KHPQrp53F
WMm9AtK4M1PnVkc/+8AOVZUgsg0hOgWeLXCPgAcI+35QoQroQZBCWinacp/9+s4s
lxnbzkDYCnVsJP9ritalWupA+y1NWLRqbU46HumPHHglBYtKaeyyt/xyJ1mCd6lo
6bWu//WL8l7M+/Ivqj0Er1+YW5/AJj7JyCUWG0Z12vqYoZenAlSYK7Df6GvStf2b
qYRVpn0O2LXCF8osaE/WPmRJ8AOLxfYHQ1tvVMmL81H7B5TXPBl0wcE7WfzhRDTE
Ixjc9ITOSrH2GlMoPl7Av41FyW3BllQBxS3tzaijpzkMpZjt50HNCiXvXOZs/hvt
bEIFZfJLIlUA4KERhyDtgdEjvMPSxQoXJlHjjYYQPXhiO5uPBuq2W+cn/FBdqY+V
p2SpNjneWuUjLdGJrvuUIH4m65PkdCdlf1xeETBPavlhCulIr4jMiEiV6wcg7/f2
TQrXpU9c3JxTSY2gKD/H+8sHq+CqMTGrc1TYuFKcCb9QiSqFQ0GSiDTPKL+lUekT
4+HVgQNJDDwF6PKqFpOakfCk49SWMXv1KnOEpnkU/shR3knUvOKb0iw8ArLqKcIT
vx0tMeJAKn+RVIYkhxakCGhn8tpaTc4LGWDkx9ikf8AJ0Iu6/73VX7tIVgrGrYyA
Z88Bw8xEqGSjm2qfzRPCfNfReieWY2SnhoHGYzhzLZO6C9RnCOyDtPdWYSEoWe3l
IGDW7/MnFH2BcJZm3vr/Kv15OTRnGORITa9zNZgI0VDDq31aoLt8L+aA/73eoqJ6
9DRIEy2PqB/PnDHW/Fu5Jx6rqu0Pz108FWnvhnDCG7QeDHod0sSczGB3QDNSIVL4
vjAh/iSxe3bXvs2iZjuCP8Hdb0qjdArtt44dVkAvDGR1mMqDT6NbI3PpdvOxnuWW
TyDpB4k8an+A7275KkwQMb6gE/zFP1q1cJKJjmYqU7te5QWyMQ9S4/1SifGEIliF
V4meuTpJyX8VJa7Qeu85E8C1gozkk5mPvUWvgOVu2kUSTrSsG9ptc9+k41CjeXZQ
TgFc2j2oMnGxT6dSIs24hK72BhNOlNyQve68C17urSuWQHJId2bo8dz/Lh+49/kQ
0LOIwGjsba61/3G+h/WhBK/zL87SKMG+KCG6JarI310KqMBN4KJcHyqEG+m0KDpT
y4kZgURITEs+emDaGdolszuBaAVZiJu1MdUWg6vzIAtdPFwkZ9ARCI9gbXL4unGD
TFBVYmoecGt+GMkDK3bIibJvy67eeaL6o5ocQzshxT7a7NsiPbmWhrUw7abnJ+9l
9M73X36gFaCrVUsAd0aAUtBKKqLMTmcK4fT8fxsC22LfLB1v11I4ZIa7b/lD0XMS
WVtMaBkAkFbCYZIYYrKStW+54mUo+j8Yyo90nZ7l+s7/YaC4ZjSG6xJ/iwVyzhly
7YJ+MjTCQiRI89YRhHXJCRPTLHFZjgkGJkiyexA3hxRecDk5HF5oxBPhUH4jvee+
hzdnwFYFiUkCMOVIcsvrwPEZKSmxKKHn7C79xpJsig29VxXsogOEI3wTpin5TF2z
c3Ybbw82u2BMCXoxixDKmTj6NXyveItacPHNQNLEQacwOXTxGNdhOHxzC10O5pHt
r0p8BQc+Qp1LWr2Hcs16CXzvlGOvZD8mrsVLfCkaJm61jT0BfIL2mfNVTJpM8SXR
ByNjVRfftBVJsCsrYfTuEbQYcofgBo0mKRCtczPLs82zklFTK35ZWfDlieeo9/UU
j4Sj0KAW+G+LSmoDIhlMEP7JIIbkbEFAGDMkJRW4YDuVY+XSm0yn3BVspvvTLxvN
FiM/L1L2aoByhaWBPTjTJ9SfkW8acO4ysdvaOxV3ZMqUfB7LV8nvyDegdkpZ+VUe
CcndvU2vli6Z24AorZRChckEP2quJVwW9mSO0x9HOcukoOZ9yJiA4flWil/uq83x
wQuEid2EIz27ry90oW0yuXeEanshjCZsY1BxO99PLvE6/RMF1hYa4yTut4juY7zM
d7qQqHuIjGr1Bn6v3kIIK59tSCkgTrKpwp/Uf93ytRt9UiCiUK4uhcvMIZt+eHPA
yxouTyfRA0vXKXwzZoveV+spi+MS9WY4jPxGZYBX6qgX891T4JsO+ajQ4BDYVNLd
YC6Kiv01DqZ1U/O8jXdhqQgoPWq4WBnJXkG43zfip9w0u8fazmE0zqMREOsPY/J/
icTN+noXLeMQI15unQeHSmVQpOFW7UpFhoPDDcFDgSx8+GCjXGa/uWw2PpEci56E
ccLlP13W3lS22OHak3aKnigf+XsLu+bCwBhybCkG4hJIsSK+3mEMq+vL2TNwCTqu
+NLnJm7ymjsRJGDlbT1xzlRZLA0ApiJRpXF0HbMX2Hj2NTtMGBtHq/j7w7xm8rp0
wr9CMmPru/mnbwxYxYeG6XjKTSucIYvwbqVYe5H7+j27eEO+P0yqcFiQNEYEhMsY
D5o7W1T/YpDMXlVf5Bx8qsFm7IIoBGK8mtpGp9yGJdrRf2uFiCci3hXvPPyFwoJk
MyQ+8bLT649JEo76rJ16m+r0n/4faT3ypkrdbV3cVKZPgGi7Zvba3N4DhTXJMPok
bjAqXprQ4Wiwxan2f3yR5CudCNnZMRu/eGLUWj9ogSCY36NfrxSOZ63NmDpWaHM7
KkBlslRr4elXGZFtTgVGs3Pvn8YLs67+A5dKspwEJtK1W03fd7so96CtrfNtRxx/
bHC5roP5Ez0rUe4qcPyn/ZZcWHvTslddJqJMDg3J99rsdZWLC1+hyIC9oOytkPmE
cR3J9+N0R24pYcsAY43Z54bEGluqpnV6rcd1ck8uVh7Hmg+Wg+g+rzqbosMiKubv
Oi4I/fJ5VgdiU0zj9Eamkx50X2nxC/uav8AOfKqMU01WDAfGiGci3rro8/yUOtOT
LvmgpzH0q8/Amf+cxi0hUzZwYYr2MKo/e1FmZOvvGu7TncangbdQJX4d08JsDV+O
s2fF4cCKOn/9/J0lxexBaZHzPlvONpORu+mDGjVGYso1Bi+OB1TRBfzzNnZP7N2C
YQsaeDk6hmT0QSmFT2oIeQMf3usNG1yKHCsexb7axbz3jGjnywTsuMy6quSlOEhN
uuWVWSd1m/nsnDtJ6jN9lxfCJ3HLnCO12XNjrJPn8XqFjKYkofyFmi8FMutQ+173
z66x6oFqeuNzV9cG2/BwC0GAcp94UeyRZgd1VxmqIbbDZUnB1ktTa8X53Y9NivsW
P9CSLPwMFeAP5lp33Y2a7g0u5zQRZViWyNKNJrgy8ZCYTw2MJQhkUuqpra6+X1eW
LzsiP9jgUQppuNJgmIz2lt1HeG3sQvpVgIX6wIueYDWAZgb4MWZ7AL6W25Rmox8T
5SizUwLTSdBBF52lsMzaatFK4KLEkCAftuv70PzhGewTmHEiJIpFhFjkkl0txgSf
LzHe43wTJ4z8gQBmSRJetUCZ4KsjFxZDXJPxxu0v3yTYgo9El0gwvC0m38qcfxkG
c6Gkqj+V0+1b0qLhbSNv8zbNPdQCeDktMN976mTge+G7ZwnN7SGiWqxzKf5i4tNZ
zLu4sGGcW/MCNhhz2d3RuQKAoxWTtNRZ2CqQorqb7V7HQ5UNd6kGgQnZJNy2YCDR
gxId6cpySRzXNK8Bo3pL7h9v8LgNLdjrwTYc0Vizijirfy7u9F2TkMwOXqkG1AYY
vz6rKIx6T+DKsoe7sjJ47cw/5Xe4/2h6VAv14UnmlbjuV2+N4ivjD8ji14wH8D5C
8DbhHo5DvpbHfja72Pnoj9WydgNm6BKy0afQD+SJWn1TBS6ob/rB06IlbXGx+g7Q
rDVafi/f8bI0NPC5EY4Ukc20OlfZbMbYSeCjsSayeKv4+/UqcvbUVgoVJxppdis2
Kg4iUmmmWBgQTIk9jlZvBbVbMfYe8MtJjc1xR2rmBqXD+zbLYGH+6NcDir05B/5G
6O7dXFgcs5H3Q4koIvKsJyZr0wP4yozeKcfeOv+gkY4KLAlRNiUY0PjLGuaYtPu7
V4P7FPQl4NIU2ehREQiVOo/gAyXQRa6JM/ZByPrbkcHio8nQzuq58qHdwMNnRo4D
xAi4qjF1oSo/LZWgoghUWa7LJ+7lh6UJDsBKvYwyRTVV12eKOaUW3paK32s/mdVN
v6yXNyH4uiKS6ks0Z26PAifYHrU4SYkcwYyvK0IUA3oLJDsNjRKuQcHRzKiBeDAe
16E+YKD5KzgLyM2z+aRxweSIHoBAdDUARaa/dIfRkD09papP+BbusngT+ymG9+Zu
EfxD4g4ViuUCxJo6LTwbHmyM+GzniiAr3UVYlY+Kugm3i+CyG2DADaiPxCM9OzxP
Z2qIv6h9qc8HmfGby2u62yUCmeTlELMxZZaUFRKc+h79H/C3flEad16ShckqYvPq
ILoTBoHK9gSqrbtfeklcNgmT1ymuc4USRHQ6MNh0VFzGM5vX4GRLDThPftlHheVd
aSTdMEgS6sZNS2WoWDqzyD+LIO4YUcscbRgSFsP0WP5v2swP5kytgXlPLIfSl8d+
zisZw10+QGRf6gq+6wXzd2QWpgMTCjPAp4cRSQHhDGK1l/4GxVX/26JaXg0R1RHq
Jq3AFKzfA2nqfN1HwgZnYSEWgu2lbOSRiVelgGqvV64tnPvh5XIl2PuEHhVlE5Jc
gK/VPCjqq7sExoIArSs/Q69l+/FFExAFWNOUsl+YfUexFrNvD3B2j3vMVTve7Cq0
rl8c+oRYowoPSuArdJLhzVPaMO3V9m6AzMu9k6Wb1BRUutf7U8UDtLe3XTIGbCja
bFn1d1iPN9jGlFJgpPSZXQZ51buUd0mR090BOlTUvsHtCfXRX01nJ75/LRyRfop8
EbHHMFFPIjs0IJZKLD7cka8ktHOM8PXg/0j9igm1zfybAU1Z5bj3IvuIDc4Q+LSo
Dg4HOvT0WJEyfGafbbKZe1tm5N7ie8Z1p4w5SHbyro0OaVi3ZyzRgKp6xRsOa2U1
35xuagsvQwXCS96iGkMgwGHlAqePgX+F6H8rJa2PO3PTqQDZvLi/TgrG3RPVSVFq
+FgmNhg4nWfB7iMixJV89kyERBzvAMZyMZa75DLVlAcq506bBLV//Dio3DzxrYK3
p9GUuxtV5/BrhuPVCnymCCmIj9tAULSL3i8MVj5HWJQ0iGxvRZjIMvq1k3ZgYbSC
fS9W96Gs144UZwzlYeLMqx/DGPKBbp4Osq75DyfZ9gdbN1VycCGeo0V3mqP2kzqb
Iqgfi8nsKTaDKqIlfQkCBLkCpuW3EhWbE1JTMLUqIHaUITBQoVe3STpM6UfVNFEA
YuSJuyKffq7xip/WDmbRbwyyWGtgVd0ctFUyucuAWd5Jy2YD6yU1vOhbX6qHwUbC
uLUGCw8lav5sncGR/6koGghjU7S+BmX4Si0dn78+CkTsxjns8wyDYfeFmLFoXJ1S
UUH229+fnwrCic0qjjXWLaZoqqbJFDji3R7zu1ygyqD8uKhDdf93wjlmXcntf2tf
Pb9+D61N2dCeooIlG5agn6Y5EA8N80c1aKTAJ4FwB2Frp/sVqRiNDZBVZTuv4SjO
dCOrwEVxGlSiCQdocz86+M65kQLKOChMVjmZ78+cMyOgzTyBOl2zpXLEXUFCoy6A
jMV0OaBZbttDfh/+gpP+j7+idFcX3eBlFWT8ttEdcgkLSasUpCNUOu2xn8ssTmHt
XrJSMUsqadrLaM4Yz9poiiT+Rm0MJb/33PtNnAgcuAATbpfnSPZqIuZrHLfw0uxB
jeZRVeFnnuEXfPZ4YHKdLnGE0CEYNp0RKzEOVEe2w9O1RIFfSKaGGcOHOrvROZXp
2bLwWJU7RNcJcqcX0km+g9jO9LqKIDDsBuoOwgAWzUybIpJxTMdfAnI6hdZwl3nE
9ZTlfZJO0WkOpmzaWoM3oyFHGx9HrF9xtoszz/R3asgJJxpryoTsTipBDQrOeLfk
Q7yTPUYabtHIymRxjdperTqaesDpfbJxlyQg6lcKrc/Tj4zW9kU5ruFCQLvGJ44n
baXWZC4pk2p9qlA+61fkC17klxLaUVgKyW7p3hus8OH8Vg78X4CnxpaoWVdhc/jM
NZ1sTRGWxoU+Yv0TaNtkTz/sQ+hnd6mmOky3kCj2eRYNdO+/lHaQuvwktGz8qPDQ
IVNElbk6aMv/vUhxWTmAf7DAvpUZzTxiOsHRs1NOSgMLuS3o/FODlgj1Zy9XrAGc
7OPewEyHtG0GmTym5F/HXmwM6kVUdajllX7Q96S4yRZnsQ7eKiEAjQIDu5Rpqykj
XDS17pWoG+CQzgDlSELr+rxCk+PGfemUV6iQVqyp1smrDqOFUqN8LjebElZBtvS1
sjrgJ4TNlajFLfFr7ThMMgYmcZWOs0opifO2g2mUST27dZPOcaai4juxoYPnS8rP
bn0UcppXj546q0S1VMHYUSePaYvWVeRYjIZI+aXclp43Te8lslUULS7YdHpwIKQv
DL7V35hxsmsUfj4wNNa3Di9YO0n4ddIbWForI89XgMnww2TI+E/GSEsjDPZ5rnaH
h6SKxNUO2Cqhak2W9uIuoHi1Ql9lC5LfQVeHl25rN65w324r47GRtxH8EgsGvP5I
vt2LUpvo4FxZslY5jNWHEVpZgdsmFSFZMJQbS7s33DRaxDY6Whh3tOG0oY81DbOc
YNvcwIy3uAnpHX1/D2eXWf+rXbd12OrlQimbkUijq96tmSfor65KDeKLtKdbXw2Z
vDKZ6j2suOoX+CZvKemkzyE362kZcv8osMaPGp/RdC3USr0eeHkN0ipzYkNtQ7E0
WTeV5tpQFADrPY9jHHyp/lAoCbojkqwwZJVm7n50NtIqHiIgphTpAg+PkkRZy4Bj
KmF4yfLR9Jn6Zqa04koWjPGK1BNrCEJMyxe/eMsDc6nO9RPTesztbHwkxL4CeZ7d
Uhg6ZNNye4vAhq6G8B2XUWESAuPrF+/MB+S7tW8QEsOu+yI5rT87jL84Z+WSV8sj
rOAgm6LpeFlngXGIKcZsE+Vw7B5szyVfJpHOrO0JYOpIE4tO/Cwe+oaokmksk2eX
5YpLHvQscE/R0XIgiz2PQQB9TOO+C4eN8kUpyxfLhlxeAPJ/MoMeIvrxeyij0eSv
qpzvNaYh3NNY05TMPVAFn40jFk6DJWjZjeoluxFlrtlnFljPpDg9OHjrHU3fsB/u
cDKupnSdgUkinpbPjIxFYaiIFu+Y0DqjgQBt+LWHeg6CuaZ2JVaV/uAzFtxHUhC6
T7Mmlz5Kbx1T/NZeOJFEweM+QFl+hybn2FDYWe+f4ZQiQmGGKkstU/7akXgbqx3R
fDbV2NhBxgZhh+ekIA8Mh5DwSq7A+5Dx/+jv88qCMXRCD3fjUiW1B2sCirxLc9My
cnVOV0Nc6eeeYkgroNREkGNgbkQU0s+xRKvg8n9xaJP58z5VhxaKcXddEavm5RV1
sJopUNia7PfkEOUbbNAp5aVJJINB6f10YzWT4iAt4/z851IsA6cQe8GO1L2mQYsz
h8UYPue5Avhap/MFyEBA8jE08RP5tV2vq1a385ge+w+tETKZLvziOQQ2k02T+3OU
zDdqAsMy1rEuUVkpocS+OShU8EpBWJZvpC8mKUemYZ1MyhGkhm7pcUNhRk3sCdmc
vdJou9DhYrhLhJ1tD1UHwHGympWgreQTDqD2L7MtibvvHDUdAppVVdRF5Dzzi5pQ
5DghlrOfDdFbZs46+wgAtrgKqPdfUt72cu55hhRO/33aERKzguSuYGQCYA2Jwi0/
WT2qZXpLOL1+BabvGfBxNetdOzdqv1oCiGfrCsDWz6ySJ0JQLdnzXc/TlWeIZUJ+
BSOQytoHyRGkQE8TNXNDd0uHYaBBiXQG9gnL2KOyzppwUShkCMFnSWgwkjXT2MPP
l9pdeY7FgKkVBHI8fyfPKCNZZsraFwee5fjP7HUKA2RI97qWoW3wtpi6pq6emvGz
NdLcUdWWzHipkDenYn4YUeQbFiiKj15IMLuGiBKMjToL13BSRLKWiH9grF0QlrZv
IA2tNgophClizw8Du+AxTMZ+Ox3+n16RgK8yVwPLSDljTD9Sf8WIQ3bT/bOdYdNj
Y2sVGqjga7+QYzP5mnCSS7xHq2MHKeeNoV2e6HalXcTusP4le5v+IrtcfX65NnWc
Vg2GtLW1rdo+1cNkONJkzPgxc0q8V+mZ3x50P5V8j3jZh2ucVwHzAQ9dv+Z1mHZm
XSRLdfax76Ntv0jn/7XofnzcLRdUC/EldYthp63qcWVwT2Elv1ihlS/0w7MygCkX
T6uRFay33TkbHx6zYmfp7C7f6p6a/qAuEpE/LpLQku8PdPa5v4uyl3dhDfgSC2G2
hLjA4a0STvjWZAJ7MRsKdT5Q/2oO6OyD5JDrFlyDLMUr5UhHGU7wK2pA3SIbim5d
TPn0ru3E+zVxuvrxkvC1KNiiWJEvKgT0uyV/VMfYscemXajA37MNKTr+nuPuVWQ1
fDRWAFna94ODiTVXMnHDqI1dlAnJP2Wy8+WwWUgU5ME+0efAsSUEKWYNpclPfzcV
zH42R6yBWfdhcxq1eCB3kuuZTuixcNt/gSxRklakI8LZDoz32ToaRikIxjD8yUUh
Rb3vY9g9pXmC0cKJgzezE+ifgSUTwgwuQ4R92Yi3Mzt4RWm615yYvz4icklwTkk0
QsHLbsSNeSfSpM24oxzYtpoTKa6F9WnOvkUaZlob8mnPNpCrJZY1TLV8kLkNDiyF
mowV1KfW76y5ZRp2zoIQJRw/3W1C6TV6l+2hjXAthfqd4TMDhy8MbFSBm5EedpXh
oI3QiI3oaDwvcm47Fa8OwZzRO3nuAzU426x9dvsrdGcHwZVmcI8YYjXI/QdGhoPP
3JKOoKt3NL5UgUOUMKYo9ihqfY/dAebtV+0TAvfx9sQ02CBQSjbrDjA+TGVrfOmY
SFuVcW/BgBPZnTTwj8/zhcAXsFw6h2YfLLs6RE3dGDNclAidj0vTcQiVuMPoM5es
frA1IYVgJeY69kJwvuFKUO94gbLKu38DZssTWpSvoA3OvNz0vZSsyRZ6IZkEzdwp
KW8KPqYw+Ix6IlgwWfXluK1tM74sd2XT32eF526iPBgp30BCysFq0iDd7e3Szs6I
F8nNFoYfiGX9TXBhFGAMX5jycy757ZYjprdeRd8KnHxZPfE7jJVj5VjeB9EShJ/A
GBuNLf9e1Iw059goW6gmOpgsavrpMhd+888oGwWkIKXyYiUX5qTqcnCnFtHV5rnG
7l+zXrJSLwCg6vJShreq4SwN/7ymSNB98pePwQM72x5JSlsA5AeNaI+uMpL9kL+l
lvNTtLow2+u5LhporINp4HkDfoxf+yzURke9yC5icLTi+4wt4D4Ue/K61irS8TJ4
wZwnGBX1YM+MYXUT3YnJYOtshbYDqEmOYgEYneHHKLw8blYAvfP3ZvAo2faVKPcv
6EXaasENwxw23lpQJoMwoTA2Fk6fYnuOrwTcqyp0WmNfDRszoFcfxuoH3vgkcRzz
Hyn8bIzBRrzfk3XaypT5u8HO1dklvRGb7Lyd7XixrRoatOiNBZ2JUR8KszQV3IPG
6pSks1NZvZ78Nnws50+nkVCnvStYfoxPJPndvSOJ4CtzbX49iRkvcKhUSBmnmmyn
4EIpdcI1y+GOZlhLjoyhq/rfFrqNKRTI3sRPuMv29ln9iFY7jpVFjm10i46BiNC/
4cuxRx250YYSVhZo1W0sIXX9sLxrZTPUX0RnfuAam92Jxq8cJlCGC2J53tbgmHCO
QUaY3sKZyl6633BYbm/pjspxdBfQfcZ06OsGCthHGytvL1NuZx2UlmPbkjfue6ht
pC0jEE+ZhkhJOmvFVC6HAIMbMTdC4fCgmOl2D0C6m9HU3l7XVNYaXnmD93eA0/Oe
S3otV6PU9xCHJfDH5+u4qeae0cMWXq0QIENJTU8xrgM+a9ClEyIB7vYIQW9Yo7gJ
XzP4iyXsHyiQ4Cu+xkNzJ3DERLixSYv1s4KlkFlM8ttq9HNlkWya0NUOM4FJWgug
KDSF2rxpK6jMNrhyBPZts8T2s17FsK6lFHhKKz28RHS1Z7aWCBmNjyPFTw0dSBE/
J/ExNlle6ThWy9NVwiothMmgmJa4HowlYEpgiUUYr3bpbqlw5mhvQxdUn2MJaHkE
Vt62oUHxpSgbkU5s+7h+FPINJMpc9RvfCORJJd8MVq/3IvYqZuBn3sRQZ6MG8pOL
aSjBdS0TTsyWE4ECBlt1b7OFevzBTnDvScqJHI6k5LiIwvbSjelwUzwPiV30pJO8
vBFq/VOucd2HKYhsFrKYnxmf8xU4fFgoO3FOYZhDoQuj/16VR5KN1azg5VH2zfdr
5brQ0SFzWJgC1rIdXq+P1Gnb2u4q3p5qFU81kEQBtq4Z/QVljrBgdaiXTjtN1Me3
thsTIQ8t3anf9BR9srGauBBuEdHFZ55fmT6RbkOmTrfR7EE1uNm4XIm54QvpGJbe
DIWODgdPSB0WzdnG0BM2tJ/Tcbv8/M5qxUW3Xrq+ASbzQQVStJg7JsZmqHgebzsh
ld+F7ckGD9r8lKXDhcx3pYhiSaz78fa4yjAY1EfmGqgHUefFMh9ImUeNrIOS7WKU
9S0RZn9cnUGSYD8jjpNVHdCC2WviWkiBcxFi6FTG6iN3C3Od9n21qpscPN5aX2b8
FAmenzi89KQ11PJXWEPQz/8iw09vFzZI4qtnwHa5V9XGQhA3S515FU6ouGeAH7jI
ZkBuKoe3wbCmaY9+7eAx3XSu67036kEh7navNP1u23eyA4AgN17JbWVX3Q6DQHAe
qIteqd1uIpXM6wVTWzoP36kxhG4TGtFbOZGhCA4t4hcKWyVA4rNxh4dmdzy+4Lwg
Aoz9qDMhpL5jUkTls8MVOsYEu9zz6rdj64LsIjvPJB9PsBOS3tKuslqnCIuoqQ3Q
Ytzg/Eqj3ajOqu9J7Qy28QDwM1uauugubUVn/yVKgBg29lGNRMFUIY1jcMbgIYE7
gFTsOBplfMzpiVR3GIRZROcEM278PaQiO82I54xoMKgrcSgxFdvEYtWxk2CCxhyq
tiY1JM3ELocxWVCVLjO/V3/jfXPJT1RpdpNVSzTshD38FjOxvMw8APONfrRPEVgF
lIJQKINwsBMPaEiR6UlvpP331Qrt6NRMxEE9bmTlqYGh+/IhqYoppoQpQ+woeCuO
TGc9zR5U6IT66fAlOr56QNcmk+vNPB6W0T/SctnbccRZv9buINSy4A0P8qk5CAqp
DRNx49ZSs7cnBUCRLJFnMyBxTXqS+3Ow/2Re+IKspor5LrJLvgCq7dak1fyOk8p9
D4aPqPeir4U8Hf5Vx5BvICmdyFhfpnkEBUBTfXN8HVvuqbpxW++/hG4ptpHBMWSK
GWEr+zbJ/YYAOF914CD71iaosobtfzWR6zntqBYJ9Wq6Y3RTU9BtDh6VWje41Y8B
aw3FT4CTR2wR1IfGirHTH21m10T2Ea6LPzKUsNWn8yCg46fAZ7Z+QRrRj3+sooic
r/Zf7hI5Xk0wCQZd9lSIKRaDhFNjlWe9ZikV+SQU90aIUSxA+0C3eOhl7gQWw1xw
yweOEFODbvg0SXQkdNVmqQpUb0S6JRQSNd8MzqeOUDgF+tH3Bx3iwOErv246ZuUC
gUTXohA1LxiKL2qk2YwAiRZO9V9qwZ0JghIbU0xhX6f7xNl3F7cQvpnCfKeRa4iP
uigfTO8A+L6n7+m6gyuojU2t9LrhLWZ1PN9BXkgOH83b3AgEnBeCA0ZC0WWKP0uA
GrMNrTintSnC8OJlHwKoWjJkQMIWt8ufsX53QJ1agqOEQlLtjnr8f83AHGZsj+19
ywzWRNknuEOTpJ01p8JSdrOnisTjl8NXV6xNm3TyCwtwUhNw9aSkEpvwwXavD69y
fEgAgpOHSmmr1taFB1GKX2fsXw+rLT744td2V3uDkMK/UoKO/S3jlx9fNLkBmxwN
gpNKV9qN9NcW+zmKHCI+RGxpA3cJk3ofo7qVSs7kvAcZaXcBekZCwEXJM37jv4xC
G3MTCzuFbjPqevttlV+L8+icES0xRrxIANYmAV2Wxk7TlIRDZf7AubA55ca2kq1B
vXpfv7qurPUn/8T1kdG2i0YQLPHgkVbubmieMDPH+xhIJnhICALN9XtW3f6qSHbQ
bmTlRos4QogdxV10XSzQZX8W0ZNWA8nq3Kg5WE3o6R6kFhYGpdrejzg1Qusfagq/
Ry28q/6av7m9ujK1DctQ6imLQQNLDX8duutvwsoYWtSJiR8WgX9IprpXa4SjBNzZ
Vq20fz3pWwz0ySuIhaolFvzmQbqlxNe6ynmWkwnZwmdGW6eoRErK0jrSTDByB9Gg
/pIcxiHa2XmWImkp39w8C3yj9IcwZgtAXw+Xq8C256xRh/ybNV5RIDvsYGkcyEfK
WS/ZI8IbR8R+4+t4Xh4Z/NdN4X8mkk8csdl2NRWbs5wy7eg13tNTOYEswlcuHPFT
xgjYTlTf0lzo0mDkAa2Ie29TIsH4doR7Oq8nAR4Va8ovfBofKuOuNRxg8GdJ4qtX
9sZU38zBFWzfRJhsFMF/+NXgtSmfmWVluRTvyoYeW4NnHNKyIqqh8BebAPNfnG4M
RYxhs7rMNEqMuClAdZ2ljLXbiaT4IDRhLv8tVWwffhEYwKnwai8b5HmTGTSE1icu
sAod7quBAJ6dZUa6Z7rbKJ2TsXUrP7lN8dckqWkrdeZq2iDTbuFBx6a3Nl302RqF
AefbDOkXUlDSB0Cag+bE/FXFzKUgtDCor9xlJQ3EuYy4xwh6sdeRE2xBJNnnLOBg
Kamzmge6cQ4Lbow9YtN5MOa0GN5zgWAxvfX997svOnyfJg0gN0sYp02J/oSrU68B
C0xi0uByndUMsFBkZ7fzujNDkbgalKFuZKw1SD8Hesoyrr9krIQ3fwj4eZy+ADX5
v5roQoJru5dJXdyX5cVhV4T5GoiYbzLM1ayVDavITt6hk4HyShhSwK+w3/ZBXKJo
jaVvRElMPTXDG/lnWIiNKEDOUqlZGMNsVSb0g+bq47mOR18r1CYg/9T1GSmg2aOo
vY5C9MR7afhhaW/lKZG0X3QogyOw8fyPrs+MoWm96WkPKYN5h7sHh6ipLO85VbeR
AcWqOcvdzg6esVzri2yuYTGuUh1L3u+z7vyxdEh+kbc8CLZcPOgFXRsk9COTq54V
VIH8m7wBCFAcFrzxtOXi/LbRWJUf9XsfcGBzj80d8Ez8xdr9QTvC9MTkisP4RMq4
U08cOUE7icJYIIOu0HG70Oxtaw8tGJXnvIDsayREfsggjfpBUOArvCcEE5cFeBey
XZq9Fe9Q75628/0R2yICvYrUpc/K/12Xy0xDPygx95eDb77cjqBWOHEt3VplHWWy
HFR/uOKTbe7ScBLdNLTvpCd8GoB8aBTmIj3RaBU3dRue7nTOLEr4vasU4C+KVJfO
x/KNCWNvniY8GxBghslUwQX/RGmiuM8Zcnr2JQgwXTItmvU9iPczWg2SDoonxiXC
h7EWnXN2u+s/WGUeGFLwdaWcjBJbMUp5zZsD54Xdo/oNdFkrAgbX1T5KEiBqYQc2
5wonondnwy+PCNCrvsY98uGAfzgTNXzXKAPjWlu25sEHgw9KUTl6jEQVv63m/MRo
Dbz5XtIH7/j27OpcqGUhMd9Y9UWJ/CXY/H3wSXzxVSDPoQQY/HVK1N6rCUCMWdzM
jSVVgjb0Y8XCsUMfoluUeesBJeU2C6Pn3KoiJRNUW9sGnRpelsLOegS+PMKNsUks
awhBD1VEzyDKcYV6U9PlIApfX63gB2P7QSDzWGgfmW7/896062XpprzS/4GityED
jAjBcz2Cj0BZrjFawk6oubFmVvB18Zmi6+TqOQzpqARYT6Ys0rN32/vpb5w1oDtV
HPGdDQm2mIYsUD0fPySq47qbZjPfTG/0UEvorgW3Uc3MdvnRRQxN5rVki6cmimCM
Bq9w2fOjkD+JHg1pZCDpbAIW+abzrs+leJTl4HYWomCyFCpyDI9Ogxxdu61SZsxR
PyZe4MNh2hPP+14NGK3JdbIf1kW/Gk7kEzXh1V5vTg5Fttsp1jFGNtGSJx5arriD
ONajRfV5CHr+9gtz72qK4MHuqXz7VLOTVlYYrclW4joy+OQBtCM1bJEbhz9dP5HH
/FJMui6iZovzWFecQn4rXkIBBn9cJpDlGOeTv77ry9x2EEUptyP9n/bESIJHIMUi
nvXGV+KWUF5+83ajYGZ7K3+wsHWn4a6ScHI9jV/tBMmu0jF+9lgdO1BKScJ4yyvd
sgtln+a/Z7esvOWlDcFS6zQpVlSIHa59sOgyg65zE3IO+24P86C2rFlDZwzJdiXk
4Hayf2z4sb3NmTvJm4M7i5yGkkszPF8JcSf6l+dPUpWM38vNeOgTDVBDTV0cFXMO
hBm0wbraK34RvwpayyzLR9Xpx6H+caQN9wPJB/xc/qU4yyDrb3RrnfE+yhSnDepW
n8FiMPIgGr2a7wbfjy1E4NX/D1uT+zd+9OAUjHruUJTYIAonF/1xs3ZSS4Cxmyo1
b/Hxjq1z8uooy1al94ObnS5VLdirfDnfdhhgG9vqavpDL5FDVYQ5Xq26/ZUP9ysk
4vK9+Go9ddV4x18vL0AtGe6qd/uPIGgx+j5+BLxHNCb6ur0XbNFmruur7kW1OGfx
HU8nmbjEuAce98Hf24leyR3od6C48+omZEBhzGTJEZfXVR9f9J4ZmUMkPSMihR0U
t0Sss09TbYQ2KFlLvLx+0KT3uqQV5iB8KlFOpPX2i4Kx+8VK7V+hBvWFZPNBt9LE
uG35zb78A0+5sjH6LH0RBIyj1U5phMiDIo3/ThVGZxB8tz2rJKoDRQ+5Wm7cbL4E
dd2RwD/pZwKP0MSNu1nnqZvwWKHjbclmW/D7P70BTqM41FFxh8YPYrOKDHM8RqtU
nSA2Tf+UkVnQnehNLBz1JSKKjUzPaBdoCI8Zi6S4Jo0a2oTQ7d8tIQSMmeSdo2SW
XbY92RdpWK+JaCONoyiEO9SBoX5EzjTMeZ64WMz+gGfPOENAhHZPJtW0jeYnBcsE
T4vxrLR0Z8DcZQ5TmYgeGUDiwFWzh5MNZxfBsccImm2oFWQQhuXtVZT10hjxMfGx
o4hlxKrQTlMzja4gSkLCxvXgOK2I3l/qnAY+gBOoMrYjXoCsRRrG5Ad/7KAy2etg
HL5JFGZIcPMxEx+EWXJnA2uaft2BWwPTd2z7pj7geOkejALRIaS/AUnm995EbEiv
/Hl/knPS+TkygAB3k+z2coODV4TILwb73UCxXSKW2wsWfpS8fabFI0tzQjlNNqAk
i20c1kvV3W9HY3bilCL7nVhiynd7DiDdgFDxRPzI6VI+apP2UuXHr8ygndvOMe7z
Dlohx/cuvOXWXO+fWz2dlsFoMri0aM5efZkll3npZYZSS9vIyE1DCKWyYS1IpEHE
Yi9CxDoWMLQ+a2YUiFsiu5oVkaF9Tm6DKYsOqyT9xPhjwtBu+VzUYojGZpLH97k4
IWzyfJP5srVgfUqt2iGkcqltbzbmEEjHXjkzEqhCSkw+7lW6rh/PNXBcjXgbHB1E
mZN2yeifjpN4HHFpu8FgpwCDetV1twdv4OFJPln9GeNVu43VAKp5rAhCwXgQ2Mzm
naNvLS1LmDFX/8pAobngFm8keCWeY/Zk4AqmdLNe+hlM4ngoYpnXaoiAiMzpqGa8
55mMDMWoD08N4eZPfEt5H0KrMjch3Qyu9UjNNK2CsKvmkJkV8laIdIzaByRu0qAx
hnnVpaQIMT5fi9jmBrMZ12C2x8Ka6QEREon1tTOzCgW8OmcyTH7JDbwhqtxr+9/1
ptjq6HWuTska/ryaCCR4Nq7TkjWwVfShCz6uOBSV3UtkLSHGi6TlcyJ9G2XrwyTF
vK4AYFEpHfCA3ILk7arFrYIICG8vzp2R5EBJc/11OBBFKhc0UIcB+6txDRrawtGn
vPg/HcqM5+llRcNaPn/FTQ82RDGZNzrFQnJFuHC0GHp1eeap1XLL6olvavNvReKQ
X0Pgbxoq7FGucvJcsI9NR/OGp/Mb55GyROwnwVlbX2qbrDmF7jSXONaI53Dvw6ya
+uAu6nVM1ozqvBlWmFnJP1sifjsYT/5hMUOWmRBRaMBBX3pMYHsQR801EQmyK1WW
fE+/9Az1wpa+bCsEP3gPqgRGoUuCA2wUSIW3V7t1jyFwgRbda8XyYYsLIpk9iBGO
8kET6a/gAIASSP7m+iHZ9P3Mm4Bv9f1b6WSMwxIIMpx7h71LUIzUuK0772hP9qhs
SB/v8FONxEaYKxZSh/2fuVAi4/ljx2atczWE5P4huywNe1y+5SfQYzsZbNi35/CF
MgcWaVEjtQenkGlqgI/u/81OA893Xe6KYDbZ67p8jG6hrhZHit0G6LuRiQhsWh7h
jLj6//wws4chFNRQebZIn07AXC0qTLVjX8Y6CJ5I3ocEcNWDlDb44EsFNKtXq9V5
gR0C0MyuRAX3IzyNVGx6j7WXT9D3yBoBO6NqhmKAsnE2G884RdhhkbHjwDY8J9zG
VdIu/9sHJ5MU5WWjpcfFwfcT+kK5To4/vAcwEx+isqWs8gl7PrONPlZ1mj/7j87A
zIkwlKndJrdA8qxZkBCnXhuYyA+L729ad77KMKoBwFuq6Y2a6PEOKJVIcrgvsEKw
Iuj6oOyR62fqPZCJRcr4kdd9FafN/przdBjoQwuVpoMD+GHADV5V8sRV9LgQTNb4
p6ivt5QVbUgeG52eUO7KCSvdE9i8Dhtc/8yuD3Xe7R6qf997F9V6QEAO4qgxMWfN
dKFjUYRUvejgQLXKpkx3CCaLEHyr4L+gmcqjQLGBP6HO3xQUdvI/NHkQ/17e0cyV
b0iaAVyce7KMYNcLXxyOPKWZmdG9NOfNo++cWIqpqYlQ49od0jL3MVlw4Tej5zEd
n0PFsCCbVj2cMleotSSbuOdCln417oWlejmp9pPvEwbLnZEvi9h2f9tfE96J6Kw9
+FD0kc/w8wAGwmso9/tTFg93PRrdLTnF3Mz+98AFMOBTbIu35w5tHGsgOsaO2kaB
cQiYy6U69W76PHWrH5NdhnUNrc3dcDEbkS77YN6FqJwvLnV61lNHVT6DHDZxaflh
hSWR/QBhGdm16cKzlBFuYD4rJOVAy+aM/t1reo7cFO14uZjkdphXNJnUJeAz3F/P
s9jUK8BWJkqXv3oXmjVMS5nD1dx1vcmQyC2rqjChZiY9ynGgEyQA7XcZuwiM3FO1
09mEk1bObu0vz2+7dc2IHibvYSIOB7JX+IuhxkyZqeJTy28HCzRYPrAct0JlpCbh
K3PwiVUQb8KQv6Ghh+HBPBa1DOA+JPGhYf/zC94E/gchnI116MXyj5Nyay5k7PCo
gKJqXbNlSUQRe/THwMpVtOpkZHL0OmK4E9pzNpAO5l26oe0S4VSfhS6hj+S+iFMa
auj1mDwnRCnqp8lh1gMi4xm5m3CNzlJ7Rdcv/zHL2WZkGpNHxphoeCUg4uDGYmPw
fAI3NOW9BgqK68wMsLZrAL6iSl1HkcEvEwLqWue1Z00LwU+reg2LwAApnBaGuC+F
62ef6g7YYEpyrlrWB6ePUBhCW1+Bnrk7q+80HvkbwMOXCYE8qnN4AmKDKks9ljWG
d8mrCEEHNFnj0YSnIPZLL9yJsDMh+WfU/Uf3JLf0MMUPVf+t0SuWxGU3XOxMJPZe
WiSubtOzc7xPi79D4ozem3vAqlrDcoyT7YdngrxuOIg55YomwPOP3umN1C1dT3v0
nszvJjFMzpwDcsO26AIucDjlUABVrFHWY7am07L7n0frAsg8o7bPuxknfNmYKua/
hCnKZo87kfvmQsuJg7VqDEBsckwVMMQxgof/itF2jYzcytspA018cMqgF6j/DLC6
+jbbkqJqgNmjgo+zXX6S6Y+MIIm81d04PPreNKryqgQbFnCe9LBcRjTVrLdwYER9
d3QoiZEVc9JZkyr6daCD3+rgHPoTpynROH0g6ZGTDH0yM7MDr1yelrWhBfXcXxkE
/sFxiRnh3SE3BOAJqv3m3Hf1nN/8bKykINY4d/T1lzUOt5Hy3NezU2kKPRk+o5DD
abxknSzn9nalrqU7sjbJ1PMhG4sC/zGN+CBgDf9ecIqmReFSDoQ/pJhKRfb0OQ5F
y2plo8dotQVNV8M6f5cTr0Xw/FdYPXCQ5bItczBn/jz0WHJPkrC9VKEprh7/kyBx
y4yMYRaft9bm9pmKBHuhVrTxTvmHeLrfKHxianI6f9uTl0ZjUg6wyKnjeIFeQHKo
uLvP+eX/zgI1WibQ5XOzUChWeoy62N0wXvb+b8xHrjoIGveUYiGu+90o1CICJjV4
tVBMUXl2kPmwxE3eQO51+s19+X3cnNU+N6fjYRFFMw9BdqYaaOEYWNgtvuT9+axs
jDVmdMiUoqAOEIqAkr6enMpbo6WPgvZrcEI3IGgI097MX4ohMJIciFKlaLRJ5Kbv
q6SpYxXey7/XHk+mSOeIqhwwvKMVBV5HGnkovqr18qzHOKsp+w1ukUSnGDM09o1+
wF4Yb5w7fdEkEwXYEibN42GD/9225g8oQKn1uMLjWDsvfsdKl1Z8CNhG8fzazVVL
JJflCtKcGZ/KXwMcTU1SDxoGs3gZOcM2MFzRXerp79YCaXZsEHSf05a6mXD/DaHz
p2HP2UfBEfqXM7Y1C6jlsSEsD7ls/PPfo600CRXqzHao/mEJFNSXZOr1GnfYZbLG
fjIvHmrD8VVJPeLFNKNXEjwHbbD1ZeUpfKoDPOkS9XFkzLsFeCbCMR5gLKCsaR3z
l16i7+ojayaHQJk8rkTycNLoA9JVZjnKgO6zQHIrOwjEBuPFF97/dxcJUmRfD6Wl
ewmAr1+ULF31JVB8mQ0erx4/uOEF3aoRlWCm+YprfhZbkkV6uEdyLE7fJZo/HME3
ujQmI7ouK6KyvAE7fUI3H4xJkbqQvJy6/IHmMlAw8OyFq03sjM6fXBgRq78YHVdY
8Z/QeS85zYukdrf6evTAzdHxugyRKhube6insQzX45yYhXyET3nB/AwR9JKo0olH
MRuEtNrC1EcVMx59ublyvh/YGHXsRl3XPdq9mIzisKbP+Wlmf4qzWo1bc491OFVF
vbFJfhoKQUQ69GfGZ9XEyzr0p2e2v35DE8E3Pis9STcZ3Up6Dmw/fjgyS5eH8ICS
ER2BO+lC+R8nLfjE53cue9lYCzoBerbr3Q5qLxdvknGhXY33zTFGLD52JruLP8S/
QW1aoDJ7QAfQb3Jn/GxOvLYeuzt9LS4FcbgEH+vRvVDDfn7fMoDw7ZwpX7Cpu2D8
qqhXi4qeHnqZj3pRmd+wSZk9mi+9SvJhcpDPZgZLS2lJUD0gzNGYJNJCaMBJf5h8
m5m/vPjCC1tgWHISSF9bW5JxTLkw5LLtQ8OmWfSxy4Panlxia/1NGMDHHICwoSHD
jmbLBQqYLD7HcPlfwzOJfo1SUwOpGUbcioxDG9edzpZ+MrQ/P8cm168E+R3kPU67
J6BOVyJEBRIAUqxDdEHYtq+uVVdqk1cGRkMrTYRJS1BUUQ7/lmRLyJ12ahhCbmHM
ziyAq4exbGbHfew1TycU9pfaWP4T1RVd0GtYGzufZq6HgcJdgzK1w9x8QlvnqkEO
PY2qUoRJ/G5ALdGjd/uUmn70E+IPPNpn5G2P117ztAXcdamoLDipLh4oGIhappZG
oyAfEWgfXvfxqXqj1xN6q9qFadBNHA1VNuOinQoIpi4wp7B38rxAqhJUQPNxnHeX
REfCGhsKutNj2y4uMbo9kseiE3AvXBy0vVTkBX+Pm4puKeLbdDg3PFjKI3pGw+x+
ILlUfNtgCHhlBOJqMr034XJJDVPMLw7R+fsm9jJTcfYrPmDKMG2gOkF9hcvCC6fI
zjHCjA+YFmXqkuOLp1D34+JQGpSpyrOY4CJWIol+M/LT7QA+czbJUB9JGlX4R1nk
aXe5bgzh4Hjld0tcFctBJoE21IlgN+VOOTge74lGO4ae6VQBfoXT1zo0nx8DWBh6
DZLIEj7JnU7iBJnFYZOaS5y3zEYXR2sRPXRxyvOYB1RtTtCtLSD0/Ten4KrUHkeX
XTaoXMgLMs8xeysyZQ0VO+0kxZRFQAalhqluDjQQisP2S45bCTo3zjlqkvZkChMk
co/1cnTHzSO/pBAjKsRWZrRTCqiODd4I2HP4OT81Wcyfw+aPVV23IvxzYg1MkxlO
yeOGCkOsebv2sw4ZoQyTtRdNxjJrx3YeZ9XrcVb9kXyY9mkk5cj9I/+H60n1zXVO
3g7XlF9+2x70EBetbTGsQtwC1l8Gg/e2igHifVmwwLAJLVQPagO1WfQYxXN/xMCJ
MlF5I8TkT1jsQ2eybr0XZt7puASOS5ygOt0Dn/j9Bt8ZkPFZpd/+uMr3RNCjecSO
HufO8f2zK1Chd8iz2yo+bslOkxYdGNSsiX4/lobrJpxGYEi72yLX86CG1yTcfmp7
YKNEE+zy9q0cQLJp/85GzzcKvOO7fA5+6tE8QTQSJGdw6/R+3/by8rDqbqy43o3/
jErw7Y8Pcs08zw1DhYTmL5jWtpt+pV1z4uD6+NKvNd1PbFVrYX55ziaAjv4zP4yd
prz26BnHcVuDo04ut1T38x2oS04Q9W8u+1PVDERzNWTfdEC9+pvl/s5yE6Xd97tM
fuud9gZvkzF344xvmSeiPksBqvcDH643XAzESkEF8xT+qpO8WaK2OHAbGvuu+74a
fHh+Btb3YFRbI+nBw27Q2WH2+pZblRxe5UfcdzYLHMqsZ8j/Q9hEbMyaNbfzpgch
8DmkToXIphstVtpGFpJNJMNoomWIuVDvLZycnBuYiQVzblVyKj/Wxxl+RA5vdmna
R4sYpSB6OF8+reYKrP7AJN4uvU/Aq5ORL6kCsiLLt67YmB7jPkbRTX8/mAjzkFHS
ldke9KShxbafjnI0D4Gi/OLC+db8oKNAcMLh7GDiH+8p+SPbk98Y17yvUrZg50yb
NxvUsJOJe2ucKT/ZPrNyoterBPbTUOq/wsvHiylqaJAvooZzVyYD9GsY9nrZESXg
oBrCU+GPlVA5MXiNJb4NXePxbNCs7wUHe6O5VW45yUZK+d6HVuV72+pj/tw6Gqg4
R6p3j02hJDZaONYYMujziwBMwxB8rX1e6qvMh3uQncVGmWN9qxdA1zI6l6lFAjVn
Bf12NECuIjrvvzev4LhUpUNenrhtt/dVSwAgt4QQiRD7XSWhid2e3yfxUuW5d1Jv
ipFNn3zJ7BUd82maVGje7akQ6aVqvqNX2HIER04zZII=
`pragma protect end_protected
