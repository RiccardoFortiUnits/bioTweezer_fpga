`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nAjLyO3EDH8SSN1+fTZZu+W7ckafzE0X3qOPkjSyEZgSH0Yojl0YCxgdfKsxUS1y
9XDv3HuR23BVJu8yOcmwLsMlhJh6gvUHUHbPT3cvC+fC1l3WfEMqjeHSs/ZBGthj
uuT2zHyCQv2jRQsjFGzF1EnutWyP41aJkHQdLEhkRwQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
SXL9XjzKum5HBcJe1SUhpeAmgri01V6n7RqTP1yMolO3kxoU0SOFrcujF6si0l3m
kZIEL8oJ2r7hFpJTltcVv4tI1r2l3/FYPfLHxSne32ah+csElVEF5R/f6DznDi7v
gepy4WXsWOH7srw18GoCd1m3TRzw51VSaLunwPvqbIOXmVFyUlHZ4L4jj8pRZ8DH
qSbsYac7GvCNJ1Nx288kPMLUeSB+XrZOt1YqhgFFlnzgenaSgIh1wt+eft7w8WMR
F/STaKnGbthEGcIlip+SP0VNr3gtTYjJdDDpOLOrhAWMVxE8SfoW/tVrncZf5+XY
WmcBlGH7NGG51Uqh4xHnWa65c5QRx9RsQkLAz8ssFqKrJdpsLJ91YOYCkMjbp0C2
hroG55mLkP3v8sxQq9xrrS9YHWKT/VTEHnI/3zW+LHaPENTvWa9K+fQuHQ5wmbjX
YlaDgjnFdroed/ikVGYK9zliHAblptmNdl5e/A0sZupLkB/6xg3eHIioKeojiEuw
qcFuwJGXQxqBojpW7kgLnApU2PybQt8BZEHuVzhLqvB/EvZIGUtajvr/vqdsDFoK
KihAcy8hFE3p85K7Y1UiOexMsRHBJGGZ6PutJP0HSWdGC9evd34tXo5b6DK5KhP4
Vje0TjVQ5+SgKyu2GYBrD9MgZ5T0/RgEq7wRksWaVlEZEZVHefRs6wYNDrl82cyl
yI5h+zqdW9j9ZhJfBB9eoB07A8dQ8uMNOs11MUu9GUvG5+h/EPw2wXlJeQf4y4cF
ZZ0c91OZXab0ZQ1U0Nl/5uToZdL4vPl4DzkEhfscLXF4FmQPVCBy/izoKg87Jx2O
cYuu68gs/4nnnpu5N2ckdzHPbctb7bfOICgur/68cKLMHRw0ngvCdfnsndFKHKCk
CG0jo3noXooz8zZDj0BNQnwGOALw/V5bUPVNOwmSw4Xqdpd1hsNvagKTJCYE8REW
jtvgVDCHznF4GvwQ666BmzhWK+5Dg4vwTTxUHZxHJgNN9gteHq8/vpu9FpCBOAb5
1w/sdrfgT0/3HvUPeMNaOeFfalXxJRt2+IN6Q3zRaqVlRT8E4UkKFfCV5QqsJGqn
eFMbzL5gbVvcgAm9XDO8yTh64r+h+WhYznmzgpKp5VJLwbgIN7M1POEg5XEembnp
w7e/IsXz019JLxIa79J82In9CRDaixE7CfMV+uIgstD+Kv0W3Hbf/Z44k5NHc+At
fvb4tGxnv0S22iPcpbwp6uCl2Vb/aHfMfaJ7660cEP9J3RmzTZ8Z+ScAE2iBcF8W
uyOK4ze5woclTj9HAdAXTTDUvzs+/o1cgJm8bkkDrAwwC3LgS0bkPIqekA51VNwd
QLihNnE2q7aQKv+TOKrSn3o4OJKl9zyzM+ktdo6arUXNWRXiIFakiBx9GVy0T3TM
MNvDmtchrj+O5hlMGSfpHsw1mJndVK8HyKJsCybrfMbeYRXfFWtmOwCv+T9Zhalw
Hxgxkd9EMmMoIOuRU5jBIEVmzreSZf+vkSrKsihrzioEWItCxK8jeKc4xuvb3ogG
XgFAWlOSB7N5ILcrGX9681xmqV8MNcfoNtO2lWOIbaVC//pUEKGRic53Fka43b13
vQW7sS+P3hxTNcQjZYhNQSZEv8l3NLh0LUQoIOPOh0NuouK8RmUd6Jr7rlGF/vDy
5shhD9BxbF0NI7kZ8Ml2hocdueGqrpiw+NUtZJGIB95eBwtqYTVS1PzQwjh9TXEQ
K1V2SF19c36ahO3ownQZ3vA3JLWlcexpftd0cJvxusTU9aPYHQvuLQyxb/lJi679
rHUgItPnab+G+vNWqz8TS5jhN3FQHW/FR//IYbb6RF2r0o3gIFfLz0x5b4vns1sU
XMQ6mymRA/171RVE6hEx2asefK0aoE3QgP/GIkO3GhROdL5iVcPqRfXvyjQHd4Jy
uJDlBZ78hcMaCGlPBdM+6rlmks2EwJA6TiOqe/fEPi0Isht364gE+EhbvHRky4q0
TvGTj3DD4+9sSeQCWVcTx4LCGNZuEQAPG/fjTZ+JzkCyN0LZDKFiN99+hEAoTVuO
2Wia67XEIIAlHvQh0dETkc4bKcWS7FgmOlny7SDS0oF6SbVzdeyBAPtqhOYmO/mO
mXBj0K8Gm2Nuj4uIJQtcVqdQI35H/HudGGUqynUEDwQ8g9jElMMWPjl61oESNxhm
qqDwukn+QVdjsc7aLLzTthCHMkX+JiLkOu5uQWYZeCUFiN49u51MBtNkWlAcIS8G
nRaCr6oE4uR5uelD4xO8BiatL6XkuzoRKqPlG1NFkcog96CYB2RofyeBC5VXtpFX
/df9hr+gPaSLiBchzHHGIsq2TKZLEoeotZM+Y9c4UwipbUUtviB0aZdwSOvMlgaG
WPaiYqIEq6Plu3ME0GFUOOlvGo0a4Yt4KDoYQNkZIKb7ihsF0LTlREI2y05/rZe6
g6IDALt7wnwZ+LJUQbDCgvCecJUsgRU/IxHhvZ5d5T2LsRDjCofcyre3M81DrxPG
u7drtskrBmGLOXHVT4Y36BppLlyvmT6hEgYpUuxZIICypxlRMaPdmWNiwG2wtwvO
82T0dnwCmpdc4/JWOOjA82+xOK22iokPpjyy03TJg1CdRVdxEpuidizzbx/UsCzf
RoE6hy4qpdPJVAF43irgAiK2bCPpc2UNVUdn4pqrjJKtcndL1DGeIGYDjhRiLNYv
PvLmGBZHfoqYGN7SLnKvvqpf5q/ZbAA3PyQO+ZzfecnGEzi1Fe12HLUzdN/Ksr0O
OyZzldeMqM5dv+hxJBH6XzF5i8zMFM6ex6I/6Cn/xWbZ9dI9Mz68ozGQKXVFVJFJ
rI/qLkrlK9cu6UW0TmQilJJ24CAMQi55w7IeK3tvxzIqxDRhNbHaXMMe8U/+LrU9
llnmIWnOzDPKkxLSYxX2o9daJmbm89csLC1rW0P2LryJTm0eFjFVapxFZnoWBQ66
FWcuwdA1VsVuX28kCIUhUe60q0hTS3bNd4+JDYeauRBsl21/DQc8FYdbTDclK8qt
Es4j+8dqHcU4qI0x58W4MA5yaGq+hRF20BqKgRo7bqSIc1DrRiQVMBDU6fJLQq9L
4W2AlgYpNvqkS6nFr3KYEGpbj66hwAHTpJnjiQ4aYQjHIBDMy5urTNz8EosF2MV+
WixVLBpozdRR3Gnpdw70LTHU3roIHLF5lisBTiaSTW//ugKh8b5LZrpK25fNvax3
ikPpR6p2PYWN1nEiGQGKHlZUIHtbisgXJ2DQzpJWelztq29c73YW04JLrr06yCy3
95VkzG87MByFWvTp727dYPv4dmEuFL+TBP+lbt6cYK7xmpFvZGwMhMgml2FNomJ5
ROe+RSzz/dvqcbppzdTatbjLWBufwk6x4ZV/Lp0Xz4j0djQ9VP0/fN3wP0hfSe5T
bwjvLqXa969hc9t0XEqTFNWFnd+/fho44mIu3cSc3YbfBzgP+lhGG152KQIPYZkW
VxMkJSNy74MKvdj3uco9rRntpiNk106SghlPO7M9UqRpwRXytPLRkaYPy3GG1aOm
biwe12q1I/hl1DfgRBpcOvifAg+QtWPK08CQKcf7ShVk2Ap6HLF54AeQvV1W5gbs
eY44hhfaen620lBtHMguxItTtSpXLTO8cfMzmzLLoT3dVs7D2ZlQ4DkvrUv37+/U
FHwXoK3dUxc598d13DTXo/idUIbMDOXskxK5TZjLGtq9wEWvXrDRkasvac63IbsS
tlD6YEnb2tbYxjrVPJwQWsumm9KMLz8RJM3aRnpLqysCdW/PW7GjLomtX2i3N3Kv
yKlEERwBFRZm2soKTMqrm6oH+HC4J6Pz4IAKoWQQLvFxmrfxfW9Wd/02YrrVBLfg
gXqRTcNcyDcHn5tNeal+mxXMhjTilGhNOlNO4lqmPt9sCXUD1i+jBiOFGoyAsqz+
i8Fye/9RjOxC9iQsIRmQe5SMLMXKVb3FX6b9CZ6s6n7J8S0Ck4mZ1upul0YQlo6c
BSXJuvWcOlHgPw97HLHdwWM+8TIdL21tQE7+WLYmPHZ2OQFLS65A2toKbgZAH2jm
ZTVYM3JkljgIw6IuRBFMFeRtncd+txHBKa4zcWBDlDDiQydLQoCY8wZ2Sn39pk5w
qXboUkW2bKq+9hAi8CD0qYSkV5wf8L0okp75rX6+ObUNLqIfrRABq19BwsEc94eD
NUXiRZzQH4pI4rC1ObgxsR5sBT+4czZCfsqsb3Y7uQg/X28Mx5Mx3hI3grkzO4Ri
ruWSpFp/0OmuzFZnvO899lAmUWt3FB5Eq2pVB+mzUwKvlTPvGUPTUv3DR433KLVM
g4O61eiitJvL70MjIzSihblY/c7Bdmb+F0aAcENGpQTrDtGmSYzxvr6ZnJEq4DCa
FjCpjZs+H7X+u2bVaU4Y4ZAcDX96akxxNeSEQwqwndcnYYRDJnPRxQtcvJUH7QtK
e2ckzt+R50ypdXW5S91QJ4pPdKXi4009PrMKqilaLDg7vAmC8MWtiWEr+lQ+9Kmw
DD7etV1kyBXVrr77oBGWJVollwq6Mlm2RW/ibGAHhaC3C8DlZ6O8OmKFqFrVsz8G
5VCjE0SlQ1m8CKSLJ1zWuykSp3uQmVwqAzfIWTEwsFBx71zFClUfOo3OEKKgAA92
V5tc3/RbHtD5zXuVC2tGFVlWP0gHmIxIFNDOoFIEQyIPRs3bJpJkuwIfOhS+WU5x
REKPp+3B9YasaecPzD/FyQsgw3Vg2M2LFc9gbo+oLpeAjEE4vhbBprtEa1vbgBXB
03IlvD/Q5ccNdyCKYqsNgNPdU9jcDsgIA/W+RMpZe6QrLxAomk8uRLNk1FVb7txB
C4DctKOc8Kn3TDkiLnCYuRzRQFCx5l1c5I5XQ4jS3Sp6sSp6svwPvELEzAuNT+YP
GNKWgsJwFfXX9Wz1tYn0qbH96xqoHUboBKX5YUmtrZ6CNrpXCyryiKW1u6UfmGA8
FK9qoK6yQ55IUP4ulDEBG9mptsi1ZVKJ1JtvykWmhPTZjW46fhikD4LZpeU45ooA
jP8uRTOiZPoJEL3dJVVVxKrYhB8/wSpOt4d5cHhx/oFFXtBSKZOR9nwdSTgo53Gi
36OI+ERR66nA0DcH8Y4Ap5V4LNEPxDVgLI9Gnj7rhcJ9szQkYRy+KlLWbvcePRWJ
lKJtlTiYPgW1gO7ceq54g/n5BNp64GPYjIQtAmVTmLqh2NwTjh07lL9YukgJzsXq
vPxR1xTHai9kudRz9PLvRDQkyYiYgnJArz0WjLBeyoX43wI0pKips1oPlXTj5Fit
zrkFcZTQvMb1Z5kbqD759nLfVWhqeucc7zaNL3OCDR+lw0Hfgqx8UcN1+okDNf1O
Soow6Iy4ypEMlGiCE4UnqCmsHYi3PYqJv0RzxnEw2euPZNyH5+XeH9kfzaikSwo7
0dWkEFQYwykKSICi5DcsF+fv0z6RkfBGy8Va5wARYyigqz1ZuvIJSwzF4nPb1Qc/
wSQTr16UoHpvoL9OVqhCeYE1wV/99FY0Ze8K3rzAjxPX+H5RJjOUdgMRRcspk1W7
e6IEpIiuqMezV/7GXt/f4lIygbOZ9IDRwpEFktmTdJwxEUUK2BBh1DToyZ0FgiS5
hP3dlXpCmj1oVEBzQutUSZoL+13TLJm/RvlQqUK72XThJziMdMblbuxE9JDvJ91y
bu4ilnZMzT+SSre8sKt4mzUeLkFKEwGgnefZmoUt3nrK/pnQRX3YqXkrxO5zGE5h
rMq1yKN5Z/lZqrmj1qupYLIwi95CVEnobo5hPTtbAql9nDJRO406x+RPd6rWtyBx
K4gXXUU8YGpJa4tRv+sZOiLqlY3e/Xrt4oyyXmH2wDV/92c2Pm32Wl3cC1cqNzqK
rIg4zzxQxYCjPqEqCOmGuuZrbYZgUgwg55SL+wCTKPB6HEWOhAUl9bgJSS4ibYky
s+O6j1mtlPSfPxGOgzzOI1SH5JK3yeZ4h8DKxoNp1osPMkwCnVV/SOch8QvO9TT/
FWcebNFoKvsP5SLyeEbKyTi7WIH/VHZB62jeCKY5dZZ3FY/KSBlKxx9lIOUDZQ+X
TBX5mcFETD9JXQ5pjCHjX27hX0smLf/1LggCgx9+RYIva8mDt9nTB+gOI4jTnEcZ
sPYmbplSGKKnWUB3vBOIRWKLQy0JH67SsJVCMPbyfmJCteqA6R7jHseF7Yta2ZQ7
G7YU4WYy3/eeW8HgyriJ8lSdfrr/9kPa+pKpVohGYciSubJwY54+3BWPomB+lGLL
roov3tKyQhFy0VfQa7UktdUqTRbMCSL2PefDIGo1u8/3YXcmstLAUYKuqAhd/KR4
6K54XOVEMhA6rG0CGI8izOlIlDx86sLhdXAwveD9KY0KNnYRwh6+IdJgTIDkF21k
jDUdOg6I6hD4dz0H9Xa+1PxoWZsMfTsFf29nQPTuLNlt8BATXs12NGly97eogxNK
kBH7bGn+iNKJlBFmpRE4/kQtPZvgLegCVDP+MNsPcg4x60PcG+6xOJ4lkOog7/N4
/Uq1vNUNdbXpumPVQDecT0EIRlR8AS33N/A1JFZGcs8W/XdtWGK5chTEY6Ocp4NX
7ZBBvgSXZE64WHSbHzrpc3VlN3K2c28w/EuYk4B1Tz2MZkcKOARYY621Lvlj8VSA
k++u9sAjvRPkzzQf31VYf5ZJjqtSxt0t52ZTB96SBI9OTBDrMLV/In4emgbAbjDU
fUtMA2WKDrTSTzL2xP2q/HRB4EwI3FvO8jtMc8O5yFGL5w5h3IQNqk151qMec7WP
ZxKorlEbnzE4Lq9X3QlD4Jc5ALo8A84HPOCZ82Z+C3NwBhKo2eDLPtLRfWEEWfIF
8YufZt5MLGaY+e48kg07aObVSZVgEIOWKR6axEioN8qXbeHhfxsIydJWUY5uG/Aa
RgPhh7WdrjLmrf7h9xoTNbodWVe/Zid4KEti9Q5eL7RhW1orbh6DuMsGKGAuLx44
wSNeN02jYnTSsq10ibs/6oQ1RaDNA6Jf0UGQmkIpHOsWTrP6de1c36gBkHkDBY5l
n0QTKR//RA0TGdEcY772462y53isaagxuc0B5O3VlO5P3VV/htBtwJiaGQsKiR6g
ZKycz2G6TV1m/pN26YFnpb7401v+lFxcVZf20i5TAr4POXx4wkho29qUhPw9YUGu
bOVMgAJtQMAwmAXYzhKq/9Vl3gF/1m264Im21Oj6KkrksAFovagE62YswNw7V+Mw
BZbLwUZgvDtbzjsrSMc+mQYs7QycHj3hx+fRf50sXmt/22/dKlVea+mEdFySHF35
RAuwpzq+dGJvpS4+ITnJk00cCkZxJ7nkfJjQ6TWj1k3PF88jwi/LTqSPi/kVsS77
hs4sFh3dFNGzZ4ck5LTj3/JBCOKIaWNmYe3nQ2MCsyiVdx3xekaqXZ8fMlUeveKR
Ob9icxu9qTCUe+t76Qf+0HQzUF56/08/bUFsLpCc6Ftuj/LSbfs77EURZfRkYQ0f
YKurwxICm2dQPaneGu2YMwIHTWMVbHn74feYwraGANq7DSFmEPn8NWM80Aohd4GK
Mni54pTcIWX+DEr6r8R+FiQobbBm5OsKSHugrlUVjeHuK+KokN+hs1oCwQAhxXvD
mBQRZ/5tJG75mNKK2Zz9oUtUtSglYzL7bzCVtNBsWtoT+QXXOpgjZ1cr09YxdcAA
cNAUNAC17kjLXGA6EfH++Q==
`pragma protect end_protected
