`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gNJWXhhr428pDh27EadPB8EyD+ZvI02VarFuhS9eMY1ZPLvldtBY1BENo/D/FQp/
GOUrJqXfT29tlmLK9m7umaZz8F9Mz/wFJad4VQyHJtOX41SK8dYLyKf6U5ggZCLR
Ez3xSGh4Ma1gj0sV/70vMD5do0iUL/4PRmeoK/sPkro=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 104688)
f8/ioUDoqMeWo1gMoXHzByAzMfqvaJz1itnzBZJXeFGn01ILT1lu1Eu2FAJ384xc
ljrtBy8xvcBH3ynspm+oWe0IY4iXTRtuOdA5plHeExglKk1kUZvC6jlFzPPev96l
dqC6tLebl0PU4oISZexTnqPCF9NC/7ZP++cMZbKIktEltJwOGy5yTkFzTWOpEGWi
x50sIhKJMexlkqzBOBf8F7nuBMNkhMj6GdjgDhuJrVRQQWvtcXsF4b2IWINP0odF
2XO7ftt1IM4IJnwz+OzjjPiMvSC3ucWqbCGKk6u0nTp2RlNXZMWwmrLIgTWMuCeg
JDB0d30+QTKevvZ45rZtvzokvUZYvr36x3aS0pCPCHzBklOZcpnm/ez8/zTM5/sa
4p6luvcktWvezcF5r5yUf9G6Mc1kxZNiqWx7Jsjl+heeIGngGcE5gbtywBTvbON3
vLUZa1xoIHCfwCTVx+/oA0PXYwRFTBEJIcUUERX6esqsFj3kz01hg6Xlc11BjPc5
R+7oR6HNzelCocHCevLuLrKJi8ABv+TQUiuBz1W/nFuDUE2PuYbGdk5zjqQSmAbR
2ceaHZ0OJxf6GyZylCk497/yNP+UZQOq0yjEopHMt3OwMCc9FnbaW5Tgtkj9TWet
rTIxNh8W+BjSdtsSMeOPNKzNJ1BfcSao1M+UWigfxB7GMHqOy6E547vwh4+J0Sym
joXJlBf2lv7kBDt/QnmrPZ+qstCOmUij/CpGAUblBZ9wlyWgr4e+ZlQQuIZpgqo0
GGeqc/heMJ/aASkEWMT6fHar36tmuiR/uEcP+S7HKXCcBP3OCdPpAXytzdGHMEja
t8CTjUeJA8+GRjMTKAIgesFb/rTbIJkTPucNBivI4Bi/wPCROo7Xt01qVtISgX6M
2olhaJ0F0P6A20y7RG0blVtadW4sIAS32gD05mTQ8leLUgH62dpL6uqzFbe7w5JF
FZKbbZ91hBzK1TUJScDH8i+BtDCLnbGKuhVu7J0bCUG54eNBmY54KMahoyMoJbrS
gqcUHs6KXEQKsG9uSdeVI+FetUkMXYjWiyfdu9OUbrkYQKcdwMh/ji+qpXoiG5Xh
2ZCVc750UzAMFQdpHnKoYjOQL47PEB/BhF6in2bqIlCPj04QUv08V7apD6nrDE0s
JudqHtxL8ZWVdYsy4Dgd7Fb9cJAf0aO7ArMOJXtHghQqKi76tge/4/ytwjneVSG9
GOJK0vEnyPp6ibmjP68FADylTrPaKwL5cR+Pn9ewiien9JJTic+4/QP9CDraBkoY
rJCRsg3FFlsnOw/NHi3IC9nQkb/nV/wLE7aBQExeMkgM6aauYJMkZP1pNuiBt+gL
gEPDQwtwmdJVYwfSs6op/qE9j4/4HVz4tAo5uCdb1BTnOZjCpx0dvVv6dZ52CG+r
ulIWGb6TQco+1NM5CPwkb9WyOO1iCQNTs4kmegWlpBr8bnxJk0vO66JyVXYjTgOx
wOoh3r55Z84JVdgESNQsQQA6QPTci1AMmwuXQWO7qGDjhyl7Zl1kiY7ZztDPEzg9
Pq8km74YCBj5eZ+NbhlTg2EDHw/9yv+WY6/g8w9lDB/ASXI+h5ExADwjsnh6NKIy
beY20uXseM0mNwATmjMg1gKlkTGgv96VQjlZVk+OpURnMqPOQV4NPk3qbP1QDIdt
+BOLzX9XuqZmLx0PWo2EAk0GROc2slMmksUHreGJZUd3GonohSag6cMyNHVI1KF7
NorOi60KApBbqESUqyW8TPkFvz18LlAbDUHn6lha0E/+kz49RarKHF+W92J0/K/+
/ljCg4m+8LUCZcVUvAM6fYzqsHRbWU997qy9GpXm/YRkIlXkINmcDyNez5jaTRdO
BwT+lpmlGcDPuqp7zTnh5g8gZibC1uJHIaGyiqjkJAqZBvFO83wnj/j8oBbrUpxz
bdAq+PKRcSJ6HxGdi4EKYHweWlmGAUEGCPKgzzJD5XgF5VltWOLwxj6w1cewEjSE
VIWaqjsVCG2onqvdw+zuEgv4pNI+Cfbus6JP8WABf9zL+0sHEyEOlykXM6zPTvS4
kIRXhfjERllXupvfIdeQcp0AVK/YENxQClJ3skXiHiT8Ji/JX1ZkFr1ltq3gOYyN
/E18ozRsVe/qhkto83Y4fKHFN4s/iAki5ORHuhA6miLQtmmt4Dzin8yDVXSGw7WN
DHlmGYeSBTddF7tvfYElLDjSE+QHwFwrkRDvafILxGPpX7hYDy3M/RjQllea9Dky
Cl4x4vXX0GMB3K0KYcFmbyM6/kDMzCQJw4cbcFqkLIJz7D2nasxzCIqCPWP6ffbA
KprELLztPwQWPPzEUUT8TZqECMJY3qQ/M1Z7zgNuJidrzMrhe7eeiebKf3fETtUy
QwX3nWCk+GWDQWi/eUtY9TO0BiV93c/6sn44PkwzeODTJrDa2EDTlgiFzo8y059+
33RGorSd5LCfGtUHQjLgccDtCW9Q7d0QGsHffKOepT+aWaZyQtSBAWqHkpu/m2ED
iww1Y3N9W7Q+3jH/FQ91Vm2gTBFgnLMqVGlBrI6M5/xe7C3/z8BtzW1BVgpbfdAY
adjT38vBsz5MApdK/Sm3TpMwWlNLbJn3NQPK5DyQaEKzzQwP1yBKeF3lljqcU5gD
1yQjf+Zt5hDHznq7AoPlNnnKqdlAJUh6By2tp4ZeXROatt2vI7byoVydjLZwNmpW
xk2eCwkqDyJ1L76d/Re3FCAicu72YQ08qI5vhB0gQtJPJ4hcWnITqcF4NkOOlmmD
kSl6yP6//9ON78I5RG10oyRCwQc4jeTVNxoQxKoHBSig5ZphEHoXToryUnaeN7OU
qVcntBvgMboDYvgOvRrDVMZgPXSpj1YnCGDfztAQxwXKM84OjMoLPb3T0mh8K4nG
+zvAbW0GznoBOwQEqR9Ff8iQNYxW17qTtncPwYD+nGFFg7rsiC4gyGhRfH/nuOa3
piZRVOlBFHW/4Ma2OUmJI0FHNp3QmMKm+skpaeMpcudu7PxvH4DHU34p7tTKCDSf
HQmNbH8QRXw4RhaZaOW1zTpjNgQNq5RffmVDtRv4+YJQmTZuWJBLchRawuOLctrc
TB7ygkx3HlgR9VKCB72SWsI8zEsHviuqGPQ3LSUZdWCi+3Iga/bEgJAUXQX1TgwK
cQCL0ddcTFIrj3DoZbl3+hxgTx+gsahLvjuoxa7miawGpjkLsyvg9uQbRGpGQqqo
3p1ThuJeT93xGWB8/UOD+qs/Q6MmIfBOf4KfZpv++MXGdmtA9U7cWPMsK6TILlFx
H42+mZ/qDl9rkGjW4P54INaFPzd52iVKuU0rbF+LDrtRmChNovDawGFVRpM7/mxR
iN6dkzdtSFfee0go7SDUEH7MRG+y08/ddMTmGY3gXXYxcS1pxidYPTWg5otzXe1F
6AIgm2U7QCPFg0IYy6Ev+ACKQi1D9u2pvoQ2H99APcNB+qSYOU1piar/TjW1Bqun
pu/gImY4nxRMVTzQn+zGdCirZRqX54DSXniONbgUdajI86JVrFUfu0YJplrzX/KJ
l2VUUVJyTe/ucpONfEgunHw6m3zZxOlEeQXO12Oxpe0o2iikKQUNYg9DRAIprKrc
LOTMRx0nqgEWvte14R706Vm/SHx1kVj7E1cNLlR907zvoCZgjJMD6FLpikrHujqy
E0bo1h2w8JHQgm37aEiGaL//LRnlqZGSl88plQso6nu0putqfNoBjgS9F5ab83u+
oN6XKD7IBZvVe+gOuDkh/18zPuwsePMwt6KAD8oIUY2Na7Vu3n5GCV1G8phX9jTH
sJx9Rg5eo70HdaYUEvWyHCeRojs6uc77bCqdpKE93eFCz4pNU8wnX/Kh/eYMdKZA
zkuPEvT/JQ6qg9i1CUhrsWOY4+a+a9aW5ZiMf+2lozoYA8APJLcyIdpdsssRsid1
p8bsx9fCljWioLKzhG2FD/7fbnaGag70twAooD8i0Y7un8g6jwCTP0HJeSLRW5rJ
3oE6M/OnpNccDRCsLaHRC7/bcbc70yYVrvWZtH53mt66TGVjfQl19OhQ+G61VOYT
150+pffyT3pYV4krRVnBtFhNa5CL+OytjKMKSLmDABcaG0+aqao4V3zANhOkm4a0
mRNbONfPgpwFKa9rt0OffaJU2AbqECiyxm71Hnvb/9DpSjVr3M2fbNQlStSuwe7E
OW/ewbyTX3g/V2EOcFI5KS5bLJRrXXHkHmUaKB7oDXk3KZkG3peFFUnTAmwMIwSz
cLSI55PtzoqhoMhDMVlLnfSXyXdE3Gvjatum71BDF32QgLTk9JepL7KM+3p+MuWB
s2IGZGcAhfeA6Rua0AAWO3hmbm7Wr4y4qvmjjwXI4xYd/ncfm/ek4VT5Aey1Fd+4
aWRwOx3ntIviem4yyj9DkCYE1bN9ykOtgnHgCBbkFRIOFvKKKFF5GvViDJmaOIEt
F57Ab+Wvc3ctEHbY6fvPJ2kI2WfbEO1TOrGNSMP/LPBTVHfT+svIbnw86pNXevGf
rG+74YrHJb4RkOsXubE8o1pcmCp8YDMt49YiPOKvd1PGQPwQpiPGBxFl1Fbu9eg6
5e/yhNCbjaXnKvvijufJgOTGkaXtaOWbLkjIdUpT15r1VHpHMNaBdw5Yb0HVCtAj
TJXs0HD9xVmr4pqvXTUuLSr1VFHdoeZc1afxJEk02OE0vNiiAT38Pb3Xih1M90Xy
Mx5F8X+TYrJUGpyrp08F2sFY/9PdewiGSxJmLbcCAdagYLWR9Yt2v4VXUfLA5TeO
4jjVqtYq6ZXEC+aj8Lv/CLgDhrU44DIR8jBH7Dfs3mXZo4jqGKFu9+QMYD4PCvYt
PK2P1Heflhzl9gBIghXSzj+EBS/xbnIVmuadq1hqijtNU8S7y+YJ/eYa1x8+TF7z
QXwXYKlhB+A6+h7Ol8FN4FWafBGGJ/MrY9hvzoWJWLWEXyAx3rVdxXtUGHGvL6gw
RRmkA9dcxutaMHZcgvvnS0KJaUWRSFXok8fFk34FuyGkHfGMvhnXv6n+FPI6VlNg
PdiCaJcU7yptnujvRREwtUVIbJRwnZ95yEfaOkUyjKekuVKfSOObQr2MiBJKcEG+
C+qrhS0JPjdBOSUz1XICdQ4XRkYvMyVnsu1XLNj2jhbL2eK99LVr12kkk6XpB5C2
9s4E0r5E7zZv1qO6sTONmTzhlXT+IdvjVgG/wHYWCRDWW5sFu/tSHJrzc+CseYuh
K8p7j4KP8cQNBC5wgN9VKWhg4VrEe6GrNwNk1Rqa0QywHyxCIlsnLe4wXJOQDVMj
mL1N3dpRle13SkGRVd1ntuhMn2paGxrkaT/VmjbhuG39NqUNjjPgdlwNUZYTpCiN
rjp6UE6CUUUVisuAIvWDoqb86BnGH9dUJ1br1ydwFZtEblwoq88lDLrL5l6L6vi8
9+7e0G78LY/kuRdJueBr4tsEZZH7EsVlzJUeFEQHuNjqlfarRDb1f23RbZ5JLl+j
tM8Q+zpuV/ohPkjNie8mxcE6kDkAX31VBKBCmyPSATINKmAzO6TgNalHPfCrCMnc
i5YO9gRZDPAEu4w0HAjvFNc5JWxr5/HUF7pRUN0YIE5hoFrxkTkw7uLfcreuJ4ez
TOCmUDOLX3Au196UEeLKfKhv56/aCKhNDdQMUqMHW+y2NYQ22gEF4IqoJdSakfaD
2SFVWHdnZAIEUT+9jmG5aswS6rjJvIC31Diiiz34PddXtTGHEh83MKxbUvCFoCE3
QF3OzzKc5qnikC2AswMu8I2iMSGGL3h9TVMw7SEMKlYp4r1EZNpIwau6HQ/lQz3W
+c2Sj8eHI3zXvSuNh5eecuAjdMdla/Aj+BK3uI9DNuoemVyJlDTk+gn5jo1aAbaV
8u/o7m/1CBFeKJ+03fkSSFoFojHg+aFU32Ja8Lxao1YwK9MADnK8sUhWni89laIh
fC47lDcue0gUMJJmgh39rU5u00F1L/NA+U864OCdB59UhLjx73rCgN2IxpYWD894
lRZwR7tUcmTbmyaCW+0Z1biPWscRgb4+aS5LCffKsQDC7EIg+EuyQy9TDeztCEQX
oB3+DZeZ8iERlu9XUj+pA/YM39GHIRwnazpFYJf1yy30D2iaRZkBOjhCzBiwBz5M
zXU2jrS4hd2b053xsok/3h2WAeS89lZPOTDx7+4G9eBAsescum1sCELUVZLd1Gup
wDQW7/LdDN+joioK0/zACmp7FODyuCk8VTzFWDyogvGDyEHLXwYLwdDO9Cq8+IEq
i6sRRG4a0BoguCgB11TsnB+DzGeLaOtrlyr7GjalxclMZxYiN7j2JWhj+4oPsolR
rWvfjH348ewl/HnBGiaP49R2nXLuT2vdq22DD5tMaXNxD1NJgXYKI1ApbsIIKusH
uqI1BQsFN2Oc6BRcwiYzVNZDiOtDNVePGp8BUuAcXetCdSr3lfMvqUsoaNPTj6v1
5GLGKW6GJuBUleNnv5wh0H9ghAg/QvJjMcDB/d19MhzIEJRbe005ieLdcScmpkS1
bE95f4ykODAExXzUVZ2Uqf9WVx5AQx71g24zl5QkRg4C8dvcKW1YIhg0LLGLr+pz
f/l2ikKK00BXvwN98jvajRjtQ5MwpW3xU1szc4gfo7Hy5naeFuZWvy8mbll5+Vyc
AEcADC8bAmnzG8K8AEJ2Vm01UiDMyjujfc2SgWwegZW5XNlo9tkHJc4knTqM6k/1
/xUavDg8RQnBpafFeTcsmVmGYFWnKISDFbLQrb/N/XIyB4WPIANsQpUkqWETk4kY
Tfs2hOv8Swu9I9qylQy4aR3C4XuXJyXgTmAZQZHwI5/sAtxCg+yIH2bcQozypClo
xcQqYnZY05kwfoV4i0yWVjKeoqJ5vRmo6IuUIACFKvIZPyZBcYHVnI//TEkyY5LQ
2zV7/m/Hnbeue0MhyEV+zV9+yxyYaS39Y8vmm7/sPp+y+gBdmV4mW9UH0VpHWAPq
pMUTgPu/9n+Rxl401BUsq1pY61mISb2/n6UYg/0EDnImp6p/jVmRLQo9uJmeu+ph
mlVqEBKSgNcC3EhhRZNM8oloxwr/kawsL3ILbesbQo0+aRRstq0QNQXzVjVLb1X2
lnYXnKPr3Gzg8yvvtidX6rTMODsKVDDejBJM7mrFTns7YOcJJvCiUq8OFnaEV7nV
ZPAKsmjWhJFNgefQ9hOcfrcYPXUJ382V3CNWANMxe1K1sNzghHaJUQsTQgFrYsUb
O3+rruv1FRVRcv3Nlee6NLOSL2BiAuD8dUWDiA5bYwdz3NpolJUcCa6XTLebX8zb
YEMEcpMiRNcDr8UNxF8Y1QPaslItgOlcbjdnGh0rgvxc49UM96yqAIh0oK40nfgK
revE6EwU5CYv5s6aIOG9Sof6X15grNHqQdH9FskAOwl+vT7FJ3bg6Aw0p349Ait9
NNwpsU1WUTGJapNTOr0vat/8mJqz6c40VFyA5P/qJZ/nJi8x6wpGFGT6Odk6UNXk
CY9x51tg1RNAD7NqHq6FdSUL9zGO/IEROJx+iLckrABjSJbthlGOLR8o0daWS7Ss
VBWv8pkqwv+1z2JTMp5LYCaWQyH1DpbiYSwEk8pxt9YJGc3UjK3WZ5Lj65DA7c+0
NVORw6ipEuCXobfaM/C3Q/FF9aHxI06SgIaGDwE+bCVOLd5bIY+0lG6E+OAHcR2Y
Nh2lbkiVGThpOfhgFqyIfkqycVsgOCAdia9smuVymjMLO5pHinQ7HZz77svkedMB
Yube9q07cZabaR1Pl+56oRS6MrbzO6eliYlt+JB1bbodCe1YYqJoAulqhbGk5htZ
zbew6XJud/5bj611C0GxiuK6O/DooW84GZLaPunENg63m8vm7Wx344cmXmi5sIvK
dfoXIpdK4yIk9NOQ6z6jfqJl4Uvr9aZyhPIAXF6M1a5ip1QZwY9gBB4x58Wsqr1U
NEtuzh8vhBrf9n8GKhw9xHdIJwwk8hgh9cLvRNKvD60LGauwAExZfWCdh+TL+q4R
QHiZaq7zEnHj8/V3xOSNwH4hPSq2jGco0ml97b9weMs9I6wU4rp+ps8gVekJvO5C
hf4SgljGmE3qEMjhwlhmRiuek0bEcMTb/FS1ClaziSzqULhoVnU2iWvgDOLiwpYc
1URUaNHAS1Iw3s/GvLYlAWB8TbQoY36U0n2Y83Vny943Wn592UlxrsLfj+VIISpD
XUK4vurjA2v81DjHivsmjHNpE3+oYdEPGWptbUfom8kXFi8ybyC+Z1s+yuEOCXbW
16/uOwh1eItTdlrkqDqK6iiX24/xFMtpJqrwWRzRp8xTGzGdRsqpqRlNFAfEz3Yc
6lAtdsQMi56SQiNdILfy5TaRiYIfmxe9YnKssvH/JuHqGc1ClLHTjBthzVJnMxp/
HEjxicz3ESmqUbw1wXVGcM+aoCQJ6GzRpZreS9ypFtv/Ijd6psvLdu57EW0ZFcii
C9AofVSTgyrVSngHJix+gRPzrejRIuvzRQHx9pvV1RsdRu26Du0UqYt9bGza1H5P
ElgCy94cMrN1NGlsXj6Px0B8FgJrWtwDZo2/880b0lkqzYs+7C7K4mRXEO1TlLXo
E/bvWEbUs2/Uy/U6CM/FTx/PCOWILcwqiqjamRjFrRxf7PIw/6+N2Fv3djbnHe9Z
1aKYzppzhpdBe0+jQ8wFLvRtqz68jDD75YmgqYVSbdp6NVXF55O8GJZiUg7blukJ
ROeV4CglAsjHjQzZRstIeiNtSqZmVi/bnVZCk1zTYwWysxiwHorTrTzgrFn5P4F1
oB/qbxECqAjFaRpE9bWrE29pqonwlpdJS2uxULj+GniVOdneE91bdeDuMBwkzqEC
QW+NPM1bh1mI+UaEHp8ci94TQxsP1ws6kD+yPELmHwtaGjr5nsTljTxAniGtBU0j
w3AbVxRius9SjPsvdP81TkCzTwDuygKBCesqoHOpf60NUx1b8XSNC7p0S0gIGDUE
adKWoyrhFmwMak69N0aP3CM2+eJeI/bNLVV/SbchKUvp34DxiWmdnDnkRNvvIW/P
sKSY5/2/fzCQQqy1yc1bzYIl/sT2GuOOAtcewaEhPtDDdGmkk6tYxcM/P/4jeN84
KMLSlRLjqi6Do17g6uH/3tQUDQVQrSSbKxkw4CfCOI15Bs/LHW4zk9fqCm/DDN7p
9El8H6qnGaTVktByulr0mmfiIGKQEFjFLuUZVKeWN4qid2GshG06594igAjeHl+N
f/vZpq7PrCX7Lc+W2U4cTkac72n3qYBvE3BNdfEoRNvx9KZyiZMZZoh8zJxW2nY3
w2uEMK7vskgGjXW2rKYYfbyYIziQcmLbb1Vn3l6leJtmWsFpa0DdePkY1XGgtVqC
CBahAiQoRjgs95lBPu4YMn8Fpa3bcoRXK3xGogIO/DXZAHXpCVVb0HfqWCwQX1gJ
BM7178662LJcJMxWyidpW845baZiOw0oylL3dhzM5ZTdCkDLXjemu8m3EKwjrq1E
s608mzUTyJ1Udu36EeudVbKdKQKSf2vrjUYJM7S8bTgTTtqzprThe6nrOcjWrr0H
v8/8vhFLryoylEAKg5wyrDcpV/bgrxTXJF9zGq9I9QgCKIiXEbJq5SXAyLQ5L9i0
NxDkHQmxS7379f/67FTFoBHyJLIkeMRNItK09ORqguN1KDSELotD7UYEpAGcoW6H
P/DhMiH4ulH2RjURsD0dyIl5o9UrIRt4VG2GF6CiA31z2JX/2DLKDxfjj3upY/yq
Ev1K+XkIRq0TZBsbQ0qBiaYxJVrQDEzbmL3ZEjydjvEQyIyoO2+1U4vYTAmdjBbR
NakbHl8P5seQEfYE+Fg7prp+0ANjt0nPv8ONq9O+LqVH/jrqd8dqCZa/kz323EnF
NMBCRxPzCV4qqFbrBVrfXn46lGjrGuCCepRfgXrnQwVrU+lx9i4mofTLSFnJxKsa
kthaErunB3cmph40G/HtFIK/+Lo6lHq079Lw5u5V/k0OA6ebulrT5EHfNdjG4DUm
zfF4NGD5mfeyeOmNeNlRLsqpq0giS+Op7KA0Po9UaNEvVl+fTOYjKbNHgPEdTZqJ
a14yhStZkKsl/liM/Dlc7AWFTcQGhKPbHZluZweiSuMEs1TjRYt9xdYhiFdVVfwI
6OSAbGcsA9unzjGbNjCzRqnPyqZdVKRgYu5vJO7c7KNRw3HC6pJ6LU1WWdUvYwbV
Xt9ElO/5/8ZPaGQHTVxblMIen9wiHoxOdp1jQ0R2b9BxQOW0lpiR5wuRrwH6XN05
ImnC4FR/hPoytmowVPmUV3xw1QRUE5q7rw+971SDxw+au+3FZ/N8kzItwn1rgC2K
OUP2h6iTwPv3DBAjhLd43gNDext5Qo8+7Mi8zsaCFmF0JPYBudFAKspyQDd89s+E
n9tUPAokTL19U3MKK3TopbrhXLtA/5p2dpgXFsxmvl4X1losYAkpnP2podICsFEk
Sy0ErdWdWyg+71gkqTQOWdsxEmpgX+ngqDs/84eO0ADqhdf/ufgGfD5h4mYeEvs6
maEYdYlLTaYUDYK0LwnI8UTwKYIIVDekfvw0YwqJxG81eD6hq1tCS4koYObDb3Lp
GhHier4G8looJp6xxrgWtelzZnpF2l9MbhIQDwDUMQlrc61wx4h48H3zkwUYazBF
AMK0vROLN2Y/oEzR19ehupUfcKAw2oNGH8gxD1+/0tStpIoijP37IXtK18symRn/
iiOTQWgNLYsGPIbUZpxj8df5LdiRr9vaIBifEZij/O8U4tVPIbHtWD6HFadGrMUa
7gclnRCkR16KCzI1DbtuDuIbuJl7n9cU9F+v936jxuV3R/ZwREDe2z4xw0e+DMl4
emOeBtZJBC+Mx+3zM3QDhzFzTBtKHtyIyCBqJhfHNox6L3FaXqWFA6XsihbbqxOB
aOMeRdDjx29DAapkkIOKkw2/KrFcm1L6t5EC2HjLQ1VoCsUkhfyRI5zDTm0cnDcS
Ts/d8YLuQgafbyQ4Itrh1j85Y7mvkeFG6a9+BVjI6237XM2+FzeOohEcaf2GfNaB
IFK0CN79jcJjc6oMs5yMFVgtoRNBeKPh2MVipJLp+FpAPz7zC6QMIpqCPg57jHze
gWabY+thT0MG6G3nU18yvrAevRSq83tMGRd6N+xRtCGrLSLCxvvf+4OWo+5IJmyh
yb2MYddh4IZxnX7/VfeOn4ETCUzQlbii+Qq60rU9vNc6AicZQo8DanPWKFa2tUs8
teaSJGVraLJ+8IBUpGiCS6vrYVU6gjQgPj4jdukzYHeZVGLbG5F9cV9RYHtIwHuJ
ECSoUQ7J0D3yNwpnj0pehrcNFj7ESk3G37e/7bz3NDTdcId1x55yyRgqoWCUrO4C
loEnhUYjv2qrQD8Q6flYxvC2tsQb4ZkqD6lSFqToaCfcoXuFemscuyqhYljiA8pa
fr6P4P5ESLsSUDr+P+XVbZS721ACPmPSXqvfyMHwtwFRIGDmUpmf67iMZQJ7iUKB
EJNJh5wYhRpLH2hdd/BL8NEGCKr9Mpr4LcevSEfZYjOd9nRpHHadL20c1eduRdHr
OyrR5zFONRxUzh5MqNjknSt2/1BnXXlztsNbrlGpC6aJWPqYWnTil9DqkpyjLbXo
0GvgwI03BA2A1Gwt7HDGm+iR3LdfKvJ3vBPyBAjjYY7NgT4zlrOx7lLT0pPYWJCh
bUavFsIMJvBxFbPgt3mwP1EUE0deTKAilriubHqfNtHt2jPmzRYmCMtqHGz4kKKI
dCahCub0S07qu86al/ULcp9kSvrGMQYXREq94JtWp2JaD1mq8kfi4UvDFzJx0RUB
JLHoaXg/fL797+vI/6mVFq3fxPMsofqk9VxDD8HfVGiKfEb3LDQzwZnOvBEBWOp0
RMWlqPS3WgMM6vE3kLf6wn1jtqSehiU9aIRpMqzc5x2eSzT5+gxaiaaq+cj5EFu4
dZeKxCyqJIniGe8gLQv4NgE+nM/dee7NCMfh6mkbQ7lAqudsl+fYRE8TWPRCym6Q
hXpfOj7coZG9DiidF0Ssn2NLkS5GFmHuejMm5/m3eN72Op0hcEVzrS2aY++0zMgQ
9q/y0aJgPjVaOJdVOFT6G0fdqV3iP2sFoFzPuU+ZMI4rcZGhFwZHGbjXnnxgkJet
Ic7CnFOmzr9V+PX4mzPZtIy6T96TqLMD5DyMvlegVeoAzq2t1/uluCs1rRC0lGCV
hB9JSPoyiZZbb+roYyTKQZ+V/AILbCdQBwzJYoHSkUqWvnGn00d2y/TfEd2a4bbV
Lwb2dAGevvlqpBGWRDra4GC3N/+K94lg7sExC2qwGPclyeTqF6ioZ87Sw2OO3JJB
hT59y1ptczJxuhjlziBV8MxiOYwib0kXjDqqlriseaSofV4eVntFXGxM8jaBFYPK
Q+dVcDKglG7MRc8z6oAcjLxeON/YAZL27vOiEFiqHgCVlm9qi9m3o1uMu6qNQMO9
Bcs58X76r+84Ldwtn/F+TQmPgG4u7Snf1/2qgiCN1DMH6bVvh4lZtxZ701APEtYB
FvskiS/v1oSC4WvMg3zoV9yTDKJBqcGHuZEdaHgzX9ljWPQp7J/eoAn1hioS4skC
hHqJNQ8HBwkVFHC+UVtwFLVceUOjqqIVKYKzTd5vK6Qvr2uq6qXXQaepw0YjhpCj
dBU2wbPKx+B7OH7deEYxU+wAcCXBEbrdKeUYh1E7rsTGdnI6bQLveq2ux/zfo2E/
WktlvOwb61j3Inkfqx7qotTlxIaRe2IuA9eeCROhm7re2T93sYx6tza0ziXgckXF
te3baNw6leP4ERm8CziVFe8OyOGmhvxvHybAO8kEJUK2URMuiFxEelMg7aQEMpi+
bDGM2CvCGRfmIufbD2iqEE7R1s34uri+3/Ug54S+HkzbjNWkecC4jwj42qtWeJzB
y8VgzpeT+4gtmlCooQ+cX5FogCpFCdn/HMdwg6FmMoew67J7nAxuvfiEG7SjTKzl
BiCezKMC3ljfaFqgW3/iYKCL1o82UJxwKYqG0yFl2+8DyHnUqKFNxCt40uAZIAlc
OFbFoAJ9E27oQdIag1f57n5aDMqBM9uWR2NFgsPEYRUf6Cs3IpDsrMVnOVjylknz
BYVDdaKRRC36/53TMSx906+oX+7bLsF8PNTIznFoobC9T9NOFbjO42Qw5AjV1kJL
VJKelQvvr7vfi1/1cA7rAkfY/XROBOwVL9ul9cUXxL0qQCjgKdKaANO3zKBncQ5j
fzz9dcpe6/8ZGgHzp6yeIFEHpnxMO/XCtNxvlVEDGWgZTVVY6fodeiDZiV4lbJkP
FHZZkDZ44i06+7NVigglTOFg6A5kyus8t4mTAzznbAwW/9MicEWtJh4SRmLLKze6
wweBRq6QaiOjj/D3u8Wi28M2tHblCWVvOwZsXIcGRRJNZvdFtcMUJ1tF6XvVbm6s
FVvkcA0CbPo9VYwPI8mMDtZ9nHZyd0stGwrE3S4ENYSGDMuDRz/Nz6rrk2MC/sCO
FPB/jUllD9Jz/6ZJPd/IsZvn4lvSuAnsANEGZTyBLjw5rf6uDBVJXJGcaG3AGiiZ
xRIhbC67ALdDxYLwDjQ46qsRx7VuCHlUB+Wmx99QCGoqijcl/BAfJf1t8Ar2R06D
HJzwbx+sneaYNE8jvc/6t9KokZeKdyhWRsMITwHnaKMxiNr2UCrXVP0Iykl46U3S
R4zh3w5Ubo4mHehmlABtqfykSTyo73drEp3/T/FBLRsU4jI6RaGn1hPAa4iAYQ9g
fAPoCMY92gFCa4cXR2ymlx1WOGnakybCk4w4ud4YmUvdTrf5pfRjDAUimv8P5nlE
ofEpTBzGhppNuJyyK4GHH6oA4fqMOcND67lVkslf8xzJpicvCwzlb/MBsHh7Jttv
hb3MOP6mHQJ+USlazim7vbs7fD8GBCA0CdjZ9xgFpK9w6AkC66cTrwugiAI5mNGS
HoXNMgsQ3m5rXoLWbIfzccc95G4QrVRSJlwucFDSDk4zaXFnL8LR7ZdzRUkt+Hg/
RfgoI6KPiET3DjDZrdNfs1DQ+96FD0SRWPI7ubYziYNUMCvzRreYRIN5vYnJYhSD
+1ZoBEjdiVRkfH5mo8d9diXiScIlf0uvmNtPctsn4BNZ3vLFsalumW8E0cd4OAKZ
fZgKUNF6ervAhgneBpLnUz+dwm5uj2IJgMODSHe5YlIsff9NJ5cUWtq4aZ9Mw9tQ
TQlOygZAbNxe3nBk2ZfVNr3HtlPmpEHy/NqWCpkvoMGDsx+5NWBGUDNtylIw75bR
BPzvuyTA0RE4DXXofnaAXlbWV2nO8CsD9H9gAlQeGFh2970dRc7w8du4mM7UOGmy
I7YwS/NhCm8Co+3j26jRHXCHxlYpTd3kDR/ZoR9srx7qJrxPTe3uIBWHlDD9EWiW
AmnKwZ76FGcWkfF6aTML9Wus+mdGfVxqEMhkM75nZVgY0tFcFv2cDiaCwgAPWSN9
A6QQH3KqdBAAHD2GgpZc4iCEcWeehp7pAH1uLkXXOGljwPK2l0zsHIP9ZSHOmrH5
oN1ON6YdO+cbRRXXHfpjC648F3Wtn97Wa65ycv8DtMng3YfgAUpAAcwGNYEFcRGR
FwfVcbqAS/+7sWRqN8wxLB3bF6dXK+xY2VyPkq4hNi4dXtsfqgxCEX0Tu5t9R9an
ZK5oqb1HfODUUnFLnnxcTETI3Ax7kXoGPTiBN4dXZYiDJEhdUntSO5GpXSvmCqtB
sOOLBOL6QmGwe8AG5IVsaQE57z8VG7igZf0oA9bhifZTB+ujIipVq8usPjxfTZpO
76GwTSlp7kUluH564SVQPRWUxTF7HolPPum3dFAehWIFshC8lOn/M14DtuB8ba+6
7HdTvLtOzw5XwLUFdcjB8VheNV6oU89Wnz+/hPpzYsOyO2RufdN/W+QGQqYK+rgw
nEBZtSSEtBy3qShseUMtAGZCIhoFZpLBD9QzEh3H88aQj66WsK5hKWcgLSo246on
BjisOumLow2mnmqcDbr7zQXifyha7xqIorkQhN50Vy8CosMmUiBGnv2YXkgwiuxK
FzNaeeyzZxy0msHmZl3qryTiQO6jQJ1DKq24jLwDCX64bDXOkdgbSl6Rt4Le0hC6
IQkugRhAw+/a6jm5Tsk4ejxu5BQZ6CmwoQ/sXak4lbp346634hYy1ABz7Vnvt8VR
S9irZObrHVa1FAaWjpsJIafgLAlurAYgGEUggB8+zCPM0WdVb3TuztdE7dhklcW0
5Ew1r3jvGDha8gmmOqe50MCDFT2QkUptj8eLugy3LsCBRlsvjPouDR4dghXA1pTg
kpXUr5m14ehundr99kMhQjNAQQ4FXp9L6MJHcF/KgwR5XCDxel/sMda131TqVHIg
49cCdGV6hX46FnG7nTGode74qC4OBmm1MHD0JnTrHbOq5q79JFX+H/GWypiMD6XM
sBno8LsGqqQCu2UaYxtXBK0u25BHjGhLcAyzo5DFFXSKzvMdhaKIwTtCooDX4NQF
U/KPgd5h7BMwAREl246YKMdPKlwfiePihrqlXTmzC3MTuOlqfd+Uy4RH37Crl8Ur
3LhtIZtfQ+nBBnBX3HkSObgBTMzoROFhD4wDtut+DvsRd6AYVAvzEllNwAKtKEWV
xbxIPSAGqikU0QdYDNTNx8ypV/6xWBgClO7hZIG+T3CJ3AV29uF0zqlE4dpksUvU
LBbkeVG0w28C/OZuJK4PudMlPHuNIlmswGBWtSQ01f8222Q4D4N3XNs0m+JPjtuY
R0a34c3HzSAT8k29+THgkhJtJLrEJgHYMPh5gOHVSDzOPu+4JMO2siNBO5aak6o7
pPta1ED28K1d7xTTbDQeDAOwxr6Pfa4W3L6bFZnvTHP6y2FzdhzJhdBJdul61oLa
VSyXDuYCJQNqz9Z6bWj0VZD4NV/6OYN+FCd0WvCaGIPbzqRX4eh7McQwHEzR9MPq
U/XRQjMBGB4umdJJ02YwooKlSCsFIUOSBe3nA66/1lo6GTzEQZdP/5aw2GDHcN9l
fizzj/HHdMM87RpHaVX77zzZixn2t1gZv1Ld2gMalGL8sLpQIuqjP4RO7XFl148m
1wgpF1w2Y0URfvcPx7yPewTJSJIbm7xWcd3hDHzlCiEtSUuTQWkiZ/MKdkOjJ07J
nrstjLr9Cg3nj98EVFa3oX6zDexZ1nptxjwgRyV/znmCYI34sEhNgf1QhIXict8a
gleYkQkSmLzFFu//EX2GPj1eQBXAldy+p2waAZcn5j7crl+ROkdSgMw/y9SHljsU
mB4d+4xeJEfksVXhTxoDTHD+YmubBHSO87YrGE6jY0tmCJgXlYxCqFa1O+rWiDnP
yGWhByORVBSqaxJ17VkDnLR4alyOvgm0R3KR+Rl7KK3dnajORoGeu+xnywZW+aZ0
7inDypD6R4s7uBBhtaT0tklHSDLvyNKTU5OcuwDUTp2CLkfsYVoQB527lh/6L/Xv
eCZx+nEWB69hUYxbAKv+Y2pL51ZMijVnux0Xp5i0hy5DwPhXcU4Fbb8xHybm17mf
v2xdQWDCoCWCDajoRoHXCG/qPSnESkv9Po83PtdtV4oUa2Iysgow/FkpzSSahdd0
5uZUD1cebEwnphgdbljAzQEehQdYkE8dlGOMs8MDBOVsYntmchf9w9AsAS+zFxhj
RGfje9PLkuNntOAq/Wa6VJLWytUnq/M6ST3d8Dxul7t9bJEVdWV/6C6WUx3UM37f
lNe6Si8fxl6Wys45gKbubnLhd9jCfw2/Gpl8qOVrgAgEb6E02E9A0YkbfYjxfaCq
DPPMuDIv07I351FDrWTlZ9X0BlWnpl0wLgoieuabHmfham2mD2R86T4ZgN14/HXL
sm5yzoZwH6QtFdkYph4UzAoR7HVDtqoZXuUT62TrkaMVbO/0LieuM7jqjmxehenk
gWtthGNOUoIrrKjqiH7d+sUxRV3WD+bF3dHtFQN+wItMed+SuJwWY9kqlQBTnu+Y
yuH2uPiBto1+WIWG1cIILLZAAN6KpOOjBt49r7VCefE83NfimNay3DsOPInH5TLX
fTp7IccutxRhUoybkazjpBptjerFhin/SjdjMPUKjfaM+R3y/BAWJx601UO6D/j3
R3XVIneOeSQh4zaFQD8bDAzcQdQU1WNJobcuMGmKqZ5Lx0RKYkQIz5LthzfNRS66
n7CoKRBEPApbGy7V7XFy5IaubrL4j8V44sBiOoj8jRnckxbTM2gn0tLrHxZ0JWIE
ilik9d92Z5Ro84OOAc8eAQCHKKHHWUD0QHWoQ5mBGwue3sIZZiJzcqBEY7tvL/nR
P7v+m2IMHNlfNnrWTNXdkJmTJwUOQWsUroHgnJm0tcQBXMl4aS/SMI9QSwY7E3KW
N43IkDDKP3/TCDnmAPjueOTNxGNJ+UR5sZaa36P3oP34TkGsqnSjdV5ENRjkWHW5
9VIHbtDNHZZH1uqw6y6Qtlw/WgLiIUgkbzrszokUQJSZy7+oyLGTgHkm73FRqYtO
akYm7mUUh8tJSIgUcIVX84LGagGvJ7eKrjM1Igsm18Dtnq+VkSnj9HL4v7yHBsd3
GaS6+GLg3ePiTBAq32F+/BEydowkJbNfkXjfOzjwz2o7UX0uappJxjH+oMWPxg0R
hRWDJP/CnJVMbsf7U7MOohNUvcb/dLsSJFB9fngTNyfZgbPbjGdP+szLJH0oQSxx
/Yl3PEoyNLx4goyG9oBPRpHkNq38FMtWhzZfwGVfLrUrEG46mO2OWM5k6drjx+Oi
EQrjwZjwM2RgfvlMhvvMZSAOXmRT9YwE30CGPkLNLjBqoYIKhM/t2jArDn+EFqO2
Ulu1dMAU537ODFicuJWkbZQPfZ3Ja26bu0vtYkRiYLuH0307wdOJUQ4QT4pJ4SK9
gkqHaDh6xU9oq90G35YDUy5b73Q5fWTednzaRzNWVbtXZ/JA1S6uNZd7JEbC4xHM
cMF80H53K6ypzhyJzimdF6KzLckt95sIFDjTTvJcqezJSJNjZNtY2VeDHUx3VVJ5
cbjixT9szrP7G02+rKztsFOAPOl8RU5VSwtU9SjUaLg7jfnw49dSoaWdMuJZnX5l
t90hkZyy4L46PfZ5I6IKrDKpeH4qd5UwzLh4SHgCBy6oEU1t5Ys2/iDOOxca6UEX
SVHkPtr3bDxi34EutfpWQzEFBQpahuubOQvrW3vYAi0KK8+VfC5+JWhdaxgn9vgZ
O4OMUSpBsFxGoZ7wusaMm+5yt3JS5e3bYIyPG0+TXvgyjO01mmRD1n0nnsY6Pvw4
Qb71XWx+p/gpA93PUUCoOV0e/Tcw4G9HGpr1Lsmmskej+j50RVil7M0Jlk7ftFYE
qq7U9NIt8wn3X/pLCACfCsj8oC6uxgwgOjtPVGHLgtVx6hnR8M/WKkbcaCL8snJi
TkA8mZ+4P8ckQNcR4C+dUFpN5i9NPzepcx+7g3aLeCsiiSQRVNs0aj/QdtRGDShu
25GROLVQQSdsgNWMTHYDOzT7bO97Q5bhyembXJbh1yp9XpT0zfQ62SaZ6UpzAEMZ
PwwhK7tj984swSbxqpDdL6aYOvd7s0U+vT/4xtY1w7EGMS36Ux4C52p0wgdFyoju
koqYlMIWE6S8h8NCywVxcijGFwYLS/YXSd3fPeS02g07sNW+WwIJQIbX8nxV+xfI
aq2xW3/RzavtVPoc8iWhDpnVE0cWd8iBworcE5YMSmM2QESx6EXg238mbpGTCefe
FNZ4Qx+ju1fq8iSZUdRcaQ033TEMabz38Jb5Lr4ZZgtB79yug4oREqKJ4kIC07Hr
DQ4MO7vogO9EIOsXWxPiU6etLhg6STsArYwwSe8ypnh5urclVAEZ+Eu4GjbimOF4
tpjCZS4uXw+U/ubX49bXovNSRM97IIs0hXMjiofEIBAm/pXm9IVGxVwKAdNhtMV0
E9NCKGpllfW+iLJglBm58RteQQuybcrIuXTArHDBj4tha699Ddjd20te0MIXWzIC
rkYXGYtCIhuyXcCWt2aZqZBBbfN1SC9EbFBRjQMPpxTrVYkYeF14PzGaBfIZnhyc
ZnpoEDQqnG6zW2iuuBQuUbstu302qocFQZaT4U8AbXF/ltZcRzUnaTmffRSzsxgL
XHczR7g5JLbC/M+oWLyWjErzeu+K1DSSZ0V7IHfOA00mySp5WdRxd9TVxjsSU0sb
YOswqOJqJArDE/EgexAms8jf00nRiKxtUPsX3zXFmd3kEr14DUgG8T+567pxyMvp
pWOPDWJmeFzovSzLuUCHf6zweuLRMbk8xArR/+vM74a+PmuB23VNwG/bSyK9E+Np
lXffqlKnBgaLmQQtkoXgGciFTYh5sjc5tZXMWY0IgZ0BsXQEyaxQIesPvDVNXC++
1INlU/bnAYbyuet9ibGshpjU6d1pJTqB9C9EuSMCZfWwMI/M6oTeaiozpMoBM2Yj
8d6URRmmQrutwGivyoskkM4uX18Mj0U9rVG+WW1CtcK4BGaK9hMNbSo1ubjmruPI
Uhj8rdkWOzKIiLVZptgYlAGZMjZ8hfW5e3FWWfvBnTLBbcMjpCkEke7G7UoO5mgm
IUVD0Q/iVoR9vBhgD/Ie3VvImZOxrVvRSJ0OSq3n+ycH6lh6Gh5t7vzdldWFadKJ
p8MfEGb0mFAe8Hk7npQEJkLL7JuieLeg/egjGXP+wgR/D4xECxgkuWCa4Zjk3kRN
pwEH7jlgSf7Q1lumaUNRVKWjocKmYa68g1YfDGNvWGdGCMeB705EYxz1Eifc/+g1
2cOjLBMyiNUemXNQiEWttebsr7NNKIHm+vFbeRD4cHy8aWGmf0D6N2pMQyV9Heo7
U0W0E3v8vYFgmgwZnD20JaT/Qgla3tW3M/ajrZzd2J6wcwbiObzf5iqOV7Q6r5At
k/zLTMCU4zMSgQ/2c+0BAGvmW6+eoCv4QqOsM6MqQmUGuYBeS+rAwREGVUIKWM5k
4grSZcbrwnk1KwF7e2VGWmGEobVnyN0RpS38IzV586RjSh3GOMOu+piL2oSWGGMa
iTmHs+SMmowB+ctCClXTvGaWiSku44zKXud0nBSuPtBM9iem3m91Q/lgUfp3EYe9
5I5WfziKAhSdvSkztKZNRNw8hATTkiqRPxzOjRM/Q6BX9BZG/yhGH+ubNfiEz7JC
H/agEUFd3uyWhNK5ixEN8XBN5QkkTj4h7HmeByqOfozkxFAIGiCnjiz0Zq2pXXY+
6ZOhXbVjfsbpHA/olq3uCHTiCR2mLGq/F5ftVS/RLK3Au1kak01LsE0WWoXvEYOe
hQvsjcFQZR6ajQReJKa6BRgxU80ETVXIBLYmdUs6lGZrBPjwOZlmOQe2718GYMKV
YP6KW6VJT9xoXCJi/pWfilV0eHEA0NMO3S64vtGmsAgWPenWIsHzMCjLQdcl1ZHM
IfmWc10cnJmReqJnb2MZAHl84WR/aBrCEq5vgiYnLLgRjiQgmZrL/FYdkD1cV7pq
Y1rBnPTGUcE4FDsmbpQallYFslxWCSOlLs8LER9/8MOSBe+boV6LIDLH/zp/FzBk
t3o7TirmD0scq9zmgxONenurAeay2NKG9F+KdP39EGi3hI9jJAu28U1IHZTQHXFJ
LvvhW+yhHiIlu9bwoUioZIO1n6aLxKJlq5YVUYONWwxsXUH23+eJt58XzbNX9h12
UBV2+68Ika5gY2dmoFqPTbhVl1zxZNEsq/9JKX6l5cGEM21zp5uWAkTVomIKzab6
+pgi1JyFrkHNUnoVfeClzaPHa62nhnbFO4tUCr0SYRv5qhx6CXT0z9KxltKrzdRq
BEEjjK11bdpRt2g7wTGIsQlLzFcOs4Hh0QJlZ5v4hOZnKGedEqbrkexcKBnAtYQF
QgVAEju5A8qvcMob3r7WuNd7VFiaVIthtBtqZw7SACc2NtYPdDwufFoCTcXZNFmH
csmINeH6iSj2rQ4BxVKPONNDzzu8lajq9mlOimKmpOnnD2XGl6PIYSv8ttRMbEk9
2qNdW0yHLBeXT0iizSZIs1tTuGM4mM+qTzsbPM0CWc1tOBNz/bCEZ+6wLx0BWbuQ
hPgBaq9/DYGOdzV7kkzzCrkhaX40p9xgTtrAW0XjtgnSAHVnZjSKVOG7vo7tsb04
mLkG3SVowhjU8H/cngDBYJwW2kIaM2wkUIqZJUWT+nmkeTnKfGSFq2Oo/RX9tkCW
cc/t5aalaayIkbD6Z0d87m13LEvkkLWU2gKfjIJQFKVN72Do3EOhGyje9yKf6oOP
qpdwu2YLAz+oiBum/VILLCNuMasc52mybmN4XxTSIKQQ1cAFzLzYKKurEkjEwFe4
XfybtXQYGL0/HnS21xEq8RjXYybXdfBlke5iwTi1u5uveO6FYrRkkEyfPDCURev0
IFBkXjl0gXXeqeb3D/i0Pl1vupeWLT4i5lwuyOJoGlCN9jeJSE0f8oM/byqYz5xS
gFu4JhTwI0a0YeJocL2PNd8aED04Au5/7cDwmMIIPSQghfP1rllXjgQJGA/Dojb0
Rt0B3hs46Lzi+MivaCv0CQ48gyDeFgZ5+Gg27TNdQNE1b3l4lm4bmCX+dudEuz8q
I0DUzCZSgPMOFYVismNpNU5QlsMx/xOOvp9Y6UlzysSRPhg2S3Qe/KQa5RPSK9jC
sjzK7Vd3wOq8MC8cF+EJW/2dm30+g+3l9BjsgTNJaDMeUq7ISdyJz5eFGaIQEKkA
RkOznMGl0NJ4yEf8JgP4MIqpF86rxqiV+/L+SKLUWZd52GIzu/yWzBfYRcrv9tU0
/pjWJF54jP8GuuEE8z4hHXBuy02O3x5nl2x+AlgWXK07N4CfCB6v55D52tlm9uwL
HGAhtqcCdDQkDupy/5QlRRFF4JEd8K8fnXykZtFn5a8jF1Liim7ozJP/bPE71QyA
VUA7gBLzCBJfCCl+oPqn1jhHDPU0eXBkwUV8zHzcBrzpi0MljUA8XqCSRKAUlTgI
soi8K3a4E7Zv+P57/AyrY/SNYM9TX/6Yq3/f+GoGXByqSYgoqrNQAbbFJF0sM+4a
C8Ker17eCkn9nYVA5kL7kE9NsIk1G9qYw/75cBypoJ8jTbxLJzlcbzUA2qyDrJDB
tp4jM0QlgaDVm230VIg1S+DfX5GOZW4ahwTerUodCK+MbPzGAHkgIligZS0DFa+N
szjX6OWjmGiW4p/srhq6WVRNDA/VlfVpNkFo8uFMfQm8RBuYn4xQJp3aFCrwWV/e
RfqE20lngdTslOVwgWz8GDjiFs8dNCHE5grWTywOeE5n6oVik/v4GSuqDNVghsPK
wclhiQHzxCWWai3q9b2s7wK23VahrGVhqIbHpH8jkeO1p3TLQsLai/Iir9ExldMA
Bpg7eSPC3zse4iPyOoZc0nhAGiFFKDCkCuwTjpXWmexlUVaUCNd+S5+V9/5Svo+2
1AZ32T/Db57Q4LM0sejLOHCxACFGE2jo6HlfdPrgjtmx1vmmathbKhCUTKKHo690
O2VuC9uB1zGaxQXn19UvU25gBCwDFqp6NzPlmebgWLBia4tLvOShiI4qzRvbGBzx
NwLkRmev72l8YB09rLveaeFnIhiLX8Msccn24xwfJzz/29qyD6VPgYIY2MqkwBkI
sJZ9i+hqwwICtRClkMhLYSxTGNnqSDifliXlIm6IROp9IRjsD2xTyjMa6Ql5t7JB
6oR2+5m44TjWeury/jyd8XgDE0bA0iA3x7o+j3J44xTgRTlkPdTDID3xmYvTdP3H
21Y8294SL9sQM3K3UoZKt//V5febVrWUCHr0ioPN85ys8+EQ1vefKQ3+kp20pVNd
X+McXuyXNvVzp2blMJplSDy5deA17eurCQ7OJ7Wm2N3yirYz90jPdmlTR8N0VlMP
bV/rTWq9XFfZQ80lYDYyKoJo8qCB9Zaa3oLjSgAaWe+FjD3spWRb57u09/oLhZOe
4puSqs6uaWgG3vlcDbOrfyWdI0D96M9GDfrs4u4mPmjxnDoJCmOnCxmOE4bAXWHz
pBgV4c2lqvbekvG1dkM/6ewLOgcsZUbfEJdChL0Nl0ob+U2mWClv64MeR0kZhYK+
+RZqD1QaHgxoPSwIo4IOWb3AixDezIxjXZYGqXkMp7XvqUHKjPq7BgQLgauEw97u
OJMki9CSVv3qAGIHAR2KrcSYQWmUjnafH6PbO6NY5zr/QCk+vx/uGMSkh4wDEBND
DYAanvMsu7UWjt+VDjUQkZaUmNHwHzjvGclJ+v/9GA7yMVFUr/KY8v2+N4rZG84/
U1IcaUAYYJm0Mr4oa61xCOaPfTdfH7rLcPmJRuc3PflR4QZk1hh8I7XSKjVTWLi0
vUGSeRuywExuxpXs3wX3wlzxvws8HBHID+mCOc2kjFtVnB+z/sWIbWWHQHXSpHGm
TbNX3eseXX0k9Bzsf2Q/MZI3dxF6iRjSUK6AG7OMQ5MMx+VBrIbSKk+g7bb0UBUe
HntBoS3eK0rvZGgim64vIM5cUdKu5bU5SUemQ8LQgbRSolujNm0DqcZrTY8SdMTO
aTaPCqqcnRd8pKO/zAcI/GOYWSXag4OPWIOEwpcOIiqByEqSS4EI/xasAKHNh/7U
joB8OiKhwpvbiiuo0WvPPvIn7/t5eDm7yI0gLUs+gTeeHtB9KV3fHHQ9ZWwSI2nV
k7TNxw4sB5oil7c4EfD3BGmP6iKDnZM2g3F29OHvA5/HAo/tXwwU2kKCgJrvzlbn
PsryGBk8peP2dTg2qFvzHOCt6d5j/rodughUayKDUxOtBn1XW+8AsoNAzqXYOhSn
LKz6mBTda7gEKNEEIZ64vD7VYlAEyHy9hfmki2W3g59YTjKnRbzCWsGldsOrbEpW
GuvBxXxCjgKj41P/lcYnKePO31T/a9cZ1KGXNx0YbIXL0eNSwyArqONMc7mt5Z4V
tu+ny3hcHAc8UmIYZs/SAoAfyTzR820EdYti2q6n15ONrkTNCOijj8nyqYPX/CEG
BZUjWVAPX3T251pQYQkdP8VMnCsdF96Zwn/47EIpfSjSv4fOdyqBBbNCRjP+5gg9
lI3/mBG9PF+SY+wxW5b1O+q1IIO93DM62dJCnEtPToJpivl5Rr9p5aTvtP50R4ki
EVIdMwC8u2Ry6MKlz8+k9Oa/GVQbU7WMa2hj4JRkBeQeI2BGc7Hs1LCfw0h0zakz
QSyNQ/oaJkTKnWpMW68glECtKVqIvqYDLmwsKFA3coJnzTWS3eGhvpZJX0R098FU
jDB5oCD+jZKYGJCPwDSJX/RUdWbr21KHuAut5Q7LiUj57kUH9m4Ib7GyL4ZK8Gh7
xg56ywD/GNsA7dBzVHwHekAFnzpXGoVTQyYKteCevXPvUJCjMzLnm6Es1L8uSVEK
r9iNHktb6OpxHHn7K/59zjPXdsVKrFveZvSqCF/xyUnXW1z83A3tI6xgr6vqwSNu
n667OV9Sf5ba5XKr7CXtB0CztlT5OS8xrsAHP+ldNXAJX+mFpu4CnBe4WTeqa1bP
syau75nuqrKcs8L0iTJlDjFLs2dYwER+/dxCcn0gtdukG6AW3Dv0T4m45l1nfVX+
MUj2ay3GEspcMJ5FL1uNrICKLRshHA+Tls9+cvF7DB2VobFcry0YekcwwNn6gGRQ
vQfFD1vmlT482QHeg9Ljmso/V3mMwR7TbfC8rk9vTRmmzfdn74WD2G0KNNBS3Lxg
BSfnLx8MYX5XxJskyIzIgL5ll1OagEzjCwLUvzoVlKQH341HaUYf74LxqEgjRc7j
cEsDHlmHdZzULk32WILVx0hrDz9O3EdEJGVqT4nBl7TD7PxA5hoJ1l9WN+2DbYbJ
Gp1l1xFZabg1pLZU53y/sO0iTYFpYt4mexaI/ySa2uto8glfU1G96ZY0PJHXoyKw
frtMIK5BD/rS50zIB/spPUILSrEdovULjTBIvayicEVbtF4SqKJTFroVlGNAAh9n
CZcm4jL2KVwitKeSZ/yv//OGmq4cs/+0DJChxtT3/bIFgbj6WpIrLIBtw/OepJhY
eR+g/b0sLnNSXDs3Iw4trLz1xdtzt5jloHOkPAoDB/glchZcoLdoFvEDo81yhiQv
SQshfjWVFyTKcViTdaj3ldVjpS1jcRKmqceErGmpQxyNgAQZCwRnrGy5DBXNLCoR
lnRx0grHDXpDYdnLRnOBN46a9gkwJZ8jWKU6kMhh4QVCNpCbSYz7vExmvFsNNYPy
6MwdbEecUKwA5kbmKGvEnodPPXUBsaWUtDarU3fdSfwVY2S1L0IWVjNsm5FanBrm
qfbZ11rLddzUyBpdyEaoxFudb66HzNcrpBCBYDhmXzMkM1/vBfU895Ek0bZqte5K
BNX/Q50gNPkIz6qpRVFsNp9iPrVF4uwagZqxdIvxDxEGpejwQ0VJkIJaqRn5sWJ8
uQGlGrb9p/6c45cyyMPRBh6IkJbBGfowpUazKdRRL7idWN5u2f20nhZudqWI1Zhe
WFaIP2lc4TF8gRMhGK2BxmgjFxSRpLZ5Kb7PEQRpFyGBReJNOrPY5gsZKeeGU88I
owhREOsd6yYF9N3PrvneblorWzwOfwqIDOMti7pdGaPVEg9uGKwc8fnAbQJFDCjl
riNlw7DQo104+3GITXjwSk6spDP/p4fwN9o6vSuaUBcRLAf/IL2alUqrXFYyhPGY
qc4jo4yJnUTJmPoM0hSyO6pLJ8X+JqB7IdmKcAMtux4i4A9VrtaD8Q6nnPfX8DKb
0Hx2nNi5Rx4V+3BXsraC//OKhYFsyCgKu4w4A+aPwih+sy87AY1dptmKlEyMiRKg
zvoKaGrsQL4nAHrPif3GWiMbE6ddJwt5zoYPj+Jm3uQjUZS8kV66kGG2rtHNjhNe
KlHcCk8eBi/XzEm1CJiSHgiCM1rSTBtfTsvf8UpkiYOhOxEuB5NSJFjCD4LJTUwd
xIYg8STU1Cfw1DQV3m3CLCYBrkf6ND7ooTyv8O5bZAJ4VmTp8HdlPFIXDWwdeOaE
JhFp5eygjPS2sOGYbqR8pXxi0bQZWYtoqCptYW0i6tx05DFOgLK0UoikyhtKzXrl
6Ukk0hvoMMf1XRvi9vEGX6Sy7mOGH8KEaVz8kQIq9ixpOUES90gqa6syn1Em/mAt
Se0Ywa1wVsEK5on3cQGXTH8PlLiFJW1Nwg8lsUYyD2c3VLv9CHKmc7mbrHM7EetA
vgC6PtoZgvpy0z3nySHQ4e1jZ9LbxvbzQj/PmkAyA/NaA/paxwOX7RDDl2mzl3zr
59aTi2zpFY+BZqzcE6NU0HcmBFv0vmLAVGdqyRc/N5uUr4KS1dKYI2ZMjvI7OBQe
GXcmUQ4gtmoCI3mD2wonC0yertznJOgpo4aD0l1MCN2HZ93TNdkYHjhixNsBgA53
D3/x+XmXcPFUmppaNdxRiEvE78sNqqwF8AB8Ir/SmqiYnh2VKo+iz6U5kTo/QZvG
qMLwMnfEe/WqE4WeYFeCOan9KrrgJaa+XuG1rH4KZ3qFb+PlSDD9OzYFJDXjEc5P
bYQRLzuoLrfzIGC45xElZfHlTuDJH6DaECjAtv3I/VP8cP41VUj2daDDG8QAWIJ9
JmYggPk8EMDxVsKF9NZIaM5adoCMRz9xj29dt8Pr9OrdafIAIvVjmRDH4DxMsmjv
KoaWLVGRHFVlqFaJhQ1iiPWdowgL6fkpsvmIzEbN9jMr1xfgDVGKO6+qwEvDZdBu
gwlu7g5A8fbk5KwWf5e1M923TGl0yLqw3BTxbRp2EICLl76WbLx0bYLZ9aA4EBiL
bZz/uI95AyGD8VRz+hZRI9J6eNPOCRPHBHEVrXpT7naKX0w2WzMPuTO95kmcgUCL
VAFH1IhF9kRxcoibP3d6x1YpGEzIScKSUE+DeROxjofJeSS73ooQ4UV4lSCB8tJc
W+a+2xiDHZo7p6BidSGelmheJxKqK2M5XojnnONCWO97kx31e2qF6A5ekd6FWkBX
OWLCYGvY4oHEzRSXs3X9hStWhFbhByHGx37tVCHLFVlaBhjJ7xdPYNL72uPZ/gcr
GAh4xt7kpxZcPfaBG1iTY0lUjrD8limaZzKz1/Y0DtcVBtb/4v7eOxs9UQwvO6lt
LX9OwpnbEX1Nlel0xqNchZi0pAEaU9IH/uyz/0NYUBYaMpH7bsuA9yuirgF0VLB0
CkXDhnPferUWpZ9uRw9edcSTMtRhNHkaqWh9kH0D9k8BhoUxeaUdUbZ/D2DjsWUP
I4obXGToo03dZZtjIQ0EIxzrhOb2cSRRa0OaLDoYLGDQTK+gwzghzhjdqDN6yhIz
M9Sc/zBZP4nky6+EPTrqIT36I8nbjJvyaRpa/KehSi23abNVgW20t3vwQx7wPJHw
DDEDVL4F45mTJ1au2zXFuuXyOsVyvuU+GMzIkrB1JHg63cg2BpHZHaObd9sKdivC
hanGF3z2ovlhg2wfxv/LWNlam1I354k73OdaGwOywgw41Nrob/5OQcHU61tqrAZN
oGI8Y+ucAS5pMFhyyx3pMOyh7V97DxVCHmDB4Uas8V9htzwkCKAHv8MJtw/yiTF7
5ozR802SC+v7nGylnelcjnVwwUOpghvieoPyhxutpRs1GCdmBLR8iryFtlsC19pu
aappLLKhB2QV0JF9eUKH1xac9xsqLnRuFRZ4hTSZMmAnB9ZVTlXa0fduZqaxUJ6b
SQTRRQ+roohmM3KlxPynHm5mNXEtOyuumBasjXD+9z4GAoDJhJQJ3l+uscSPNN5w
2CXfmys9gszl/djbot0h8YFNUEmMT0vYLGGYuWAqa0uJ+KDdYurh6N9pnVfx0sQt
ISvwlx4Auma12Zccup12AmJFAwIu9ngXgAXx466whlIIztxV75wm43NF+yP7K6IG
aWhNCsrIU0Df/CWplXd+kZLgiU/DEwMgBeTCSSf05oi+O/IDUNNqWDJPzyHzVyGs
WEFyz+je4LAvPWryPWHnEpt5X3NYRMOEo/eJ9vVa4UsCEmz92mNZOjlu+RIWWS78
GMkM3EfH7fyVjZ3uuvEvwDkiGXXsgzkI5Et20nFSGMIcdFoy6L4N8ed46OrkkCFK
CMdx4z1CroWn8hS4Z03c/fjC+D9dEe8JDzm+sn0BUdYlvq36Y+knjLJFqoi2LqR2
v9E9ss64qqC4DIeGiL60snz8uNN+QDyeb5fCQMiC9+BG5rav2m8yKkwhwaUpCHQ9
e6uK2Sgzf4mqmiFN0K+9PsAVMTT1WuAqUDd2GXc9BeYB61w0HNzJQQ7uE6sg6rU6
kDm2YXQ/aTZMXSHCbb6BK9NhBy/t/ljmFgefeg15PrPHti9nFASsdM69JBOspT4W
BWwBt5eBB45yL93HJdQLmqDkdb3hFuylVKkG5nj5+zi+yoh5HbhRzxhJIY4fH2Sr
xxQjvCGUEAqbxyy/nvTPW/X6XULNNwOUstak2sQdg7hX3IqtQyOkq4JWXi6yplkw
xY3YDeUlxPX5wtAdXFXXBzEzUAfGam2eUWsTH1ayCWOnke/dzzc9449ScCB51N+d
lvES9jBUXtV3FiLgkM7UKCcmEYH1KsmeKRvRq7izuPoKqlZACNFJvMuhac7HjvTr
HevFoZkrPCNJXZg+zMc2rMqWtqrRDjqflkzfqyBqfCIKj4qF4CEtsIB+Ksyo4Hyy
tQ/Jd6QZ2gQgjtOLuVH0MS6vic9v4HRQjUp55RgknXctvqUoluBGJrzxaKpNewKJ
9QT2zqykmbl8bpF1kQ5x2yoZV2yjLiQHCr3XbI3MNk044XJrFlqEwntKGHlFH6Oz
CO+9ffUW67wwY6S9zd8ohl3z1FJf01huF6uFaCO3YUPVVcOYoL8JmjwIBlle2Dns
KDPGG11PmFLbxCBzcbueyB8hqZ3S56bHXqRmllFuiD/NsP1Npmtxn/T4kfs691P0
Jc7JJ2fbYRgEA3CMsLiHZ2OzXXepzyfM+Qy9IUfbk3tVlwBfl+ZaZsaH0WzQl+eR
84Wq5zI3hSMjY62avtYlk/AcVLp67UBt647gpRPw+fV90DB95U0FNANw0QUILqQ3
seHZfXadEUbeq4o+NUsXovHf7hS0xDYqM4fKNnBXpMkCjQs9HQR+ENgQluUGczIM
Vx9WFHVjY/zBBwA1Z57b0Jg5wJkfNEvMrgEuQMkFnq4Z98sUEC4GPP5qdWI3UJ/F
IS8sA9GSSqFViaDPEAJIOxFjosX8IFOf/+gszc2TanbEoFNt/oOJc0i6eTIX/ZVS
z8D7ztBU0MtOvGA53iGoZGsbPeRw3Xr3SAKcoUkDjVAPUCKskgxVKq8GQ631FPNu
5X8KbnmAw1I8GWVQue6Bmrdj/4DGdc3Jgj6xjkJiX8K3C8ldJz7bZMEeKuUGRohH
Z2ZOXt3fJi4ZHAVBM83JV6elZBpgVJmZu1SY8HBszt3wP7J/gmZFyz2i13NFlwF2
ST0QUVI3wByZy4lHLyi8bLtCKdlMFNe6SWdJhiAElf3lLoLIS4b0s10l2K/MWgif
IbiwZdLFqvbUYDh2GjEFNJow6Rzxelq0afwxKFvOW1/T+tOVyBSqBZLBjw6VDh1w
btDTQOrXZe/jUq8tOdaexu67ztnv5p/Yn38uKF3IhRqDl7o63wKUm7fvZaiGtmeW
n697BIHSio6ioFfBjdphV8ql7yEzow5nK+nD2+ydYu6oXfqO0FMCoFOc93rlfBhu
ENhmwGsSANTYt3YousAylV/0qARHZT0jyc5znREJZ8nO3weTWK6ofH/52tgjJ3TJ
EALgjvdDZRBLYRrTDy5JlFO1CZWyNIGGWy3jG4Tf9An/DUYeEr9ZPErF/2jwANNJ
h/WMe5lvWXxbAEwP6sVi3GD8er8uBFxyUKvOdx3IIBTZEXv9gYjPTvsPVXd2NuKz
Ybkt2UZBTRQmvIfAOf6S1qRWX1TLYb36AZdQeSvZvKGug/pmj+lDVhn37BZzJtg7
n004TwSzElmOcjGffYdIfWVRJjnzi7wjcellYHI1pkK0MydhNRpgc0CHYp8TacW8
3QA99U2S4v9UHR1hDZBIHsn6HOtZWu+cskHsE/wF0XE+w5TfJE1zM8sU49duj/kA
Ap4Vm+T5PEgRmRW7F4+DFXcuQjvqgUX3TlzrsSS7J9PUYnwWfFWV7Sq7eWyGflLB
qRY2nScWD12wLXylU8FhWE5MG8HqfhLl/Jp636gsA7QQO+NqL+MDNYhb1ZRtaRaY
+TrN2p4Rh0n0ACGkNb3pLBPkWB45A7perpTdT7lMywYjfohNgBZMEr97e14AJSHR
8hojzDkf3S6m6xSlF85ob/Nn5A1BDAPDYnDiYEvQWd9AnIZk32r0KHPeZnYNsDH/
R0r66/qwlnMDMJC/ehpxHj9doDW3GxvIhJKOeTi8InoDRIXJP8+UCRHa68t7icP/
aWNRcLLqw2i+MLc9lIPYr5LOsnRSDpSSQTV7joeGtbi07I5vC4hM2TKHLDM7cxoP
ri4Sk9SV6fGUq3oKHOi9rVx8vQw7GZCEjbEwo47ikW15g4PPeQlFMZit2lwJdO5g
Kcihm4Nin2vb9qg8ucYOQOSmazvF4nxy60OAYzgO2HkEc2L64xoydnDCr0aI+Em9
62tRTUF1SA0/dgVsLBu2S+X9s6NoY3HL3n0zLd+5/5SofM6skEJCUXp4t20UOZz4
8w8XcmpDAhcjLOmgbHqwDB31DkYGWzNNGbxEh0NoIP4kBTlHfUy90POfZlQfTT7+
GJRGZFg7V7oLD5hQj4fwRFFkopnQqMNWk538pOgyHjltQGxspb907w2QoHHZujdY
awLrCKBNDo5Hn+XWzpZt0QXBN7FAKmnuiEfbLuxBrQ4YzNE/8beiWgbs+Yzr3bPn
3V/uU12ob0WX0zXNgq0QZOL2haYLIBywk8wy6VfTNcln/VSUGYOoRhF7968ndP4x
5VErT4LUWaCTuSaX91HIe8O1WLi6aQIbL50DSlfq7kaxeOG8rVl/J7DOFRC/1miA
Eq41g27SfiDrU8lBlVcy0hiQ9rqoKricRSYpJqOd9bHEVI3AJLqov6bLkF6VwXs4
nZ0G+VjsgO+s0QUFXOrgBmmPXl4EnMkSl1O4TC6rV/z1wLNfS2BmWBDvOVa9YPGM
DfMFTnvKmRrDMcBvhqGyzFERvOJE6Ny37HR42TF1mrWXUDcoedVPEWTCFlufS6tr
NLKG2zZ+wCLh4E4cASIwsI79yx2XMjx9C10gc7ClCE6FNjZH6P4TF7ZnGRrIqRh+
IuMzIjx6DwkXmdAMU/sqbSM59FlhG2OiT7T1aHOj3SAIZlti8lrGNMo7zTxrqy9d
LlKUmg8k0839aFhLIk4ugPdna5cd46scr2LvMDzPVcdqh5fFy7WYbbyKehl2hRA0
z9vTzJ/oBmjKUvUTg3lZE1iyf522HUR8KeZFgg2epT6hu6o25H563ejJBor5unLD
NTt17O3DdpFCXcnCuz18bBZc/aHLK/nIgkCNT25bYoPfSt2wEMQq/A8VFOU1Dp5g
BJmkfzebodutq1/1Xma1We3lvgNJl7rZiS0X2p40HMGuXCx6Y4/Lyy5Jdmf++pki
Ata2JmpguEo3CDH3nHxdLTD+RBBkVOAKd74fafzg8Gg6fm3oJwS7WaKFSQupewa0
08dBB4wffp2baEDh5FSrvrI7FNdphVlmF0nNcF96KvtdHVjfdm25ZxSwQ/z88GUq
w9K03HaCWec246xwsKWgwCfdO8BqumKqBbI+gSCew4dNhfcWntTQiEbSNq0KaTO+
SOGRZr0oTCp/W2JTAg0LtjbWCa1y3FsxH6f3P+01mXRavdhDMZLByeX0UY7satPD
yHbiV+Cz/Zzxep3SJRaOhCNEPnOTlljHMkPnjonkl0vMWZzKq0wMLVJ/F5LrmXN+
eXhWfjxh8+YZGjUY3a+LcXjTb7NJDf9kPZmCd1TTJH0CzXhqjxlrDqcuvNY+BAvv
3lImYpLRjoeGBkuwtPQp7J/iM6BXhr4jjvmAqbqd3HBNaKL4uoDnTOBW+dRfLgF4
W7TwZ6Qt7BZ/QM8vJtnbObAesXF7lL2eJ3Jx96ISYOmt5310m0yzrVKHyDJzylYb
z1UrSp1ECVn16kvqi7Vdxe0SR41Tf1njbm6KkDc/feppY1P3NJlHUF+RjsQTXdVK
H8Rd1f9TZJt/nPXVo7fRxJ50k8353tmPDRdBXlD6Yjm3SnKh3def7zUSfALnQF6b
/2CzGS4dgkXFAZwX6TmXFUr8wHoCTdSANGg/2MTwlIY3p5TayQmoTiVh2ceRw/bZ
ut1X2K1+m9pb/ZsAwcWVskwgISAxPIzBx000siRWzzeKSjudC7piIY5TG9vhbwsy
Q4BWNvtOcwbnJHniB7Q7YUDRpf5h+GHyQG0WDGwCEMssw2N+Y0pSVKU9komlYQYa
5glidA0RyXriyMLKcJSJ5iHABNxSIyfTAm7NnoTIDkPVANOwtdLDb3qaPYVhnW4F
ycb+gkshgVYxIOpxIUJ93wlbjMgm+NUw75wL9Sz8mDS0bmqtN59UadkSc4cb0B9I
KGpL9LGhf2pabLmASTfqthzJgBXfxnyJdaS5MJWWpfSqPH+Q50+ka/KF5RQ25CAS
AajURmrhtYx5Z4Y20xF2Rpdxa7qQrzKIkLSvWB53Nm95c8z0UmUD+DhXkHFh6pgl
7b4uITOHrvm/RHxOkcBPb1PCxhKhy2YhNb49FGiJeyShQgJ/7EnOwqaKVsYFJshB
U3NW/K1+q38527awby7pBhAMYLeBp71FvQt+wYnpGwPNbUNS2OLtIMNyHlVHtRFY
r+37qhTzxOfEatLlFQIQ6kB3ZpVPhVdenrzbDSkZ0WAvnXelEFyZxQqZWAUhWAjS
2x54+FsJ+LyxD9tDJU3sFX5iLNVABaXRyWvnflnJhFI3Y6GhixnZ5SHnVkrI4SNk
sHpRDBMf2nwkJZjlPQxj+UNW4f8I80M2WbN1cgJzmaZZhK/VT8F5lScLiKo/tIJt
UMQSGBJJ4p7oe24l9Szrl/ffeZKm95LizLEeik5y1WtR3mnFl55bcPCt/8eJ1cU+
rXpeoUvJ6xEOydKjeRbIv28sfulrVJEJPiVN8wVUs8eWjamqFrncL1WB/ccCPZv3
xvNHS1YZl46AOUkZD2iBhy9uelv36ciZkBcIo63+/yNVVcMJ82bX4auX/ZfbS9vw
WIxxSrZ66LlmrZYCGVQGKGQoSqs59hZ92qK2wWvhW5g85v875K2fdffFTmQPWgU3
zm9oefvVT1+6z5kVTP5QofwifezTrdIoIREGJlIBIW8dWQp+spF2NZ/24jfYToZ7
r+xt0rV7I+eqBbB1YJFVd9r5owq+pQczuh4XLzmLsmpkIgdp0j0ShWCOtiMAXObz
YonjkOp8flr0VS0ZaTQ1IheTU3L3O2GScVJlSH9fcnRpbNtC5mb50vYd4OzN7bpz
kLxdx9Cik4ki79bKWKeEOvETSfjt8/r8WwAnU+SMJAVq0LhptIq0Q1T5qMbeTYMp
Mb+BG0LxhMNylZPV5Rj+j/J4rt3bakemak2wEW5zwHWqLH9ncoSud/Djfu8lpe89
ivhknhUa62tCBt6ZDXNPrkLvd2TAqjW2/iAbTT8CYtpjc0zMTgYSZJSKnGLV2Tm/
DCasm4U4oLSfC1hgJ7QWHIzWqT13D38qmdDdmd8UGnEivoUzsnz/VWbhnEGu4LH1
Dl2FQSLxObnObdkt5nVawA4hnS+PbG1uS6cbll1QkZ12at55odXkN9KxkOYj558p
vODiA6IWW3J6JoSP1Okd0OdQQJYSSi2oGP01lGCk4i2azQYRE2qTNgfs3NyVD7HU
1WMut1+uHyRMeQ0nIOuus9jOb8b4tu2X6MFrkKY0JxevzzkyHJ1at0Of55RvVVJ5
/BpP5WStaUfqKB/BDiXrwF2xsECiAwqYXcXaG8TXhRcbBOb03t3L94LZumg8Xwwt
VdNB9nNfuO9s9yNFUO8G88S+7+Ti6EntrJ3U0IXuHdhnAcwVmZAN5s8SvNug938P
FIxgilXLDibFZx8qJkrPdWs7Xj3XukYPejQJ5Vndhfx02Wmc57uS1j4PfsJ5i5y2
WJavfkxuXl/N7mTp4EhocykZqzOXjg1V5KDOp/nveBRaQIoEMp+zwrSZnk/UUYoz
q4R4q+/v5YulupEOwN70rcbd4je0MZKghsCHSgcHbNdexlHyljkIMBGcMBolxWo9
oETasUk/cXPGILJUw5pCxQHqots06xFxniXBHQ1HO5nrwGa2K0OusmxfWCQxIfRh
8svKlS9I6QpLCNrhAL2XVTO/7QUwYUO8vnVI+4TzGWhoncY8BC7UEHZIc2yb7q5H
lIOsmMfPhrMaWuilm/ppTNs64UmDjmTVBG37z/qtY7A0gZAr7QK36+u5OmnkRDB9
0V8xfqu/MYrAMW89efii2NFsjn1QYKbjubZiAPrXdInqDcF3ht12aecoYfi4IP4t
ftBuX4wnDkmHfeusPYqhqn2DqRDFworBIJNlHwb/5jBAUlJEhegQaeZ0Wfd2ej1V
e6PKWibjBLrt6PRZoYwX4OP7MDvy2AgTxuwMmIH+r5hjboXPhgLnsxWZPrLyS+zV
jjw1qgIz9SK8MEZ+uahSk4DRrG214yc21PzJDUGTckSgU+19kl/x93jun8ZYPoRJ
PgcjAUs5QeRLGDEAu2/5A9roO/5t6JSDC+Brp4auSAfCTW0pJtxdnzESN0RdzCNw
/YOX4i6EDpmz7loUGR8BctJj4knIYVhAwfZjsLrhkhSTOOtpzppT9x2ZC6jJsby9
NamaberM8ChAcdsYG6YXit/gk/GGg/rRXljsm63HI+mEBrK5l/SiAoU2dkqcMIGn
12nHtS1B4n0n1gZng0Z8UthzgWPkwdVnJserYNG6Eu3eBjkytQqmQQrgATYOiz2v
ngGxBBkWSgWfG9CUBv/qX0VHH72hKvc9wLQrAI4GYeZgqpNSe2iDaA/KoXQwSAHi
4rb3qeTFtaOddGod14H/kEemwweaJnWq9Vq4Qsb739gE0WxBl0P7o+Lrw4dfCtHs
tsBRSLA7f7q7c18UBnd9Ea0RWoiRNuKfN/W2ctHs/Z8/q1VqzHCYG5p2Q2P+PF+b
DymIl6QHzQFgwABzhf0kMmQbnCt75gJ+aLRzmRIgMoNZ37644rGOSmj3+72f+41V
UYxlA0824WPnZ3cFBJLHxuacOlOQSJkdipYcPeo5f0fW7wgtZ46eCEcyYZPpmHQt
J7UmizQZqmpOQ8CO97YBxJV2vWsNzdFZUeOuP6LMetV0ptn+6HvhkXcYgBdI18tJ
1U2yC5BRbuySMehEl0bY2QxmZRTrNyFvC1wNwB+FtQhJlu0n2DB3FvAHRo65K0Wn
CdYhCVDNLX7ZLzto5t46Z4vSFuklSiANzI5qoUi6hEpqTTESAOja6xUpKYVl+VCk
PHiOOWX7XzJDZ1+ofgJ5CFYGVGn50kNWvKzsvHpA3HDT2LUOg27N7p6XtWkZIgT7
Agzjy3ThfN0NG5bynwnO/nniHswch1IyFbQSEioJJGC0t9PeC9T09Neh7u797d2I
VG08AGuO079SkT8vykEvfbm/BlK6Y2MbZ+VKhN2pMzIt0bzl7SnuCJi+TtXnR6nm
uyr5gaLCFXTp2khAQjoy6cOJjjatVUcLQpffBSDwryBwTqRGe3y+WYQHMkCLsjZm
wcw6493RkFJlenaINzkx3MPkLqEWwq4XY9jYjDfMAVNX9jz7FaPaLFIGlV2j+o7h
8tB5kdscIgm8FkWfWIYcUIDImc/wAJ1voL32Pvuzlw91opzJwTBOyXgqHyAoLgGi
vxYm2nT4TQEVF03opJQyd5t8zr1LOiYoi5t4tTrVhfISYmEJvvv5w8x6ESt3xtMx
bwZomEQi20nUeTsYYJ9HMlBkRKeqa3EKRlpANlpzEjynKOlHGnGIGbELMdD3QRYD
VWEoLeuEVTaZb9tQmhZT3xZHGWtiRqLRLPkZwuCHRdBHQSkzFlM0gDmXinM1vCgn
myruEu5L1Ztpl2MUtAOKD5mI5ldnmWEwqKcYSWG/IGUlJqUmyZKOCEPWLQcSXJpe
d+3MPNH7YOW7XduklnYn+kcJKg8G9Mc/8Px5QQ8nPcTnFA2uO9VDVEHOvYBQHJE4
Pz7F7Yn/GP/QLJ/tHqZk+v6XTQFeUSf3ltUykfo5bRdNgIxUmQVAejZ6Wd68qREw
ptZ1GyBRZ5ro1nNrqubAxPJ7ERp/y5uVsvTqFdfpH6pdCBP5yTtdIYuPqGkKcO2Z
Lg9hwdB5wQQT2GyKXz0impNpEI5z3Xyh5UAxvnZ3X/eAjPLsZbEfFouIGWmbEOAN
eL30IuKmLDKbhhPw8BeeUuoAsDaZUB28gk8caXUBF2E5M2GNoCxbj9lnEa6AIdw0
9dxAPaotlC4dwEJGCjUUyJShluYmL87Vv4u8D7DQ8gulHMxRrV0TvICLH/SbEsm/
mx+4l/cFSbEtmw1xnCPt50Rj/RB/Af+G40OeEDARzfTwJrT/YwXczXEq/yELInZv
ipBv4grRVbAyOyYrXXO107sxMBZ5tifUYzkC546xCMvgeBpq3YTg+0Yi1sONQqy+
OCiwOphk12FYUEluHVI/vrZOAq8FoaK6R+IuQq8lEZLHKLqPB53uTspYTlMRlx6a
ra2J2RKqFQG3jYHYpkE+QR2F1z1FuovtWBGHEM66YKzIhO1YVhhRr9CPAkoY/gze
ExuO09cqOYXCpZaPGH2CXv54bgD9olHuBy0MpPG00xvvM8TqoZb34CARmGr4/Jhv
lqyc+JG3Eh2ajf6GS7/l+cAJ40hUZ3fVv1zcdS2H2drcQDPCGIoDePBltiXDFaqH
8bLKLT4f3ahZ9+Oq/fhLzSDjORQScAoNXJjt/b7okhw23e/8zMl/DMQoHXKQfbGM
Bo8mDfd7NaulBqUn+abrUsegJF5i+1oIEgpDa7zsnZJKwFfObIdfOzNON/FSltwB
acMOUQpMIKUQ7hpoBxA8mbuqlnyM5RKTvT0L8Hbyl5chWX1a4uFD2PdeP+DU1+4j
AUji5smgaldAg8l5RxXfoQOHTlyleTP5WFQS7UFFkp7NnfL7gvR/KgAkIvTbT99S
rVAMB5COqqfRKd5V2uq0QafV6D6qrN52J5bgx10hF0Td9/mk9U6ZTuIvJzVPowmW
DO4yFIoAWRVVpBxnke2BoBz2YN7UDtN5O/s/IFSdcjkLFveKgedI4bmYpcqfUjoT
84gI8ORnwCGFzYKcWPRyk19lBEQFjPIbM/OqSZqyJpo1LctjyLaNuWkLN+BTWrQy
EZDxqonwEcqTzDVkzHLPd/sKTwtnTN3Cd20RLEKwHObjna/ip8yuW+WPTGjVaMal
zHSuVxL/MxU6Drcyx5W1Ck4p+eoiPMgzOVR0260qqbv86k6T+FoHACbIljf3ox/O
DDIDv8Gl6QDLlmyozereQEnficC10xBdu2hWdig81ZGfH4eaQsCkMJLztog6A6tm
gUW+fGhoNL/5ngdQFwWyTYx4/ypL0g5wwSv9lDYr1Nl400wsJNKc1b52wNzHzyB9
TiPRLqrzjuC0DG38sxu4dr28FEUJzDGZWFlo5Ya8HtjGQVu4S6RLjhRUzFkiJd1C
r5lCrOoIm+iCB1KR/Q4GxTG8L+8VY3qLVVsvgj7ddU3KirlGaK8RuCqLWAd4MEjF
GeYwZClupa/1K+zKI6R+L1UUToiLG3VuBD8ne4dorVJ4jvFvVmJ5pDg0WLRVazPN
OpohfoH+PhCeKKPZ6lwn2E3nuqNwIqIO1IfZjZD56ZBGSBIeJ1P5Z3sLCMDNWiGk
gkpxzc2i8009GL5x4e1xn+GfWVDheCZAS5F57yulxoJSk+gxAGtH57le+BSVvepL
4vlToI5KN1RoYFxucMG93A0VwnYh05PlftseGfGAPdyI3gplaxleCSVtryOD2iv4
RH+1F3JWKFiqmfXiecjKKa7G+GEOsP/NaHGuu4y9Na6AwGmyU8g0/rgHvgSWSKjk
ytSRhAJAIvXJD9vsLAKtfByacPnlUMnRgmbeROVl6SDmVpL7w+ZZhaTU71EN1QNh
OA63Os1Cc12D1H5C8JCx4QCYfiz05+frqyFn8gvQsDfx6yhICNOoGMyb6Um8PJCT
UPRZ6US4wLNmlHyRA+yLyJUHZo9eXXM9UQCmPYNNjF3ZGwd/Da37zg7ITKw4RTgF
QWS6aX7b/ROGhgNHLfqzPKkICew74Ebt4GMc88BNyq7MOoGc6UVH9mCOAzPLu34k
1kg3YT0tT0gCOxdzSxwI7cDdamjtwaCvsUzQOcQM9W8TB7J/zYKv0wKjw1FScnAQ
D//3suW3jy5qv0F/UP4G7mA6E7pFyASXPpekFvc7zlMDPYhZvAY3SgG6iLGSSOfq
xKtRIYThLZ+40ACgFsbg7bWrGa4LD4mCwosJ8cLNBY2UJOYdUq8NuHXdeqN1AWbL
vS6AMFTUbKn79PSB/HNxrbYRb/p3vADElQtnAqBEg3Fxh5rsh0yi/YL1yqhuNjjQ
zHeOIgfXCCVSMDK6PIal5vFcUd+OszhTQ0CZ6LTzRkjZhE3IYbMJfqsF7o/GC32J
439eqttwilfEd3X9QPrmrpZROBeBUcAMLk7M0x8wJzBQloseZWlOabcxAVrDij7u
4wnuQNJIhaW6EC8G2t+gAM6u8y4UFYVAxkZcmz/YsOw89wZI9fz+K0Zh8VgjQYQN
PH7aj2TRQet01SqEli5aR21/gwua1kjjcGHJYNEyHZj0tIq4bP6NMhCVTlR7Wxk9
hzlJd9/U68B4NCScddpSBUjx+/0pYfxqt39C2wCCdpm5CTv707YJvk4m5T1rubMt
53+QOgt4zJ0OQR0NmBYzCrb9opAjluTsJ0edm9bN3MvTo93ABN9fBYogDv+HakXB
1+PVrgpEsBxdSP5yNqYOvuVqmYmNk9oTEgczMcdNrElUplqr43tUFbLzrOei+Z1Q
YDhbSzwFaB7IzhBtw2FkoKkn1z/28HiQkOfAHuGXE9GfZZ78s+wKwLbXf9vliHF0
hfsL8orh+ZmIS8G5Fttvdk364OyVKCG6cElemdV1RizL71GjGJ2mmtVZ3VUqR8ik
RA8lwZiIpW3opUB2eQT0dkIUIoyz+iFBPK/qbl1iyOk7vT3Jw5YWdz5RerzEF+o6
DxB3QzjAAsyszKUJSQh8mpZk1j1feyxwE/1LPNqUE6LPqZQPrYpQyEqrb7ESJSS+
Pn5f3OjfWNNi4plZjbk2PfmIHqW/6CNYUXZ+0KypFTGKFYRi+TIL3dDwYavQmSFA
DALpClbnJ1/mJYOQ3XWm/5yVhpquImP6cqNm82FT4ChbzTZ+jtk3RZ4QOyf4iKW9
tjIgSS60QaYNeXz/uim+y0iLzkW9LjExtUQ0jr8ub0LYJMPKR/lDJX9gswNeT5+Y
D3pETUFtlbGPkbirxznjoK3WNPPNZQMPwVBwym44SPHSQ3Z3fSdpFfRvy5X2eu4y
Dlf93BJtOGEiJ/GXapiPOD/f21yrdP+cUTZjGSb7v37yA5XDyrd1U+tNlLn1jWn1
e2e6LmlMrsUzowThXUowXhVTfmNRaMkGP62FgO5NxC9mOpvAhngjj6VJP2h0Aduw
dBrRAGE2EWUcdTMZUVm5Iuipg6f4uXMd1VyEPX9RT1aMgX0Czy5fwIT6wvPgWdnI
N7NT0MO4mHaB53wpIluG/iBuCjqxIwRP4cimI5qYdWStOmz7KAsdgNITW+lcvlRL
D/FlmGaXi5SQrbnG5dX1aNhUZQK0mVbZzaXjt22YTEwYQLjKElTMCPhjDPV3kzL7
3i/kh/zwICzBVoyfyVCPTV8OdkBIPjPScIYJ5Cztej0yTmMXvSnrh3cBHhHQXh/I
cOuKh9Lah4L33KCsw4iXV6Z3GxXPoed3wfHst51fcKIhGJjsO9zIaeaGfhM1Ssgi
Zh7diCLn24UvYr2EbErYDf1JqXCkOrp3MFi8r9o8zE6tdfsz42Riq9ZzYTCRDvu1
lfP4vdGgYAaEIiNdfC4vGCeglg+5DZ9X4zq1rArRgwXoTv0kpKTpnnhK+TDI+/ud
dLM2tb1Wyvcquf7vMYE8gxzbln5EMSkN7P7FHJsmq7PcYTDiXLyiPFMT3Bba66/z
ja+cPjw8eseIiVFBRkdS9TAWv4NEvj80ifoMg+O012KVfvKZOLLkfvPh1rCQKZS2
6ThNkFsL0WWdGu+dDgRaQ1lkzZaVGRaJca0IIBLwI8m/AvUJSD9h4NUeThyqo1Z0
ZqXfgDK4I3K8/wf8dOIp8EfaSAesJRAu/cKGmjRlRynDVX4ezDMq8THvDnxRJYG8
U9z/DWJBg68o/dwLDB4RXOf81rGuNxQyxVxZgMght2S7YoqIVeAdx8C4cNXEx6Xb
hurVpVxgmlvN4oR6radg6D+8YdBZhxxTYaXCqE6QVSjNaCk7X/OHTtT+Y+c44plP
WKFrienHH7T+zVbysN6ByYctuG0UxysmNL13fq8/J5EV2qWT2cnXVyMjLm9kX15A
6mSta5d9LI9gZqe3SQQkWSfDLFA2mdHbM0wxJENn2101/TB+82ruSfqrqjuRfZKW
RuV1pn7jvY379JUICnK0xFunoFqy8Qw5wWKDGagTd639GP+il8anhGQhd2ZFq84D
BNHH9prtHqU9OnoiLGkN9VG7QcKCUhhyJE6goRPmgur2QMXNXRlHylfW72RjnJN6
WA54ELJUMrZEGey0gmLG3HGCEsrISWmsCy720XvlABftQ7q6rfVlPLNChWMbXf0W
09Tfljv+Vh1wIcLzeAA1CPTf7o7yTEPKpRtH3B1XWxK+Sthfn/GixCznPUfo0efg
+yimtNbvhEVpdC68XHybCoem1AzoaVNxlFgwHwQ1BOGTOQAO6kGA9M0D2MpC4OtY
L94He8BFMtZF2C9pnWfT2QYKjK5zYb8fBOg0QofdKcfs3SV5iS2Q5GUc8FzfxpFy
3xlpNE1oqlyVngHXGZQ916uaY54WqwsG1O8COonVkOBKygwy10eXJP4R/grpT4eX
t/XnFfhLmgeFSHVqVJFbbfh0eXcwCYmR9N5/5a5an922xbpfocjffkjOBdawEpVm
pmz5FQsCE/zflThQvaJPh+PrQYel2OET5FOrFQVXAsQ+MdhRFkjtQ5jRi+l+oy7v
j26uXk4Lcel4EjxcKnBdA40DKVPdfulb7/2flMgRNMKUSKfWmmpfSRBSXi+tZYbA
wfEkkXOSi/rIuk3jPubd1SVfUMJEt5is+HFkVTcOmYY3YnT5tBeUCLaz7IToLtmH
GrnXAXmbB9dMiIF2I7mD4VpGib0Fnl6T/Tk4ZRGujufZfH7PxJqDdqceBUURwB5E
JZMlmTGEDDIdW7Ld77NpUyk+lQL/IjQQgiOcKBb+1MLEDMnd9c75HYCAcWxm7IpS
S3DgpN6C8j1r1fqG2dR4c9OibY+Lc78lY0NFmKRI8JEn3mdGybZo2g7gbnQqynI+
rjJaYNd0QpXpNQGlK8bKRjAK202o4ScdknxLDqBndg7pr1I2rySaSMlB6V1+AYpC
AHt/R/iF4u2YltyYTxDEIC4f9qwNmSEcrRUJS1I1I3LNposkynIal7dN9sCdMXy8
D9myW4G3DJXtJaDxof2VokNHCNKRgsmfG4F81Ds+iXVnNzCipFbfXrK5T6qaFPrf
Vc2bR0ifVG8YPSgcomk3FfZgdamsJ8qnyR2W0Jcq1NeChFa0fM8LbVA3u17Mx2B/
B+TpLC9ZLXLVfqZUZ9IFpSW3UFk+eYRmEYr8EAVB549nWMi1E4DuqJGTeNPDvYDQ
sN9y34SKXeybTiGe1YS8Lyqb3D/n3HaCH1K1ZjzNeuuRr7C+HMmflJ7QTmQXcGhp
ciSkCaxZYpjwF0srtRAJDOi2y51F9oNueG+wVSA+5BZQpzOcTQHUnoCtPjXWrWYz
uoezcP2fZ3Urpmgxd3tdnLB5FZj7fTARby/o07/Igfr/L0oYq2HzHTyfF5LFknJf
yE+nsi8Dfso/ksjllMaBMjESZG6fSCaaHVsDHOKh3zqQvNMcL94NGBuX6B5Bpttz
ScEe/HKrYhdKMU1Pv7vfhIeZIPbHpuCAGX2aB+5815kxCnyyvYy9ywOmlEzj2aD7
ea12Wg6LhdI98pg4PyWFV98q5wAp1FD0a4A3ytQXJ4z5P1mNYiWE6ytPf9bXTgMG
kSfRCfaU7NkNHZ86JN5zIxOXlLZiH2AHsMtS1sXPtQ+qF1/Z12ytr8/dW22LzXnu
ppPREhbVXsayN7SvQMAwNtJA/aY3GidJPiP98iUUfynreyjNiRgpcCgVEHxaOK1g
NDAmxw7X1BAzzxpQUgUx6t8HOE6t0QEqytIXnhbDuJz4UBBQg1XoxGdupjDOlofZ
aHuLNTi6m3C4goXmY+Qo4A/dPZM16FxfOscOSrzhkoIBQk8uhuortvgytdSrl0eG
r3Ms4RaBA3ZJTlPl9slUpTmbwLKqo2Ql5n6PECCc6nXr7nPoIRmg3zWbpgFCDyCF
fO4M+cq52p+QG+cVgqeof4O1ueioPxtOxSLIyyt/6ESJUTszWSLdJ0kcB/j5A2DB
vKWKZfD8uenBJUEzVCKeif7WFmExAz1tLuoYHLqe4pFvk+bQNP/U47Y+k7Y21KF/
G0yD2jboDM8J2gwycDa0/OQtplbrGQY9fsp7k264WI+BVSw7CyxyS784o22jk7GZ
2cuae7V9dnl6rfkU3UFQQS6QObTMqL4uB6+rWBlGRPHyPUICPwrn8PQ67Fbtb7yo
tpL40hh4/GBrS77okNVHAlnYaPf5ldm1wep+8BD1aULqyG2ov6kO2CObcjuLELD3
u89EEOLjVI4TBukvdSoQKCmrETE2uVZbgcw0ZZqIv0Z6rjdqpWcSmjgVPm9XQxw0
cVZrZGGkktesdYLNUYnWeq+xcyummNWqEj8lCwCjSxOj+ssQs2PQ5MP9w17LzE3k
nlOgEHJAMAO4xDh+/t0foYuqu80XkcnBJqL2A/XngiCCEOAQiJrtjqI13wGCmuz/
Hzlh4nrva90POfmKJZJZjTApXfoY8rQPKythCt5prDSvqlp/RtfuQaqMHNDSlMAQ
235Bec/Vxa0fDOvhLQ23+n0BTS/+iFUzpl+lYkfcNZBoj5fA5EN38BipPhpu2XOT
vHcCWSVaSd/8Ooo7lhdhiSvJ8JShD3txgca6ABYVJiEnQR/SK0COAy57Wny8JNZS
g34umb7Gw32Mme7LfnTUQEpLfnmE5W6G5CLDGAg3pQt6TACtJeXN0f2RF2Q5mpCd
2zjPvR+5oBwPFnebBrhP+3iGeWTWHOvU5o5T68FWYYxqxmMXRHSEItqYpFr0YBcN
bnkSRjnWvwzQoI4ycA7sribW1BZqm2zDXfr8LBl2INLMu4bo2rlNtfYrTcZEZq+k
uQR4v8ipiH0pX0WwKu0/s1Wd1eOM3ittlyR++mRC+pvYe3f7roROyViJRHAD93g7
vYYQwuoQKuq7QzNW7vjtaGdkDsY3EyaAJ3WXfSMZlHaqrijxZ4g5hl0pSJK1uZEi
dTtGhJ76uyvcs1dM1eSTv6rUBBuGdCa5Bwf6u6eNletytb9nLtnVI5vLWMET+UcP
pz4xXfqaq4HuIsgus3F5pGmRlsbJgWWSIjnueJbeUjoOU7XRPE5Bzeet2QM4mGZX
VbaJlZ3FQJnFOvVyzFJwV6TSIe7KNmHsn4+UiVek/dJ5PHsd9lUERmJFTqt2i/Ic
xtH6Re9yYlT97lHorwDp6VcBr0q9F9tDrv/XqICO++tJ+dZHTqUm+BvM/Mrsk98i
zx8dk21Wjzxcf51MfI3Y1lDXyqaWnMn5Zv1eG56v42LArK+2CBemMbV/2SO8eLMz
eCVcq5z/7N7Tvo96qQHUHC114Bp/Vt/lft6cjCkCA7FD4rOVO6jDeOOU6MN8DVq8
wu92MDIWFrQY+CLT5jzGzf/fHwrn4WuegrWySDRxrbnDifTy8gBvrxFcNjSL4/EC
x8v8OZqelJqAn3xBMTTyQlcRaR0PJIL98OBQ6i86IUCWfjkNEvCa2AysmdJf2LZF
Z8CHeidpd2EfxWNTDrlalZnIuHNjf4jbX9yy9Q6FLohsZ3OtH2EZ+Yiya9a/GOGc
wsgKeXGnQA4vQEaxKwIQejzQBAZOY60lqYo7JODXAC7F1/hHxena2uL2rwJSVmsq
DlBwxPO/FdxAUtyXSUX9zfBgMsLax8i5+OFqpjvWReLfHmywF05XMXuNNPjmoeYv
NHN6y+UX5VETrfqXSGLpxF1Q1zLvCiNsawnXnapiRVGT4E1qIG+NpzLO7I9t/Pgu
VKTn6JWDFQdR0U3EQVl3zcJq8DL5z7X4UVUEC6k2OXpbHiIm9LlxHL+UczTHSRJ2
l7WlsphHwcTPoBnCGHzIQuw7ITXHSiBCWpc5vVdHqlnbDv4F/S09ul6wCKFGKXcs
gNVtnP8X5QQYXGVXx72P5RK8FjxFAHF5nasB5VaHfbPOThZu0RdTCXplt4U8ZzqL
ADDhFMDHOe37P0j+VkXgwZc+CYQ0VtRLmX1mjcZFG45Vu7FSdNCOnQYNR3/ff4WR
EH91X1zgxWB76cIoW7CNcKCBvVa7gMnZDA6ey3GcfFLrvFa7K5hJqGUyWEB8hdNZ
N3NsRnYspXxgII2BwruXPhkx5pbb1nMZ6FakBnNLQs9gebJ+AlQLmwDTBKYPUIfk
oobUoakJmorHh/TA7cTwSwblkMPA9Rxl6PnauAie8wRHsCziqv5uQEjZ6KXRVe3W
Md3cjtTbd7u267WBPArujHUicgND5VwuUsi3Np2mmuZM95uGGsCou12V0WL69TX2
mSLC1lN07hYcC4yTTBurWDZsT+98N/n8vDPBXmh3oggIndQzADBuWR97Biw3sqp9
iwCNTHYXxcG4PZ3mVYhdEwajHBxEvyTfBGkqEELKzdcYU+AvbHLw5sJvvrMLI5Xs
sKcYzy0azghHsjZN+P+peFG9Wp07r37PkGxriHwwaQMPkPV/V4hK8qwXLZv0gGck
axchKees5qE6EPGVlOL06jrZh1izwQxtRGEMNIS5Yln7J5kjZkCUcuJv95FGud8Z
+L1uwRYRT6tWREUDykl45pz4FnzbSWhNtW8xl3R/ImliazE6z7dzVmA3cXKKWzRj
YYE4KGLxi++OUWg07wUUaCuVry03Z5914o/1W/9NfElbNTvFVjhyCP8rZcxkAtJ3
uclCNn78baMgmcEZQ3My0W3OnEuIR+1o6XkwXK2ChMiN2t63dbqIO/6J/CsK+536
2NwfycML5j2a1hp/M/7RXuPHsDkdLK2zHrgVfYFM/Wck1DFAWqQ9RrZFsaaKaqcL
/8bvDMWyNLw8m/LXKD9GgYXzULs7u3KmqjbK9jrKdevSTct89Dm8xtjyaRwpnomR
Dj23WjchnXpMjnmGf+MKG92c5p+2V24XbydGvJml3IhB4obOezU3+fY3Lo8MPgoJ
Vqlkw8Mrs6y9nqp+Qh+/cXJB7BGau2CWszIS8wwyLlgOwlJNoL93dRvLzQKiujN6
YpBYzeYB6M+/duG/5avLanB1XVNhgTaczbWwdjyIgp9SMEkIXXXoAplxtzPCSwej
IkwbsvLGg31NgDu45zROCU7nnSwVyLPWAblnHNze0UN1TFmxUDHAQsxTX6CVytAP
7U6fXeK45XprY4Bltqxv7845Gc2kZ2roASZhtx6mo9D/oE54kicDZqfpcVtJ+OPH
upqNCmBYm4d6cCcmq32x3ywbLcSOO1FSOTQvPtHXJVFKvIuIGXC9AvdO6n+sQdOM
/BOM3gI10kJHOEQqkwR01CeUDE77zLPgAvusXzLKcEXrQBoWPSrww0oFsYtsm3Pk
lj3SbImuDfQNr8pUWx5djfxU14LsCUWDG3hKTpzKZDNQ8on/XGAXd7gluRb6W5dd
2Vt0lKLgOiOv4TpmjnuHahAlmn3CMy1m4xH1hKrN3R6VVw9LrfzIMyjNtWmpVDac
k+QV0WWXRnCj3GbddVh9BYCWNYzquqjOlahMaAaqOgkDM0DQ+JVkBHi7TUFpwj7P
amcAi8j1rE5NLeRlKsqjAo7DC503yV6m1ZcM+V2s4g5h0DgopqZBvR85RSg+i+iB
IHpZPl6zpyrskoOifBAxt8MKz0x2GvV1kaLR51Xi6ISrUfglw67jWq/2WmD8gK2z
ieN7Id5kFU57s4mJq67S4f8ioisNY3KgbT/bJt+tLe59tPMoI7FhPkNBDGOD8xz5
rOujYn/92OFkV+shIOH4RRUThjzOQFFaosKohTSRs3t4D/mxrJn+JCc4Vp1YMU9h
L0UoKW+SqVWqrn8AUPGMHbr+EqnPqud9lGHaxaQB0laGXlNNPCWEffgX+LWMO10U
ffx7dOm7LjvVLZlHbzVJSWsC1xFolAk8hpVYn5C5L47KYPwfRFVJ0VDOZTEnNEDL
rYtUvkBhm0CmPESXz9RwwbAX8tJg2EME5P/WgWBxuLxTxvMyjPpW4Qihyw7NZSGj
W0xWXBewi91iJVr9khEiTqoQ0QXJc4PokkRQJjSy6kZh0mVunxZ5qtQCicKIhzrb
fy2d+lY9X3CYX3NAS65ht3F546BgYx+LKVR/BY/69e6duvvFh3SQ3VwLUyp0T8uW
8TwELsoJpTHMOPardnZP5TomgGCVjAuUxPc8IIcK5t1WzgyjZSp5Qux/Z/kNb529
OK/QvmErwFYbJNB0h712AYlbZbLAZ1Ir/E9chp7GnC1UM3e43Mrr4dE5ohj9Tp6Q
xlTqRLsJE2Hx2OOH9GJQ/7lU83+Z8bdMlZMy8n7qxkAGBnAtYF/iT7ZBkYXguXGV
O3U6nFEoCj3lz9qfm/KaqgsGQ1rrBT2XbNKam/XYzsWcSO6C9iUbqWV+QxA3Sd4Y
czlL9G2jF0Rrpkd79UPJ5NkfUNngIlFAI6Vr6RcsNykUAylVDvEgb8bPyjd0dRGr
+lj3dqWoh//TDJAnN+sp4YoDWhIHpL5GyY5Jz0NSkfxirNLc9rFfisL7z+lwu2F+
pU6P3N2hanwgrZ7U7T8onMxJpr0DEnj5mL7JRJMsnFzkqmSMMGgkBFp/vsPJBd46
SSfKpNb1w2uKcZh3nxlE7dnjEVV4vbf6BloL8vkgbYJVsyPAJSqID0HrA4kzwRDz
5xhP36vuL5Rs9G7oZx3ePFr9njaPRvZIunK1qKc+afZ8SaGutBTHURsoNjUTqbJR
JtHfM+sqALiJpuwuUyEAS41bOHOKoLWmwhD1F9oDdbqSozIlyx5plzElCKpSLonD
OI4FEG14/l76fR3UOH8t5BJTiYqumapetbt7Ey/dQ9fCZKJYoKxKQShwH7RpAlFv
Ptmqxb3TK1NpozbCTt5cSMARL2rnAgERgx26DgLFgILPyRpJzqS7oCuRiPGLfGod
CUUrjWFOT7KmSs5w4GrIB3u40DmkfMf51kc8nO7qW0ku3JzFWgbSOqNx4Fx/30ja
vupwdBB+P41IPQ/vmXvYiDGwVITq5ctnTXIkfHytCbKOBwLDR6n+rttcR8fYCOec
9+44izKntNNF6D/Z8NRfyEC3iosMg+8toTkqCg5X5P26k/WF5CBAI5K7G41mql0z
Vek1DRlFfo+Aa2L+77zF5Nyg8u6d/RjGhCYg54gUgA/pxo/iooD3WOPVE2EByU96
zlBEH+llIUS0Z4FF6FnB1abYWnUi983i4AKtIDVLM5LR/W25qALjHHVgNxbWW8aE
yo+dtc6odWrr3kLmZbjQgl7a2lTZ6Wl5xD5kFO4+VUU8eGjBEU9yryBYNzxT+gfr
svOpZGpd3tqyyyNRsT5Y55WhbPtz7CghkXrxgTdSghyimoaBPOJOm03DdQj7IRRn
Nc60xpzoBU1ShBbh8EcOYxVtSXUq4jCgG/RuMrx0C+tIohAQ1aRLY1FyYIX4hNbd
1Xh2KgUPz2FWjCcFnkAtEU265jYfN1Q/PoCYxNs/O7y27+c7xh91kKUgiDdbzwkb
SiWeApWrJmyFWID8aLDb0q3cPlrqIjQ7W6HIo2YgNSSXJFD4HZNmNE+nLHsfChSI
SO6no+BUt3d6+DCj/er/3vxPlDU0gVMtRe4tfC2Q19MTspFGcljC4RWAb4ZU44iy
rL9Pd7AwmoMcW02fr/k0J2fA1x/9FwOsBmbpliCdUwUY7dp/bNpPfLoMt+hL5HS3
NKzUzo6VUaWqc9C5A6cbhf352D+bK7zQMhYcDbE2LSifT+/b1H15CmAWPoCLv4hN
BIarwFYDRuvfu9ODgAUAPSQempciIE5BJN/LAe2KidJW14TQ6G4N3MiFZZ+cu8pz
n8YumNhlpe+N/yAVttdQuN48qlx2mpAxPv6T9LuJM+TZgsnc/mn61lxCm7ppFOwk
ovo11LbFEAr+Q+GSPu+7yYiQy81amkPk/+5X0wjPB9S6WHYI1wGfZJYitlnjfojs
/up0/Zsna3lpUuZ98bBq2wwF/N1drH+IiNi8MLZ+xfi1/70KXYQDrvJoAZItHMeO
6a1gX8SYzYFLs7FuYUaWQwQVSIPZL6NGNPTihgnUd/Ge/WEtlWGeo7F+5TnDyLJs
kLCShedvibDc+KQG732ArPuSc32gz8R9OTdScqkXjw1ZGioIkOSgW4D9OYWG9mUb
h5ecTGczemMM3nM7WF0hGF1rokcUCWqiBtikInAWhtpe2wzjs+PmopRLOmvwiN4X
vHp2ZQuL+KXYuaKEWkZUMadG78xX9OkbseDdwS86kSUBFqH7M8fDw/2MRlrvanI3
ZHcK9BejvFbXjRFGaUGtOTzu0hVivi1YOwA/ecNNhYlQua+P0gX20OVp9AWdaoQ0
QuIO5rG0K7EHNM0LWmBrStu7DTknQjoF+9iWI/zjvnn5oLgrd+yhclwGrtTv3/4g
7Bt0i5D83+hpbFNNd+VnUEqvVsbvkxLcIWKcB+25RGNDqtNFbukMNTWjdKU+uqmZ
jCziYZ3AeSCKc+9X2cBWLPty8NVsjKT98QWtR0VMBOBgon/dTM700KrnLvrcFAmT
rENlpsJvlRnpFXqYkmDYFNWbVORAMUxoBFH3Iw3sS9k7vglZwastmWftAbV5cP6z
Sh+fA+SLxHAkKezshJtPvfZ/HY5/WQ073w8I06aYx9CIE6wJZcVeCwEa4meGg/eZ
9T0kkaP7QPCerH+sHTJ3ZmfAJIyWl+Bz1O1b3qvguNjtjM5PHyi1dG91eKxbLPS6
V1mQmroKrCD+C1CN0w9EmlcXMU7lKUrh2HyaM9zamNg2vKmKPVh/COlNcwJP9xj3
hUyfpN7T8KoLfsiI3u6C43j78HJlCAA6vYs8H8zQuGfq8Vy9DaFVxEtQHRnJ4K87
TYw2lu6Mr5LOH5Mcwk5p5hghdChppEQ7ErtKVrHuEuf8tW+3EL1Bf/z+pxdPru5d
c60mQtEYPLMllKhjkqibRQDtrGeizeIGJckogMj9f0JWEr8Ep2tW5H3XvFuuSx+H
NbSXJ9K96vREME1/N4E9B1MRDxlOtfOVJbgH1pH9WEdF6U3gpb/h+mnJyH1IqLHM
IXDuPdQ30z8uPm+57W5r1S4b5jllCRVL/OrvJJas53fjLoIpcRxikbzl8Z45PWMh
V99kapSEWLpUNp7vc3YJl9BJtsh4iFWDFr1PV1IcX3yEP0QGZV4nwArEmd9wJsNm
k+Jz+V0q1X/a4l2UIiJFQN/mF+5hPONiJDw+5/fNFID3d4XrUUYWfTd2ANatcl/6
MSsbCgLL0l0onkYLT4Am0OdSaQ9JXgyHejxke1p58tX9w1oB8QwnhLY3uDJy09GZ
Jl0fOJA/cjaKUBn6E3giXzOejhrSnWh/46cemHVAI34BW4rO866RBBdP2EqmBelv
JuHWJiYTk1c/euggGyqtgVPqT4pcoF39hia7F8vuD2ezU5xdcB0fw0sfTWgoT58s
hcCJmCEH15FWSyTMcEBrPizMy5EPVCtgBAdxjc0vdYnkHvRm2HolWUnxHt3CyM3w
UJ0Qb3dUHtQyAOd34NNSJslnLQgsI44KSUIovKG0yGKzNTCZgPT+P7q7Gbjo79PA
L+hb//fCnMBojfRciiegfdg2P1TiGnMucHWZvPrEiGr/96/o+a9v2QbaTabMEmtU
8gNBFpl2uAVgRpbzqyvGcmGpjXfaRRzfYzXzBlynoyGjHlW7Dftlra9kkeaBWhmY
1635aQiTl/L/rVswGPcE2XnOhwm41AZZmTdLxMveiA2EXgMASV6Y94kZ3UFjSUIl
QZVtoD6Fj8aGRLfvh8w2VC8KG5nNdJUeCVnKNrXqI4uh3mH4kF0ZIRFVHn3d8ZJU
UDLxpYT8Zl3+MJEH3piBksMUg0PHlk0tkvS+oygLwjA13zKK8X+z+HLRTatIkIib
fEH2LIIaMGneaQIM/+HpL0V71pECihw1W+7Fe3py60isD+Q6RM6kLYegppY1dCTe
txgGwkWoa2H2yXnLsBHSmfImT5Tole96Ap7UVX7OHikxMpF4Ele6ehT/rFGO9UlN
H64+pEWZ7GK1eyOVuBN6VGfA8hanqYmizKDfhddy+caxDoM+gtDXf48/hDn0M2tT
yzkfRq05/2oFA4OXGuySgiCd61XQIuFoMYU/fgfZY1ykIBu2h0DLjOi3d49nDkhL
GpulW5vaJcLzr7bRrBeyYOHNIDci2rlDXGYsmrXxxhACBcaWQSNh+vtOQTfiQ2zS
WBXFx3e6qp7ZXBfejMKwfmodHnFgHU4/9FuQG0BSU+fPnyw6f7rsBrHbkdCwgg4y
3TXB9cRrqbjTi+jv+4NK8YyBme+5/pOOQN/xv8N3THxHBqy87WWi2osTBAsB1RDP
a85KtB8769JWTS8CE86YfgXHnQVfTQz4rU199J0+MiGAIN2ujAdTtukatzXqhmmM
+L7NYK2vbWepsz4zwAsucp2CW3c5P2wGvAf+PibRCLzQZG0CYIhqa/Sztxlu2uLc
qO6saHY0gym0gAIa10h9RKLnoUuuaB71bORvEZzWKdB2khXaeKeMQyX74Cyh/ENi
L0ISiCK2ddbW9HiqliK373IsZ+9Up2Q2Yk3KHRHvdiCC49BD2O1jmLRLuY1giEtc
WqwI1+p7otuvykEiZwYeHL0nP+Yi9PWsGBIiohcRdHoljjUJpb4bAciJoA8Bm7GZ
K2bXX4hR7urHczY58U0p43iNycMySXSb8BIiKch1x2rTCgvvva4XIwFt1ErSn8Ib
u1DlTnlGXon8Bw1tx/dVYeK8mwgmMCtARzZySOdXLdXqrcfhwmu9/LaZGEGWjvyE
PyY/0uYM+Kktcm5orurXezzoD7dSF8FzMEplM9qH9JSoEz996EwIQVyPsphYhKS4
7tUVBupuq8KwvA4S1gxPqdvGafZsbN/axmTir4ZEWatwdk+y/5+DHL15VhJ6A8hy
KJvynPbh/RdlbcTsN2bLLsQ2NzmdiJV/hamiWKAEMrBFkn2LMrEYH8Ft3kjEtyYJ
25q+3Dswr4CqmTQV5KPqt/KjGzAdDhz9IabKUfO+aK2lkjIz+Ob30IZB0IhER1uQ
kDime8oQQT3ne4/r5EER/gl68YKgBxqCZJffeJ3W0+wYVqAeUdbo2qCm26/pTeeq
tQ8+DzS5CNZX7U35ZeIeNj1zaGm0k7MOmM71i/jZMSu2xp5MHYCgJ8vpMNt7TRnV
Ns2SB6J4or/3WuSH1VvUio+QGDWEuqa0PBjYGIN1jIthQPXHLekNE3oVIU1OdhTE
Rji4cuyxY/VveNR7fzsEaZGtvAvqCUBWnNMETjK2yxNxHpfl2v2Y+NBLhkEXSUSV
z0Z82Kd0oyfdMYsjxXfpwa//ZiQYodgqf/bzrDZ1nloV5k6ogLdHdrNYEIPQX3YH
Y+I5kytrRBpAitT+qe9cDsG4dc75/Um+WVk1gTM99qnH6XPlWT77JwXAb0e53Rzz
DTFf7yhbKHPxRUvfEeXMfgFbI97MWXfi0OAq61QiC3pXNrpVSI0lh7v1UQ07Booa
r8tWblKO8fUkTjnqlWnCunllEjN3AfJmUkula2nDmiSbn3aoIw6JifYe96s0pPfQ
nFXUzrTxa5wqIqCltt7ZPJaejRrON9tZCJ5ct0OpjAXly/M2dUL2pDlOg6/a2V65
EuTxxOS7eXzjizIHjy9CglRYW398fzwPuIh0s9jtxmprXTLg3IpotRwqPUK4K1Qi
ww7PF78ZbNPNZhhPHZktzvWilhVofC9K/3YZ+yV+BpF+bfEW4wK+lU8Qmombw7Rq
ZGcI9beGMpyzwj8pZ9R3CND1ygTK0i7QjeO2bQCUxGq3J7z7HDQ6sG90pioADMDU
SGc+sIbaFCV+Bamrq1ynU1vQaLhr8R+IeSLpyUSdM854PmtgmeUOT43hVHuHf3v+
uXW9nPED8692nDCICGlSuys9rKTDDm1PizwYtVvwDLXX4d+0DHtAH3W6cXq+hKfh
vpuUEA+/z9n5ucpSMmx70vJvFDn6/QQjmXSU2WdqD2FX/SGqNmOifz1tlU1KpGn7
Ych+W2hU+cnDX3HTrnnRSpKhoud0GTD/8q8YFUGy9Zi6IpJ8Ar0ZUF4tYVAawCtN
sVaYDUHaol/Y3HFNrmYHkc3Bv3P2rAuUO7bWfH12Le3HbgBCbce8VHTVW/RdwVnr
rPUp1kHxEAAdBPaY55eEikbQPQdpuHphYyBX8WyAT5URfPVuj4BF7+KgBaBL8OR3
XqxAyuDaDFjlY7hnMblDnThSxg8yUO/osjPEkx4WJjsPFlDL80Mu6CFlna7C88Ja
74kAGokwDv2+kInzJFy3UG/cHgASE2WtOPoQl5avyrrVBIYioQrIMkzcdRZryLzN
3eSd5nwt2Ke/yezGLVX8sUF4O2/+OX33Ym3o0xu9vkYzEvpmBCITYf6ABFVJ2Dev
biSUf4gexfFhSOCp/WdYOH4UvMiEXITlE7D2fSonWJln/3JvfF7k5DTfFYkFnq7S
/2cO8qvV7Zq21YNY1ka70I6nhVdN0Y7olBbEiSUl+LquDlr5omRnX0o9DjHlGA8i
RJ5Y5T5XSBjvZDqXvUoobf+/bPOj5ecKcUGdnXqrmU9FqigDUTJ8OVXDy29IT13K
4btqCBZLndciXrFY7WCCHB6XXAAndiapw89ePm3BhnIwIU8F+rxy0MC4/wv3NMTv
xJCzdPk3EDdHfP11RXvfCMecdjeCf3+GtqTpKLCuGxWkJfO/LPH0QRwa/B/dgu59
O//jcTj0ELZ15njraqm2jgzJCeZ9LHRuvcQa8D1FcVHvhpyheL4h777s4nzIBbvm
m/YHx+SrREgkfFP9GISt0i30vRsbSwLU1HlhHZ2V66z64/PaK3/9HfrJrYcjtfVE
6fp6JWqjpibUWMeJE8xoL2uzAGIL6uGynoQxsvMN4QYSwiD8DTmBQsyOMYOvsosu
PVTXOZ2FwLzNJF/kMPr08yl0JYjFzp/Gb9+E8B6rQYOZRBmpiYXzXWpakMch5wew
rf+gCnAxAo2TnvJQ+exZSThXIOPQXCE0pHX1J5aKOs68a7wod22OfsPdW7NapFIn
UKxE1lDR5/KTS7G83PjvvjeQQ7HxBE+WAI3MyOeL+vjM3wjUlO88HBwtbEkEWKqk
UbeX3AgJJlsFZA0V9zpKfASbWySCbt5ZTx58H2WFSxOwt5XDIQlsDxcwCTlVbFYu
Ftil/undBcnQHIubENnEu/+C8PD15aR2t6H3Qs7Qyu+tpdbTcnlOBh0c/NfyGNes
JIvhl3oGwF+cr7IjVVRVQkxhIir0KhwUQNVkyuRihDPrDIJCnRXxIWe08DNhcWJ7
8Zr0lhlpzztVaecBCUP8eRSxVPBb7PpodksEywoVP7uH3W21bF2WMErkeXt3vf87
DsoaQgYrib72fgmyvYmzELlLUvRW7mFZ5AcG9vo+vGJBh6hdM0awv9oO2Wydb2mq
CkwQ6ssPNz365F+IZo4oFaQO0osJREd4NegBCw2LApRHercm6YHZp8GyGv/noQHE
ipUlbGtWTQwzpoF3vuJwHACNp8yXIMYwwReelzCm9IRBHz19/zewXYmTCQjCKNCA
Go+rNpvY9iiz1rvb18cP8sI2SetfA9ne6ZtXoGOFUHNo5zUpHr2r1Tn31p9+7Fg/
zmu8E8xoq3Y4glRRt126BX8IisFqZt4joRrDL14EHzLmOku+aCHUvvulBUtewkw4
Qv5SjWIZewmfQYYQDkoaPuhelmfOBQ9S1s9WNYHcvYy/M9Cz7dZ0AuN0/GwHiomz
h+l9IGiflnD+9JEW/7x518JWpEsum2Fiw41WOjUc1qkRs1gLMTgiC1CU8hYOKZbe
mn8Ryq8uKCZJB1iI2oyo0Axi5qGJ6aHF7B39kIDSfmYyykQ8qbee7D+MAxkvejFS
5YCo2BYtTN+E1f81i7W2RMV04TbuE6JT7sQtZkzjGWIYR8jcteNS1iytTqfHSvnU
NUE8AbQ14FQiLsBtRZnRaXfDlF5SHxscrDsGLwCrzGiq/8L1YL6SDIqiBBvzTie6
cslj0O6rh1jqN7Lgnt85USE98cXwq/mHYPKJtJzos66wApUNVbARZuRcBCCyy4Fu
8PDcm7yDZVtgQAaKtJHVDFWEDogoH993xP2XkQ+2Vd+P1DRBljvM0kp+9q7qebOV
cYFFOF7oZjykCdNq6sw0smSlUla4Y1eZgmLqNqgHENkiL/YebfHHU0xQiCyKFcgC
ZAkYI5V4ZFJbEt3eA9f/ijqkLi+JFSQtpMFkdLsyhtCJuJsWmMO0kGN9P6CxhtnS
e5Uc1Yv7FRe9Y8Ve/jvI+x1VKpkxubIGyMdCEi3c0we4pWDMW3VIbPCE4g+yJp+O
Qx7PlM8ZFu94xCdHTJMYSZ8IAxJG+92suhy//L36j61S5mYU3bjQKWNToCWeeXOz
ZDZE/BAnKPJgUyZruYrK5zsVMlW1VKhZsICC1nbXzmXpSS4dUWOL22PKneIqH2Z5
HGSUPRts1VdYYsoI6L1D0cMeoMDiN3dmqjv/5699WDBELl9lI25In4CBvNHy/RCk
MCUUaZL7JQgAkRrQvtLS+QCzDN82JDr1A/tJLkFsrpAHhx0nfh3yYSBMg4iwZKL4
TMwletNOw+NMmtLHOw0JGhtm+TRf2BfWMKilxDTXI2CkqgYpWngbGfz1TJR43amd
mOEMCBQq1/hd2DN4iw+PiYdwUa3vggpXuYUSqVGAg2B82L+2xqYwE4O2RrA5cXUl
AAjimkNDMywZBVGRyJAqaXcl+Tsetvqf4WFIxVaqb9C76t9XLA+tPfgd/01ZSWL7
lBcA8aRbVRpjJtN1x8AWaOrDmy48fJzm6oQBy5LiDFQSLsLtzy81Z0870agPDJfc
5fflVg0zmv/XQE9jmriKArjlOJlEeX4znFBZq9/rTqFyCDn8y7kLib2eSbm3duic
o4h/qh1raxs5Cu7uROfdOPdLPEbZE18Hqwc1cB6iz/ec855sNMPyqonimVHcxoLh
5IRB1MyPgK8cEdd/swqTu6aBXqu3uN815zziE1YTt0QLshK2MQuzcSwn+asLggMN
dqK+S+pZUVCZCGrGAxzZ4bPr3s/3cyXW53JNqZlWlsh4q+X3ZOjTejoxX6Mhq/FA
Ovr3euKiOOGnj3TEi5qyLW4aYsoP0Mhh4c68wj4lDivpwWjKePRog2MhKGj5smeG
KhzHdHlmb30H2ODzwmPqm3Q6GFGxPA/lagPVLjS4XTTQ3BBhxO39LiUyZaFBwLS9
CMN+czEXdBX0y/nb7B93Axik2+OuwcNBd1bozLENZMq8GIoAYoQEGcXIHnafiNzL
DoNJPChYzMk2mdq7BBa5g99SuQYkFdMpznpQlwC40vl61Z/rkhsIIqapDKE1T+Cb
p65WjDnIeyb7XZQEVrWXnI4Hje8SbdOMuqrva2HFTKUM35gOMnFkk2ISdDOzJKhL
Px74FBjIZ2a/a6NQw46o3XwTAa2LFEXc90Uif4F45G/52cjR6H8qkoqxZ09tUb9x
Kgg/bAlTUPdq7tvhLm5P2SbPRic2MxI6DrZP3QSjD2Ei/uG5pw6BdKc5O1t0ama6
US6PSM6FgkoF+juqgaI+FVFM9axlTekEfJOu16h48Wb4G8+W1ECG+10me2IZPHZH
veNtMsXUsJ6Rl9w+Q21uiUyY4CtdCSXCOa/Qa7SJd1AWdVaMQW9B9eRMmx9IyRfV
Go2mYJpay3a7Ct0N6ikVrPzmdZi/bCj9wqcKQnLvKBkWT6pgGL4c8ZR+w4bMDAFb
2AArrAJkUMgSMlWOOvzZgifW0G0YjB4hiOfX0/gY+S10yckH8F0RLbUj4Pk9+65g
p7E3f1FU/U1+xvdjT+M+G1vny2x7NJh84B9H/CBFGG4GBnXjEkgmcbB/Zdd5K+R2
y79+My1kSnAiLZW/8MPFOnb7lG0gZ2zgYrNhhMcURHyKanBOpiscDTSecjvBjmY/
tkIxDlfW7uxj0mXlWO5JhaeoaG1pG8jPU7x/z0u73C+JsYEKEN7sKQgXtKd5CI2W
jLHmXAD96vTntjI3d/j2n1nOs9+wrfTi8uVHe/7XQD4GBFnveKZ1c95VQgMeffmX
lCVGmsHPc3F6KaRVQ+ml0xETVvxoogIcrsMgn1qhhbYMxA99T6rSyD+8thJGhYTt
Jzz7kttsTxukgFuLhcGxsFLRpQjNhhzzQ1NQPopKEtTst/YbxIUfc5Oh+8jF/Rah
xVd4REJFsU9hsnU76KJC8Au4GdKDJQI11etN15/+cetb+xiHSnjGH2C7BtDUoN2i
WFrLLBfJ6qtFx2HQVL/rNRH556h/z4bJu3vQv+hhNdEihx55Sx5vZnAlw1xKGD8o
1E8LzRfUMzf68K/xaRly4y1+h8jBdOKj2iDdwnLM3NaQmNnrerPbOBle6Q/tdrDZ
yeASEDX1Be61FZgU9bL0um8Apxs4bNPBRsp8bO8C43c/B1EUZsrx1TODFSpJcMV0
83IR37U0xYk0+XOKwnpAlsdCyyxidDDpf4uRKcQeTvsv/lk7SKeiowd72VDoYHT4
iub8wv+/HrLU9UM466JhwdAIAZeuwj4K5GroL4alnvX0W5Hr8iTOUormJr+T4E/Z
ATuHYSUN4TWLO4LuzC4bJV6YzStQYJ88I7luNj1TlGy/vLORh+UMNUbVyjwvXFLC
zIWGlJX50ze/vINNJ4YnM22nSMeIWhWriuaZDIBzLEy3DTDk5V0yUChLLfzlHshI
H9hZSBE8a+jm3yB0zOIcpolwnwalHcv7wSg+8kMKeeB3QkHHVIkpX/j5BTNATZkq
60r0kTm27y70dibE2z+c6It35WxbcpGE44ibYnfi7A599sYvld6D5l/NRqmOGtqs
Iq4pRJG/UT/KvLd4/jQNQfyGFaSkbZcKuLP+G5Aao2G+q5bVAmKxULNgcFOb5DOv
QXCf3t0MVSyD/iIkpeSlCugLTNAQzVXRCFf4UPe12wEhtAv9jk9/+Clr1iAVdkVl
x919OEUkz69uj8R7DcAJTI5JoE2LL2OZi57QJ11niU/mCgFLnyrNWvDCuDBKCu8l
yeBG/+AUES+96/fNBD4Z2PONVdpACTyZ8L8HAflCcRQd5Z3pUmYZ81jAe7Nk6YC9
93z1T3LO+qJ36JADngtTOPDP2nsaYCh6GRWDWpzyDVGPGb16oNjBz3RcAtiXk6lu
3ZevuGxkH6/0qEBQ6ofBi9F/GWEBV5JDVcXfhF632ZHMWVI5SzYVzCcMGvF/qnin
IGgHZNN29EBpPPuhGQCwQAZ+BYuKnv4OX1q3HA4wGp80V6/seVqWsT2H80BVRZQX
GlB52hfBkB6s7lP2VIphaug5nEN13qhAL1SGS7xL0KMPCv3obeshnIHLcbywRdQS
y9fMR+MVH1j+Zekx3EjVMfhhvWNsOJnBQXpYkays3FnSLuYqHvdRJE+Wy030aqcQ
J+crvD+rbuXJh4dS7qW58gDskku557iFgcMm6E8XqpSpaewWxxm0RIj85mqKuV1F
h7GZxHZXmfP3GFUf0Xsw3xttzMDgxRdTd+XPsJFt4ax4TQAEdLKjImt0oodGMph2
IJETnyjifMNxwZLlgx8bfKul2JGCcNV8OWZkgkxV+L4SUUFE2pGuCPMVYoEcmj/6
MBorv0L372oNOfJBu2gCWkoOLGbP9RO9lpRt9kNAoMreXTY9rd7URUYHTyP/lrbR
J2CTOv5uo1PqSIwrS3B+srjQcH/ZMcLRus9fuEmGT5IvH9WnHUTSx2AyFblDgR1e
5m+w7ZdmNXVf8q9YKPDjp/xt4I3b/8J//pyi9Ge/nn2ipp/jjMtTY7u91jGIoBY+
V9w37oinV+b+oNoSa+4dgGzevCmAdb+aH0BS2QCwB3Fn0VRxxZoMBmQ/Tfl0qw20
aiSb1V4D6/oyureJtt3eoeejVqvyb3x2/N0fZXMkHXmxRvBcLiUWBsgagXohrKLA
3fqHiMOD7tzqkq3p+yJwEol/SAk80bZstxmbFReASA0JbqZwwwxb9PRKS8/GG3RX
1rxUqTrxQo6xcPxJf43imIgNdXzNw36E0DQKH+FNILxTfcB7Y8HvNTqsYNDg/SeI
tBCB9QnEPd5aXUklHMz1N0ulJLw6cuOE4CPfg2Byoq1z4coSVYJQFUbmyt9iwVBk
VVLcRjI94+/zpeijJTAd3psMYZwO5+npWxXNrS2Mrti7Kus18oxTChvivSQVPeM5
TKmuqaN1tgHap5ooNNcAF9z8gwuw8ozlx0tQmioeyb8x9v/nINdutedDg69h17RC
J4ujjoeY/2DKE4konOvNxRTN4JBvt6k+7UuJtz0GsP/RsLfows2PmoTy+SHJI++b
eftJ30/fmrd/HFNhwpSOxKGIkWDK22hjOe4fd5+qA9Xi3NXG9GkyHYetNx0zeGIw
Rii9l2sVbXPWSWUgXDrqxhBkZB3XytKtvPf4QCqubERJgAf7RGNEh943J7GrQxYP
5RTTz5gJFcveGk5L04y9XkVK9+FD8Amk12gaQlGqedCboqhJ//cVuSEBal+rjNkO
v0no4pXxyvpLwwqbc2Z7RzEg9n41Fw/wr4C74zJgqjb6zcHk4377itRyKno/X4qp
uImkTJW90M6gqbu6rJfioGNYdnICWLhF0qzaZDZURq7P6e5chCPYGzIMeH9q1eO3
kVyb9pwLStJ+B2r/ZmJb1Lj/yueAo7wU8sGyZGkjqz2YGg2FiqvIwRb6RxClWf6T
K0x7Wr2wutHiXWs8U1qKVfAwElCR/FTuKcWHnhLHrmhtLTvI2OmuwSAQffL28/sb
OauGD6Zsa5+mZ4GxHP3i12touE+f4gcxU3s/IESEYPQwQzo570aq8FcXL9n/uhkJ
0kITf5HkmwEtQCohWvJfdGEXBVtmuYLVZ+hnMPe693GSeWW5VMv0+Xov019skEfa
ovxkLZns7wtFHFu671RSo/YqAT8JFnqb8YtglUigl6yrXE1tIzwtRab96csoz8wt
hVdLKkgrxQhL6Pa7U0dedbhH2XPZGoyKNwLRFZgIy1IX0kawhYWVYq+eBdoqRGkE
UHQLvo/JoEEJU2fSBi3ChV2f5ppwtai8n9QN0hPWWNfA2z8hvcqLvcv397Z98yfa
DebYJANDnp+1uDE8FTldPuSebqCYS/kAxSSyE9gNprGwpqHe1gC8PWsDjfNbgIpb
MIr6N4qpQ1WvvBe2rRuXBCj/GSe7b9H3TZKzI3ehdpBmMfeLGM8G1HfpunqIhIal
6iYL5PoUcUixFW5/waqZ56pHfSbGfm7d+p4cUhXHqvwDGDoiM2yGd90BAuKvjTT1
GPxZzEaOy5TIoB834soOBcdD+4aLxmBhpUPASa6YrLIe5ppykGluE+CYnHYGltVZ
zaQ1wEkDa+IFM44meCINCh45DGs0A3x8Fn/ec2ci2/gDqJRDRt6WLzLPeOo7RDgf
GLYSNwDzhdiChZzpJLDEjz5+sWXXxe3vvvSSJen7wP25LAqdDLopX4OQVzQxM/E0
cOFdeJ1L44CBHduu0f9wk7sN/1inmknjEUuvtxVqgPWosPhD05dpE04HvJGXTzYt
awDL6p7Ma0WeK5B6ogfX+UTiN36Z0boy3fOkfs7HiV8W+CqXDUxNey7q5vArZf7Z
RfQeWLXcuNkiM017wSZDpdxcaChArknUuqq1rjBGYkA12u6n416JMLlxyEoX4rac
5QXlVQP77oKx00zLd+PcX1rrsVV81JWbKrI8Z0Ha8wy/1qnOgASupEX7z6I0JY+x
lIq65M5z9bioTFKGOGxmdn5c6S5/GhRzt95GAOrHk6NYc7ERDdQsTEiuWXcsTUcJ
TC16NC0CNYtEwYIv1iKQ+qFf2SCOU4ZWq0Q+maW5/NWlWECcs87W+kaGvDkqfRb2
LNhVucRfCFKC/EWG7CAod0roHqo/Q6ttXadcj/CtaImK++PKQ/KXCuR5/HErCV90
9Jb4BiF8FBe37ScKSBUQybTsuMoc8TdiabgzulAESxQIkqKITPODTupl6UsW/VVl
JIjqZHNpa6+E3hk9a+ZGFzNzeoXhh1FpzxoAm1RGNfbyaLCJBwN/ie4IQJAL/78y
9K7wDQJW5m7IFKNYjIdGypVXjdGi1NJ4As6OsoeR8s0biqoVca8vujnHVSyB4IUG
u3TbWVMocSG9felq1a1/P3lebBA6icLZ+p2aTeUNGU7rAHTY3DOQk/JnS+YJzMhq
7quiKuT4TMgEruw8n0jxl00GnDDmiqNZBMp/mgy4FR/cl+WWwoZxPZdy6i7mSiG5
CbTZuXejFYpcfjezOhDVvyf2COnDlOtnnMcinteHAZvCpLQIZXn2VPKhdXnzwZBT
DuqWbSxzogHZjL2cVgldtw8E/14TWNPS7YhcDwCwt8yYFmEKmfAikmB3SZmZOdeF
1J2DJiHQ+TA8xFwrQe7k9WJAtFW6/ylk7JkVRqpUhjHPcS15ciaxUtbNOSe5kiZC
YAlvqR+fJn8mhwtexVR2xTQHBhMj6wmEFMGfbb414Ks+9NiI0MwO8zkXUPptPKgC
Ls4MX1VvMBLS8Oi5JjLugDLaDAm+eKryfzZo5cpFXDjglexjh+QPjJVeAPR99zpv
IZ71h5NtX5OaNvk9tI9KoCsDZG7JIA9gq0JMcu8XHMRC1j0wHnxpThUUiqLlH7mi
mriMnaICe12jDboPoKCokxlx5V3dlJU2G6883zXyRTxone4ctOIXDa6oQoWk6D2M
03dEJ1KKAZF8B0XOai+FCywx8bl89hXskckBr5uIeW1ApxWHivQU+PVQNTpuZv8a
L8DiGXtyE/lwIKDv6/U7s1TFuPnRtPGir2O6OnyauvxFNWrX93xUgflqxIO5tE+I
UMD6F72l+ifLS7wdhcS+nbOCVGEzB56dSw4u0O07LWG0IvLHTyI26O27LOUywZV6
YC1FYQjnTU6lhOrh5cc8wzMAR2cCdnb2D+QknsQap1lyDjeQKTagHIrPz3+Kb9JA
I+eUOyAl52mnj5COZ3Iza1++oFUjIwcpBzOEnttu5GouVmVB5SDb3Qlnea0eNxTQ
i72peuuIFnW+pDu186oLIygdnU/oNdZbb5zehR8b9uCKQlG2B5wQFCbylWYvrAH6
zy89YaoiSP+e6wDmgT52TsaGp9KQy1TLo5jUY8smETpDDxWnzLbxC8gneshckANG
IzYL6/tWHEKp6kIefPYQ7CY2pRNz00cw4seO80EIkrW12kdUC9F0Aq+QAgKlpMJa
3zWxaiqvprIgtoXIg2hZzP7nyG9cb9Qfh8TwdUBiWSW6adCbCElXpua9rtNKKuGt
Bq1L2AfbdMQbJ1w5hYka/3NAPG/Vp9sZK+wvcxTI3enGtI3Ku2gqK+e2jS+esDj9
l0aVFNBHCSKwlkOYl5+Ws+wLR/gWq10Q9T8pr6bZdsVAgCVdWGdbEMNnwYCPdZwk
1iHHSOhT48esgkUFbW14P3hKB0hV5y/h1/nlbQvvqRyzkKnI5LTEWpXoONRlOFFm
wcdN8zIWmdVpjIQh5umU2/h50GwjEiMKU6YVz1PeXvUsrh9fxfoHypTuPpVefbGT
M0VzUcBqMXS+l37/MjATAyk2bDJwcZgGX61WyxGVxRBXgAPJdYuc8MJkxvAkRy2W
T4JQYMAqN8dluAbrz4C8Tdo+gd9pV5iJfc5cBaDMouXC91CVPLP0EyYnZev7us69
eLgKfDn1b81i0OuBHhA0ELrTNoFYPAlaPRjg8W/ShZLhc21Cr8qKMrZgxST3emN9
ImzUbRR2fDZ2RYkLAf1xbgkhEiSjUZFbp/Xj9cHFhEnucXqpI/U3CByfBYgZ3Q1s
F2Zy39CnMopiXw/1WmYvfrQQu0YdZgrD3f7e6XGBsxoKtjCVjIgQwr51N8+CUpbg
JxcsefnMjWpniRxUgY7wBua3xC1wbYN97LAozaThN9gru4qSXoL+hM4a3ICTcjZG
BamzGJ0qZcMgC8N62yec5UfyqiuRXZ7196AAG5hnG/xZofVThWym5xmqpTayCbDG
HX/jiOcxWxCbwfIjGGwwXWVBAE/3ZxlteQxis3TM2VlauagxD0pNMYAqHk+G0ggj
YhU/9DbDNo+59j2GGUYaL32ZzFY8tCC4hktZiTcuM1/cipMF1SPjfvW3gIiWFF04
G7ofqzuA6ETAs7KWRN06wdxfh+avUsYbwVvfH00iZERIZDH8NEx2MhZtfL/KJ9ew
PH/4/14pb6jszNL96HxqEN0e6h7zJdpSDxhhoCrmWLyj6g6Uxdx1UVhTB54lYLGT
Sa8dWebRQ1kYaq631YmBx3r1PRzKixsP9nzBgvTUGEoCw0fhh6Ssl5FbDLH11Hqy
ZgoojBzgopsycLlDDIFFOOAzO9EJK2MPHZ9nOmJ4bSZlkOiCZTjinU4RH8KXL1Ef
yV2eoRDHW6/H0ZOgX0wTtHKjwgAz1+STncmJNoFOJsm6ndeV8s3yZhqwghlNtajW
mCw6Hs4V4NYCSpgmr1eoAQSIwtUAhtbrihw4+CSmM/M1wJHV9Y2jlSmuq2DAcmA5
+AqyMtpUd1G1OsIMs9wwaXIitmtumw74tiFE+0W1VpvhQG3y1ywNcFN13TgeYxCC
QFMAV4mbHsxzEn2u3xJvIJlbUzcZCaoyg/y2WzBBemzu/wJotkTKySHztXzvctVT
Xv8whAHZQY057Q+PtqSnT1lm2FjryG6XDquCyZIXwjwNBnAVwcAb5mTQeLAE1qzR
5320KomC5S8c4Tvut+qPi33H3MsO3/0xTFCbBBQLMEfsa0mnd7JLn0jSzFBpbeZ1
KaXd+RgQ+FYfQNN/DhvsXYBMtMECeVRS45HfpLXCS+ToLzGnASEpuRsfHYhVt3S/
s7n7QjMi5CL7PKpNC17eDlO00ohF0YOsyUQCOq1un5AsxjdPamxEUWytBEEQ3sU2
rQLLOOm2WhDH1PUkgvUw3JDtuntLwQiehY8R8eMFqyOJIOPddo2SI/UuDGc4j/Tj
u+07raohu910enttJHjpc8fsjxRh1iuJBraqbXE+ZQxxfnr8sHx2Y7GE4rO42Obj
vBABs+OiZzqECwGJ82k+eNgXWseMPNtGBe7urP6f8uco+P0oxdb9h2ijrpoG8AGf
r246nD80BFC3hVfWmySmHjdIVoE3T7+oUFpv2oddq/pNDkv7gv+S0eGkoVsG7Gzy
q4XDxBFo7o9dDQmB01FSoAOGZVOpcRThkhJz14aFFKsEs8MDSijdjeTrPlISnY01
qF9OMaxCJ8NjPPt3aoTwDYJdVaDP0ilMBO/Nht2/LK9kHuBU0xcMEMRzpGNE+qSG
TFKqArLnWxP8m2JzFUOtHlldyO10KtVkUINfsjorFFFR2T2pDVWV8nzgkxoJToUj
Qz9VzIx9zwglx+r8+93S/iG+GsTeUIDKX0J//gw2JXtW5HP3AtgeaZGSkwolzDsy
lYZlVkS+Wzb0nfGwFBavjVpzU/k6u6UokN31iJ9JP8RpNuYkcnhgTsiy/sjmWjV9
VecPVFLSFK8WIthJYTPMowtK82ZshT7kXq/Ex0fvMwKX310m4NOaKDKi+vj4qjmF
vanm+YcugEZJ0ghmbPzN3ngBMXR0FNrlJr5Gyr4CMPC47f7tHx1fYbmrxcFYe0IL
n8O0s7TOCWP0Cs83Icm9tjoKnmcl40f+gwWPRxJl++OmsCCxC0XFzUi8gEe4FHLY
7q2LgTm4fQU6ThSqye1mZtpkS6RIlQJCLA7jS6sLoRKhdbocQ/UpeG6rT1cqQOeh
ayipYGyEEGf950AgWB1WQvwbCZSEUsUMaLoz4SBlvgQ7HjCBS4fXkaR8RyYhF42J
HVnV89NNcHm07DXC2aSoDP5OvpQ+soUC5G1Yov6Ue6oLCMAZ9wOUXocVFdPcjZJJ
HmFS+z4LkrDOe06QS0bVVDS1CYyxZBYpbIB0jxaOTRKTVIn5MMdTf4LT9DbyXOfq
/8NIgNwamK36JsCSA4ZR1xWL2rOTeZl/IILwJQhY5f63pXyeFmKaOWVl1+ghjeJJ
OIsRjX0Ysy1cJYdHNTGCdxrZucAHQGpRsl7bAycvQ3kqiop59HiU7aLq+w6GtFfO
UwULW45dUfR89iOqDkbxqk1PvMGLB/xw1Ig4JS1ogtGFWEH4wJSvgriLz60A0yxT
R3BzzvkPvXBVZ5Xbih3PdKKkSo+bxdPdy0TKstNgOVYTP/bPo3qwAXGzrMVfSVmC
y46qVOQrQTdyUGthsFMJkbVbaoK7SbMH8665TDZiQjNb5mXu74NJjf/OhfVHJBOI
SnhXDtD/5P2Xt9x//htqEdo9976gjn8V8aTvVdP5NYGzVCsX0bDzGc3CnvzJrWu/
No58kJIkoqvVT7ONxV5kPo6kr4X3Fxp883SD8528vY1jep3+LgYCSAME51v+1Z0v
l0Mah2w9J1KgFzYzHQyeAIV23D11eyNnwjDr1VLWE+P9Ixwok/7njlXKKc64hpbT
bKKf0raaiGBB5wxEKM3QXgc25wktQ8Ym/LRyn2MiAmERHjNxMNBcfjrAi4p0pw4O
vclFXgRMoVCvF4YDcA46ndIlWE55Nftr7RCEriyda4QdiMcv/1jV8d5Qa0dvw3rp
PlTonEXggjPThZKggX8huTQQjUPUPJKWs8h8vE+VVlHSKGoWXsNjXcuIZj4PBBIy
9uJVqP4WazTNuGvG+E4NBrEJov5PjyIU8gJO3tdVv44Tw3cMUaqxwlhDK9oaaKHe
tKDNjhwlCOBEQLGI95J/9tmwK7ACWrbopM77LmnDd+jnzRhb0x1ShQyfuqZtFsPV
Vpuwgmbct1YWILIsZVuSoAqxt98zu4XgTl4ZuACPVaRLtEYqHR/lRkx4sl0bld8q
jUYGZ7oQYm8vMO7wzSpw7MUlgLvfogwc15JoOonBddj9/408dEXhWDXezZFwNqVG
lZhdmEk6108YkHWF/ynt9CUgYNIIHr9/Wuor5iYjau+GKg3UV0RCpeaWKSrGvtRP
W+eTuMz9I1C5tf5lwDp0HopweabsTiRFHWBPAXSia8XQq4f3m41lLTNWaVdVRbzP
0TRj25lMsSNB1Ft/ENFJCkkQT7UZ+J7lnRCbi41PksyWFE/wgWCI1v5K2PgEGG+G
JFhQpqFWkZNRt7VqUkbwis2aAwr2l97m9EToAV3HGchrlt2rRbP2Xw7p5/93iBo8
0wVXDK9ZqZjTvWKEfsn6h07WO6SiBOEbQeZCEOuqb6lUS33ehcopeQVSkVBILivF
xwg2TFJ/D3yoZG/RPPC99NVLGd1BVysO3iKEqg9IgjmZjPg2M61NoN9tMeI5g0Wx
oUpiSWI01dt//BcjISPSH6q2Bmo/ymzBoYDHWmXLaloBmBtDlOQool+zkv+wtKT/
1vHjCfw33Yd3ChUMoXaL3BxrusnyCRsLXtcNIbmtbc2pzjXrwlhurwiHgKK0zhpu
ZqbRUn0vABUoU6Q1+sR4YXxbQEhnuHXI/tMiNtFqjiZCaaMUZYX9rPWYy86IOY7Q
8S8kisXbUURZBwBueA5mvzLs5EzvkIPA0EQWKxzgpZHY+J0qxv9gW0IQ+nNqYrD9
MAZ2W0Is4fD9HSvd4eCwM01ry7O626X7vGikhtpiSix8EfhqSKk3z++BL9mRkDo5
Li3LpD79cZBxgAR7LxqFWo9kT7JOxais6JMv1OwBePOzWFO8S2WvlnalwckQRpFp
2YDmra5qpHCDT6OBVOLHJY1mTE0h8XKObHmDb315Rg+yjiqDGhc631kpOtqE+gY+
M+3he2E4bXDWnC0Q39OUAkZMWoPerF+L1WX4WDJHvjKnr4oByMPM/zpQ42Cko3PS
iZ5qHVjoEI3DU25MVlcGWiKfHNNBnkazE0oHCu8QdjLvkBbd9d+7n+sCxFs4XLVq
tHDDBPo0yZU32BRVcERLAdwW3yeWg20LTXIlpvNeUsUCv4ewoUwhRPuVqchKfAy/
pCSQpTyc70LJGornREzvneJ4utOwHu02eGWRnmZeGPZb3nUo5Bcx4BynLXHjZL07
+VIhFypTg2TXm0nK0Dx5KQ4ccQCkmnJSDkKOS2MldcvRK0R/UyUfqQsHlklyl/pM
tD9JnlKRzbR7GMBM0j6LnGb6Kt7xsSqnPu+Wax4cx1uziMz2q30vO5GAO0eJsMgh
vjTjFawMpBS5sJhCbQvEHfNIdcputkFAFlSr/teklB0lHC7Q1B06bmwTn5QR6S3S
w72xaEpaqxN0SAu20M5fLjQ4iyL5r4cc5nVKNP+I/L6cO3qSx6sgUH/za18OuRZB
G0cjXjM4a0W6WJXt3BsNmkRvJJxyLvaIqzEHoX6kJ3s2dqzAS9CyxD3OXLTa1syA
8vmxFeCjjNyzsFWME6rvhLln48iEsdQtpTBVtIboFCPzL+V6l5VE5t4kuC/FTIUt
2542tCo4CJwn8JXmtKmUgGe7Y9UCj9DnC8MRlkQKbMduTWuW2hsvZXq2RbHl8+S/
wMjN685ME7JGet0r2q+gm4GscORMXPwFHSBwzKnGCgP1c0/+f2+QI9G1H3w66wRH
n9OpUPqmaRTFM6cYv5CI37GUj4wYoeofaJ33rR/0EfuVNYbsfjNygwdQtU7+zvZZ
lars2n+vg0aXeMftWukBK+UjjxJM5J8KSLrOWC4br964XUQcaoIVWTTX1t4mbP0t
MmM/Hr1amnUksstqDFi08V0v72u2MBflym0I1z0wq/ue6TuSiKxCustdUb6807lx
Y2RNFd6vLe68ey+vYO1fYrq1oM4xi6WkQFN0G97IFhH70Wv+QBLMrmROaCQp1hFR
K5o3vP7Sv5SB7Shf0JbMQWCgnQrJl3HFnaXyJaePWDTcrwm0tM03KpDbVHcqcKrh
56kKIPv0cxD+5JDqlLhqSnSz/I+yH6X86Zsz6lEA51UZE675nss0xy6HoaiMHkjO
IJ8inEMvp06de364zprnvsEf79eh/wqgBtejf7cwjZG1G4hHrK+fovELmh4Xyqfs
h5jQxzXf1njJSfV7ahwZM+HIffFH/DxDXBoY4b8KKA2KfLUIPhaP02Qacfj08hfK
wZw70i0hGkKh4asptqqfb3Mi6lgrfD2p+I6TVznKqftREdjsFJ6KF2IDrv85LwP8
Nn5ZdhghtRxMnkAdaLMkjGKc/orlBc0WAb0f3j6vvyt/PevVN/Qb2RBGEq/jkDW7
Gt1WB4ziOF3NpqoN9fvJn5021zU09QulGJqhoI8Tk1WfkZeHCK8hgOJQllYC5liZ
ISb2GVpllpPKRfKak6JJpWA+mkjJaRcd+lK0XHveWK92VhYkzEa5Pin/IUie/YLt
YZa3cI7vYMzS/g6ZLfcH1nJdW8Uc6DqGc0w6WEmtUKCctk9Fu1nqGUgra0PqRcd2
S5P51YQtGfAGP1irF1RE0C5qGvZ8zb50tpEBnWscI1ekHtVxR1cVdworOoPCrScn
MM4vjoDRx2oqXe2Nc+YfGqafL1MvA4WtlpU2iKTo4jAfUAnjnY3BJyoMCpsqReNH
L3pSzFzdJ5WFhAgsYBcggRdevzE69WhKdHKGFu1Z5HClno1MiKkKk3ylqzk7hyd3
+JNnPwNVbuaI3KAHBPh5FRmlgIXer0sSlCHppyEQApX/hL7AJ3hLbI+ZL2y9zCu8
cjKu168wRTlA5QriR/2xmUbVqeUeoyyAo0VarPmOB4YuXY+HObZIaIY9zYX/ZwTA
0Gqop9aPiqKL9DKRjnlTtC5YZvNCoRCx6ieIqiVkalnrTpHduBH5/lz+2WOe/rQt
Lptfr1i9ZYA3bfN+mUbilb/n8S5v9TjL8eHaqD5u8W6p0egin6LJoHWQaEw6GTGL
H+2PPCFr+HzFk+jsvFiTCM+t+JsypBsydrobCnZyhm2jczvdp0JSiHWG2XX5T9EN
rJVv5YGNu+Uew9aYV7WsvTiIAv5ytCO/ye2L2v2mzCUDBkt4+jayPlgqdCHsDsOA
kSO284d8+diCJ/J8SyYuG2tSJYrx/lbasPUJ4GNA2898/TZ4qkrJdfcbXjo8zbeW
xuDB4yj6UlqnP2ddb+QbJ1eDHIshYZDvdupDGrTMXQhBUC+VGnkN1CsaLQY6Q6Wd
Xw4kMl3UU8+9FUOYk2N3Vm1UH6BHd+9t3XUPjr4d00ZZT4BJ2NxZPLfqGscJM/lH
RntuwX+MixwBYGZcw/OC5b20w7DJOjdhnIN/eCTr3wV6x7n8aJwSs1HYbRqpiKf8
Vb6yHWlV+WbO8mLE098LH4bYcBqoa7/0F9H9pgvq5067bOJxJ914O6mqoKx1c2KY
FXdriBtpBaiRy8gYogIX7T++nmbRuKwujmsYYnQ6LhXI1gvDMQOqjiGOyGu9dVXf
mNNTHREoMoUGcKc2vCZx7WLEaaJLc+5fFIBtBT3TAsc2sYvlIgs2WBpXFeer97x1
Y52lYEgzh69V3RU1ylFcnuSsIxNrKS6UyHFWPA5tEWysVtn1Fq+GlJzifVMxjbPy
TyS/Ew47I7fp606qykCTdS44Y2MtQMa+n4knbKX6gVsymu7XNwuEI7LPUSycy8uq
nxei0knYFD+Aiw66ozM5ea/9rjfsEi4KsKumZ3qAqzKSOolC5fqKxJMkuzI+tJYU
W6vuQZeMARus5JnSB7reeXeEPiurliTVQK/7c6jvlp/P647CYWKEM6braqxZMBiu
eAg6h7vbn/NJBPezGpIuov1bN4SP4aL52XeT032qu8OQCGpqbmnf2H2ThlT6F4p7
vkL/rYz/jDdZcG7CE/RhCYKCcHk6Lez9dEvPGK2Ytt7jKKbrUoMjQ43A3zU9jl3H
C6jnBNO4JzIxfyZ2emSEzvSQ5fRW37/dq/+iqZEjUDgT6VZ/ysVvkTOafG25S2FV
qEjRkB6klbjw6xMdqPAqz1u/7PKaYnfdsr3fFJfKN4lGGAcD7pzhd8I61QXRycEu
aAEbkWTJFSDk8pxCSJRzW+meUUvdZlpMXDSlnknqJOgBo89gh1byDtrwAt8QgS9t
HluvKbGuI/6QcqSxT5thIjoQWsy5S2hcjUM60CJhe75wTPNWZEBfj0uk1uaoTNsw
+qAzHpTn+rLJKhMx5yNlLrO2QyI0OICq/D1MH9Q439lVSEVFHZ0CvQDwox9mdYO3
ItuN9J1KpspzGfeHxqQRShfiPJwiPI+0Bs/vL6HLXaGQzTMQGdeLKLiLuJxapcJd
vD2Cub6I3YG5vsaeBVGkzUME/FNV/l5j5bSpqHXPQqkaH0G0a380zNvt5s4JnsHU
KCXxuA+UHmd2Zmmv6tn/qzbiO32kLBxygt68BL4FFx1X7c/2O7Hzp6nFHWGvUqOS
AhhcMP44Gp7zWqOezetE84rVX3zCOjNcZcj6+W8j55kowiBBXujQXPrU0EUpCwyA
3rEEw7HRuFYa8v1ML1sqGB5ikKaYtVbRSXNriBE4k0GZqhO65LbbcwpWv7A26fOo
Iy/x2I7c9+5PGGwjfDsmKvAoftyibBW0pN2O/s1ohKdsl/SlSHNAjS+RpqGPPoEo
PO7c2obl3+atq/ng+YQdDL1jgW6ohWSEWOmaCCrj9IyUy1fAO8PQV4vo2UUiA0Ls
3slb8mdmhbiVyy3uk+hPbneNyh0vXqj7tHLvXTkhonFNZmKPx5MJve+dQVsJqCKw
bjuEdNXaaGO8kR4z836aJDVwJB+RR59iOiJvp4dYRC0juTsF2Kiksu4nau5weMu7
v3JhE7YgRJOE3egB0EAP6HzfpVgpLgR0Ph2R5F0d6YZjo1/1QTHQJGV9Eds3Tp1U
2lDt3H9LvFB20zpViDlb3VLpO1XQ6mY7ArdxHNcEzXk3nwOh+OVObk1W/Iv1Hufm
cZWe9yU+DrXx6X7Ba/DH9jpVYmlgLth3iOsU7am2Q/CnbUs+lXELx0iVzbFtnPgq
/y4vSHVy5vmHYisOwOHlO+JDvMKVDD/b+OaiSK6xci1A3M8l6TY4hCpt3oUjAi3N
W1m+n9lpolC7j3ND5zh7/8YEZyIgH+MdpgO1DuXoVO/vjGxiNcAX7jFYYsv4Z0e0
dDaRhp5IRTiQbXNicsIUeJoIBfywtKKBgc9S3CklSdTPyTOdlhGiPW5qH6ozlQ9o
mHFrvRmpKdfwhX8hVDvtA0wH1/iH1rQLs0oXA0Mj02f1lAKxM9Yg/FUA4DusJxHC
/yYRa1Q5YgmFxwJoU7z4hQ1Y27v+xKuLoA/cmxndMh1XhM63jMSPvjyaMxtkMwC9
l9aEiKVwHHvLPVuQhZieHqds9zjmvaqZ996vL+0RaawZX/df5ZdMFEJNpGJEdWOZ
xkkH9LSJaTJeWDoFnkqgKSQQNq/kz+TXMtzMFpoUpjpIUFUjvQ+HlVG16SyUT6ew
+JbD4dE/EYoxLfsvvl56kyjp/JTBxAq6aW4wfKhYuPbNxFuaW6BRKBFoUYhOSmbg
mSK1PWJN0JCBCMkXFCljGph7gOxQAfYZnew4SZ38JQtir2CKUUqez1ADnCgTtOX5
DWBDS72CN9BbjBtKMOSleOKWkz0ERrCyHgWxsc35gF1cOETPX6p/AHHwFyjsOedy
VJ4Tl8444QmShhExK43ycwMkLauy+k7BZr2mOVNEcpESYkhJegE22IUC3vG5oR69
6DubTn7WSCkfgtTjWyP5CdSgGKoOOP18Se91eqfUBdg1OB0R6yupNIZv3UuXleit
VFwBDDZTWtZHfnuyOs5LOlOz5MgKwf7C5HsLm545D/FzVvk/jKE6urtcPRZ2QJRW
Br1u8a4oSqHR88q5Xm9bA2WKjfXnea9Av24n9QuYYaQp59A5wxF67ZgJd0fQPuR+
PJL4l4DeaXv8H/Kv/JqVGYw4btiEP3XUBePV3msYIeIgccF+QC603jfKV3euLExV
J9HM+6f4CEgRYPNSjuoB13TZ9wpsRBza99pjG0r4HhCj2n/cioG/Tw9qRNsy++KT
xDaO++MCEk2+SSCBhKI1bJ5P+jzKV6MsXrYvOxtCfbS8hNIZdqUXdmvYAaXxLkNb
eL7SNr/PsblKf9ce3YykvHerG/QP+w4mnOlqW4iUshCjZXw46goQLEblWXI5AEU4
BSxC+eon/Jk+Gl7NUHkONX0KIaSXl6GJFPBW+D1H9Iq1zVcHiC3F1Dcio18vd87q
Qota1cW21d6vKYexk4fZ+NaaIRF3dgaf/M/v9DTHqVgjNRax/DJ8eB2BAtae//pr
b3CSaamPCvGzWa+EZIamvAYCQ4F15ahPFNtpVkYaD5/7wxV1GTaLnFQ6gO2xGpS3
QK46fi8ikCS2Jn3Oh6UsoijpapMuaKZTduOWGx8bWfV4uP6YpASIaCMxW3/bgdWx
RGVurSQh9nzN6zGAs8fwWGjqwrfH3YwWDUUXX+MRewpfsObZ83b11GTu8o4Y1mce
e6THXS49i/dx12z8t94dZNztWcbSIO3wCos9/66jCkrkhS/vWbjw5rW9Mk8ndO8Y
dU/u/4IfiabxeSU0DkdmDXOknGDy9aGF4JPVXhsvD0Y+nq/jyKHRfHJ3gCFuwL8I
nd0SEzSCgLrgMjS/W8/OdHLKKRVhzwDLbK1fhPfo87zPVvYit/gbRI95WIN9P/je
pr/dpIei3f3DqauyoqKmwBKyhww/ScGW7ELXxZdUm5QlswvWD2AYFrGr7DgGHZ3y
unK11r54j+3qRUx116EbvDilHSkmdS+m6McN6+wnYd30PvfiVqO1xd4YdUyMlfXq
UM9oFl2QT19Dc878ElEpu0MS/dhxu5/BPEe2R/QU81Cp3YZHgUjE4uhq1ODOcS2F
sIWPreO/k6qc/aaw70jJxCwbFA6pWm7aBD0TuVob8A7jv45D4kHGu5DmBrHqvs86
X/un7IcUrfvMjoj0+tA3vvmIrcMQ1hZ9z9Za1Sje8ft+o7onj55dP1T1hhP2IAMp
a/PQxONqO9e/nPnalbC+joRfdpbD1hFnhbtJq4/Tu+xvOrACzeocHlIcRerh317V
aYv412Zac80+k+NdeZ/KeL9i2oYLauvf7ug/+SDuqE1MmPRqohui+ybGbZygP66H
f19u0dSsa7Hn5ATOB9/EbTtCx5YSjn1d4GV/LQ0bEcEEKXA7d6mTiznFTJrIgX/l
wVcqoR6kyKFQq4Sdy9s3XDhXV6+SmAeJw2Y9TUFIPmHvu2GySnArpU0dA8tOwbAX
Ru7c8YT/aa/+nDw2/EXsJVluInS6VPKiWgJpkWaFG79VnB54xI6H5+se1PVMWVMb
7ZkU7nCX8rFqmWy0XrcLwB5X6FePIQ+hEfbzVVz5zZswO7/GXtJMnWqweYcW68+M
mG5J+hWrW6JUgV7ErdxjYklFX0+Iu1Y+yH4V95wOjhFjW8cswVifano8JgAJr65M
Q05PYIpEdJnoZxfOny3eq+yHVUwkwumxbdbOhvL6OJaqFFPZDM1rLoluty2UF8GP
l6iWoE6AqlhQ0OHkPeS4ra15Uy+xukF59sFol845RPVMLfXFxDofOaTXpPs3cQQZ
O6BvdrVU5NeVC/amF6FXf9GrM75NIuyFdhimXum0b+3MC038y6x3KJkFgAPmfFUE
m3rknmmIXN0vd3zK2yTdgP7S56FkdAG7Hif62jf2hxVfopwXnlt+xpXn5llvGDCa
SsUDOl1f0pWL9Qi0pOr3zQ1/hpIGY71BVpp+gQ1CvvstGJX308G1Ny3SGUmGFJ93
cSaxRz1kxJ3AML1WWDPfe5wGjcbP28Cj5TsrY8C98XwcdEC4CeHYdGGrkVqCAzlh
Ltvi2Sxxc/dhkMSPLqKNg5xDSL8n/opLnMs8vDYaCuQAs8bzJ3Liwl4i+U+4S9P+
UOLPhIDkfnnn8vCp/lXpQh6jGDbcvseio6gECv1ZR3py63F6WI4n8vL1E/l2pEfb
5U3Fr3wk0BIQlwQGlBa/fDnEVYutlc5C/rp4jUu+Zzg+B6CV7+7YWMdXyh0dxRl+
XU+zM1uDlJTKRNhtu1Twp/QvXN53B7f6lP8isa/kY7suh7k93vjwdY1HdPHOvu5y
yveZqQ0l9yCRLuxJ+/lejXgA5MpTMEcJTXiwzvozjwIBN9zGQ1Y04MrKm99y0PrR
1APsvqvWSsXqiZFmIud7a0KBuC8t+PGSxPPFsMIuIC1wwxl5aCggOu++zSeq/rHT
E4ABWYgf/eXdSJ6zcCiGDF6vn01oLc0NKlKJQMcjcM/FC1daiAlzCkz+gxR5CclL
RdmeFP56MOx506xib2mzhhQW2Z6PEqwO3X40h827Ir01CznlggPdRNDjTsSFJn6o
fJnWqC112fUStto+LnWqDgRPYcNrqIhKL6Slk/W9aPs837keoAJQMxsaaHqXOar4
471P1zCiX8ThOkwzVWZYqywok0aD6ib4vcle2aUpcokPDOwcy4WVNJcxQ+2FMzBr
bMiDp90Q0+SRDaL7Zpe3OuMegz/1HQMFi7gePsfvTIg4GgNP+3xh4sFjTzYGYfrT
xBCqSvlweLWRPnwdVhvZbAY3YFvTdOgX5n3PbKWG5/0uhXf4i21YZy1tjofTc4Om
xMBBquzlR1pZJ2u+4kob+OY953aQIKFnlWlIY4A5Hkij2cGG/r4B5F01xNAeTmbx
fXuYNpahAutH7spsYTRF9gKKcLKQUsI/r9uEFwPPYu0U9TsCI5OM/AXzKu0eJZbR
OfvXSxUnBs/Hh3iHGD7cwnP8gSk78C7LnxM2MmFv/NmAzyrJU9Gdwm8wABvWjcs8
4jEjxk/e22Wnlep88wjCoJjWXo2w0F5ILYCB+3QHnuDeOug2nsB6C+qIVoa/21wj
63jh0w1y4uR9IkwnKl+F5TCd5iqAEr2ph0JPAA2PG/t0XPSti8ZNx95UkhlEdqkt
L/hvGiKq39tr5n472ae2b5vymsbbkA/snmq/sYV86FWPJSmGR6vyOBMsCYcymohW
BdrDBkPfH9VHMgwAja8f3/ArOiPtob9gwFOTt+MwKTo3SBWQPJZuRwTHqnKXX2dl
8Ew9CpAgylwjAnN4S3e4/D/THna+doQmxEAWboTBi+tZii+XqmUdxk0MmA72aDSH
uI1GdPG8R8qFx4k274mtjzcDSw1KsCeaBPCfbvjJW4l3OfMrXDWgYBs9kf5uxaEQ
IOlDz7HIVcU8CMC4/5HmHnBAo07Jxwlph2S7CIMGwQxN03dky3JEGtOViTxRkcws
dMbbX5ZN2tC6V6KecfAmt7SebciYes3eeAtKadJ1kLy/eAP5h5EZ+meMNFQZNeeC
Kr/zdCnrn/aSjx9KY3dg5DNWz7CNkUSwbUlnPsp6RLGPZKKwWH584EbU6oP3qy9J
9UpQO4kuEVlMfaGV3UDgO0+QpuabhuMKzTDdTLcM/uKXXuz43/xOSWCPlSmSQF6e
cdoMKSIM5aPg+03EKzkfVcW82dZR4yj1IVoMTuTmu3GoRGIQjrs79IdRVYA18O74
XIRb/C2mDxzieHD5iWGChm8Lq7p1eYg/v4qFwvSFXWrabXdgIv2jVYKbcIq9eTJE
yklcRU6caYdzGGO7CfpaRXAMIe0U47Ecsa8o7AshWN/yiiGSY4/ZsCRd9BYQ7EE+
dgQC773HDRytQShB9USJOTfH+06ibsvzm90rAIu6cAmk5Kya+414I5/WfNXqshAL
QdgYB0g42ssF9sSBc5UryZkIl2jFdfo0QkLsuKCEML1emOR5Vq2bf7m8jGTkPwp1
U7zu7oT1Y8cflhOL5M0UeyyABQFMtXzUrV5AfMQC1H1zIPkpy1XKtTGppWWZASmJ
CsMoafLEaSRGO6PgPxW+OYa7jBSEAINhTC8JXWRG5d6dOFPH4zf84lCqB+s1h2Lz
bp3NmpqbS36bivi1/yFIZaR7H6N30jg69JWkEBDdlbWI74bj/tZcuLe10Wtwl44i
j7uMb/XsZ42KJLRT8+pc0ITDgJeBpoHicNbWat8K0/FIuxkgr02TEh5PqViYqR8Y
3LfImRpICeeFqeyga7pG+OGkFep/jXk/OPcZ8Qfla4r8NvDnuAEuwxVdzn93C1s4
OMAwhtTa3BQ0BciQSPLLDK4aFjULvc9zcx8FkTmLOMwJ+2OuGnaOyPANIM/NkUPL
hTV8gwA5FdwpeeZfiDf6gpkctnbbgeICwGfjmAd48bmp09pt4favbl9+scba6Jib
HI9rxeqOTroEWlJSeR5lN/6iLH41jcfZcKBp/FciGU7NN5xHsZFjmURTF7J6Awt1
Ve8M5FQmxkRztvD5BvxpX07v5BWy/hmBwLJbFVauuGNuRDlYmPg6WToK2qg/o0t1
9Yn4yLkN2+IQUk508JOnuXe+tSJvLN2JYfu2ipeV/BH8yp7jR790eNgu0XsYUHQ4
vRgB82W2Fh9CiRYxeGbH5VoCmmL1Q8S+eqE+nsgXHri9jke+SK/PQ9pRSOdZbyjG
rLtM92ew00OUWDBCFOkoFd8aVTZP4vi1/0NOS5zWE9LtSM8Mu5Nqrmo5BlsAFVlO
W3c6iB7kKyYLh38sinBZL/Ts6x+3hn4mERdhk69Mty9r9iAsHSikssRo56eVQs6O
ozlMru0aEVjYqvF75uvbfEDepwkiorkrjCrJrfWLxatc5ZjojkfJgvGOTGNwgFNH
zjq6ERUlJrRQq6r9u+P/He/2Do1MthqYsYLgOrKUA3+gzu+++E0dpe3YftPLQk2/
fxONPG9FzTSJKmODXj7hcOjHRQl8ankMRugfyHsAW3v+qKNuguzHA79Y+pRPUHBH
Tq13KYm/ZY9PaqW/kn/cySQ9L2u3SZw7HDxw44S769AZwNrU1BsbRCELRPWYofl3
gAcbcIPQ4GM8iry4uMXZEV3dmqQhBwQDaBWZKyra1rLN/cSrLBYPBOfNfxHcn5TK
+ETmcd3RQl4gK/7SQq7ZJn+Rjr3Q2/8gGCQCR1NIN9gBNO6kiz+CZ8lmTW3HrUxQ
6qjO1h/G0ZQdwRN8oKb58ZeBmtDyW8+SDDp9H2q/8rvZIP2OoMAYdZnk9Mxk/IIe
C36JtKXamHOBizleh8rRTwZ2HAjkcIk3/RtW7QGfehYMa1ZKNYcN2FS/wdVGFDpR
3dtIwd4pMBpK6JL0OzQf+Ci2sKYExiSvDgsr6fgVhCKfQkBInANJyahpkiVSvUeS
vBtFEK/nXs66WWJ8kVb9JmgZCwKlCuS3hH1lir3KAPK3hyvMEz4SnbiQ+EsE1Vd/
wF3D88A/nR/Mmh/QhCM4JZIXR62KH1EVKYzejltIOIrwxwU8v4A2kRRDwkYl55U4
lSEFSFOA8Hzwp8XqPkPj/eXact0MbYrjSpd/xADWPA5HU3Vy+afg3foJ4KfIJk+p
NILJxygqTI4OYONize9lRdPL6+CLG8b6l74XwCf9cCrlgvE8IAh+UAN9+zFxlbpG
k+yHc6wJ6o4tynF1YQBrqeLqmpVOtJeZ21qupPCLVNGT3OVSuvByLkiLG6iaE7Mv
jfs0xlB7L39kgitB2lPuURwdRc+H39GxK0GzrwfDHQU/IUfHO3zh7pE1l/mIoSoV
dhurDIInTaJx7ySEEE571/5ZVMkvtB64Rg1UKlLM5ryklgtdrzKfkX3FC2gITS/b
5TtyYJmGegfUcqwPBHyH+ddUFwlRTFzrubApauf/ZoSCtk11AkDXDxz8PPMQOMR8
05m800F8FT3qRSoxHdXJloyPaUGWlp0LNkTLHJhmpcsQhTEFcFlmYtKUG2+Bjq+b
iquFQujNV+oKrWuU3UrxaoZOpGM/J3R3/54i6epx5lO6NuwidOS1XInJyB0p1FYP
jKk/EIZCocz/sbJ+TwF4KTP5QgHvTlcdz7oXHlCpzK8GQxFGGqY7oUTkA7ukae0l
I2FVnNjc8Bmhh1rd1QtUYvFSJpd/vG4IUU9tSA6QzGCVAVeelPBW8z5bhWp23jAo
ORdnENOBRht54L2AU5L0bYCIQYf86fPeNthwfuvjHDH7/sIzcqNeUr0HtBl1xD4R
9sVaH3gZAxd2upwsNBy9PkwtK9k1COF3gkrJGutTDViOmDHwJxlNjDOZrXJXkVH/
m86gMwdyZPjIlOQuZu2zE2iQBCznvYH2/yHvOYVxAIMaUqXFotAJUltkKbS7L0JA
/2X3PYhJXPY5OUt7Xhx9mzzICkDJGfZ10RmRSZBbhSgPDujPX0U1RQRYEBHVdUtm
qm7nTMDwATBqEuoI9yxEVFXI96jzCjDSboU7eVuZKAndQrY7qkP2u5mMWbRfHJ4M
6qYjTM7IQzfDnfXKsgLfvM1e0DIAiRdHQmmO2cadm71zMn7QsyB28crBvUk4kPna
tkRwyuEt9HUtuRyHO5HwXd08l/9mMaUnIPrGQ+5wSQwSw2Xjpz5rQEo2HB/U4ECW
s5ttKXUmy9YYC46z4djyWs00ML/BQ4GNC+wc54JPIe3IQDQpxiCczEGk+U8G+rdx
xjFX+jxcq9n1naOo5o87vMRGYs7YGyAnQH7iKK2Q0Cl61GpwIVPNQL/pzYZ3pN0P
AcWowrBvO74/8Mxjlnjkapbl3pQoUpX7KzfNj6sSd5gcLtUFpQ0680gkNfBrm89z
nN44pqms+843XcbeXfrkOAqZParhXjYI/U+Qj/nSFnJgJc91+FCo6CQJwBF8z3V8
1siJdfnd9didIk9qttccz+pYJ7BJaKZ28ydtQ4r/CJ0bC4OOhYyJbnxv0Zk8dUZp
V/tm6znce+WbjCyLtyYmdnMS44TmTvNiwTWlJrZogPkZ8fnSRi+yn7EKGZ07qTo7
zrabdjzl70qFcYeAZFFyqn+xKJqqa+v2e/UwgyMfIxLk7ubDUt1mevCB4p66StGH
IQKqW80JHfxbOsCyXJ7RqJpCRQzKSIokjKKSd/PtdLzsMMIYzmkfExrQXpATVhFr
2X3g3uDCwLeoEB0ijPBsoURotZcJczXj7usLCLO/I2BL1YunkwXqIB7BXRkQHW4V
LLJVF4V/fcpHoT1X158XkzfAcKLZHVeiNgMKE7Y8M06gon4iORLL9ige1MKET5Px
AA31M4six9mVdkQ/5HkpqR2gAe+WDo1afQBVXdx/MBBL19MfR4Ozc/vvq1pzJRgM
LBiQVwL532MRRf5YaYmoYsFDLoYyJ2YJ5gHHO9FaQxiPpUQAR2WM+Rgd3ZHizRKs
mjXFKPL2d8czFjr5qJYzBwYRFbMZlzX+xJPXCnRW3rmD9sl0wLYZ0x6YSUb9DDvE
sgELVZZ+fXy0bD60INl3ZYIBDHqkbiAFyjjwxBNLS7+Imy2HAupN8rcoTx3xzPBb
1jEi4ZMYwb1ihHn9EgXFrnW9rb8R78D1zPikJ6LDdeBsnxh1pGbQ0vBxpY6mJ5am
NP7cn33Ntvc5H0T/0TrMAR2s5OyNR/XVN2DBH1VC9bRWTi/RTKrmnF0kblshqWLY
FxisagGBHE14rY8zOI7D2thCMJfwl4IONrSuTyZ0MGfS1llm2Exlx7AChSHHPrGg
UQMS5MgXHH36EyJrGavv0uJv57eW08UIuHi59vE4PJLlOygBVbqCTTn1DyLhXfYl
E9gEnd/Gqlioe+Ny1/KuxTEDIuEBXkQh4llteDc8AJDc6gyhH5z5o/qyBNM9NgUQ
kXNJabRAMWG8sZfU03Oxl35omjijbuSGJZiS5R8RhJwT5JOfnCEBMyP1o9U0E5W9
MMghY4rX/Wb+06JpOwB0zJC8CtJUwXNYmL6mQswcUkXcuqNH+HJokSBJ+f7GKSGn
xIbfAFfSZX6ppN18zZ5lywLTtuIh5q0w6bxVfH0wGHG7URcdpoJQgIqeUHyKJVAC
cq0aEhEEHDg+w0J8XFr916UN7RUguv/3/zK4i9H1W4HNxiaHS2d83o+S2+TtsweQ
VN8E8zkuEAA+IHVb0JgldP2C/6Rw2ooyjQM7OW6v+4cVO9+owovNCOngZp49UA72
gYFL0JrNxYMM6UwWr0YZ1p32NKGGUy8avGNImcCdSSma2/lAEqb9jZ55xg3jgYDW
OEq0grX1Xp5XT4y/Fh1CnPSJ+cNLHmSaqlCxu7cJIea0cu/+HpZ5gi47ebU6Q3pj
0VfhZPHv1pHrdhnt3XgdkKHo1qtgv9hCNS+NxG+POGMke4mcabI2AJiM5HpRM3oe
lcTFxJbBkPoh/xHm2sSvtbY61i5jXF1EeChYjrohPC3T9UQ2p33hIEAPv0s1pBMv
iQ7pfwnXnoDIeXPt0vNtLtr50XhQpAJwG+3LP1Nw8flJAYXiqdSJ1c0Q7Wj98PjU
5cRojfJcRfwU1Jj9JrUgGmRxy2N8lvZRHa/eNM8Kmqf+mOAC0lJfFOE+82e5Died
jwLhKlvZcS4ldDfjNdL5QitHD8CEl0i2j7U1J3d9+1TH2oDA8+TQMYIXEdNObju0
Ce1GZCItYHZXvOfp8GLVsjDlbfFWsPZFnIUmlGK17ShkwFdup1oIbP6ElCHxwfDu
N1H1PDiSbXRTLsZ/baMgBXfbq0dH8VplIvF/F/v2Vf0NROyozIX0bre4ZOkBm/QQ
kqjyvX+uCvP3QaW0whMlGBHq0pj6dXctKo3m0vzbDMuUmqkXRlkxH0TW9gmeUkmH
l0x56utmt0vWRE+gMIOFqMpoTf7/gZ7CBNnOBIlhmHnMXKmaaiw/xBIVqD0g3EJa
r2YqfjnNpU7BjDXqjYcNEuwHkx/bAilLUp4VUZxmfeKU114LbLjZ4zMdV0dRertq
mV6ftqQ376sF4zgDtqWKBbeqSjHH7R+f7DOd4w32BoN9BeRsbLR1KdXcp+nrblAd
vdK92WJ97pFadrpJhSy9PkLFBTbno+oZE2ZIcO1rxtCP3wjY+ePTVxnIImSjdNE5
g1sFoIjkpkQvuYfAH9twPo0O3r/yVjXZeKj5yroafQqRBNO/XECwyzMLdeGnXJNN
tq2n/bFdRMu4t8qvWQsxRWLTAhWz0+PpQ53EwB82Oeal5GIN3F2jf2TTpGv+ujie
zAAPfJQzOYgc4jZn0/L+f3E7ndDkuyuCRDMBC1QsTHPY7XzxW637/b6+aTfZxS64
A0nQoW8oaNoBK3l2IXmvCvP42+D3nVvax2HT6IxiiguaGZ/UsAGsvcpI6gS6/IFo
mo93IKSrQRpzASY+pUPyXhEA2rWnPDTFa5zrv4I8o9zWocC3IbZIzgIEQ9E6AdlA
mM9pOj9bHOP2fTjUtrjY9R1ASG6Qvy+1m2+90reRsoxtje6Hk91tWrLzrjh2/tlf
knpIhh7vxjMVl1oPOu+0v10kr6p6nwtuFQPluH6U0q+t8rTUDsV62mlbLDa2K8Vj
y4ZaJ5g2ZZsKQEPPvVsEXlcQKyrgCSFpwWJiplZb5j1sdOttrXX0Yc5vWDI1jUf7
Of0QU6/CZLiJ6e0z+i3aHmjnnVXsOamdVfme/sZcvbVXoiBqvPaNHPl4HBWr65Ft
Bax9YPbrMLHrU/lD2thkojpC2hS0CaIK8fus1Ny54c1o+EhSmA9Nndrn4s6dTtjx
IRAkxOcMzTfCl2yYXXVrksHSw1BR1WljWz0y2UGesVcxBAhPVjp4oznWj/cf9i2R
fMeX/KkCP0c68XZJK4QyrI55S8eZmdjwLlH7goycHeu7TzVtFszw4WuMJUNQkZF0
t6Rl/dMo2f0En3wEHIxH2ndOnHiAKhnqs9OiWxz9HWlnYDk1J8H9MLI1BpDI2JRE
pmwO98coImnlwBwNjVsHgVhrz/+oP7iVDJMQ504eU4kPNE/QGGzXp1G9Cxu887Su
qINdp+3u1nIlXCuCoRoaT2I8ScHwBVU+cF1+iw+ZrOAYzGQo5mMh6py0pORTZJid
ctJRDYdT5mfY+yRIQcPtsF+BByLXQIcHktkmcX9joz6gFrzxe2DB5FREhUlX5CuC
eHmIKhLkArwQ1owsvcBhJJhgMkFjmdcMAgboyqxX7plQQ9jsj8P3OnvDWmZkh/1p
/2RXbZ2yxDq6fuO1LQ9JxzgBoN37wkvm3zw0Kz4ybiyvozDegd+O8AYFz/z9nnUk
klPNwdftS85Nv9oeC+26x4YvkxFspY5BgKKKqnde7zB3elfrNZW2VGHG5fAfhFmn
4VWQDicE5T/Wj+0v3I8ULfUQq0nnpf+lKqeeqUIXqiWvr1WdrkW6n6xuY9Rqy1Uh
xClRXpQgUF0sGiTH80pMieJRuLjlYzbMoh/YYIOysH1uDu1N2yx3BGuSWpg/1+T5
3AgWKiy042f07WD4iItp/fP8bJnsHu5883Ds91N49ZlTLwdB2O0Wk03Izd6tMvRP
FKkWkuBdSlaRfUqqG0lTgUj2806/Vrxb2jvSABPuYABhK9Z75wH71/6HSvQ7Xeub
7o4QV4+FyBO60aMQqOuqQCHiWiQ+tiZHBByKKUeY+IIPlXo537Bcw7EvD/ZPHYnS
fj+Bgs2cBSUlbsHKunqb1i4xRsQdRHwTwyQM7AO+ZH6gSF/nQb38tnssd/HaOqfE
s+Lh/i8biTcuz4SAp+aHMQiz7y3CLlMsGqSMVckGyqbyWyU2rGZSpd+Hm+nHHKaF
GD/JokpknWUM7IZzA4XBf6+IQAE517NGTKeC7nM/XjkGrCXM8bRrMjtE3NBf/fNb
QS6iDg2cWncWUD8V0yg3795Iyz2FJxR78XAu7mdRaPnmYN24gM5F9VBdxdiLbjMi
3MetUHJwzY+jSrgSXpN7XEpIkkVElfnJDAboSvNmsUikMV2dX+GCOGvvwXKUNrR3
GwkKUzPn2nJ726Zi9kyGFDb3QENpp2YIB8dx8G+gGnzgKleNH6bhrk4bSANS08zq
rGXK11e3lfaYg8UpVio3oa/+/xzEkxqzqFUXA78VrFDslPXStl8gyBRxNehWIDt7
NlSAjb1YE4ek09UG0JIR31L8Owna4oocPHotp9Jr563LNknOcQPijqgPe3PJKXMk
lz4c9FbxV4ng9mw97OooZQntgesD+sonbtcWV/vIKyAhr8EFmHPY8ygC9SomcCVx
N6BXkQ0YQzWwZ34ZrKLX2Vrqo2SLxiFZJYz2sf4PANK6qyPjVsw+NBoGPSDlU8Zf
NvmKoUpFmsDBwXU+4nwKjgo03FZItBDPJMnulEP1QjH9JuzSJLO2Q9y+xWDIs4DC
tlrPp/tMnMQ+wqw1pZGBfk5GitYZsOgGbzwvTDd5rL04jwBgSBk/JexsY9vs/3JO
A9pzYB7pbpDR1usalGCTjMlgNLWtbxoPNiR0n/Hv55gn4O6wPCmRE5N+t1R/2RD0
GSc0470kWATMCivEZKTzqJ0XtcZ4SniWvShmhSwRTRCSFLtA93Z2lZps0AsGXIk8
8x2oSrOFayluZ7tvT2vRvE4Q1Z34F2v9iSjw24eHzeS5a3zyQJvPNbCqHxjAmPI4
NCl5+NZ7V7GwZVmmUtF2sp3z+37d2Pv+mSlhqBxirbiNuQMoMJuuV09rHb4aIbMp
sFjvpo2nwYaDMBk0OD34w7pKOlR+NRS8E3r7zty3Pw377MuDyWke4cXZ99S2sQvM
2F47x6PDiKQGAqQ1TTF2SUNU26QE6aaUDikWkv+a7OywfSZURuoQStzOo2jvY70Z
Sy0UApSsGF3ZtUMTmmT9F9rfRbXknGI3/2H4wqxE0gt/8Gs9reb0VJlfqcgrOYwh
gj8dSlP85lwKsjvv3tra1yTA7qDzEadFIGWVJ2LPT3DX+N9B4n13antWBaPVWkPD
3W+Ox4bX5MtdZ+ygc8u6BuYEuDdBCauJhrPD+pg6b2oTnbgGTjLrw/Fyplk5D+tT
PJ+46L3KCeMepcyTZf8ykDM0izc/2JmJ7iCZMxgzHRBfd8tQAUSG7+eq6o5OuxPx
6LKoa2Ps4hIQFYkillk3sx+ncfipU2/PS866jReDAEVcLaZnIHoHpSJwk6b2CegF
EooX9Z3tiku696oPTZ5CmgdyAOeSuAlibpdo6FH0e0DWY745xd69Z8fDJvjX7+Xr
FaIJYyzu2oMdOLYUrh64QpfjOlgSyaCukjyMek/J03ZjKBkCevpslEm423L0XnAo
kSI1OspQPD0y+DYzP0dN7WzKGhy5gR4iLUX4jaU8krOwpCriEXVpnubaUplDVES3
sZiAA5yYaBI1WlfmPhP55b+U4JEQUymNj4mU/3UqTW/KxA+ZdVHZU/arARAV5WKW
oeOSgp+2bTFb4fzANrly0XRHJNspThAPd2IqjCPfHVMfN1J13rw0KEJMrMYp+Aed
VU746+Im3J54dVoKSaTn8SdU+CMqB0jkFlRz1NNekghOyRc8RCGKUKGNLpgLQfEN
SE7tB1EsjvObRsYFbj7sFAqSMjmlqkutXo0tjDhsXhxgPn2660lLIiXy+LSCPTqD
mqThIVWJaB6fZVGqehCxv1Gu1kAwQEHioBSn8z0e2iYRHbwkZMGrmPHW10F+qtQR
pQd4PDPMItOmDwADMewdthMVAQzO5LeEaledKoVtxYMRjtIPTvRJ5lJPSypRFo33
nIh58uhdCwnX6G58dWZt1SRQg5ZQ258ZL9u7OYuQBJreBf6YjkB5lpAnujpUMXOX
CMVoGnUiZLtMOH7DE9mjzmO1QJs6L28Khk2ehQ1k8tGPLE/irksQxmig1E/AQubF
Dn2y8R90ox0QaIchMbLwcRTkh844pgEMMaaR9fMrWJDMOcqunB2bNhOW7oBxTKrD
E0iQ36ORny/FMCxTP4f7uR3ButHzk4mFDdhTXDGumMhjcGouoCBLXqib++3pn0z7
SFVVLa8fZGlojNh48PoX6daFE5ZY0OdeWltPuIGO/BVnZ4MHI1QW2Fa/ELzd1Cvk
3YisYqadYqY2kytV1j54undpjDlMkS/byaLlApaq6Sh5eVAOuf6qiyh7ge5uDV+k
22/SmvgWWA9HZD5CUT/Wq1wivrfUjaZqISF9HhJBDRy2TBuzUQm6d0QDORCKGPd2
0XfOr7Oh2+GFKb0IHH83CBR4shg+10y/z7U34cbNDfG+WSEzAJdGb5jD3x7zvCtD
tP7ehy8/qMZQtgrgq/bpGIOtpL8QukwDvw74wV6TN45PxW+084jnXYyqJ+/KCZDc
rcTk2j8VRdRjv51wkayEozeGEKysdJtlw1xkttrKhj8rUXcdR6DN4u2ofdUI8yci
MSGw/Yleek7Xgr8S1fdTHfh8V1cHHJWZVi66CFVbPqK+VIRU5MpLsADo1Pu37ra5
/LnwFdARpPNcIxzrLId0ujEZ4I+2QRm5d3CKmVp+y0eCH8DyH1PFU+jtbph7MaKz
LJ6Pa+qvQpd22mHaspCDW6dby+LVswqG30etmcX+2RYzrVqD6jfPZGtqnVeQiQJl
AXtzcDzOswTwKZIC2wIPCpyTOrJNFlp1CzsKJOM04UEPt59vKRV/A0SDDl1Ph9PC
qEUOvVTyErKqo0IXiKoPboQMapVUCCHT1Hb1331Jtw3JnMVGrr+bIer/gf+eKbgh
xYuw0trvSQ4zPOKA0334U9TV3u5wMTtUkKYOkHJF83BNmbrJcH19xvlZv8JdAWxE
YyzDUgX/TDqouHPLOforDFidl3/rD5lClstIavDCBqnL5EStCkmi/qYv8CGYR3dN
3L80X94TJ2bow2jRa0ZGdYHQEFhRWREIeYzaP4rn/95qU5cjQnoTQcmzE/60FiVd
+BXX88ivnk5+LZmlBPyPezrvJXmdon6qMSbpqfnbeL5Z6G5JAyje2kFt429/Zrwx
gfQtwaTThzopYN/E9Y4LyUO7xeS9U8KVBMoqfaWFz0C7rsk4MfneCMl1uXQqIOeV
64yyR/ZPh8DhYFLDCO2y6CxMAalOyLZczGDUXPAjGPNB+kPFOfxcj/0BCh6UxlH5
GoJYKgEvvEaZfzZzUeCAvIEAMDuu8nSD4WxTlm3KsvIInnVcpRanGtcL0Jr76FoU
kuz4YrBCSaoL2qPJJ9NU9aKA9uph8jcngy4uCw0gzoycuwtpFMUijasVPNbpHsL6
A68goole1eNNet2fV44WoPH94Tnjmhv1Llkz81rdSgb5gIRgOOAgDLAzEOSEB/0g
VFYzntCfIqVR6DUXN6eb1pTX+HqPAvYsPbTYdDjekdx1+Veo1e/vkkLT9o2V8UcK
/+lk/xLasICqNAWDl/4oaSl/m1WpehPBLU7nNVX3wgeVTf274uZ1qDz1/mKjWXOh
nFQvRO/955IEW4+ESIdnQFzZNMj8dEHmLHI8e7LNAtCJzncfa6zPe9su9pWKJdti
As1GjcNr4Fqi330nZ4gWjy128D/vWjCl74d6xikRKlHOXhhMEkt6QYclMVO5NDq2
mjGaq3ccXX1MNDEWfZSErMCVzP6FUqhEaAkUHkU2XhKktnbi4bfEMCyvkEDWpEEI
1MgqopSLa5O3egRsCu8nnV5WqIOaT4hMQj/jyJfTAtPJzG4/c4TYwcGNjpHiXxs7
3AlAQxJljFnuXiCyxWMW4OTWR77rqrh2ErYdUK8w7sKFzHveed9RD3JqPNRxgz+q
BkKugLCj/OfX5GpVslJ674DqCSsdSwyLjzuHhAaymUI56JX/ceS942jluVM4BmQM
xFJBhp3Qa2GpqFuCplezkinMSxJ7FoU26wH+O95XmvcA7QsqgODcWT5tjo/itYn1
oTzL4TAwqgOa6eLf2mceINYIF6ONEdxzcbRAwfcv6SbGc0Z7zPREnfgnvGGgh6bJ
DDr1EXWwIoVGT8cXKmFs0vaH2H9m5XhhxOoHxwyMJMcQu55BLMv8+bl66aXAyrqA
z2D3o8bB5vcakHGW097ZWO7fPI+ABH/GOpYeRysw0lJSuC+s5LEU7CRXoTkQI2Nr
asMITtdzHOCDWgXOck78o5T64MU8xDMeH567qE5x1JUcPAD9Rjx/qO0IXSGUUGTP
bwEqY0MW2XW9czCkvNoqCazO0IB4x1MsM/ZVz1TUuIDylFPs0bWwWzfF1ykT+Opt
VP7Jki8cxo9j3/d3T3TAXeaJGMLv3K4r3f5NV1fLOhy/1zweic1zLpanAuzQq6YJ
tIfhyr7XhS9DRPbwnwAtaukPPtGwNJ4Db+kzE63agKJoVwb+f69w931/DxSd3vnA
3lwYjwJemRfhQpapVxRlroM8G74oIKtuwRfpV88YaKIW3hx/IS3up9dF55yp2Bp3
a1drt84fe3xOd22fCGomHCbWS4U5Q5hmMsKwdWEB1MWI9U12RsEii+kJ33s36mx3
98q80j5zufJPHf4EANq3dTeD4k5ZIwbxg/ceWeU/n/z1wdLNivmp9KgeN3mTzO8V
w8ZjnSNKf50mhzdpAPgYuXYPnn906tmSEa7MGnoNIpdRuHNuMvCgvFBDYDHBVV9D
S8q8MYKWEzDLhIYg+i55modcri6FfdLhtQLxI7XIR9NwAhyzgrnTRUYhr2phf85m
3MSCyhhrbskqGvJpUjhkahZxDkszDqJ9CDco0OSYOy8er2w9zmFmt/bprQiWKs4W
+LHbska4IH/qEDSqLPBDJj0D6F8H56ji5IBoS2BQeFSKFmi18p4kKW9xNe9WwSGL
A+QYcf96rasD9gfe4orlcLaR9tCk0iHm3xfFG7NXUpq7cggHE36pumyvbvf7iS9G
XkWpSIbhu1YTX7Y0TVLjF8MlGqP9AaOJBavT/UwUa4sRwDlDzT4c99coKurkgqRZ
UWM94TX3NcGluv+WueY6M3nGjfzRIu0gGCwEUSt4KjBPtghMVLXmBOW96j0ujVwp
4EKkbtLLuqXxZYg52oR1Pg9fV66kPmR97RaP7w9sjOSFeIYVevVeNkGv2Hsekijk
NyPvgm0UoK8+bYPIwPNDoWmxOeQDyj1TG+25bc057NAbk1FjDLAxxUMeh/RlMFqy
W+CD8UZ1pyraD+Uz89n2BHZCp1oVmMo7CotL/6IXFDaGIJR4R0RHYFTm5BkiTwfd
bp7rEpBekLxe20u5q41ddNprPXw+35BkWJcj9QM5lnInP/mpZyVhAZ2h0ftPAde0
p6niXSe0IYbUKB8cuotlyBeQxk4FD9fnCRXB4Ulj9EvmMoEmN3I6JVigeC+z9GdJ
ksOuEQuhKRbtlW8tCGm68ZgN6wDQFDhLp6Z2mcmLrxcZiFQTvNJ83ghYXUiF1WLP
7YyDkhL1RAXS8TIEiGRowMSXhjaPOZBKNNFTVhH3dsNJk8B/51scYG1pO19QzH4t
0DIOhhHKpV5fj9JU7b1P+xmakx915cwLJjg0RpDLo6lGl8keH0+grFp6zOStCEAf
1mXG9b8MQ6BLXSoGakPXNmcNI3lKSpjuwz+Lgwzpm6mXgG/SjisRN8CweJInwEsD
VJ5W02cPrQd92u82fQtFpGXjWjpPGBjLi/nkJ5/KiL4kFoFJRv2bmQY0fiYG/zKH
rNrFgOYBD63fY6gp5aps68gh1NlDviki9TUihOcKm51BvcOJxIvZX88mQixCKM3S
IBXJA01acwbB3wbRi9S84mjoUhLr83LL3fVGC2h/P4YojdzAg0Cf975tWDgGUiXo
CaJ5gLszYy1i6Jctp0laJI77SZ6mr23WyveCKRdnuQr7HMz1U7Dr6jrv85w9fS1q
rsEd4gF4iCJnAsZ76qf1Jl1IRJvrmLEYAW8VBHjd/F24RyYAlfUyhVn18sEJPqk+
3MM5gMJA1fZ5h6bEnVs44O1go4N3ExfPNM6x6P/VqGgISS2mn5pGS1+DXX66R35B
6+2Hi9tLu47brFj4AYJezOydJesyC3ciElaVBCSvuBkA0LCmOLBNmGDoOC+zk0ny
9guF4z/YzA8lMI7gLD1JOmBovppAo848M1KZ3rxpjhvDPdwiMT197IOPj4Vp7DsU
TgQDEvfHM3kMFrQQOjU1oMdjfsRyQet1cWLuXjpIbk6L2XHyw4fMCBb1/dnwpamo
09lST+LhOObSo12JVahSWgIeUL3fFakY+9q6EX6AtlEIaWwb/+Oo7kaHKi+KjPWp
QA65IsJcJKwKQXgEkUK+IwEfA5cx9Zv6HjVH+hwlDPx+VVoyxlTPYlZpe5LHTqcL
7hS7p1Zq3vjc6SAwEK1rX6T9BnvoJoWmpuyLegl/ImZIL5ZSotya4svJ7CxHQwfh
4BvubwaHXnU/O8QZZzFdJZIyuOUbdHyxuVhUi7t2hqV+pd/cIT/frVW7R3qxnSey
b6bjX+eyfjqj9AR7vqs7ogVSeEyV6vpKd53yMtyxYQAyyQ2pW25qjVgtvRxJTvZl
jUqWdIeY9SOsUQWXKzFNNDCd7Rp9eG+K7RIPdgp61x9H12flNx8AQkKrxL55vp4B
ZAsBhTo4lqadLlOLOpQHis5PIWQS25ww/luVLMS73br5bAaALyhx2UvFDLDP/3kG
Q2lZd47rmIH87wXvMwB4JAFIVSwxo1nkDvjXL+t1cY6RhcoaWQ3T8Q5J4k+mpqNF
1paq7MyD6ho/aUd9ZdsK8eiuNQ+BlMfgBc/EuqQBzGqWPRZkZNqp3T8/YiaorXNN
JTbJ0uc5ICILi/ux1gkZ4xqQJ2sdpDz1YZ4UWuz/rlzSJFIgLa4KbJtSSFtU48Px
7c2z1F2Uo4XNw+ZM+uZf+pmndpyfHkXNgGGJYJWCyInPamrAScqtr4qYXNrNvpvz
Cc8yKS38Bl31TxOJlWdpXaImSLQStK3beL9ut9dq2aiO0m9gNLCmOxfCrN7ziGOT
X5NQvAEipxm8oVvXhMK6moBmEYneG47QlQ4OV7NQhVyj/sPnQ3yNqHYdX953J63x
9CWzFeEdvt5r70qcwvHwMN684fayp7lmgpalhP+D7fbV7gXz+JeYYJgQgjqtjAXG
UzBJElrQnFo33WUy9T+JwfH75wgiqlaSKl407rht8Ik/839I5x3E4z+VXOC3/UJS
srxP+QmqH0QEHBJaK+7z5XQIBGhpl6OWWnOyPyc0gaR0TCGYm65xWbEsaBNyyOhw
i7iNdURhX2WoGuWx207ak9i1DnA7KiyZzJXIvC075J5z1tR2wIVN2lSPuaC7JfQ0
ujcHsXlHzA2DUzvpey5t1NS/awjpj/6RhgdNwCd1nbr6MupV/74RkQBVbRxsUUXd
Sw4z42G2nFOAA2pMu7bsypKI3N6B1qPyFhx+NYw4r2Exv1m+AcGhael3PgzW47Np
2WMRkWNoydU6jh/AjQLYM6YLT0mFbd8hL1mRAGxgXPkrNZlSOHo/7ADgk3p3VcQl
G9qi1pDUnJrXfq3zvhsQyFdQZFaxKxlv6sYjd1plckol9D2BFjA/A0uE8v0vdyQG
BYNDo3/uymQkN0+XgyMUNlA8dm2bODihpeo2NEG7+JdER3VxazF50NzPIATnmw4o
VhcbtqB+tDLsHB61E4qIBgXb5DeGW6HyJFTQ7F6fRLdyqcpPufnpJS15SuMtWby1
UzRBP0J+fM1TSKPxGhwLmOfWvqUqpEOvslJ+AYB/9/j4LkhuHCu3jcRtpUB5hlpY
kDdOSpgGtLh41tDxMhYwSOCmB20ViVdpPnj3fdDjdnx4RWzuXH5QalTwVqnnprMO
j5nZFH6PySwHlzA4wK/Lm3F1jB+yVRBw1D0rLF0u8j6q7DUV2KBge6I7vovVkzfH
Vro+EXTOhPXZutCQaMbnTzbTzLlM3t/PWzpl/vgr7M3Q28DjwsnKpAUxBP1+52Or
ghdEso2BTRaQC7YBljQ8pd87CgbZmT8g69QkWtLCDlWr8vEP9m21AfQd77IbCP6Y
+As7G35HdK0fAri7j4JaItMKoi5Zx+EzqZ91ayRy/0/Fmt5TtWNW1sglpcCmY7Po
u5X2/DIOqYmPVr9e0sMNEI4kixxhNqB/qlZvPRkYlxYnk4giuDrniGoiNoXipcf1
phVYYCarba/92wHzB9FSMoMgZEK7xpR5rhTbqEgU4mQcAubEjeNAC7Y3W53zl1Mk
NWFFFebqAFmOWhlM3EYaz1WWpoXWAdaDEIdqmgtUjmpKYqabFixzkbnwrTS1bELX
1szPLUv3/sCwUll27Lx3g+qRi556G0IQ4HQpRb6xoupKmcqe07oM+56JxCGT+yGb
7kZybFUXjI7utWUlS3WlHSOPrSJQs672sbHKYeoTpV/zWjJh3ricH9IIaXreuPJp
/FR92eewY6Fl2QiBt87rpayKuttuvWbrqBIDwsNiPTXJOm481E++Mxkq3frhc7DE
rQuHqGo9PyQENnFZT8KMrdqPKVmG8SSIZiYa2W6Gyj/wlhLQg8cPz2vJ6lY/gdVe
RW2jNKkaghp/y+01+FVj44l+n2z5dwmGvTELW1VlOaJ04P3gmkIsrt6qmRr+yXDU
xxGJK83ANXLj6ofl19dk7217+l+27NMU2X7TvFm2x265AWvOEQyAx5GqIuKdRSg/
BVFYp7dfzYbToeznlQujmvc3oaiN8u0OOIr/oeOez69RQWpYWJa95h6gB7XSAaaj
mni7FGE/sqd8Pd/p2tNSk5uQqS0fXmV2/SGHNeI09VeRhQfqCz4CJ9T18sjG8tlF
IwBeXgyEGSnh6MbnCo9LFhB0qqRhepELa9DokAcVgn1oqcUnmLDYav5BVt8ie2r4
pUQBuwS2CeU52ImxJ7+OSXV4N9Ed1aGCwVtX7r6k8ABP8/IBAT+5OdgMhNgrQJz/
UtSJiEoAGAMqCyvZU1Qv3G5USmd0Xp2ZxnhWKtY0QW8MqHZs2F1i2q034BYFJnfF
ShX+rtNkqq7xqt2cZVWgkG0Cn69DRc0U2QhddkLhfyn/4kSrZ++9tPZXq/XouHIC
ol9IV3+jrokd6HwdMYNJtnIsdooZh82iww121TGVHDvJMhISTyMQjLq5Hr5Jdwwe
2QviBmaHV9JEmtHXTgX4mTgkTs1l3FXVXhBB5psbJ0ubamSR1DKr13k3LCmvNskr
b+nTslkgQMxJTxDCuWyHRkvaswgIgV8BxgyN8RUBWmDqR7Z/3BEmmO6Xfm3mzZ7G
ALxtvGh8y2OJl+ch7s2tw42rf0ArCUBknmnjXM2V3f3dQqn7bxRslYnMDAyZxkJ4
y5mU9ZWpdoLd69iJH8KYWrmugXg0vxbzCw29+QFkmHk0pDxZ95qCIXchcttRxmOZ
wqdGo4LH6b0dTxyJfmd/zopMLdis6S7ZePJr+22pUeStsytPOKzP95oVc0OpzJAv
QH9xR3W7PSYohM4NZCltZ0Z2spdpaEo5xkQ8xp/n3IM5oKgr7/hFbT4TLNFCLx88
mKDXHJ3ng5A+6PdVCStobZfeLYGEYcYQAQxhDcLHbxlyFTnuWjuXd+505wkJ56jW
MyHdi/ueAT37MmZJwKdF+xnMoEsQGh2p7x5mq+Ey0w5+1mXa5peYRNHjdoIdORfD
zVbkK/akBbj9s9F4ljSIRQmJ7EHYWyaukzFuL7zifKDSRfWpgC2NiXwTLWOJFvfx
7JVKxEKleqE9EeXCoNy6CQpcKUvus+m7KQl2SDfYBRV+840NgljfPr5PHQG+5Fv+
ELH0QP8U0Yy/0Pgk3UqwygvMCp0uixFfnoDF0HdOWFT1lqLnl9+kPd37Q45wHJXg
hFSJD4HBtyHaRQ6yLVN7KvEnuUZHQ51suliuMoJ4GRXf/n2ChFd6hXA6UxIeWpWD
Zg5Lx9QOWM6uxRMcj4UFq8zkURD4qcDTAxs9EP4ATIC27pyCamF47bQMXXt949e+
NALZFCzI4m7Yjp2QSY2h7zGZDJXw4+MtF2Us+JeNbeEBmeYSapqWKbRhRjCoh343
OWf52J4ko9k7wXM0QrPehP2KPiJJbPZfVarlsYH01IVCQGWsBiAqCIBmL+2zKoeU
GQQMvYphO5uF03HtRV1ulkKtEgkfq/ji7B/bcK0R9OKmFtFb4fC3UotaLHoDDgNG
Ki57Uqo6/9QFhzIciwuiOFUVfs1BU+Qk8Jr/Bmceq1lwZ8aa+/KQZb0GWxAejm5h
ZSjVpiCAXUMu6yY2A5YUZNPEA3Prvtthay+8SZ2OwLYWHOMPCMxNMy5xSCExYnlI
MqZJe0KlA2eHajX1MTmmxRW6b4PToTfYXWciCagjbxyDG6kFS9wilWoxPug+77QG
DFCe5RFaxI107kHPM2XwDnNFRYw5lnWpIseXQOdfJgO7VifFm9J3c5ra2vMFKFiA
HAenPDQqE4k/MVwq5yTFCXei5s6XZVwZ4GeUDRWDsqe6CE0BYlLMM+fk+Xm6pK9M
y0wRQZkeXHM26Wg/RZjISlXuYQr8FbZWtDqiueCoAS3A/rxvtz0ZEeTuKPog7L5R
qs8gH1WMOgzg3gLw4hz0yvvdkbPuN5R+EqJxpC5CAZwH8Pd9Ma2Sl7ONm3RClzo3
RmpJ4IjLmcktxYRVvAOPXt2GdxoVf8FHfqGacKB/QbaB+tuUY7oe4PYKPXn2awQ2
UHcc4Znqugvgbi7E9n1YgsU2FbtL4kXaqBui8cSCfSgLIcza8R6Y0FGrUWCkp8gt
0H+UkK9zkc5qw0Oh6cCKjiOgL4/gHmxV+xc97BiNeAmj57Pt/ACGHK5PQ+N0zYIS
7z2j8+dnutQV0H2GYA8yXrVPwPDX7Hlxn6tz9miPTrB01JvqDAkfn2opnZEQ4ThB
ZgAXtRFUX5pl1ReJllc1XJvHDYG+SUFZXjGo2nFBhzAS/WFmKb3aQgGih8jjCGL1
xUUV/M6KS+4X8k6fDTXd0ackntgyIRQvZ2ghm6CxLTHpidv+zyqYq86zue2/RSNi
rwxQYwhje0SajsmNiVs4436bx6AQv9gU7aDMXjiaMFr7j711o+aMpzy6I5FoINFt
5XU/xfN6hZaPS2L5uRJKQ8dkl3OVBod/S0hhG4BaAmtlwd60RW1gZweQMWyGc20n
5ubNzMEzr56fAaDuwxZSr8l6N3BYyRgpVKlknDT+V/mZmaQ8QfhghuZyOUOd4Ovf
61xMn6C8BexVEMEyrf0zOpx34W5BxWODPP53vdQ45gR7c9w3xnJC1noG7uC/5gD7
hVeUedqO91gm7mEOvT5RaK4gU994RV+7S8E0HsEH1db3SfxBEUhQ+t/GXBbc81LY
2yL4asuetBhdBRHLTovwog6BA1XLmNazXJc3uBGLDgMkAH7kSTLxVAzVaZMmuPTt
zFDHwtjscIdp+t5Ws5Qi/7JA1iND96/jIQpt/ivbdCQ6faTKfpncWqGZz/CNrfkG
wvBt9EmHAtU5APHopJw+GvqUUDN/vXnF2EOwRD5gZjZtOyW8waXXxjiQZcopSVN1
e3T4W8FbOI6Nehr5K+sZ/XfWK1dPwgIy8F6EqkcnLAuKV1jVgTFwktg4dWlXZIor
3EyfPOfStKx28wH6l3CcG8PAuucljyNrMgfrOWKLp2G5igB+zNuSxDGfb3LynEqe
P+rzUsmkI74jb0cGHtW/2RKF2mzziMin/3aHpGIrZOjd0vKwfQQFikNfSSniH/cV
mSfhhUsNgv2Es9/Q+7gmIUqd8IZtE4B0xV5PyRUpvKCafOxMfFxri0VHjmWwMabP
qCQrtv4QIBhjftw1AkjSXTVz/aF+FHRCgk6lOC+qy+JyR8LyJeaCq16oNqA/yAFl
RWILZ/4F+V3jBTPhPQfX+xXAZehQy5iZH+QXkF2RU4O/AOM04vv6IhQJlRNVs4Px
1JiCctrdaI1TOaRc04f+LUxRx2AteraAVZvhpjx0CoDVO3i0fxhTyq5rYGjWTBca
m1xJFB8pfciJYhHT7EEoUFY5eVUUZCJNW2l//atkjAQTod19hCQCEVXFiZ6RFxdh
gkaTIcmNa9fa5S3a6qoJ1VyDWx88BIlwLYt6TqscnjYXGKulpOwjHieSGPp2MPot
1NKoEwJFPY/1QSp8XkvDux8laL5xwq5IKZbNDspQxJyuisUw+cw742B2fDVjUWCd
vw8LyF8VoeyD+UCD96nhknYoH37enku5kxxagKcEFNnc2I/Xb003W0mssjxgemjH
bn9HyCmrfY3YQaxrp1F67tTAxQPlnxiPY5qJfAWHZ2dWgcF5IugKrfFDD7ZF6mmn
WXm9leiWq7wAnnrDJrjMysNzVOaxHeRop3Fa8hC3jfAMirJ74Rgpao08AdzZ3NYH
5yh3uQHiQvNBkAhYlB8vER2/sxEliGZp0rJatTYCtKKJ17KQBWgboQf2R14ocK6R
DJlDMP/rZWu9VeIJD+MOMX0WuJoCsP63vtCoGJrh6hQDkM+rDGIObtQu02CxoIpv
AQ3IN5C6OPcKnpRqy7h/NMpd9oh+sm0/2d1MmWkbdCOfqzPXFNA1z3hw5l8ncwJ1
JwBSEiRODJLCjghABF3OSSETxreTmGICBOaOljki1nNp7PUl/3/mklrMKLLdMn4h
jaWZSmuVdIk3e0seGJ5GCqusKu80VI5kO4GY6lbixTP+Z1XidzOjMTraDCNW7vZ1
lEUz2md6GDIxAlEMcPpO/XgVm8X3FVyTbAXG6Pm6G2H3bszvIjnTKyd5Frjow6+O
BVuJTeKxoOr59Qd6a1ViBhJ1HLcaDj38cL92ej/axa44HwQycMK9SHDGZ6t5JFe5
Xv2A4S3t2//HaE5DHfSrMQ5d/ELpWAO245NArxSPQwGRczzrE/22czzZK0EYSFjk
A3TNoKg89Fo+rIn7LL/9ABY1JX9Qhaxrs/LGQCM6QIiq4rbEGLKfiKcX5CbMME6p
JbZ92MSWwU96ARAj5ZEIZyc3sTtEZgG5+b+xKyY5pvdTtD4T9T4vk+pPiNRBQc/F
hpkLDoSavIu+8doNHAgZj3DtPW9izxXOS1sJgZXluCanCMc7yWTFPgVZzqoF4AZu
pafMcRHmsdFYCA8PBm1A5xk0l+G7KUiGwSG9xeTnxJe/YBiIGOXuO6ViCIFKC2C/
Na5/+pZxP6L/3lv/xBJldbWgt1IKUxn/cAyHCtkSijkWf+dzXij/aK0P2fCHqira
MzJ2e5YVZQorL5BlQewW6GGwTGK9TMF5nOX2rlpayOy1A506ASoXXc9PytobRmtN
pEA92Oo4XG/Hf62MVkw++U2DWUI7R/HHnTOgY9fcQU5jEeIzmy4EZ4ehDXCSfrDm
EJiZiItbE4CdZsFxs6yzG+UGDwu+v18RYTRiiXHRVZFNP+cjyNXx2pXy4HlyOfMp
HuYM1T0m60WwMpiS3IjLqIIPUqQC4iuGU51GBDsCAV65pzG7wLS5kmjR2R/WHyNW
aqCMiVdxBASHVHMFtf8CAX/AH1EqgTuttYI6WCB7PUnrHvUx9ptu/GwvoBCEOPyz
CcCe9y7Sau4RZ9PRfJOQwoqfUZcbSm03RBOS/qdb3NZxNdGM20z462+/viKJfky6
2i6PMzS+j7ZDry8oyKnDWtXMgSpN5HyG+ouOAuhwKeQyOZx1ZH9cAQ23bgUl0Qff
Gq9LPPTCliTKQQeOjBCAxOC//OPYXnczeEoqxSwc9Ym2Zga8CwHhA9refBxXWxuc
/bOU+YCxGyJi7Sdv414wWb3uNj219ABeypVnbHDy6ZOWSh448jzhdHjYEUDCTzkj
RHN4tAfxULko1xRxlvQMb9LxqPlPqNNLCFDgyEpxsuni8jeI5vaT+18JyIhYrv0W
+vCwAlmG1PPCCWs340VkN+Fwd0pSmcBtnNaD2YyCM6apatMX5/rgvoEGY5fjryWR
LngsqnnhBTtvd+55hFCO2wI1bJB95BPfKhPnYTbwM1pB6JwTPMqeABBtK8wU7/hi
rPo7E2mb+QKGRlLwt7l5ChnnnPeWBNoWVIEZjhKBFkC6vOKKZuznQcjhkLCCt0Zg
SKvHWkn3vqcn1iCXuyS1C3r8P/I7j7j2zKfgrsRBQINWjCeBmwLwiuVfQ0oIjpUQ
l1aHogGw7Mjho9UKnpfix3TVsgqWIWjU3FVwUZrCtV0AxlTv3zhjGA8HBjMHsXjL
2GHXQkWXDQqbyy7UVc+eMCuVnDAzL7q6VpZdJ+pS8bcijdUibwYLMDfPBgpAxpUe
TiP1KaISTKWDUOl5i3peqoBUDQhqBwwEY3HPwXfGeGh5Hs9ut4nXqTTX/UBAZInn
HZdsMSvPfASFKwGDtyyQvZhgcMx6S1QAT/H4XxsfhjvE2gq3L2ycWm5QCi1lnkBl
g9j0xYlmmRzew/BVZ8fJAGLkdUzq3WSl9EYLELH2wv41/WAbnXE7CqmVNuay3Ljo
KDLBWK0+XVMHRxvTqnaEN+4NPDjSebLWvsDrCk7OSvR3Ne6oMntRiiuptj0c+Hku
3D/yKbgFlgYyIVNX3b8w3Afx07d3w2ci7SvalO0izms/wxjMT1l1ImvA2i17hrW3
41Zr9uIJ+W1WxTCSLXHjdI02CUyCKszm0YDFWUBy7MFx3xgzqH6918D3bvCr93li
jQ4ngj1u83JREcA6wvTcBoVnmUAvA4CKCiG+GxY2vBnujsE6SuSuy/V6WhnxyN3e
qNDgyYw4JNcaiT3YoMQtQXdWMTpesyK4sDc/t7jNVCmyQuzc/bzd3FhL4AhZI/ar
uP8qyIlTlQilBgMFNnjm1+cVWX2odrreEaA23PwUMHytJnDHbW826LfDGwhaKysQ
L7I3Ht1YLwVGaRtssggRp1OgcaD2hy8EdQPD9ntXy3xFIzxszH34AVWodECuIsH5
ir8PoX8hqEox8qUYyTF8IPftUPD8q58lSZpy6nkdN+e2EO9DkK/8up8DvZlIi2Lp
0uTAPY29tZTOnw4KNkSVx945UTWqbO6J/rtrmXjE7+ObrKRVNEDeFo4ggh7iHvWo
HykhRXjodyoxBnxZyPb65inreFjAmUcoB/I6xGTHj4A4kt3kAKEw4d+0Yho0DuYy
Q5xn0Jk/vOCmlJePeOGoOFmZhP8JT+2q7yMNayJq1dYPe8QWJopLgRBhlOoHNQDw
qPb+5WgglfQa+zelwSEOhqOyrL/QPJMge/uVwObJTbvmuKj2Ex0GC1P+dzLYZ0R9
2IzN2KL5zVC07hoaTkW/0vDrWYbsHQBeabYxMAEtfpeAFkJEKXZzR4wiSCez1bW7
bdMOOcyjFCCkfZvolfT+X4kssJCOTT/4Crir+EA38nua5Evle9X7cXRKKrJMS53H
igk8oMjk6JgKym+ZKnbwvmRnicfIhOXIJLxJOfnQEzBy2XR4f/fWmuC3C7aYXqoI
3IAQn+gUNHdOF9OrJqRT+gmJjm3cDGv+mA05/IHQV6drVeBeeYP2nL4loRe77k1i
dugPUAKL2uk7VCLc8iVJxjPEy9Krnvbh0enbHnyY93FnO0lo+3bo0zFeDXkg6x1+
TXD+u3XdfYDeMwjG+MjTctExd6L0Az/qQe+b5+4XwPQZQRcgUFfICJhw/ZoPZWPZ
9OUDppA1LGwBUkSLsYL9l7uUCgig7ZVj+GMpSrK/j4P4J/So4DJSZ/GzjhCntdME
a4LBodqmpCgEZVY28P2Abuz4bX42k5FXb2VaxXSdNjR/IryNa5RbVylvY1stnVzp
boskmWJFJnCz0vDnJ5SuXj8j0tLYguGoPa3DKemeRjHq2569h6VfwzXfJqw7EWm4
BmWEZQCuy6/wCXEcWlD6h4knoy1QfXmFLbcuUt9DtuaUCISb+bX4WCbv0C/t/0rS
eLGE+K3K2c7CyCf0ZcNehxf1YDz3CVvU3dgvH6IkUtpLtrgVNJmGpM2jx68KyCH2
yj90oOHBDlyph0K3UKTZv4PxcDC5lLTKrJNrEBAuzONI9ekgVYsM4Qi1QMkJqsWQ
YfOtxlxH/iSs6Owj4yLWwExoDK6t0uXKBAs9jXlVnaIOwkQnqqH0l2scQuxaC9TF
SdDUYXJcmuP8jdBPrPvT2h6TJc0n8bdZSdk4/5tyDqnGqZhe3OoF8S/fjjByZFvA
b1TkJGy5C5QdfB2jX3XbgE9rD24jBFBf3cwYbSchm8/VPeuDHhAS2YU6DbLEwXoW
+jEptEHS/yjtVnUlHNpmu+f04cGS0eRe0bPZVAHNFfo5zciWWsqasG+raXeYH5oR
yhtGhBtKsKb1xm/tYELzUOKVISecG7UpGxw3QOfFHVmefdJ9J+2s62nb6csth6P9
JUMb9xmAMfUywN+7bVdYCckCdorCDcwO+tOeBE9y3vM5Yll01FDZYJ/AOXA+Mwqv
GpUKIffsWe9/VmB0T8NppMilTnNAUOKJflXsrL5fRWvcRwJHCBT2y4iQHxy7Aflb
g0G20FUXxE1gQ9H0akXCNVcSfcCftGjxff0nfZn2qR4oFmGVSqhRStu/wSZlbxOy
Zr61rbaZ2Z6QcmodcLEwIQWwoQvIuc060Nqmea1rMSuSuK7YqUM6TgEzWs9JVeyA
1HFCxk5KU6pmtEwojevona2OLT8UYXqmZ5xW7rMWrhPtZRVCZNP6BKKEtOHkXT/D
n5472KqWFTNt2Mc89HzGmGN2oLA8a3Yc1JgvIJPqzTngXGoGmgLcwnlWbcWub7pS
1NiwmsYAFMzXKui2uW5Bj5mpjCsWTpZZ6fNDt3UnppE/v2jw58hYLOaNUv85b8+a
ff4rKbSb23mjaJtlKuemM04UlfypgF0HmD1P63mkfWeCn8DNPp+4d7CxhieX9xAH
sFN7Jq9wyJKwuroft1FQ5ix8d4nH+c4CVf8g+Ic3a2CN7PJXKOuSu+cc3Gyyi1V0
/jOI3wfSfvsjE+/PbAjI6IGoMRGfal+Yz8p5YvFRF8ShPtMx8c3nmsgJDpW8RNd4
4K1Hn+A5GeR6rCLrs7BJsOT22Kk96MN6cU459NTJHddc9qWvRfwMSwQ/ycgQ3lWf
STafMuLpOISt9MNdD5QHEuUBNgL2BgsbxjyzhU6YTvE7/jmHy1cwrsx5X1UzJP2U
JLSGxL+JBk8d/xMurroWV76Sfyv09ke3Q7WCWBj/RxA62TfYBCEFMJQqTVnWkr56
8Fic/I9UQghQUfMTAG1PkmBFuRq/3T2YxAPo/hIEMOYmtcH0NnBy1m3YOEvucTET
bpyxavgMxn7Wzo6Dxdhl6KcYG5tBA9Kd6ZsO9iWg8NIy0ozxifhxy+19veIj5K1z
d8/AXVS0opyP3ojs9LhXkXWV3JY0kj4AU+T4WTEE+wjmDbgtpJSUFblXSXyoSsRl
VSZUxXwL7RK6PHwvZ0wAYopV8iBqG/HacVKO/you6FNKdFM9+9AuO2KfrA2MA67N
tzqgdX+VGeBrJ8Fmgqhual+FLhVHfnAG2Xj0x5Vznc1/9OnZfl2mjKa/fRg54Npd
9YO3xKQ0wFO4xSS+JRkgj2N615qVxskG2YkFaz7Kd7kKHEikzZkvZH8URJhn4sxp
KI7efvr+G5XAe5hXaRRenhwIsM6hqQVZg8uLx3UKsPTnqIRYABb1McXB7mX0RNuU
hFe12Bw5kyj/IgOervfo2T7rjV5GSfQbjdu/pyg78lJJB1J+FUu+OTzfCYAha0sC
VaPwRDacm/DFgKaj7oYWvr1N42DKH3lMBEXeuLbD7+fEOLkbicHi86tWhFBbL/hG
ejh/EVeuBgDuJpGTg2CbNThM59t261vi2oDvu8/LR/pMtQ8Es660ye/6xziO36NC
P/WNyieY5y/Onw6ujcRA45syIumVhUNSOpMX27o2yGRVShzagZ/C/y1lojOn2acN
LH0lX5ZfV0ZjOBgGeRtBhtuiDb91rOxBezBBZM+MWs8lKdSKhZacQOQla7ffXdEJ
4Wmm7fgmEB8qb4RMWoxJ7rNOcxzIA5URWOJJCC7qXTa/hABsMckOtYoCEniObnyU
yY+W4FeDxuBbkUwkPWA9TNwhBF6juxlK+cp3+q7Dtc/o3cw6SXCn65nwkFFQB+SJ
sYx26KzGDtNCrR4uzlx+CF+/jIPdntSvDvQfxy545WTCLKb8xy4QA4a22BIrnk7w
DpsC64kXzNE+bzPJTRtVOg/vg7bKhglGDG7O2qdRLiLGuIPlCLD6356+4UpHI2Ja
+Q3HX/iKJNasjGtACjl9QE67HBZtRirkRwAOLvVCHMFvlMjpgwmAhA37yCC42b7R
bO8P1mqmWDeWS0gxxfmKp6FxgacN3UE0xMnBycgiPP4dnEhwgc4nlL0nm5K6U9Up
F4irfT4n5lkYzwIoqsaGkSE6GCtuJJD1Qgvs3zQrpnCXnSIDKLmnSOpJ0keN1HK8
ORDYiNqW5PHf3NyogkmWmhUT0k5XsDGIPmNY4EUnwFDrDdF9sNyy1aQtrbdkqOng
LOWticx7j2quUx5V1zZqpv4I5Uruw1JQUBErmmTRIWkVnW0ModBuo2lONEvqIfOx
BzSWSOmQEUkxnOOIsfVCXnTP+xm5RerLMMadNvkKzPfWzHc6TPLlxIskmQ40JOWE
L/SGnckC59mckCzTJ3uk5k+qpAJTt8Vk06kWKUCy0VDPYc7AoOkGtuQuOPVlVcTX
ogk1qqnXh7nB6o74b7NsJZFJndw/85uS+O4ugNhcJWu+fhWW5cmnXW6JTcAwwLzm
/KEzrYvCvQKUeCHum9ocqXdWk7jvHuUlVLPhIJktHu1wQOR2EhToMd7hBvQUCz50
nCE5YDuxXhi7YHSpC0hZkL2Ivk7j2rMJncgynOnLTyGtXPs2tuIfban7G9f3Qkjv
n7/P0NEp1wCD1HiuwW/a2HIkOAm9HKqh4fqqFnid1G2a2qWI7B1YjDBLMWDdrBlL
r59RyJtt0JN7rjz492O1hEh0yH2is4se1d0b1wvYwRdUWV0V/TpQpN2HlaKm+Qds
J8FU7tWihaxGIMhr0ow/BGJx3Xshm5/opSFJhKzkkpR0K42DuenwE45yccZRFreU
eH/Gi1cN5NlhhZZVDnGAn51h9AErIyD8+Xq9LoNhUdm2h8dV9x4g8pVPMgmwnWT8
BZ2mMFbXaQZbgjvEP0ucHFt7JEZSYEQSJIoUb6mLUyWwc+QtBrKtoRdLakGqqq2L
O6ZmlH4fbq/Epds2AnxGUDvU9kOYj87BGc7EGDufCgeErOVXAQgNATFT/igHfS/n
NxhEdDfm5JlJRTQc2QxM53OHYDKuy1viUsPpxG5ugSQl+4wBc7As7Yimf6wXI0gM
jXKkcEif/MNgTZLwtpPNYN13SiPyXsuLNjqoPVcAzWYNcfah/zmceVENzM6h+TTE
qlDZ96hwrk4g+v+GUpMdrFDv608Ks6EXacsM1/UdCWxs4QCdaG4mHdDSWx19YocY
hmAV0bUMwjb+bZPe23hPlSzuFd40bjNe5G9gy4PbrHXg09luqWKvUiPcM21hLkLq
3RCyUHKeOTx6ImztOifQi4IAuku/8XRMApl8UsS+aLSyzd1SmG370eKce1mti0J+
ug6O4ixd6NgMzZEMLVE0DyIsdSdMXlCyQoI8QcFZkX6f/cSbvvTXC1yvxQ8GgZFV
8+SyBXgyoc+SMbd87h7YHCTWLR4qOO9dgzY9ebk7HEplz+jK7pSMXu+wm1GdJ/UY
kPAwcrXKuk2BGyDIG+4N6vYhJQvjHVfA5zMzOyXFqfTEzoeNuz+20Jq6miy4b2l2
bfvDhkaS+XDJDprIvsD4z1PvaHgoh1xaMV5Sb7NONeOosI7bFGQP0qUJw4WxmL1/
9Mc/MtHHukwUpsKFw70rQ0n+V0KQzah8sQp6l00AbH+zYtFJ8v7wOMkgfG5DwAYh
cj4zCXqe9TaCdBm9Mqps/v3g6bVaU8OMXQMsnerBxGnMAV3PbmMyR9IbVADZwNii
2iHa+XojHN5NcbkXDe4emKrtW6y80foqxhHPq4VaNhhu31sHQk28gaO1YlSqeM/h
mIcsChf35fORSYMP6ARP/k39LyZJl/UhvhS6ScHaKCYFdDxbtucEVy4FiIFU+46E
fMVv3FuxZRhkeBcYyHTnbMiWqO2w0NQCrpXRziuQiVJkKOkjQu25bC+8omAHZPTx
PKgx2CRDjYGdZjaYMkLhai26VGLqBMMRXbaoQRgm9XGuW8afmXrHg1ktoYn0H/q8
3bDRbZ7ZPTZNK9fzXcd6eTmP0RA2UXcgjUrOqWbl4oSnfN0dpzQaOFGu6DUKyIPT
3TYTpBNgCIyHDTH0OiwmqzBv6VeHBTjRw24nlvz7UG79fjWl8eG9m5gTYtDv2DeO
B68HW/lKTGsPhzrpgbNT6FbbkV5l/cXFp0PlDd9iXz671ejJAW5zNPYdfpWHgtMY
fVRn1nNpqJ7EUjhrPHW17ZNQKMjT3YAeTpogO+Jp5DJUe/xp3DoSRQwLNj/k3n5P
Uvkn/1dH8KcebycSU0Tvo65GewWfmWCBWHemEKObG2DEbgR/EbTv4ooZvB9XKe4T
JxodK6jlGCIqbXxpkrKfmvD3b88Ounj91Kwj7MLurMb59usZ4JjslDCFKltL6bUg
u5O9jK+MHm3wlVlp8v5+J3w6M11FLAE50eKVFXDNEZFSfc0KdxTJ+ZbaBfFxYnVd
m0SVIr8aKJN61afbAPLMW+lOqjOhcF3+uxaLBOeGTSBfOAiBYVbFVdY0va/waaMM
xwlqaH5YpJc3Ck7QPGXRZ0YUneyptAgFUddehXeqbF3S3MUtV4++ArE8CCm5zi+5
zb/YrXNb+ah1pPpPP55+WV+1DoN3aVv34kukjindlBf5knzqDhd8DtSdCdTIfWLo
l+8xkhVBgL7w5kanyDykw3Heu7DQ/mUAUcqxxjUxU5grpz7LVOp+GQR2ayi7C+gd
cx3FW52GEPs0GJH6RqvNX0U0h0BE0YY3Y0TKOf/mwmR0BIA9E+bqI7F5PrwN9pKF
i0dAK86UDkJzg6orVV6ZbEYLsZCIzpD+Gqa81ivMXh2YV7ShAPW8PpBYT2M+QuvS
Zjfw94GppB3+AgnkUC3aM3/BDJga9SXlKtWvysaj6GmDcOIv5Yz9qP1L61PHFGZQ
0x5F3KJUM5yp0veRMvJ8lTwz5OQ0E5LBxtMyU/3AraLcq27ZGo7faKmKkCgVL10a
DfFQHwF/49i8024babvJLy2I4gimSXwew2lWP71itVMo9CbHQyy+rctJXb+Ks1G7
qzOq8eaXmt+smD+EuTTU53NwbhfqvS/XX7+firQ2ylr9f5XdgHYTeSek+TOroT8k
nAQh60Uw5S8OYLVcEjWGqx4d/NBDzgAUSLRoj1S2Q/Sv7wOqSmXi7OStF80JrG/7
E5Cbd9BowN4+kZXRoe2UzFxnQsWQ6A+k+ZSC2NY7+5ORgk6dRgDs4QtMM3rp9IUR
jF+Qmj9fkRoPjpovlNa5iJPg0aViVfgrwH1C5HmWCoKrfKj05ca/yUxyTqOYcwYg
Pf/kqF/ZCRrxJyL/vXlaI2QesSIBczRY9aTDT/yMkd72ER9Gxis7K3ZbS8hYhF4Q
5Nf8zTjctvXuVnGw7W0IBQKb9YPqvy/UgMMGstZdWLIb8OYTBlmCtjuQ/aaGHSEs
/xD2kCgh5clv4EcVzZxGMmIRRZZtBUnydpJ9+Ht9IeKnTiQUuNsfyP4L2iZYrGGc
kUyT6ahAXaPwixnJylkIJrENpE/kom/QKuXZNuyd4tCKfir7Y61M3G5nUUALDO3l
4mCbEvQC/abPwxIM0gnUXVp2nu2dOoCWsIE0+D3aYNOKPW33ZHZ5vSpPlBRXyLPB
LlpYIln+IWH9rZd7w1zKNF6S3o1My3TZkKRh1KxZgIM2VYbMFWwPUYXgv4QETtnu
CW5mz/haMvhAM/zGTX4HP4fpmQtidHQEEml6y//2ppZx1G7ghLwES1qH8R0eRzVz
PG3DLbuFzIfbCwMKa5JWpJtACVFJD5G9zXK0EwECJzNfwalMXqvUjGVaGzUyFbs5
tqfDTdT/+C3Keq97zBc+4X1gsrrFGQktUgIxjP9YInj6TfjAI7L0BqeeiGVGHgCG
5bcxOmETrQFTAXYHl6olpspCr+9naBuVSm7xy2ZJAk25Kv2B3iMa6YFV2R9HGWbU
/4ZHdckZb/cLdbqGABB7gcvi6hYblJ8yJ36f+/IiDVyIl8jUlqkly1GnbTiNn/km
pgtY687U4eZnkm7tG52KLi7+IatxoqNES9OUu0bGLjh6i7sIM0LVm31hV3kJ706t
o3bpN/bvVahvWfOFc8lgWtar3905ZjiQEhuxYYi2HqqTQgF2Xntc8A2TA03TvGZI
QJ3FLVQrhUxSi6fObXV5j1Qsm8nE9LZqWVepCG6vzSRjveGy7DfWeIM8tpZUWKy/
dGcg0AHQUG+lqSbE8OR3dbGd4axkrdrgLUntgSZBiI/0uhWBIuHUHJpsDt/1oTMu
9us3AAxgNy9GF6BA0H/Ycp7Fam1vNuKAxQnZKusibrylYganAbHmGGtAL30h/419
2EiQ9x3WA3sfI4QtGdcqB60XRvnjWmVLilkid8/AvxBJSEB2abBzm4V7BggR4TTq
vyKKzRk0c8ye5NkKwTMIsmCTpDJAASPfwqhFCwG+W3uqRL3mYwmU04+X3BMedO7g
cZfOnuCsyv3DEsohbyAZxkipGoOBaJ/Td+pmD1bodqXNOAPP1rLUlbg0xOfuKMgl
4Utu2pGr1NbakbrtqT6zMr0jPa9lVuiichmiijtu4Q/hoOulQ4c9EgWtbwxhCH/Y
5Ax4apRrJxtZ5QV+Bs5phgB65Z0CQ8N6FGaX7UMm6gUPF+QRnKuB2C/IQX5Yjy3p
+49iU+giuXyhfEqU5M2sz6MDILMXXej/2eNjI3QCA4ng6vD/0mJ7wxrajLtCAVq1
RS1LN8vC3XdhAh4dDArXfymME5+3eMVSDODtaQxMTPteIvO6FyWaJA3HPEBwBPOI
7NqzFg3eAfnmPhN44y+7+NNwjCK/Iu+YeSANYrdpciya0J0duXtDXO/Del0hl6AG
xwvA06NtEc8sUC6ZhJGHi1KqyQ6c59tkl3D3YSyDQqMJsL67rSNeFKEOgzN9rR/B
bfw0z5GC1oJahui+4VPP1297yU3EYqCLz+TtOjbiItLd0Rlf0iJ06MUBklGZD3wc
/Z5VTG4lE9xwPjOJdtRI17qnkxWAKwZ1kT/xwAiHgqE0sS7XjkEcUNJblyifSuaJ
HnQ3E0+JrLTgBp0GJR75WQ1KLXFAsW01UwLZTdsD2mDOSBAbZI2z2+/X1nNS74G8
vofpDZGzLFnIawCVTyRt9E8C3emc8Wtr1aiQn93nRaVpyoWzYa+achQsxM9CSuhi
jvxVO61r9gAhWIVYmBlULnQKUyceK0K+SRRMCgb0W26I269nu9IdMnOYLoHGkc2z
yBpsw5QTtGS231alDHatxRToY8RljnSCL8hFq/HtQatC4ge7YRi3TsfkB9w8WARC
ulTSHQtKC9ncJCrEut742qjR9ZrALBKTF4ZOJ0evbn7PuJu/dGqV0Okii97i9Gw6
3MSsx6Cluh3KGSjWr9ak75IE8pDC3xT4+SRcuUan0/X3/QY74RYKa1Et6LjHbyBP
TNZwnntSHj46E+1Ofh1GsDIXt4/4k3YjsrVtjCEKk4T7RuDE6RPIFkMAVrmtU5+o
3fFfAZqnjc8vodvHDlMCDZwyxpcIhnTGN4xwbFns2jZqPqYe6V18Hnm36DjNBkkC
jTYY2/OhI9f0y6ylj3GpRJ2MlvXx1j5reA6QcQtrEpYVjeCswJ4Qra69QqABQVkS
MLm2jTdNSos6h8MQkutIjmTWtytnWp7bSYiHKywdWpJxuYtyQ8Mm68S3ckUmBxLf
paea8kOtHw2t2RPTgjJ/nD/1HxSvjPxfEeidJTKBIvJFSpx7R4qFlaI3cQk0euzP
ZY6RWep2sEluoq2D4wIwKixlGnyRuE2CV7dAsoNd1E3ARwxyOeYeQrVEhuuixkxj
naNWW1AxJ8LjBhfY2SSNdskHRMq/q/5yAxhvjJD47SwKgZufkBVzhb7F0nM/nEjg
RJHNTqo4Bz3sz8cUj07QIbQI7qYl1ZoBUfEMSWMXdqgHU4WgWjiFrApegqf12Leg
oBswyjaURR4MEtAa53ZmsC2Msnp8ZKXUMQHtIMGnnWutNRO22ol2KylzbaCaKgRf
U7sWHdBYY0cL1WxSJxSFRFDrJ0cpRRUMKb1Sn1YATbanAiNjfWKyIZEgg0ubIPoH
wvOrQZz/ZSmEmJ2dsA32DIgD5zPLXR++IxoMnuqB8caTO9dS7EVl+dL0narFy4Uw
3T8WA87UT8BnrYYW0PmSf1iKe7nd0Pb3umYPEI0woybdhg82b47XE8QdkMFancoI
k8yNKU+vWR0pGDxPZ+GeNtNtsbLNPm0ulteNCVE1XqoGN6rNMdJS3ra5EBi7DQme
vqS6sGA9qccIu9wtUOwps2WQlVN4pHIcflLp+rAAWW4J9IuzHAUbOYs8xuSaMPoG
+8jTYxRkELVP4dzUdjJqv8ytF+TDEJzuHjJ5U2Rj/acl4h20AdHh5+xXZAOPsYoY
MF0XgxP0PISrIOyIG1Gu/OJq6HmZfKHDAL8X4dtwEfkpi7j5D+Qvnf6mZ7T+LFul
uiwSVrK4Tlh1XvqqdRHrszwODCy4KV3ENLlMtpOy7Ms9DWu37ABI8heXOffA5JpA
JYrsQgFxEltlXlz34d7uQUmTzCs+PDpIrycEqiQQDSSBmywqVBBh9S7nMD577F/a
234JadcdcqInSN2oiSe3JXFVkHTWgUU8MHVF9Bg2zEKNSManRbYtUP7kwa/qLJ3p
tkouIBPvYqZvbBHEX/ibYL5UdX4FFeopiykfPgXQN+ySfs2wg8BFrKfxScJyhKM+
zRrr2DG8pph//N+BnH/NDYzKtQOLyeezGOHnx7lX1QLGOjc6HHU7u4wQsEPP1EJi
bhKuJgOVaVP981BTptxkpe+ggRUkIOUHsJCewBm5XjK44gXo+xCc0VtY98y4boLx
iq27NEFPPtZl4AwT7FzZJbs2HfT6aORCvCfSfOmJziE/H1t8o1s3cUKtli2J1Ndd
nf55ywvZ12AtPPjVSRbsiFx56pBAZlwLqfOfAv8F/qEjtwZUnCk4BTZdgKaNfmzY
6ihJ0QwJl3EeQv4MlD+sApB7H4sfSShae1SmjP3wEhLuZFZfUqYtl6jg5dErrb8d
eibGReaajvcpb5pu29Ar9c58hcrFfo/yCm+fTz9lwNZ4PeKztvkoYVThCUIphFek
yUMjGtd8ZgH+u3HjLYFNz28J5RHqZT5ZuBPrjUveQ49x2JTUfDK1XrFmmXF0xyqy
GQcA1UMB7wDmskhnKoe1/9c26idRrmXDP+v6einfQuBnHs4afkQOTseFTCPt24Gm
dBT6BcJxUaaJWBQaCD4KoFOJDxsy+lOjtGuvCPIoUgfNXfRXhvFWJ/+N0lAdwL41
toJzxY7UP3XqKIgVfmCJUd8itOS07MWd/myjNHs7bvFpzh9RkU0cYl/tkKZaN6lC
BLDmHRSvlpxzi1vyk+NmgS/zRcGOvn16JNFY3ghUuwzZ4sf7Nen+Tc5J70oksM7s
rof8I7wW37qOoynI4qDSIUpYHaFpLqVb0gyCxoqYiB9FCu+S1QEEk9nPjmdcJH3C
MiSRN2NLdLVEs2I/DVFZ3aWsKpgAb+iZNj+eZHdJkjG+sd1MX5/LxZlSsnEK75AQ
yorp+hGSI+ftZ9xGTyl7mSeuiqkXfaIDd3tYFLhZvGeBaYtnKFYKsFe8YkdQ6OWz
zHJoB92yffSzxsuMSl3j8M1yLQluirXPUcdpKsDSOBQt53rytR7dHOkVCt3gI0Ul
BdXV56Fzup9LaG8MmS+vbr2PmefTvlGMKtUzSzj2tv846IBrF+zEcIb0Y5QQ3eoR
mLRGGSBrZl+RLcvKUcE6oIgkzGSQSJXbuvlArusdzXrO31q66Gc3c+/9z5GckgPN
VSATS92RjeRXDNMXdfkryvU11r/MIrR6lyXHH096ZDZ2DpB2upMIPw79DK14/VXP
WsABBU76vOaedq+sE7Fkz95gDEqlpbR6QkY7NEvYfcl1K+tzmaEV5KogdvkHVbuO
4uxc114JO+6LyqWD6mihmPu3ac67lf+RrcRJKmU+4vG4g3WJasOWjU2J1sffd9YN
dSeN6rzgoYUsfRUAgLEM6is271ajlKAGORuN//kF/nXzGXtVGngdl4fdlZvo2Y59
2k24CrYSg4xk9fw0DTiTH1opuAWsRcJh4lhAOCopxEgKjJz8umloZV/XpkMgaUsK
+leeCv0EjNxoWLkKIwYlxmKmFodPBmdVSsWGcTfgv1Odai8GZmEXEU8o25CZ0Bit
f8cEpynEUaB9/2IKNzHWmqBAJKM92UEQy9VnA5v2bOAe4zMfD0wk4ovZSJo8Owna
/MliiFKO65BMS7fC59GXepptV4mTWCUOx2OuBeSHeNOh+PwlXtCPOWVVPbxNd4+3
MS1wNBy+f4bLGQkZ/W9c9lpSt0N1CYNBPCPGrPsiRsUc0gVW7KlZb3yyUXInKAmK
oR2aValjPMaYkLouY1m6CNDw/NFWrzMnO0FYHFeFeqCZcJBP5tnqhWXPn9rDkl5x
Py3a0NvYhym/ZdLPSCytgyYHrRRZd+mpV0Dm7Rasbx8Kf2d1rqvQ4jZtUv4MBoY7
c0sGDgMS/UXgELCT53p7CswyiC5u9+FqfOQdCMZ+OmLSqiHa6gwUIed7zQ3tFVDM
b61y+nmuDpyGfaMpKDn0SOsZBLOP1kXdkNSLmIJslsZaMIvR77dNQCJ77suBKvnC
l7CbZ0GojqvZCtRlfECKuRWa9Q7vq46tzld/QQiiZtitaL5arOo8jHBilbklkbsU
Ko9HWaUZixCjiz+2all15yuiO3njMkKzpSnFzEM+bpyATPyjPyydmZiJuuiiSo0P
w2qqdxH3ILek/UPoKUYlHLJtQhODa52tOf2vnbQgdSdM7d0hSUnu/1L0YzjNSdQ/
oT4h4mNGe33qLJmz7BxWOxpeXrWqUjGu55H2j7IsSfIn+br1yDWnzhBYcIFrwdJ9
2eIfxbvZuOv27bI3mbI48acSHKC8YzQVxg74DMXMmLCW+TRtXsppu2XnqggH/5FO
gkLySAx0Z8t3LooWVNjy1LrBIEU0asYwBB4MCK+DGnBk8THfLEQ7lM55orCLJeO6
tY1zSowyHJzz540h/abU6TBxDMFW0W9bKwv9/npl7OGvZP6L182SxawCdkYmWQkm
pt8MYrkSM6Yq4W4uBDonJKE3B0+oobJBgNH1bD0ZNYSgst9MAqGzErClccDaH4Mf
A3Idv4ZeeC47rSD+43uF/iRP3YHv6hIcw6i2uMQ0HNVZYRcpuSfIk8SoUNSLk02t
qsUCR6F++8qCQ6YHqqb7IufuXEs90Sq80t16jt3c3ZO+LNSEyWklK/p4t//UYuUx
ojyr+9x1YsZOYuI5jnwGT8b2FwfJ2UIyivrLRXShUfn072+0iveScMb+i8QhLIYy
dVhpsGGP6bEQeD3swf91E7gcElkzJxcRE7e0P+4kmBNmc/8hgQZg19ZSCyLdX29O
txeRD/VDnrPl8e/KhMnIP78v0+cFiPqI/WkGVoRG7VlNpWdy6vMno7nvH3UHlb2s
yeMaqjDq7gHvhjahOePw1I5e5hxUmvm1/28NWUAR5PpyWfJvpfCRNgbGJJnuPagy
OYj/1BrHxrtTHtFCcoJUb9MST13MT3zXhwm4/q6NnyBviD4TjFxU/0Qou6OFV/vc
zTX5UAqcyiSCIgFksxXD/lDclQ4CuBygXoUNiKHy65dJpo2vA9CljnCOW6tmpQzM
0VL40+ldJGsJFudEQia1v9zS0W2B4G1FkWthL9o41m0yYGm0V0DkZn0SiY9iJyzb
OTOMtncMhLnc7K+pcX0NhfiSPTVfJO6mlAVPgkvi2AUr6D9vW8o19qX9DZU0s7g/
5TG1DSBCzaehmTwm0W2V4JO580telIEFfmZC4sZh0c04oPuuskOPbGQs9fyhR2L3
6ugKBDQPdYxL5bLSTkXfIF/XP3zPQDEVfoO3jQl1DRiJlCWJ8JDIoGxIranoRW3v
5lty5C52kemXS+obVcdIg7q7vmaNfCyuX1AEcojPUbD0OYbNIDyjy3aMBzD2qf8s
abCuYQR/NIrQqrxsvZYm8U84AhOX/sE8rRhKHIwtXUnSu6YtkBLRbv5iaL/sprNO
+/1NzBy5K7hH3WHosvnZpJQZgXZz6aaSAb21SJ0JPDxFQMz/uX3G581K8OhsLUUI
ZnVXjCrOznF17SQKUOL/CfUqiWicQmI2LoqKkMgdPuMMc1E8Px+EgPtNRDnWdqkF
tvVtpLnuUN6gKu2KwBCRuEEJ+3SfgQTJAa/y8IP5qw4rsIHi7p4N8sYHqtWsYvQt
UsydsmDD5QFwgxpy4Vtc2XSCyN+E91hPBNYJqUJhJfKip3EG58aYalFy3e0CxkpM
ACjHyTcD8YEPqlPEqFSUxfWke0HrLB/corOYPdQ4nN9JdXh9kll9q/APL7Nv6fHA
+Shxiwr2qHNjZ6Uu9DqyxFFYZH7pjBCIMJ8PC1IKuRCe0+Vz9S+yy9sDEzMQtHcf
muGhN2FZks1SUsbm4I6M95AjJbazSQ7xrTP3H3BhsbWsgivvQpGoSKaBYMWnQMse
1Q4qwFyPIN/Qf+jWLds3f4AcGjQsPAfHHpbHdyDO+jaYeQT85T26BCOSlkHGV8nO
8Wi1tSGXy9SMkTMHGMAU4KzhJVY5KpwszivQyy1uScG99/YpTtle6d44i133JNJ6
dn+UoJfqveYLOKfF8QGnFSDb+YHWzc8udDlevMJBomG4nRYIluUXF8INy9eW8jXE
ewbJRqNArlaJp2f8j0is+f5peGzF33eVcNZURbV33ThwF45h08HjkokAJ2m2jxnk
nEHnTjC9KLTv5hPqdoXGJIdcds3yHIl1WMEMnV9Kitexpa1tFVE9r6XITvIo79lc
K0soTSm06B6V9R5sE9iKGdMpz06NLzGVrNqOH6JdHdKR2rrC/4a570QosY7ldv31
75tjAVo2vVCQlkDxEduvqkSCvgmLxv2jic3scWKdBBO5HCs+Ds9sPt1vWTBJc9kC
hvWb+I7BtuFpuTyoUunAGqGRk0dvhIESokR9lt33AUlEChhh9xFSowmrO4B8g85Y
L4F7V3OAobbmOX+PcX+i+TltuxEYqtZpZ/HRJfHzpjoA6kCeONLSUQNxPVi+gZBF
TELo4kUSPGkaX5yD3eXU+UBRUHK+z4bIWTciF4izkXGneo09R0k31Jn5NwmE70OH
8+JxU19GRgJ5iAigUK+Sl3p8Wq2JDThojelRqkKN+up3gfHfcGNgAL/fGCJsam2e
dnaRGUAcchsDqJZW8kX8Pb5yPwycXNra+vIm2HZqVulEy4rJM1mEDSCqNuOvmvfe
ej3t1Mq5u3urEKNAbKO+Bpn1lrYvuYRnjkNvccppmELMsnBa/U9ccXZJ0ORQ6y2R
D6Wr6ACVwNXIet2MHotvgBat14IpXOLZ4cwgagyMHFNN8MP1mSMip6aaslxNicuv
RDRmrY4ukBPOuD/WlG1X95c+1N+OrzhJ/cuPjNHKIoi/W3Q/ffAF7vjGLwQ5/HNd
GCaVM1SKQfuicx6sIF8gLNTLlcBXSosVdGL9/v6ILUQv1a5uzhOmScgL0dsM66Lf
Iz7Jo58Ga/YaTbzjO7i4bO7KXg/FgCYYKpXOuqOk+K78yBd/Mb351Ag2cQYJ4o/j
9dMZCvMnMFhdBVlR+nM4qPKOngxpvHzfWUhfmZTXVLDxM+WXgO+85V50gMBQBSIp
YZoExd+DHi7GwtE8Q2h/A/+wlGxIRx0rnKywUU5CslMn3RJCAhbHF2QiihfyyQtD
R4alVLsVwJDvbHd7rDqSZppxF9Nd5+XUHzWuYI6XCzSsqRmV5ViKJjX9Oi+xCI/E
4H4YQH5gyzo1lXTDzaomrHCh6REcRG6f1fz5bBqWGAOyiUjoGW9hc7B2INsK89n7
AVuwDdaJRrdFA4Botj2S2cQlDIivfZ32wPbtN6RVkRZDPv/YnC+s7AXETK1S8FN4
cz/rZyUUFXGJtEovnj/Q1H72ZjBStYwFoo9FrZCyg0PhF3bU62GJ+ZgnuhU+AL+D
eWmvz/BefgThRc5jtxPqldLa4UCO04tmWQXEuVYIFa+zd+0e6ug/iY2vcDgbPe+1
LrhjTHDX1mfskk+BzqscSCXV0cRkKE0vAoBk9eedAcG+e46phxUigSoc7jkuM774
QUAcjv72tkEN0i24ykMcQscJG7hcSiLYXCCZMTmpj3Mzzz7K11mb3OGorlNE3r2o
dD6/qy+9FXuMghajbIs50lHhziZnAHIJvW10LCDeBANa3cInQj1l4IM30jDSRuh+
MrDWQ+cbvbcjwr3Tj5qkfX0TA1LWfp6GnfHNE1tE5bENnUr2ysL+a1H6yKmv/VuG
77umE3Iv9NpOigyltBS0LKix2ZhF2hrQlxZTfIJuulgpRdBJKZ/DrR2ROkFiZIQ6
qikyZ1ogCRExT/q22zvZVToygLX3yxwlS5Ot+TZYGY1M52kOpUVKRA+PqbNoTt2O
tbKpsz0ItWnZvzcR3OEUnpkkJxCrqyzh7HMnqWKZFe86ARSEW4Z+mRhtiAiHIf+U
HbdPCfNKZVSu45jZAJ/QlQ116zwZcmkj/OoJD+cSjJHN1eGzhlRT8oQRaTZiXHbO
bCvgerJO/f6PD8OIVOF3Sxj9i8f9BN5vkj9+rmnsU019erL6jsGAI4f/ddi0FOpi
5xJ3mzvd5KZWxruYROyzCyS4dqbYUR0L3Ez4oDufnJjYqJOGWjc1Q9n1LK9+zlug
yju2CQjX31L/pw563l6WIyUdgAuNMNDgcuztmYIFScSpzuT4GxjSD+s1ZAflqzuN
ZGXW4pIM0LupAC9kZjKif49BQdR+ZNA1nzij+1OvFzyWkIt5e0HauQddoGgx8Q5x
MDgR5uJbRUGQtQ/58eBY9FUjdpLERCiFHrux30oK8xUIVaFailTsZQmi5rR38Uus
RtIDAv4swlLxYa4W9tOV6RfvvpxkWrjg+nCEvDoUIOx9sHfdlwNAk9H98BDSdvMi
/7BdM0Qhi3Ndfgnj7xTk1pej0J0nfnHP39nNtV+x9MAdIot8nOUaPkVL+xYm4ifu
XTSo3/L+tY3gND3F3hrJwKSYhCLo9vjEed2W/l+djW4ABerbW4iJPVI393o8jia5
6KtE5MrUYXXn02uZ1s11LAtesdQZ/qQwrXZ4iqA35Vl8YYE4Q4+IgVmnZthRjB4H
7pV6m9u8JwOzsf+T9s0yfLdoTixbmU8SC93Q/uIEh3zePv/dZbMrM9xC4yt8/Ioe
XViBvQZ5NsHuu/iwff00KIjF9wtcZRefTxbKtjJ5dOPTpaJ+1Yod/11bqeYrnCfT
EUb4WAHVGZGI+SNs9UsNqO9bfjPMonatKGdtxoFtyAaIVMlu3HLgbQpgw2g5K6jL
oiqyQXOPNib90UWoRM5V6FKqzFjVnMa6AGWLJyL4IwOV5pMXhrpa9w3jCYLEv+TD
hu4ZKVoBOqkTrsl8Y+PX/kO2FJMtFupRH0zIexy0KP4T74mqIBysioRi4yWorM0z
FeMWEOgx6ZAdoalrB5mmB8uqpx7F0pJGtvF3VJREExq/s4rQhOxoRWK+O50FRkK/
cOt9lJDYiksiWROWXzko7+oA3nue/5N0wz3C44uTEB1C6n/Xk4+4Yig+Pguze5sy
OgdPjajvfkWErfrJq3sgXcS+9a9XVV+nNnMhwf+jsnlTIb7lndWywguQbQ/9Bq7j
EGfQ7koVL8hzC+KYK8hUOxJCbi5q6mzqDMfxQyFhzYJYYq1qWrbt5WKV3F+8PqPb
C6V6BAU+3Sb19gYpMo/v6fOkNTrTMoGJcCxKlDnUJJjgkIC/vo4tNpsxaZNeNS6h
gfqlgN8jN8hOwF3R7DvG4XrQRMeGeu5/qdRopyIAkUsWnMhW8ffU8ty0sYdsWysX
r9cRo/1STljn7EjQjbIirx7ZBldIUgUgbQeF7y356VFJtDtXACq0kMWvs+s6YPV5
+zcNfMsdQzQFkaqd6ibBxai+jxWIrChVn54zmHPzfnoo43XsX4lHVLnxvfELOa6h
daKSkPcnjZajB809c0KctGef7IUPpA/Y72NtU+jFvQQrmIBde0HaelJgfUnj9cCc
zq4CtOlU13bzG6wlAtpG7OFmA4RLgh6wkZVXvAmaak132afP79y1tqDo3UK4TvIf
b3IdSrz2dBjOvaJmfutOG2Deji3iTI3xUHhH2w9ti5Wqv5Jo6xmIva1f+B3Zl+tw
Ml2pCpPUl2X6QSlOcy98k+Cf7yiczCdDlxBIpaWORhbE+SeURSPkGGbHg4raa8WO
7UKpTe1lXk3826zWXpWlSq3PjorqGygllkvFdIXXT9tdlvk4sYf+i06ktYg2XJGH
URXhAdEnBvM/wjfvIYMJtzaTvvShIvRZrebYa0GPtKElpFljCCciyyFZcVf3Qh8Z
y+ye+YMwnv6GynyZWlUuOSN5TeUudPcOxQEO4OiFrRnu2Pk7p7HVryi72LWftycV
Qp6NG9Ye/rqm9wNL/FjKVOZz/jZwo6C/Q4BIIgKj1+4Bkwr/ErC3VykUTKM2CuhR
KxK1vpCDBpRab2xrsJQOr1n7uWkZWdOKiCJ/RwOnJJtyjalIasKBK+PbvSWTKGsG
CLVb2/v7ThWBVWsgTH89S+eId2HNlVDOK8wnNf8fh/BVYdcofJOhF+8cIwkl16aF
ISu3zdZAoHhFgzrl5qVGmqKVR/QFPUV+NtwhQgcm0gebTha8O+LpWaO64AD0Or3/
zPznB9fmE6KE62bf3dL7qBN7tlLP28kABJMQKutfLYttrQGQ3L1G9MdZji2+Dr5X
1vF1o1EGuZZS+5J0KA9YB2VYsP5WddTyam8FlKJS+tS5DUqOPJSLUcffAw19oxSa
q5TxusR5ZyO/92ymY+FPngTOJfiPJ0cQNmpl718XI1cJ9ZAEo3/zEkJCd/9jesV7
/1N2yxGdlpyFmTPg5Qwa1Kylfat4kR6/G+Bqi6euPhfAhp8bhVBpzlnlu7Y0slcZ
Mued+srbaWHqI+Xhqxnm4SLez9fjtv2Z34kDsFDLJw1xNxUwrVW55hgooIZi9/Lc
t44iNk/9yyyRjhxGKnfuYeMUoZ6/rnFm1mpP3ZJk6nB0HGN65MWMOOOJbtFy1AD0
/OADkFvAmQcncbzjopBvteclre8bzUdN/4qchdVe64msjMNbnUCRKvusoAJly7fK
btkHEMdjClKBn6WIY4Z/nUqsQWKRLx9FPvNvgx7EH5OUfk6WovhgWmZyQjKncRmc
4/BwFMoNIIzZOkpVq3KBzVO7lHzYbAU3Fj/93Sloq/lZ154UcRal0snM8DexaQ+k
HQCLeNYN4S3tuDlemkBdr7+F/xyHIM5Kb9ICldCZPkh2TYdFcplh9ED42RudSHjt
Ea3Oc46ck00M0nMps/SCj+wNinzxfyyyC31FrjExuB2RNq3xau7vAA/8dFbcFeZc
WIwtqe5HmoV3FFs6Q1xXTTg+obHOebD09F1eOUpxBOudALsqPYoRiM1UD4OLnSLM
NAsE93riWBTWGRMrCqLC47vUJuhJSHYmXWRB8ptkaOF1Q+hCesYl3tRBMko7OopS
zqfO8T/jDZWG9+AZ90wmhyWSqV3RJkVhUJN1NOGy7Rt2hQV51uEmncRSz3gWWovQ
LIQOgcFZ5JlSDYXSp3/FFCMTuKWXWkzalIylsTu0I6hwSDQPva1WU4qo8ofYe8St
B+jtbJ++l02KW/OSs2FDdoRJWHMUEnp149ylKXoSQwdmurGpBN6r5QmEVHA4+VP4
EL/QO789+4i8zeEXRHr1v07Zy2jcAg3dbrntc27obaAwUEzpqN/6Ugge194D00/t
yeHSEFU7EFZZlZ7bFRG7jGD7n6OOg8ETOWmDMypYwBSjER0yo5FWubGLVzGaP8um
3ZNnT0QVJicUkINQLGynUScwxA4/Lo0NMWUBMWw1M6LcpC7LnfhHWF+WxHe/0DpM
k6JuqfdM3Ndph2dSjd1TpF6DSg0/SHUnth6wZIuvahxf8GrSH8q/qyqt7+S7+U/0
mb3EYntClMR5Cio4sIDw9j7dMPJN1629IpMSB9egmtLBpEzO1gdblKd+2rBK9VKS
7ebLkRecfLh5Ou2g+QrmN8R7Zw938NR62OKREuu5sW7egoQrwsHNMljXinC1j+pd
+h1sKp35mnSwyPPrgimz2Sp1xTKTv09JkgKtGa6PM9QqL6vXaYdTSDWSkZL28dZH
YswXxTf6Kv3wr3asLxBIJrgZJYpgEo5k4D8VlhIA3I7pgFh9SahWBgHjILF8BS0s
KQRwdPY52kzZmMGvWtWpODd9ys0q5T5wsTtlXYxh7tsUIp/IjbchlquewEXEoNz0
/jIhgBInYUo0x33uQ9T/9AS8nQmZ8KiUE+g/yPBFV6sExaWtBaOXxW/hZtPKfDi4
hgj8PWqdIh2ILoDtP40tj1/trzI6fo8LrXko2PqfMibo+eFotvafsR5GQg6v+7xo
rxowUnJTkVsq9miXsqZx2gQeqkXtnjvnkh/FnAnPVI6mRHm2SzoH/7USwLkOxNJA
ykolBReOr14N9Grs4Hj3J6Io0WMK0GK95dTpmgXpqnIcw63+Hd1KYWyrqRJYy0u+
mhSOhjZG543Dn73YcQiZYrBdfA5uyCtZ6kaDTqr2IkHkFpAm8DrpmmUwVY0uMs49
eWWANj4q8X3ge9ay0tjWdIkiVms2MpmMJN6GiX/RsQlhaZ/6TOsd/+CWva2+ybG2
fIKD0duZoYBxPAuBONtq50zgmDogOKT+HzfRLsU+VXybijh4W/nPrwCi8oQWFdim
gUPT3M++d2IIWQRavpnr9FaTDgc801dQu9LwGdDj8MhPfHfH8hVpnesZimLUIbuA
COpzS6Jo2MtB+pyXV9VFtp1Bxo/JfwtG2Q5is2jDimX1P67/ly73NphqYYqny7YE
wp9BIis0Ac4paws1mfF+MMyNv53ETBngQ6do1PerymMfBzO/0TEnj8b8uvUzBSD0
MTHVE6gyxqEhY1QHJyxIvkROvHCnuhJ8TZqPzA7Zc3yMUjNq27kK+w64Xp2nOAfP
r7oXlN0jKvz/gERuDzHxNctGGgz0Ppd+OieXrUHsBzFpe6fr7p+4Ng8cRduW3iSf
kqbAKKWY8pMschQkG0EKZgnv3EIxNxK2QfzQ03KoaJ0ckPbZ7YIucsSXJIhzm3aK
jZP5eEsHe0kv9cNIp9JUqihGKcqPOJ0kFfjOKh6DLYh5sT1dhd44pqjon64laVwP
F/UHrCAjXecOqZqCiRTIKDl1640phD4WxIUJNXIIjgb9Or8PkIzAK7BmPT2zHezB
0hUivPHxPiCc1x0jDaJTL1AxXA1PhDWcQHm6tEZk7RfTteBtW6W/GYgcpJzX9qbp
6qCsQGfre/i8PHAf4FcaLe7m9u4MQrR837GxbzUWpdBXPmytdLXvRRPdf4PLm++X
wgDW7n6woMd9lQSdyo/NQIgoy3x9weLysQkkWK0qPnjeXlqvHZzwesAd35akFfQU
84B4mlCgvNWVGLxXm8VoweyC1+DgVjBaAuijlf8vtW04gg8+fjFdY4cGHNW3dlB2
qVwUKN5NDgvC7j0bTXnoVmNnlZqqEli0146hNhJG/VAcye6xCLZER0nowxOoV+uv
VoSnQMbNIfQot9bgBalLa581Bw0GUZSzaICkbMj2KfzKXe2VjOR2IICuz/RQEedU
iltqN8H06WldfJ7rLYZ2MjuGSuVpAVPwi5yni1HEIxLyJ61V7xZTj4pOkaU9/ykS
C7QDiTwG6X0SSyPeR9ZB3vbFTesdDbo31vse6YGgcPhMY+FjPYIbHwLN7LuV+yjv
0AQQ64qEJI0pSs9AJcOy0C4+cSQzA96giIwwXBRj2bei6nGLsUjHjcXUYaL36ePF
4+5P2zwC1LEsZMg0VfjZuV4tTE8VLF39m4SnjlU6Tc7VRSJCkj/NRGl6kOjxrtfo
tro2CVFk/gob7R9A/mmXdh0DKtxk81FZKl3FZtSoDgR+ve40dfG0VwD97GgRF3CQ
KXkNE+NdRpl7FirS1twmztEDzK5i7A2M//Q+uTpc3H8zpIQJy55YEPQvUSP0FqTi
FuedW8RjlgZ8R3ELLRGGZju18+AEkrM2Q6UNELIh+D9QYodg7arvuYqh6jd8evoQ
yu0Si2nXNEoLYU06mgTaIqFeMQrEmxmJn+QfkBoO1jw4FATMi47yJ7BHCM3B4GWl
0GG0NCMUqhR4GTm9pHDSfdyOPr2fayouPjp/LI0DSXZ6TeHxgH4YbY3oB+TkBKdt
TrdxwQdtmfUfayusXncJyc/LH1mZvDsvvR+VQCEewIPc+hfrLsF8WiWbbanR38VG
f2eq/z1mW2Kvt2SM2S88pDKfhVg+AANYwHHTlB3M6FwDcxTbVqSxQKG7WqZV4Nvc
6UpEeABo2xkAljyMcfFoTGDpdS+aeBo8Lz/AHht/1L5KREsd3XSGIA4D99aN9OGj
/NMvLNbjLFCAMFAHLDSRc7zLeBcEu/4aoo+X9IaZBCQNgrrq+TqOPJcBr14/BHGJ
qkoCEdqc35kE/nI78nemaXUhtUGP7bRPI9LB/kUdNDWplR91tMV/IQ7/EDzNkr+p
fBklCuthCyX5JviUktN9hJop8QOuUjkMGfBrY3PP14QX+Bj/1ksiZAQu8c3zvBl4
pv4z0nes3MSUOQ2eD9M8SqvH4+pk5GneSf0HoprqphaCyMQgVe4PtruWk6CgDxTZ
t7JpvEm54J/5wxzpEJl+b2Zm0hiPQhHojh3tug6IDSffZBynTqFDFvDWc/yy+61h
O3wJCO9JEPlRcUwfBPmgIMnMrk+lEXqnAanphIm1DzRfWfxZTmsbNrnkb3TzJZLu
T9v4AT1gD3yxPv8+jB+qfaStvqeEj27lRP020kqVfy7HZEGssPM9gdgd9oS5RBoC
mIaSGH76aZZF1oRJRYiwB5I+S80GZIxo4i4pUk0HXX1OntuZVGMJdnmu/noxHIYy
l92/p/JuzGAyyP/eEtZJGzF1nsDNMuCXg31xRuZjJqdMOhrM52XfLfYINBFNuRAZ
46bV3FccQu6hRY5N1TqciZ+z1amnTcx5j/QnmT2+S6XrzCk4cxwyXe2ODK7nfym4
jLsTCgP3T1EhphIdzx0PupjuXEJ9wyNUr0HGBNHd9Fx0By+LPTAxFASTejUWR8GM
hlOFgDzl/ImWJqliZPlWPCN7AjLpEnFGSs49hH9ZpQTJo57Db+nFqKciAttjWD2s
SJQhOiSRGWrL+7MOYMIKKAFFj5H/7QQx+dPGDZSkLDZak1OYlM/xdg7ZEHUPfim7
lkU0+ANevGM5hxjDf9+eHf25ACOCnTTi09q0J/E9FOS6XAaUQggWXtftSBMYjr5z
kyWJfvGca0Zj7pMvnK230h826zUaRncYWVw1V+hz1nsdwmr1GGJBRL4ePcylUANw
FhKxYZrqrawMSFdtORy5zAHj+x0CiLdeX7f7UElSf092HMJiYwuyZub5n8Lk6uFX
PtPQ3Z14KhJ1/0FSv12bIJzT0y4/LzGEGbuokG0jYV7Nn0Alga1yeEyeWbdRni/x
ltidpKFige+oO4eBRq8/yXznMzXYE2w7cSGNqPhLHInu3PJakiLA+Q6DhFxymBEs
3cPJE63QcDYfRHMRXqf7+MU7FUGioWABjviBQvt7dOLu6OV5FDRXndX/2tNqrTB/
IE9UE8SqiehrRet5NJGG8bnGoglv2LFOP5oO9HH4blOKE/Qrs5YNCrRxuLeu61Fs
PaOzA5adepYnWb4xxAc1elMc+QhiaMfL76fZ5q/V7SlKVhG+dkhL3ZOKBIoEoUHH
PZDgxLX7CBaXmzXpm2vRefHgXdAKls3erXD557G9nw+vHrSrADEyrWxzJPzq0QzW
qerbk8SvOxJPLDFl+LB5mpatsa4NzQsdqKqY8OQRAatgxU2DDyxNhu+COr3mKk+D
1MnmGfY7iDcpfe6s+dwYPSftVUQKg2RSMQTekpkRImKxV5Vhuk8Bhc88lfVd1fG1
op+AD7kjx6q4/vYFK79fPLL4ZINVNM/hYQwYtsSdKJpSAko2fKiP3nGtiRITwSCI
3RxM+Ba3mhED5SJeC4GPaXkzYsrv5vDVyFdBrzOYbyZqGxJopyUcqYnsO8QN0/w4
ulNbbik2Wn968sMJAnvjBG8gmEI5Jn14sV+uT17Ebso4aEnjy5d0QLp+02X0BpBF
G8tgXSxhSBEHVVF/X2Wd+xBeSVBh7HaJ9uIhVvtanWP3zviPSRsZWH8vFB0gm1aw
B8Me2rM42K/g3C+AHARxayGxnNWrkXeUFXrpo2zioiXyVOnNlKDWW/9tOsfYegIC
4JzAlr3rT1BU4hOL1MPtRF8AsOMpEr+RRpcOvyTH63a9JUkxKMDzXzT0hkiWXHeF
AuRbmx5QMLgha54AfSS2gYpCcfXGRjS0ErLNHdbiHryNHgaBqgEzprZ1FeVWvaER
FXj+23mOcrnvX0tUPRMxbjZNOXpaVibmqutLftd313I0xNzcYkLmnFUTDDq+zN0U
FBK381H9sLQRFjV0qVGa7ZVa9NLBmCTe1f5T1n3zxtI13r8T56oyXowTz7W/h4dM
+zuOQ6WMjhOJbLVmRnmcGkaThKZmsTjDh9Ge9braX6vDDPbJyUejdWj5aRh+GQpF
CGYrP5aSgA0OyAJ/PDN9quFmk00Nu6Hbl4wghUXMaI9xVUvY0PmIOQWV8olzXb6s
P7XIzvm4pu1ykmjat8T9JGOLBK+sbOFCbYdaygy0sC+Su1dMuRrq+IXoe3Z4HtE5
50EAPVU++5XOmAM7XE1KnutDd8nJL6sAn4W4Eb/AkTHkuWlwzyJsm4d0goH8L9z/
dYsrukG9JcXlYS67Imn1odUDHFbnHhrKK6DQhM29jQGBDDBGKRSYrUpd3CkD109Y
pSRYznHXDiQSt/oW8cQ3e6VcHtG6DTH1hdWOfuKYtik7RKXCZawptK4E8QOKPADF
bZ2jJGIRW8Rs+KhXv/0OtVNQhqco3v43lXyGrCf6E0PQCw5JcuP5LnPefP34EMoY
CNxLxhUxilKhtjo39cjP+ZoA7gEqYNmY2HkN6fgTlLu4s5iXIRqakGiy4iIFIuV2
4ejT5xGGfWRh0P7FuCEIt6cuxLHbq5TVpvsclSos5KS9q1YLMNukQS89Uzcy5YrX
bvoaovo5zNqeexAeGlOcVcuasXPujWl0FAfILwWagu0s4x24/67sSIUBlPXfduvq
mg6IdKuxjROvr6xSppM9x81VevRWvWBRMeLPjvLswBVXjZBnhJBXsiVsFh3TRk6k
8ef83u6wwaFlK5k7s/j0APX9362GIgUApsVYQncm5Ze+R1iBiY0JJN4wi16xa6cL
JS4IONdaegKLy5ZyGLS8UBRIjXX9XWZ1nOnd/BUBv7gedQjA+DgUslY03ZxVIPwd
wf0cnDVtg+cO7cznuysOyUnX93fZ4huIBbeo+V7CPR8oMHlGtSkyxkhkmvfRsw5k
5WYDpDmG0KZtJ+vz6DTWJGI3kE/ydVa1QdDOiVENTgDQr/1lyzLzhcEJBb4zmBNG
6bXr4QwogFFhGAX0AJ/Y/7pypzSXGYItc1zihDY7bqwxflhIAWnphkjatjmJoYsC
8y2FyiQvlXLGvDzlFrqZw9g3fY7P6RkVgHXlov5sb4aghR6kndoiMFzfemga1fdj
NvZozFDEnoGCrvlPBUEOvH58QVqt9WuZYfnQ+3/PC5MpnnjJijqtaaP+2zoaudNF
gc8lZvTxAeTxJip36AgIT1OoZdBKnav5f8BC3lPdHF+4R5CaSvyWyJ2+098T++R2
Ozf65u1J1CYGSYVDIChay1d87CbtXrRnBKJee3Cb9dGKv5AUwtUl3I+jTK70wR1O
1m8soMBnqjRtSS5cJCaSl2ayy591I3tOd4vGSscrJ+hWegyWyeq3tvLvab+fOpcx
9tb/fYBjoeivufBgK+SJo+N7P4155TmSGumzb5MbKb7y0xlBEZQ4BJBKMFEJteJU
kZy3uVJNUP++33PhL321hT5gKOynB2TwxpPeYp+SBmPB2+F1pAu0UxFwGQ/p8Y8M
RXUhaW0VVaHgv0ZefxPmtZz4Sf2j+FKvMpiBPPe0TeGiZm5l30vmSwUMsZmnJfTU
asfcjQXF9ARSL+MRY8UYMen1TJ4UhZIrR/916lLHuSUd1WqhKonqMdKPeIfdrwgM
U64EdHQU7mNZyHshgVZh/KGvcdAu48bfixbGA/nOSzgpWghldaTyhzfRuVtj6rBW
lxo5qu5zXDhJIrkH7j0a7Gogr9sHXXWX0zERZL0ws72r/WSmfNO6W8XY9V6YS4+M
z4wIdpL5pgNG4vtxt3hWBUBnhK2FTsycCqKqSnulHhTJky/+6OOt3OKXd2eG4YaF
yCVF2br9YfiWcKnoiOfuWl3bb49AoW3PcPOO768H2S/2hn7Xwl61Dzy7pSTGNAzf
oeUvCmUGdWd0PlVYZBiEntY9BREfHEOdYmqmOYLqgoDRDc8mkJUetJMtvDcV2Xtl
L98WhGmVp6Tb12WHS+mTvU1hVRHsJN3c+tT7xS3sVWf/qHx2bO0PuMKEMIcgDUd3
L3uEQk2zNsZBJA7dVxc72AK8YVoTud+B3r+LvZAFGhQ7h8KOvMJ6Zzpv2XtENZD4
IJKB4FP7TnP7sjaVdlOz0VTQXtc7Uv0wNfIqcep/l5tvqA6MDD0xzOlkC7ILd+lA
M5XZaM79RZzOMFKxtKEPEEcT36ppOPclQvDLv+eEvq6lEdAqESy0ZTfEi3USrr0N
n5Og1r1vflR7OROqdsWA9FEvVGLit1QIhx6lFQOlp5A5A+Rga5AiA5k4c2ZNpjTY
JWR+2w1JcOlQ5xjf+NVVaSaXY2fPSnAaHaeXTHdBOa7FSWgO4g66x+v9Gggj5uj4
V1SftQqR4611eqkU1bGzYNxg+5v2AtyJnRoxA9DXCuA7hbCtzlTdfydX5NyJ3XJA
KJ1aYDAHB4D0Ymd50uy+03tGmExCrdG1XF9m+Ec8lKnILgYJC0e3wCqnAaymPyDk
6M1sh5s+ZKNNodhAHIbnbyCUU/EM8oScNC1zLHXThGD7pQPCAax0ubMEMdxf3md+
5wVM3kfU8geSaGjr0yxkXUpJHMDPrm4d3VB2FHBJB4iQ6frcLb+eDdetC4WQe7zy
NKIH5+fKlYvS4jOxo/O+kdQL8+U6xPQtI+y7cMpJZwSKE4Qhy8ahGIpEMe2syzFR
0Yabgica8g4ys5NkeCGkdYfrkIZRoRnGDkpJUZA++d9cr1QL1atU3FaXfg+wq9fo
z5goXnUkl/SZXFPEtUHP1Q6uHbJr1CHb6pryWlqnhIu3lEN4LwizlkozOqr5ENVx
o/WLYWqyefukTKiYx69ps5Ropp9il32VsEq17tM495ZJd1c1WrrgudaLa7QmhOBR
GFwXq1rU7LChd+B9PF4SbXTtiHalI9C2oGg2EojrwPUTwrpyRHDaIzbaMdhlSXps
KlLKlC1NmxFQyVjUMFg6Z46G/KVuRCJ7cHwbeiRd4OeTo58591EqIFUMKs0m4buv
tCY4dQxyn1DlO0G5Jj78xRvDwFM7TgiG2Ub2hFOjXlQxAfeT0HIuuyIH61UA9sY+
YDmPy1UUr4+OzgOYUWPbQYd0tZa7GecdPXBpmr//uQS+7k/EMxMK5UCaip3dL56f
L3MHYYENWYo/gi7YIuDcKA6ammNX7anmjkDYXtrYWFFI2oOnhEih8OCq5h+yDs69
ju5mXa88ZKl5iEtx81YeoGkPVHfOytwAmgCkmPmE277nlhGmO/qKLpe89vxr4mxi
bU4rJkLy5EWNX/+khDRDLR8eLHiPy5bTi0bUG5ufdRdizYyP1/P0fKTiKqCreHM+
1o/4rAogY280cIj8Nt9ZdDlG10H4LUvvv3osjXWbm3LocJOJADkZl5+oo3MT5+Xn
bVIy8/5NzTuzSEbf2lWsCSurylGMfaal9F+rRUYb3z3c9MoeYOblUe50pi7OFEw5
oLH2ZUfn9OHvRdXeEUrOPaUJPHa1Xda4CU/WQu5ycr22kRlQwf93ApKvZvvYnf3i
zCOFy1Pxiz9tXhQizwUpBFZMfRdb+z0UT78sAOL667X6TIlwynJw47RPYsKf5O34
T8JWMKF4zGPGnGd36RfUhju8wpYai3JZxT1YfHV6rVy/BoFHvpkyzsWenKdm1KRg
yzG0ad0amjUNjH2lJnP7flPBn2P3VnvH2gjpOWkTBZYIU9nSHEZdbBmuR8PMACi3
3Wrw6UzSLN1l74VxT+2B2JdUmZCb8gctkS55ZzDbGPsX7hoA7yvH8uI62Tqz+G+h
7koZUOQLF/ezZx0cOJh189S1jipkiAME7NrYNlJGFEvXz5tEnAd74Nv12vAklTRT
QA3GesXipkQESL6PtcEUB48RzrKCNTdFUR78GfVwW9c2KJfTpRB/q91FYE9kJAiz
9A1uZ4qba5QG92smnw6gzJHL0UAw+dBExAuNeHqIXHhkjbrPEsyVeJBVZPpcU6+1
L1DeG+WjqtntidAdNf4mv3ke9fA068aBjmD8V8zHruVc+mtYpKPydzV3E5RmDQnP
IML7NRFQuLcgHfoAGPoMhBA+Up+D1AwSNiqeyT5qL6bF1+4uATL9nGoyvPzSK9li
A3qSl8C2EcNo0uTpSF4RTIf4FRtIFHjU3YvhwMEDwLjA+W55LZ7plkwbHTi3OTOF
oU/J0/up0nLA/A7N3kAiX1ZuU3MTMcACCFtGS1j+Kojjg9tGvOmn0WThVqXj4NUQ
dO/SPouWvum1noycFLNhFXoxBHj9NlPGJ++Kw7L3cfR05B/hC1YHh+jpJyyJMPkR
tRGNQtKzmvMaoh1oZLI0m87CTt3gh4rIffgTNdfavmYGn9km8cdf6ZcoX5S840Vj
xVL2MOib21pyhWVyP8EGATlvKFL2CntbEgS98bw50JKF/sIE7eV3gkEZz/+Oil9j
txyWXdV5pkrglTE4RzRJUBBGKSQzQkLcOjfp0zDVsGQWQThBhAuQMQ8RHFZimfhs
N0FkdGIeMIQQNjNBEvWscXcEPjWH3g7E0f+v5+EzDsxZxlsKb4becYqIFi9RFQQS
lQJv1ZoK0v5K1BeRu64eVOQxPyafK9rEXgY2iqVplfK/EnfEhA/q0hYepRyZFe6E
jc+7lsBOCSu6aeTOyXOTZhiPfpzROlPCjhkFdD4smx/XaXuDmEwL4NYJ2rMKNEiP
TeLJE8P5TnyGkhBTI7Pk07tZYhIY+iYgPu4AdlR+4OcoPN/LtGbVeYcfdB9bt1hg
wetuJpH/TG1WgUvsERw8QDw7YeQCdX/D5OFXb5agSBio2C8aacKU8Dsd5jFdgc78
EV81md3MD52Jlfh8wqpG+o0rpKMUSoUhdbPM2yUl2ac58mcwgBLWiKTmUiP/wWIZ
XRdTY1t/mq5Zr83xFL/8oF8kKuVYQ/K845oJKVeDeap3fIbQTNE16iqD+Ylk/tXJ
/ew+MK+QCVL9OsFHaL6oKzBIgrszWxeGa/dTAFK0ssO6D4mdnO8j/KSQvaELKCjF
fkAuotf2glRMxZR9upTgXniLz3fknlOMiyMo1JQERapPgEgNktSDad2GNbG1dMzX
S76v0ykoYd2qsBN+kewat56Tz/Yq+f1mJhIbOO1/C4EO1+pm8lFTZqh1sTZqETAB
7g93lidgc12bcz0WOXlDpncDf2LSfgaTsoonftKgS4y/GEh9YP5g2AZcOO2HcZE3
S3GfrKQfEa169cRsvEm57td2CC4e9z0DLywXX2tcfsppySZSUBVQwGlkbqP+3+bS
7TJ4eNMTkRKPe4aMrAHTvj/RSxViB14CYHRwyYh/d3VX3nv/IT8QJU5Mde2lFIoO
Lrsal1wtR1XDkUpthLgohKlrpPMp8FVXV85iZHro/iu5Z2yZqHkU0Ha0G1JetN8S
n0tlfqp8Nsh+afWifWkIIBRn7i5UDHflLXtxFHp3WwU2lNFbM6SiQ9DJyrBvp4aV
W0uq7v/gAeFpqZQhIIa8SgzhYTZbJMPq2sMQjPpgVdzwMFeDfIRMkuKccW0XuzcI
a3oEf9ScnwNMo3Gs6W3fs1VcQqwYvlNlPsZCyMi1ByGw0ULdaFICrhR/dSbk7c5Y
5nvftxMZkXqXZpCSF43V703OpMmHN8WONPu3CdDueB0CsVGbebODrPcKVg5FXuVi
xWoF1wltpG6pNui12H3P0R4kpoG63CoIHG47HEthTTO7MNhmRU9nA7Ycxnykx3EM
oFK0ud7aky+tAG6HhgzTg3Q+8sdaHuGMoHC9r63QscmnndzzT3RWOPqxkRRDM5m/
AdEpMjqBuQP2cWeRWzidtMW3QB47k/ChkdkNZDUEJmmPKPcXnXDLfLj2InVZMxDk
OG0jwkPVgSolTGzZV85T9bz7vjJ4PR3d3erNc31pUaiwDZp3AiWsWpk66qY6JQlr
8EUw+X7v1Cby56SMrSKKqTqA/z94adE09GJJLIthnZ6vHlp0AHZgp9PNU6EcIca2
sFU+JetIAPJZPE26AtUljTwimrQ4yJPK1+zkMnyA2YT/M3n5292kt1HXrPY81uQi
564hzHFDkzrU3gK7JbnDEB+Yj88uomQFMwDaPlRg8wNFRh5EZaqjzmJ9zKJVBQ6N
G4vzvW4bawBVsqE6SgMeb+xWT3kYZUjqjc8JbrPoxHiW84xjS4DsvBndMF37oI1w
TZyEJrLl6hK8W2w9XqXVxJhngV2PHcopzh/S1ALW31QxdxhYqIZ+Mq5V7/lq2glr
J8+mQ7DLz8EDGhrAl9AfcPZhoczcysaKSwe/ODo+QApnEnW+PsK1jdu3QV1dbgJw
FVc4KLEBril0itO0OTQjVXR6cFfz+xU2aSCC3ZGGzWC/z/+07/xQ5q4Il3CKHaq9
0nxLfYtyH3FTC9nPjdP2YBreD4nLF8p+yrfWkmHdaDfKEVh22X+6krk79eOLF8IP
Spx/Kbhjjo7jLJ/J31E1Erc1Titkv3FsW21Uyq/vK+GIFqaC/3qv3d5WWNnHONln
plDxwhSL+YwGDJJ7CSn22TwmUIrIyJ2zlypi5y17FwYUsFAwU0Fk2AWI1Sf8AybC
XMzgeWeM+GJz4DNF/1n9n4o7aBGeOaPKgZHBLCQWEVtA7xc15pun9+MaYI6dI7Ne
tZtbnEaR4grCKsWTOIP52TIS8B+LSfcUJLY7k9okSg5r6Q5s0Cu3pbO1pzZeF9SQ
dIK27pthlXR6bMcH/fR1NUdYD9vwu23tuzC5jatANZwL9rk/cQ1G1+da7Ft8NezF
61D2coRe88kezhUq/WRGD+CcDQbCzQ18kuQlcKILdQM1MBpsJKFB/+bJFeGOQiB8
rthc7/pebu1R+7M5Bq5Coj3vKwBdYYPkRjh989wvxS6Hw/3GDq1c4THoHuO6bDIQ
uvAvyyXs/aOaylhDBR4W81xqfCh4L4VfzvJvzn8oy2O2WgN8GhWIkcV5vP0FssIQ
gEzz4EUvdqWgUoweJMleK8xJuOTgBxlD3oD0jJvvmZP8Vc0PGn34sw61r0wuNTfg
t4NhJzZTl5jop16jPEeaGUVDjjUMgpsLu4abEzKTPaJ6ZfqkQrZKfa/tlqAYBYKv
pYNOWILgs4Bt01K7B3EWaBDQz5Vj5iUB98BlYpmQH1DDyfVQQszz7nfa5wlbzWrg
ENcIsRJs86hI/oNchI7eXBGiNq0ioiGYvMMGnqKAv20+x3kzciGKEJGHXK2S9Rxx
Zn3ABYXOU9xkyAaDYrmuKUIWbcWgh8uLgvcsOnQYI04M6OXqbPnYWOOU3pusdhVi
xpTasJUQ+QLvFVCc8zRx4wzbqajuqPn/NNg7LdfJk8V2gLMxCQqUydAI+tEyva36
1JDcUMgQNczmuFIa2QYOiEjV/7Mk9UeNtuoTPeq/r9dmt6+1BIP5ec7QTGsBfYUS
VA0FMwK1qg1MKdXE2UNllgcvl3I/vv6UAIWdCWNfofJbm0nj0tNhSKXMpkNrC1us
9yQiHsoRVmXtEqCPGy/Q4egrGij2/geoGwZK4OALG1+SweXYXglIzg+xgFnMKqfo
JV2BAOUVE7b7SYEewsxvpFS0w907C/0SjAJrs6U5X29faRFTyV9HlejyHjDI9vkw
RU1u2qmxLu1KByPgZO8QvfxhTFv8eDL6BhDguk8Q5AY6JldVcH1/OOC2dho9HEcF
yIL/+zBTatjQH00ACzM+MQVXfKeiZpkSrUjeTkFBVegsaN/WZ49W4RLY+qIelUnI
qg1e/YGLeG/lsRQjX7sMEiTBo7Kgr+8l6lmfjwqNoqyPP4ftMRZzQ1WGUpGJ+SgA
GytjNsGjvO/n+HMZWsCjsZBZfFDibRy3/c/52uzLsCYaKygAbeeRSsts/1ikjFMl
UtpgCVMBgAJyap+V3x5MTMmRxX+Fmbn5F3f/mzuDl08WdQ26MrBziVuuphy5vpoG
buNNQCwYjiYZBw651FazHP5nSnJlZy0OU+mwGNmT5levPrHz2RBvdtr6kK7gVeDT
A765/mZusV+7Wcz0p9agM7F2ibO4bWO60d3Gb0k89dhqrD1z5uMsyJaiA/mWRKOO
wkc9M8vRc9S/MlSC2esQ5324BbOWB2Yy+hZLVRJzPPIsc3H782Mklux5P+HEeO51
IQARcntz2lAhAOd/eBAVXDKYjO55hsFdJvuDe60DsyGYSuUAaWUBs3/IBWREsLgn
CNMPRCZRHgL79MuQMY9xKOvs7+FesP3r2kfyEq5J866XCqXHEopXjaSlvBCAduSM
iAJnANA+pR48Wu8Sy+Qc4m9l4+GbS6mp0mqHo8IrvvUNZDSMEyB2tl/YhFW00C3T
4S13bUD/w4wEZfEYt3QV1PxX7xvHNtUBHz8IuZAliDmzKUIujHw4MM7/v3Fj+E56
8OqMdmZPxjUdP9W4rwT0pW+cPc3gClZFk2cSidTWb6TzisrVyi50f2xGs2dIEM4X
fCtBOIZsYxdVX2SYpGLcFSxGo2YWgzQ36EJwbKSVfmcyBwr/vOPlKxIHJoOdF20W
HMyXdEmoA6OQkEg1tw9oJhV+Mcube0NuJ9dvFRR7WO1NjN18HZA+2C1ouAd300Dw
Sz1q4VTr2tIXuehZ5MrV5sjofmN8NVGVcQG2rr+CD71eTyScU7MoB+9gaMl1za/J
6vpdzTeL+0L9SJDupZkVu9Ruu5KyoYnvQ21QRm19UxGaQ0TbQ4+2SCk7+Ou2Mzmo
cfH7By3qJFMksPO3qglAzLmeJkLlPEv08Qx9qI8nU7Np2PDYXIt6aVt6XmiPKP2r
NsenXK3zhISZ5TFJe5dR6U4XIrbqX7budtbfE3PTjm6ZZ84BxE9ZfQ18XMZoMn4t
H8QTNHK33bceuMus6nuA6cehwQ3fNm5SdYhmdzcq1xUR4CAvWomnXv27TovmI9YJ
jRFhlaoVyCHDyj/FUcHRCX5uaGXuHYfDO07rcaVAmp7o/0zfIXPDWwbSEkzI0CBu
m+xY6NR4sjCCA4HTnH/8MWsCelFSeUkRw1AGYjeOyt/B7MKEMm/UXL1CPykkbevf
X944xoYJ/i6CA299BWB/VcFpWXDj7tC3MWfXM0U2UeUjnQHYocIIfkiomVeKFmp6
SfZskyqhv7BxQ3wB/Zg0yVY0+PNkxyl/UMcMpvFrSeOq0DPl51vZnFJfZDfVn8EP
kiOEPh91Ip5JHWq4e1mqBaTR13ob8hAlAtXWacfZM4F3ALuzPHXc2KofO+FIK5Lr
d6vwqxj++tyY5d1Ecrz+mQFSyHtSW0wtfCraU7hf0GvgXQ/mzIF4nH01G6GKcf2q
LxKLYUPOkkaGoNrmAeodk19MXZ/RikgEIF6cYiizGE3ij8Mg1xA9O67sXRrrMArn
aUO+iKOSXOwz370GJzh4P8stKfJ/1u9my4ZHlKsBW3ozo+WhR4MjWjcQxletcGLt
NTI7XUDI6FRtoBtO387rHZM4LQYlc1OBJ6gVdCjePbfhm+jlF///vlcUYkRJrX3H
2L09muzx6OfudSQMgdofNJf9l/Hav26BAkjOLKLvFYvwQ01mLSs5MsJ77XMPMJqf
5QJ0qJHzIt0DMY9agGIlzaHdRVHgLTfM3X/7Q9XtVNyaSjmh8lMHpPgjWwa8f/Na
3wHesdWks9GdkdyLkYK7YUs/T9WTH0Sg84sXX90m4Rf3I7iPLqJ+JRoXwUOs2+QG
5ZsZTN2clLSF9QmTDFYNIfEDaxmKtywSB9WOO6GwwIzKDSJBDBYQdKCDonXc9nht
VKSSb2Rnn+jpalgVTyMmhr+WK/8F4xYPuDPN6/h251dZPjvTQwzuyV1WvrI/DYyJ
jNbNuTs33kXHbPqQesv23zdjN+5BWIN8Onalya0M7Uie3LcnO3GwAiiudl79W04r
eJ0Pwq5uL1us15MnpfTYrG+jJN5nu33oQ7lGNjJ0fpIgihKDQyeZQy/Ldf2GV6pQ
RvXDPNfEt1lvjp9eAZAnXuJ5P+8TKT76auBprPBmrLnR6nYb6ImZxW8fZjf/YBQG
UggS/Sjjw9rVqNWUfdDc6b55TOcscCj6CDiJyzhiRHrAdNIn00DvBf32b2dM8JDE
jDGZNIsYSMUhXqaSMxXIjKwRTZRSYDy6pvPs8rRmDfPU8fy5IpPV19vTG45NAdeo
cSTBWkkb4+81ZXn8aReJqZOO74ZyqBlnVorUAU/nNSOyjGTzbJQyVLY9MKlFKsHr
zxy4R5wrV9gCYWMTS3assbjbH8NAJrqcoz4DbsvT3VmnHUOhl5a9x9S5qneN0TMP
mF12sw/sFNsUkILVyfjpxSI3ICDVwvRKAIp2MNGpNiZW60VHHyQ/RlWQawik/Qk5
EhO4j4qZ5gmNB69WCKgyGV5ppg1PJ0xp4BoIPyRA+CO7Vhr7052X7giloSTMOGmt
r05rHHcwIv9aXwElTDP5lAu0xUPRH4UqhF2GI5J5oQXNgLtkkTIexE70fYyPB6Pk
B+H6E/+2K9pX2T0KwJwMZsWMgFC/loOZzsrg8Gs48coDQq3hzszmKZGHFxik878q
coDfASfVp47+4snqJzi6ZyAGO3eFn087zMuehXY7y6ySvPsiez9AZMAwgGOlZMcF
35rgUgYmyZAGMg8f1br1vTF+sJlXHN8Gf74QddCQxpp/kMTp9m9BXBy5C4Hg0H3B
Go2k4uNNNQnddDofFOpJTboiE484bcLGNvThbtG0ZuHWd3KjBEJoaXzf15URhLYC
qAA+pndsTgegYFrfaF8f2FwJURkK1QsmHYtG1wJIfjLx0OBDBpEHAmNYWqwwdBYQ
HZI2zVaF7VpMMLwZ8S1stUe1wN/xGAjetR5bMAspXTemVrlQVROua+N9/mKri22v
rL3ZPj4TeKToHmj9mJojY8vXJN69cx7IYooUM4NebV3qvo2MF43Z3SuecpON0Buq
WcSBG4ZkiWNodqMDLaP4yOsHoUNYwF5C1eAQemhX3CyCZDhfhsZELPT4SRpwncLD
Ydyw4uAOe7TcfeEE/0wzOYSP6pwb3V2CPlCAmoYoZE0Zt82oSJONt/zs66ah/QHH
Eor+wTjbob2pbHE/k2StxSxxrl4rESXN3AjZoDcLvHSgtHsBgOOB6Nx5meu+tV5v
9CPXULtrJjEdNe/v7Rclo5va8Rtb+L/A8wkTmqChpFdO9dHhMFSe//62NpVR7Z+/
f52K/kI5OmE4EyOdEsC04+uRXnZ1IcCUn4Hu4TvnhIS9OrXAaorximJuoHOh4ASE
Wh9Vg1/X5o7sgQgA2oodvj3jEuhBE3fDAeahLq9uUoIgimAE7OT6SDQjOo/X8I7B
1QfwKpuE/hBXjJVxnUrbRjVPAL0H7mqqd3v4LPCMYJHSe3vUEclSCOgjOqzVqp1v
zpe85pecXYiuU/zBX/qjSIX5gLmmrmtdEdQTq1JZNRVqORHYGNb84Pe+2hscJ9SX
jKp/2dYEdNFC4hEV7sK05AHoAa9M4L3TFrVizv2QnDhA4t5E6x+qmiPC9K3jfOZz
8mD9X32dYYkLJoq3bRA3Na+suSvGN+W8gZNvNaxs0q1CUWhpOisKjX5AJ7Hl58Dj
7jYoFxUGJjVKv4hBJFN1fy89W9j+gT7+WbvGRK/C5VvVN7woSh0GOWNKSn/xXmU8
sjFzIh7DNXQh/xpBEBWWcxayg/xew49p2Qc7mv1slnMa3O9aMvdS8hr94Jh9IDux
6wD3sojqB7bcQXq7NYlGRmPFbb/IKx/IbIbiF9rSBhfSo5zPZHuOGQyeHiRmPLVq
pP1fLr43LSE7etWtZKaVDv5K8BU41viH80r74K0V5VEKfHEE/Ji8gA9v4xX3rWZp
vjSpcB0WNiXSBrHw2JxWyiDUPb185guZkFqgdWUJ0+HgP7zrYa/lezpFCmxkEK0T
uwXvw7bHOGKiDzJqi3G6WpeipYMkuU2+8m+V5+Jmr5DY+nSbORr2eICEEX7X/c1M
vH7K3jiSyfi4Qi3nyOVQAg2oLJ00DDnPemILUXJGiSGeSmY1IDraTLIILuZxh07A
UHk1kkL/2EXd+dnYtMKke3TvfrVUWk+9XaIH/cJEuqSOYpDzeeOSFVlTz6d/S5Jc
gEtttoT7spqKuWr2FOyzqSK7n1u2Ug+JXqdV3SVIHedZqKJchz32kND1gg/pR2/x
Yuw+R0f/zGWQ9dZExuqcj3vRRD541Kw2kkjsJk+1fzGwhycJkqiHazRctalk4NPa
ApIPUJ88A1TQRvpMI8wTxvq0ihDvbF/bGy7HZNVMrjw4+16oCHVXeOKHNpaZOobr
Vxf1TBkLuIhi09RUtzeGJeReRXkv9JjApzQrSmeL2HxHX+kTQmXqixDjDzNa2jkU
IPUZq47tiazCrWYLzHQr3YZbbziJgj2H5czkH41qd5Y3hLfOkxveFvoO/N+c2HNG
Xk6fKoSRor+TpPu8tdqO5auQ8wEUnj9UJln75V+ng5p+baEp6G08d2qzNt+Ghu+Q
jzfVlXGyBqx2JYCryEvmS0q7mDVLhQc0Pd12thnKspL2pvmdsgAA2N2gVC9T+eF3
Xg/tvUIAeuJC/Vl9MWxpHsCjMT9Snxky/qJVtbG3TjVWGAfSsBxrNuNdxtdDMOrS
Jg6Y53Fbv6w+e1N4lY5mWde3HLtLlmbdtTZy8QxwGs0pbkpai11vdrjWhA4+3voN
q5mN3+ZI4yxWo1apd5gq0xB8MxlU0uwJY5vqe/xwb6K+OEjGseMA7ClOV6bNnahJ
bWCpfMOcDU5wTSQkxbE3mWXvEWhpP7j1Ua8O3RIdnYxCFUhuxHfMH2MMnf8xBDJn
YapttAaae7pghagmTNqg35wrwBlPH7Jr712InPiRHRV1JY1NCMGL+mxYUDeYxq0k
1P+dyJewjXL/urV9EcXf4jA+ya+HLykgpMVWCLZOUp9ZAbTm3bjakStmA4UU9yXZ
DzfA6Apwns8QRxs1XElGaUF2HaH9MbZ1NjMThUY4EH5Wey+zC6Uav24X0nS7vBYg
C1+RZLEnTCxww3Jux+qX6LjTrV/QvT72a5VGjn3nbRyviNcVTOWdg1Lj/g7f6i3c
xzoBtygaQsAk0/yqWYUmbsftrpoKy33DV+JIKzo2VRuekDjRoY7JMRn4BXXbfvGm
/mXzfu9fguVOxXCgdNNLM4oUjS/yHCgpwxmJxv0ihNS3tqcF2ovqHecFj4x8Qy0p
iYl0NK2qigkJDVAytic70lx27UfbKmg+bGorKVf8e0NC+J2+Q9XHQWrRqz/WCAYm
LA8i4BKe+pAN1oJmASnSLOgCrC0TbhlzvAt9aG6u9jhK8kUOCvkfBRC2srJM3OIr
62ym2FZaHgy6Nu/xbdY002Q0hT0mfhqwjoOZXEyzlZmKWjk+pjPZOSxkA5mcu1dv
Xg71D137cJTYECh7tEoffwbGfQek+xL+FjbTCslwpyAKbJLBl8OrZmF/3dwVp97D
h9VKT1UpfOUDMjiLrLTnjuorCvU3QUCNDAXL0yWhiRNOfGbezY2Dj3AWoetZaU5z
FuI/vil8wrNPW9GPjgFbKGI5AOSlIJ5Bz4qudeMbBrUA1+9OYq0Q/6M2VeRaWvTn
Wgp7ZyMO9L+LO3U5gqecjKbGrg0oob32zlnAQFXZU1XGy+FhcbJiQk+QqtY7UeUH
vh6UdxOPWYGrVil45gJzvkfPnWmTQyjTgl0usDBqJ3C83wxXsjTNE0Mn/u1K2CIO
fZcsESAm6YlFku3BxBspWAC2wwdhUSS5MuNZdIQVo+gWI5kgSOxJo1XqkiDgFU6+
PUHP21zTccOQekNq3D7vL5cXh1Pc6HVAQPiCfEQDrCADUAV9bjy1UAn3DQ9PWQwx
/JE38qbgLzGYXNIVFFGD+YWYh2xgAjZecVVT5LfQT4pnsYR5N8vr7eqcYcQCKV0U
kzHBZ7il1KEvKKB1PWmilmOx1eeaId8Ao0YC0KO2oGPjQkQzRJoz3KXgu9D0W18P
H1h/loSQXcGIdQ+Dqx2GOCgpH8WK+rtevnfZcL5GGTplFy8XpmOXNhA3tMpCvfIh
2BguU7P4YF+lUHzSXhxJmoarm8ym2H5CN/4zxMKAuxcxf903fsNh17q9hY9Sra4M
ijXFe6toV+tpRRcrr6XSxPhZDUa8Ykp83qmCoP7JiyFku5lQX3r6Rl0im2CuHEEu
3UqalrSB3rKVEH1lcErbJ9FtRBZryenSc36Sr44r1t3JuSvUKhrP4BEhZuCkSabS
rlZNB0n10bbaFspFpFYe9i0QefoL49mWwjve7hN8kNkyBD2v9NnpGDSHbO5tdWxI
hhoO78gHvSGQkQlmGWJFzzmFSnUv5KXpLQ0d+gvEIqKn/EzY71RwXxMmnfKyOFr+
d7hEW4H/AO9xPXvTpbjENY8YhW+M88Bz8mnAI+IqhM1yj1jJxQMdwiF4jp5lB8lN
6ntOmqkemuEDxPE9IfLSFKNEG0oiv8jg6xMsT1oKCNAAyFOt7ytqXIPVe98VQeAf
q9FIoHIhAeigmxiWPQnCTraG3JTnIGEIF4uxGCYJ1DpuCqku5mt3Hi9A/Qepg6LR
xG69qLpqEuTocF5RVSOFB5acgdHwSvLcif7LpcgRID5CxZqy3oNOd/i98Vv1Qlo0
xjP37SMANsuCl96QjZl9WKDedrZPiyHUdUufRtZDkrojRpLTClPObQRHO6hIegEj
o62lGBcktGSDmlmj5k1Qzv6NEdLa6DV5WorYdBe4zzvL7iqtx+Dq9NrmxsiauFTx
/lF9dq2WnqvOeexgJ3iU9iEGGZrwzgeDJm4r48d1soxrhYoGM9kNZti9xcLXdqTA
SfZ9F/qd43p3CVJeWyZuFG452qeHrsO6ZPAKwxl3z7djjp/wkNt/pG2lk1mS9PP/
Rwaok6/0Gd3oNv3px/WiC7dqhTwT85OPE3iNvf2Wi/ZVVDNZEM2lJQSe5viQcNUo
N65LNn9WDGkbrXG4UzarP/rcy9e95UT6f6MGMaNDo+vMO1v8rL6w8YZYwIunZf1+
kjAmJC1DvGoRaR5wUXV15Ddz96KtjbyraSx9porSZHlQyKmKNDWSbAGdt7Zp6m+b
/014vJyl5HYnGLq39XqnwdIBoGGQ71m+Q9b0n98oBYjz6UZS4rOYhVL9jSgK46KI
+yAJ6Fp03Hx13ecEvsEF+nT5kSlqypieau42L4N6Ze2Nz9vOvBvP+urLogyMqlSP
IuN3IsOVJGhXtI5YihPsAm9B2Nr3uqNMZ48iCGNM+VodGeVviyvM7rHM5dj3SQU3
2osPxI6IydBKzfTDhKcAfghfQbjrUzpcqUw2gDNnD16HNE9qCUhOr83wsF8kFWcJ
6X0fGoSIAmHtVEkgjqIU02Z/IBE2ogynmPNxwLKOLS5bKmQqARBxXBwF+L4KJ2Cs
WXKmXh1CXG56DpQVoCpA7wvZTT9dYvVDZ7IwDtNrU8lJXFOmQH/Uksdgn+hO07cL
T/empmgrN9V4vD+YMtcTVBPeKVXf/ari1hK98Egv+wslVxgKtO9dLY9eeW2vy0o8
L3e4qz4IPQyKZZ2O61G7XMHlcIkW7+lI1kSVlvdvfB/CW0zhd2DERAm6ORzeVM6Z
BqRtlkhBgji9WA5+pGflwFeDoQDxMKU7ZW45TLfZ4lArZfLNwZ5KxSZmO+4gTMJM
Lw1UMo+woH0RXmcz+IhRWIf+tIBiekdYBzlHKzP1Y/mBk8gMknnK93/hmRrxhxuK
miOMsuyrYmUCwTEr7i4AF/Po3HhYIXjgMSWWZGtwjYUa54P4aLkT27nb2HNyOe1k
+dwygO7p835oI7xeAOgCEK1c9dakbgjINToiV/nDA+Xh/qfQo5EDuxADi+ZDUoiJ
241stoh9ZchMH1T1Ql9FvoRJmwdfJd6SsV8g5bIepJ5yYlWadtGH9h8Hk3KRvN4r
yWiARygRRDlhkl+7N/s2yJIdei6748jFNLzvv6Fqlu6fWW+ubrejPKc706f1c6lI
4Vr9VPNlO3sWJLrGXFvn7etP4ai2GmQ/BccC3/JCC1TICd1Y9DIKg+27AnlvCnwm
GJ9yaLOQ2swDKamguU2/a37z7VfeWy/vET/BSTo/gJrU3J4a8jwtyFhWJmtA4X6z
nThtNpzKRn5OWdaNof/kjhXUjDwkIJmNfXbbpE9AwdMuJIe1xj8IIhMA6/fjZO09
9p73Y27QF9qJ1FBSL1CVvJpiaMfC81u9xD4ekt8AQEaiZhv96SjbuuQ+kYuPg0jP
i8vbbWvlD+lY2Am6pzupCWrMvZAir2yCVR6IJZDdwKoYPRGnPBhGKjCPXmrKshkf
ljHo/lHjgCQxKyl73U/Bh8/HIMRvOjZ48qZuXPDSfJeI7McBLKio619nOUO4VqTy
UYy7TgbyP9j6hcMhSfk9Km+RBCReu7BQ1L0oqo/xkvIP0T6+H7ZaSzEXp4l5ir4b
Ww/R6mhWYUQyxctHYKSa4QFqOnbAf3fuAc3XhqmIaFHff0l03iKf26/2G4byS8iB
M6saIrirt+TxSFtGHHmKMILYxdw2ExvasaYHclxwHlbegKd+oYyzHoAKLEbeVfxD
UuF8Iavp1RwcMx0Cs6sLNnmS3Xaf/hYwdvQ3uCSQPOujxYPyy5sJ29emBYpqrOrg
W0VIqsPlAlyGRXVFqDsIIIiHR9fGlwukxHyFKsfDLGnALeSfCmaEz+DS6ydh3HK/
uF+fPaq6wWPh9Qn93eT4LWGaBpmN2qJB/LQsKufMCexTKx2un8pftmDxLOB2YPZ8
tIUB3DEOyp0MVdbyb2+XxjZAS96B1Ef4fmG2yLQIwHBqqIeWvswfWWqi9NR9mVVm
HvlL6sxbf+YRo2qADuqfUpxcpZrhp9IgxnKBSiFnJHhGEn3ojYSQnYUOTwHCtP5V
UgE9Hc+dyXzw4krSmF+Z7Smfl46emskbxGxOEhuuQPm0EcwxcSNOjUGjTVXch4QU
OLYMT0PbmakWkSnC4p4dDB78WRz3VTJurBzK9vLGa8iKn5f9D7Ldx43Rwb1oF2Ct
Q4BGa4/BjyJFtI7e/z55Phl93OTh0fXolcFQjRV+oKmNMwkWZ8Fn4kSk3BdC7MVb
TjSloDCt7je2PTmHZtcDyV93WOB1MLLbElu+OzllfCDbahArtbb+Jj732t8g3BKn
Ht1VI6wWjfVXsq1BE51YJJjH6y7xcAXhKNgoagbH7HvVlAaM2WvgsnSrigsIiCWP
Bo6/eXEvr3jJ6W7PGhJe2eECPXz98bUYLf8Fv47tuXobRPuLQchY9RdsWwvqLXz/
jacCEKXGedH+E5jAAx3cQDeSLBK0I9Gcsz4KUIqXn1N/nXIaUEcS8hrf+c1Mjc+V
7E+NGoUiknlNhiE+pnG125RU5Si4s9sDyoXvqfNfoFaN0pPwPrY3rw8uTwXMN8eW
kddMkPo04Qtqz66fL4gD0bRpl4ClTDxcBlRmUUTccAXXE4GeRrW/2LALUdj3kBEW
RgTThwOjvrUjdDVpDgEJVm4xK063U1UuzDkZq8qMVw+qPqkkAlKNS06unfl65jLp
SX9Z/gRx1m6kb+i7Ka88w0DTa29fM/U3v/GMhph3PJN3GZimWbq5AHJf25xmMp73
ArarmwnN5mdNSR7t2I/ViOzUYljwPMtgLltIj3mGjIl4hZB+EGN3Ke/i0uYBbCiq
pZC7LKpsqQCSgFT8I82m468b041sbFxNnQzyDdoDtDsfTZ0gjfLmBkL0JzS25MQZ
AupcHtQqL+WRnMdX071wMhaoce4BMqCm/CECJ8jPWz+EfOO4jHnt1JPm6w3R9kT0
REXr3Qkae/sLtzEV+tdeXTr4gIYl+EVBzLFG3xiezx8j8UfNETUM2OzkTGJzK/VY
vCdkgtLgXA3O4Jvrg0/jBXH+r1AiI62kGGBU7HjhXOWoojVODaCZajaexNycQbsQ
8OKVyubGnZbv3CjLl94MJv3AIVn6ttyl48cyldqF/9J/jfvhYkUD133+WVT8EZZG
6e/MpyniQnM678wl3frbT/Ad8LNHo/JLVvDANRG4SpktIfVaVmaH3Zwfq+LFPRma
RXl23oDESTajt8AikuZpjILf7fN2ADplgumD0UsBh2Jy0hCI3bNYDToZ8SAboakU
hRK4/XJDp6FtnfqpCwnTUVjODOYJF3iF0Z3EY4ggsVNs3P3ePtlLusMKZVk82PB3
sx0qw3ymsM8CKVYTA3A39DK4nYvAhVHOFjTee2BRhOObZiZM81RlDfrQCxLbj5Xu
scXRCiuyIixdtY+8TO7mpH5ArlHT2QfT1X9Mfm3cD6Sh8I7Ssa4aAWwrkDjyp619
1QCquqeOPJbGJ2fjUslbLdxh0aI8a38s5AW4uFon5WLvuIgVGy2p01aORCULNPOE
QhQCmKE10ckxC3VbYG60xYorWwInZZlMq/oXsayT21CUSjSYf0EPsC02cVFLwZ84
GA5cC+5vHvKdFj0NgNNZkNKfhdCiyXiK2FAYgM2TlQDbTkG+7BXNdY5SbJhVoW9o
nC6603VuLSO2dMEvx7OiihULpH56DHjMZagSIIBKLbZa0UrXet/T9mhLkSCUYpkc
syY+B6Zd1iaqmWdCc/MJPM/EE9N/OlrYWYQzHl3gdrbPWdCg4ksm6T0OzBdaRZOW
ctPcMfoldfiE9Be5tWfV+46ooH0QoX9BCS/kcGymjQKj5su0aLQUjvQSElNY8HZR
Rbl+vovwkXojKUHfpyXNMR1VlcxHgdksQpelbDpp6U3lDJ6sLvzSL8KJGX9fIOKw
ErqLLSZN6jNE4ZHnEg7+nYPy0Qf5eccTUGakZG1nk+vyM0chtxfexOU2KFfjGZvd
zsNlGrUcNo9fHM544bS3PsbmQkBcRu+TITVjsVETIDrcTKFOsGyGfKmRdmFdLZIx
nFx8PCXeAn7IdwUFc4+ZCV9seaGNr70SglEeZyvJkShcTn2RcK3ZdUtXZQCNdpT2
Q/53SddEY2Se4ou6aRytDX+hU8Ese1+Q8BILMw1TC+leNyndp8cP1P30ZQ2N/Tmp
zC55aiYYQ9E+bv0UT7lIXVlD9YL3qHMjcPRCk4VuByna6V1gc8QR3AxH7g3eoOxd
RrIRTYYg+GOaoLCc7PCDhmt/FROzJczbbe0nNOFBOQz3XOpeO3qGrFPfLrceB6UU
xh5pzQutzVTzLE1eitDGjcyEF+QHJ7pMly8hbHUr7O/BaeLudj4PNy8AxiwQXrDW
sHX17Jo5kmzmi20hhvqWMPPyAaK6WgiifO0HBEYSyRtFZ7YrHFtf5Krc0j5UnDTX
87nWiaEfV5fh3ZF/rZojoBOnDt0PD36DimffZvPy256092/XmlzBCtsDvWl9Prpx
/aBn6aaGdaT+CPGOeXQPoKUa2v4FdvnfGciSOFoxPFmhlATUl6PvRE4Z4l8lXVxK
1Ftha6agDAiQytxiKX+K5MWR24db2zGDHsy3hj6/ty68y+WxUYp4pWq497pPSZ3q
Py8f685OgQrBNxo6q0aQ4Txgl4d4PH3fttEzxhXLTASREHrVvV1IdkqrIqKTjO48
gxISGrf3M5MVhtwdXlWMq9YeqmKRIX33r0gtwJt7lT1XmIZ8o57NDCg/FY9Kwru4
15eiVxX9ykO/oUipP0Mu5SqoB4M5RAgpxw1Sbzfm4fUTsnVPG5f6shL7qAoWxpTd
H5EtYF71zmMxsTsn9wFY48022EIOJj8HyezNal8c1xQz4FlspNcBL3j+hz7bSRa4
zAhLY8mJNCSoN6MEeRbc0gfqjc8D9KcFPaL+zTrM97hFZCEVEO3OAKFIVkGq9Njf
u3UZgOEAAbvp3LAhaQgynzWkcILsDU/hh3lo5zgI6c8yLN8i1rlNvmNiMorpDoYw
gpnRLlhw2Qqmh99BoHK1mR3T6lKBwCkHk/kzEb3koCaUj/Q6sSl3uaNYfunkGjMb
aSPSjlVoZ1k1bIj7vdqQ+mwt9+Q7osrGIlWXEWR2TH1j/rdOrGFmHsf3xlH7vja9
VZMIYNZHbH++KiVRRqRii2iBb5g2Jgx7MFymXnjjnKnHCdHItDumioQjm2HvFS6C
FHL0CQwdRqodN7Yc379dzrqr1ju+kKKnbaO+pJ3T6C4ICvonaidXrqXy6Pm30yoe
`pragma protect end_protected
