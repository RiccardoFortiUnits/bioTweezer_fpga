`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iCci19fdxl/rP4Y2llC3o9X2uaucRIyDyHYH+BJLKysqsuas9xiqs7mX/ahapbR+
6MLZloi0qD7ak7beEehLHMvI4DBLE3AI5L8jIcex1CvZTCrZzkolF7uJ9j85dPmU
WHkbZIoBsqgPrtjEFAZgYdoB2unGwZeySWzRDIOrEH8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22080)
OeDOIRsWwBmtbgmruTxKbQbJ0lPxvrkf0mqAhblkXCFHwsC+kphZz9XRN5Bu7/Zi
YjDLm3pTQJkXCoK/Jmd9hnjsWG9oK4CvcP31fS/WljYNS63RrM0s82Xeoc2n8Y7k
4hTpizHfe7CLWuv4L1X7rSWTQU5IAYgpSdryJ5wqOKQnmsnY91ex3GEle9ksL/Cp
Ffz4fMNLmrfDx3ZsubkEPKshfeG6n+FAIrQlohGEXGushjav8AcTsgSPt+0vUAB9
BFyMQTijGwHA+niv3+oFeyXSNMUPPLD9w6T+FeCpxY/cyBX7O6YuD04+WDkstuIY
RT4J+iIIodraq0y2pTykXKbp84z+BeYBhENEXN5YUsEGOqPMlW6hIClYwwbLckYD
bqU4JBf8bsmYCtmY4i1qZ7ezIkuTO53VhZhoZzqnrL2l8D90xMYkf6A635PsNMOe
WvQcnGk0Zkn/Sf9UDJjPIdVrsxopr5azvXaXoJqdHQJ34JsHceYvRUjZiqBkrRry
7Ip9qmQrMRF9vSso/DQM3fhv+KAqzZe3fY3JmphOaBwfe6xN8rIIMzRxjKeC4dOK
wPzlV/b1z7i/6v0YE05AwWfPQSa3crJZ+Ax2id98qI3GCVhCInLueewC2WXCKHD1
WSQKbVo2hovhgKxoXbvnBPo62jiuniEcjFEfZuMOljsKu5ZRh4i7Qe7lMcZ5dh6+
6PeFNm694LfHKcehcHqf3dSLzfvUe/7/SAV0xvR7S4+dUGOc2QYzKj5D76t1H/yN
jvlTJzvyKLtLRAAdCeHspnG5zmkxjOMyzRrFG/QxgF8RoeSdmWUTOl6ZogVi7AEw
RoEntU4OElhJNyHdqm96OqIAO717SYY6xTeIpSnJazSLa5ONLCah9ejabzjRaYzF
UUK1/h84gfkD04cWURqrJ8tb2fhBP/Hwe5wXpRmuJHhQteCIU8/8P78Bwx7mNSGb
Rj0dw05JtR2zyL4wzEFuhx2MkZCi5JAGvneOGq0gIvkcoWXbVy61ygsG/xvIveG+
eBpO16ecKSJcf/Lx+WyYplQGONgrsdya9rXoplK16Bh+zY1O3YV9U2ENXh0u/Vi0
U2FyTcZXq1EaoKOQ07A94QPjpukl6BgJAG56VC6prUnCw/tyYyzJEvK6gpi1s0W7
eyx+Q71ViPWv5SJWaI+qlqGhcqIK4hyc2cMgKmZaudLXU6jOBBcFu5uXAdLSom9k
H6RWfFsUJbu/geknr4A/d1CEv2ohda62axREoDv6pCcugl6Jqfx5uBD5mS0z9Q5P
srTrlwpPKYTD2cDGH/1us7uo9VHg93o/1Ies5LRRZXtk3nwIyWu2NiHQPA25O/Jw
TSYxTLnLS8T/rUFAzK97KOir5PuRVyGUrcdrhFG11LOEpF2V2Ab/SOydd68gq+7F
lfiRY4PERkb+ZYdKsg3K//CujdxFBeaaCB6Ja9gFvjj/wij953UwBaU8dBtvTkhF
Z71jvPvnBf4R9qw+2iyNBWefuyozl3lQLSJetTLvdUp+9bmpyHmL3jyDbB+ba3XB
qb4ouvBUbO6UWc4XRd+2yaGdF7zlTvGn6YAbKHd9Mnu5mz2mdIuMQk/PdWh8LnW5
cNR/KPq8a5pogGsA8kcvtK838e71tH6gtfqdc/0C8UYZfSt73wprUM1xRnPiyBYV
bCIMyczi3f/Qijdl0xHY6GU9Vdttmz6ugJCMYkMJmwUFUfxMill2SwUMoBx7UIZ2
i0Qh9a415ft7OTHxDze/jziHSuDckwBOJzdRb3+U6JJuZ5ALDre+s+3waDR+mmwd
MPFaoTSSXcJKXJQcuB7y3hz0NVLeYKK09OSXvr7h8cdSvDDXReLjpOeivNcCptWP
DciSVAd37vxmfU9AfTzRMrI2tHk85nOiAJMFNmHuGTeH8vZQL7nBZVgOoV0tVvNB
ghTBxchTo3V6tV+nWi6N8wsfAchZIcqdm2aPKjSzIsSnCrQeQAAEZHkd3Kn7teB7
qh1Ru0NO+pdEaDAe/JXDhjWchpa1Pc62ZwUm0hKVn/yPqqgHo3zj55g3IdlPHK2l
sqAwMaNv/UTe4yqzUFCVFN2BZcLslSWhlasEBM6Xp5q28CeuehswRGHbqSj2UKbM
HQFw+vxDi5somRkSulcZgjC+VKtEjW43MtiYhMjsgjYeozFTRMr2M6fXUV6bwDp9
mZHb3bcK7u0MzUMUgxwH7v05cJr7kxhgZ3dd/ka0v9X775s82ksT4VenYaTwrDul
PR5RiaAOcrbwNRKJgaiZjsBDqnlBGuHRZV2YVpsIB5HvBNWWdYx7J0iJ3rJVr/aR
Al06IAxOf9eQlCY/ZU/MiZ2NqLnR3e0FH13LBKTxx2NlDsn6FhGLFShrpSnEFzDm
v0QpqCQVFSgfIk0kaVqBtoo6GDicHrCjppv1CUvlH/YImkjjztJH4d4p1rfeQCbw
AFRHNNNHgpcE0QC/exXQ16BC/2hy/eEwnhvBOYtArrTvgBsh48Y9iyolhqhBUyIW
Q6+ahnIWYClgjRP0Wv+Kjb8PTBOCgMYiYYw6KdT5G3RLuOaTs5c8R0jB5we+MqkW
IRO0UkgFGN4rWCJ8jxIriG6gxHyXOSdh/G2a6RU8NE+KYs/mKDM5yC/O7aX5TeMN
qi4/N7efe5JdIR8vxyj6huhCQd5fMAqsmMUD0m0YCYybscLecwM5i0/rUBt1I5x0
9ptxFh/4c2weveAFI9Cr4OPknWNwB87Mq/6kqYsi9NghA5rKAgYHFvR7B/r6xcoN
AI3zWI+RvuO789jH7J19iJCQNGQPNljAb1RcuhgxjIgpd/9jM9QyXPnUB/4j+88Z
Xs+QBbGLnNK4hcFisBkvVsNcaYz4VL3nB7MJEft41iIRHGkfHhdH1w/WX6sbaCVN
kvCXALgzIWPHrPTS24QNE/V2Zl3Q/3FzCbDddGxz5zh3b/rrTg3S6TyCFbzrstQk
ku5DIf4eewjfklMr1XZiCmNa0vKHRfS/tglLrLO8aPLDZCukXZQTr5JtIq+XSbYu
kWwnFtX1yG5GydoMXWJQ97T2Yir8kzq8MK2Zn5SBwYccrQZsmNA/98O6WxZaIgFz
7KxNx1dngQBYEsWWcPpmIjwUtY+OWDta5bDtHm9d8x4y1Z7ntXgyiYza9U+pB9+u
fY5955fBgSuHJWHf4PNNBGSH/sfCA1P3H3rIVtJvYg2y/Nl7QNdLL1/RMfuJhq92
l9jMUPUHAVUtK5NdMY11YnuM3I9bXrDAqJud2wX9jxP3NshgOnbHKy+xtnu/+k+Y
wM2pSliqbRvWJi99xHYp3lzix38tKq1oDJmEWPOm38sNK4dhmztFuKkr3I4heljf
m5buIgSjVSZ+hteU+EHZ9TuB/jNvV3N2RhuNziRKhLIaRT+8NBJsQ/9tFxqn2L9n
3JlK0YMqGHQul2GI61LtdbCXpYgt6UKeHCfe75/EhsVMhRNh+qciQqoj/IBlAXv7
qaxBZsX3jamVLn1JD8bkfPM1xt2JWSIJ4b1qJjbyWU+j96TfJyNM4HrnRTLzfuFX
92Zdez1M7UR3Ux6aIaDADqtr7Xzrk87U0S5+ZdT6E5BZRIdMHPi0tgtjhNwWjV/7
UUgZWCsC/11paKUHpvNxyo8t7imm0PihorhASWgqVlm/nkBZC6lAxA1oc7DqNlOs
Ibbobif3p8qFgaiOjdy3l/UcxecX+DcanNpHkQst43guvyHhnbWr5IlZt810ch1v
apl3NYWrC0oN0+3ygyeIlQlqm8S2hRjGUND6MbaxlBgf/PXkMKET/655v1561ey/
ybITGzCAuzau+gnWa89bAcHAwtM1oKSGld+s7bR/O8RTb8OwCTEUkqUWjujUvrY8
tgdEe/HogJsD1xMYk6AcDrRgPNzmYCfKgTKZWYiiONoTUcAVFYTGrgr1I2xe6QRh
n5l0WANaSe28eFQm6U+y6eI2afa9PMCIhaQ0G0JCar+DK1yNXig1GDEv+kZ5RZKm
UH2yCxt+vJ5IOiArpP8DznbfWTa2iyjh72sgAfw2wzrFgrHEEn6WpNUpOqUrA123
qcqIlpJXGHLiY+llU2FbT+6JEFpp7gW+zZK7p6hHRP5k9pIqrzRSHfLOZw4M1szO
565GmW2fGfZst2V2HKcNeShVCCTSOkMBA2grmCXKfY5EPPfnRglHYLQTvQcvc9Cl
ssqbSb5x0cLb0uM1KQtnSG+0FY8elGotTWOPjtKAZj7rYvrJJ1BfLM8DekXVKeNs
woIOSHAkCh9Gk/VXZmS2PQljWqyZGFyNKnOHTtx+IwW8jV2DgYvmeqEYDtMaRGqF
F1XwYimnU2HAkhp+ZB2W8EHMLpbLnh4W2Bo+9+bc6AGPSuWfoWTTEUkVp1FWw5MB
T/fkE8zSHG6Wc1MaUQmAM7YQWZei//Cq+dj4balyKqT/dIuEoX/9kU+smrp4+On3
UUNJlOlx8/m6rxrddu27Dj6sMsTp39je3SQOyTn00Y5WDe7O0S8Of94OHZQ0ei9l
w0puJnZOc1mdjNmmyP3r5SmBLZIX9NsGo4glESDpgDCcXsaUKVqb7Yd9lWijJ0Or
JxEm/YcptHSozRYXvbK9v01OpG1VPcsgeJ1lwNEQ2HcJ0/8IacdHAe7+nQ1sta3T
sObBNDBHfKUXcsMHJstbJJrQqmh9lTv/t59dLETNbK1bkqWjopnaTxEEzAQE9dxw
Dq/OKImAjOVG86KQkl2iqUa86Rt815L8tH4I/EtzwKH4PpREpSj2PYxBZ/4CthUw
0v36TzXO3+0oh2eJ//eO31B+3ZvULy5njCCtJ2UNKpcyrcWRrIG59125LT5WEMsi
i0ItAe03LJwr8z28t6Ppnch3p7NKJ5b5A6wXSbpV92FDNJZB5jO/u8k3p4FUP1u4
s02La+F5D5AomNlep2cNZzi3u5U4EclZ5OfUiz/JPinIVzXvUqz3v747pUe/X+is
zK0IahAPykQaNdjb9/jqrVKvrkl7p211YkN5vyVdcZCfVzwyGQMxGYSFHNzFsG/C
co56BFdJTBNDt5AZaJPRBl+SgdDYLKmEcrqU2jtNr05lgVxO0Ehc/CN349BY/evH
8gYa5+7/OOapvxG4riKSJnO3zDvb4iXrLDU5Gr7m+FgIK6LyNd6HROAroXa1aMDg
qHCRLe93MwZW4nIE2HK2Cic9RiOGNNP0GEFdhK13FdLxDTkkyFxUYVphjkhqg/js
tGac4Eu/9mqcEBrDBF0y8XS0Crn3LjXJWTWAj7hD/h7l0boCKO0kWxX9Llux89yu
nebi4znJ8mZHYzHlt9g+n0eTiDml4X9Tzu4K87pVgXs9SwMwGnhgFYQXeat5vIWy
g1Ogyh9O9Umlo8cp2VX6Nuw01vaHrB8x5Boy+YArGyqOwfvgte5Idpmcr0HJIbMB
ZApmLZHt2w4sVvsLbn6NEG8cjU9UAYN2O8Kuuim0nqEN4NGQCyDdQ2Mj2lBysFYj
/Z7tH7BZ3XtKK2LyPiZvjk1nmVWNp3wvVbcN1faflSsyS4Wl+qEvUx1kGZG/Xypq
z/v/r2ekVC+gM9j1V/sfpG+MhQ0zjlzPlSgIXFr/FQfKVaY0YJYAjcEN1cSjsRFN
ufAoeKAkBgHmkrC08WmnzvsoOIyybJE2w80JMiVdFvIroeFzMpTXQX3lyc5crvPo
qkmsiWop291Uadm11Wm9XBZqlfgj10cwl0XKaAJfK6ZPvQxhpOH32yAoJ1/Lr2Ue
v5UMIToNnVVVpUAeMNbEruFDnAmA6quQKN9/9sjABlzSqgxJnDy8p210SvX0FSZZ
JD+O5PffMP5z4JoXO8W+5cbPePXZrotXkdRuMsoFoxJCPG68HKMQ8lBqvsAv/S4d
Wr46n1u29OF/h99k1xqpDDCgmkln6HB9QbxKtCnHJkfNvdPi2k2MrYoNHkv89Epe
8NwEcL4/AKqMyxGrYbgLaE1XnaOpLTvpBwQwjoSJizrnwMAwlpXaFNMpEijHJG8v
yx6IYXp9sJVcsFuB+6QnK3oM9g+gS/Z3KrWOyFxd4687nXCMNGScF15vK3HcpLJF
fHm9Ta2cLhFvETq8iU0DAro9Z5Gt3SM52zTSosN2Ex5UwRdkfYY2TxOiK46XqJ2a
7QRBzzT1TxrmZIYrDnsjZ+yAqlaU6qG+MxXVu2t8R7ahwFXC9jE++Z0A7GcyjXXs
u9hO274D/f46jjslC96CnBdgJv28javhbBKI6ywTVnMXr4vcVxcPiZwLIpbWOxgh
PZAWF0VpNyQGGRLl6ixIxlrh6NOEg8+NEb8//kxO38J2l6m44D+23LZQkD/Sg7xP
G7HEvwDD4UrILADds5Ej7OV6tPGb60duSp6p62hiEkdaVomhgKuROViwDtfrNkOJ
WuUrD0jb4RIuWuZxkzk8EpMmn4iIdQ+cyFABioDARtto1Rzqe3ftBk9NZERJbGBJ
tSdkx+fHQBjrThcSrt8cjLEeGFYnEoOulxxY5syn0PAL0D9yFrKW/GouZsalORjQ
3UR4fYNTi89G3djPTPCCD8hHpbOESoSBhxNew9wucaYQc4og50zdjyQLtycq+Oic
1qSsV5l/eZ1L3lcF9V2CNmEjGNqnquqcREDt0ocz41vYfvHTycnYPfTv7iwmESYO
dwCmDtB9WDnTYLuB9KwFHxpgTyF2lDQWhAbfPVlewpScEg3SK0sc75VbrL0jovYi
VEoG3faQSzsegvnBVUFhmuboeyb6iRoF81aY1vt6y6MvASnzYjfTgEEwH40Fp+6c
xG1ELFI9Nxi+q3ZQloDuSCKIuPPhKbSmxxH05E648Lvuct+QB/5K30bITnMTMgv8
mwbv3HESA4WaPtejtr0T2cZs4hA5cek8CaoATSWhzQdALreI0Z0Ik84d7pMcMerD
+GS6wn9ZAaal8EPP5Pxtx/JR0E8/xtuHo2Bdq4i4tSJ1RSGZV5H1b7red4PXT5pz
qy8GcaTMLmI6lgyeAc7UbpeohSXjhkEjHkAlykOpCZdxnIZzr6oaNYusiQpBDcWn
CqU0T9hQuKWkNWR8iq+JKHl8uxwa/w0dFfib8UEyjRt3+wksg5Uh5BPNKwYQjbAy
yzqfWEz5R9hx+1bn7zTz+3eBOj48xOz5ILSGr9CUYK1a49OD0GLCHTGBpTNyRdTW
GT6qveal7+ruQsHwglir/zrVfjeyd+g1gY0bm9JRZxDuQ2zUngjxz5nC1hor3TIU
pDIQcEBn4w0wQ+W7y6XKJ5BsRc0DsEjOZHZe59BjKApk34vKxEYeXzdYJmXcnxPo
bY1ePtNXphGyhX44aLtHJzrcRZN+OKTKN3NV6aC2RURUie2ZIhzYP89POkHtzPz8
8aFwo90Jdd1WC4IldUJqBssqq8e3DVoopn40JUL3Akn/wPDOWAIs+iXzIuCqlT+k
XrkXIykQdkdCQRJI9JzCC2DQOiFhDG4YrZf5ljEE/dKtB7dhMYXkuowIMiXoBsrO
eawU21yLDd6jx9WItekEniDnOCsO3lcUq4BMMlh0TXOhd19mH5+xaW+ITtO6efcz
aT1ZrqB0v3pBM+ATG3LjeyFt9I52t9KiPHnBIbqZwVf0GY/NYxOZ+J2b7edyP4Wj
IK8XnIuFnNaIkoPtm4oFcusx1UbjCd2TF444U4da+GG8Ci1LpUFrFx0KlnLvhBLo
GjI6ON4dpZFozlSrvJNshCe62LiGqMTEdKXwUq+/F4/dCJckPUTVVjNx3mart1Z9
danlVSyT03nUtReMyAOUT/GurRkaK9APRQRpx2g/RqNtGUsMBpEH8A9a/HnSuZvc
WcMBTVYqVBKqoiaSkZvlD6iggSFU4a1zeGZNRkNGsye9mxujk2BrnQYZXHnVAGsm
uAQgL0WvBGevP8tmwIdLYMkvxuNqHc+oHGjXNJDol6lzY+i+T6aIOxwN3wn7R+tE
T7/4daf/9i1Vj0waoCLXYDAORPDFhPbuM335kb75l9o2nD5IVUl9Bd28IUzx+E3k
H2NfKQfdxL7UFFyUG8gTzGXmP/nyjlmBT4j9uKHjKEcMZLxpV8oxC/v///kWY2JJ
rh4E66w35/Sy7pzmS8ndXsxEfLqL6beUXCZ9EaGvDMd4zBfy/8IRJP8gj9yw2Fz8
F1ZnKvTDm8VvOq5F+XZSQF2Q7X8oQ3GP7HMbSrZKnCMWbzeXNTv58AD+h6VDJ5ZO
Yq6qO5NvgiVSISC5Efhwu52WSZYsdaJWvcxsqyI15QrB5DeWdhqkxZVxCYp93fRY
rJOkKdbzj4B/FPDGBl+S5Ib944vx9ESDRF2M9vPd3tfyup68fcBgQ3KbKQFsdmLV
FJKfZ6c8q83+ICfy5PTyDW4Gjji7TWfF5RwVZv/nButEOOrHueWmpwYwwRPkY90S
ZFaV0EaQJK+uPH5G+sJ4KWhKiAhhSSZskUjES9j/Cnv9r/BiQrejYB7aJ+3zPrb4
eN71CiU8DvwS5ZroFTML8QW+BpTPCxD3a9KejsTVEV+y0skMnhB1JRWNz1zcHGmP
Km73VP4jhkPuy6W4nX0qUWFKYaeumcSoOcaR+UbX8FbaN1wOMSXJcka/IDsa1iba
8BvTrXccKuAjjhaovDVZ6Y7+vtM2sT6ftwVdo1s9jRanKAjZLjFYOypjNip4m7gU
BVQLCganeSZ/bsb50j4zxnDy2PoK2sTKMWhEJGwJImSEQ00i7E/SNFejZquzgfO1
XRGlj6sSLOplEEMvDWjuqfuEAe5/432ulA7LflpXTwReL/K97fdJyrYv6wLvpAWP
+pALz53nwbsmobjPlokAU8eGDIiBs/O28SoI72/R/7BhORYIQOdanNtsMdk1xup6
R2ff0Kr2DNF5GZMlif2qJ0dh8/KE7ZFG/r/OaLuyIJXC95TuN5xRrE4Q8TzuSfSh
Hyd43pJTvrtj8V0ZwbvQc9vTPrY/sKtdsPxW89av+gAq0pQAWV/7gN4VJXynZ9Qa
cMw2v5rQivQmx73OIQtHppUBIQDmooW/7BVKRgWgkWvlxyyRqOOZ87x9cUT0v9p2
yVtaZMUbL26unwRAFvUfWyWl3M1PgMbtDs1XZfFPnhYWCzojpwLqcSezsLcRfLAH
Qc8LWlowwSmSWdidQttGGA5yx5G4Dbe5EOq/Q+Nv6PNyH3JTr2NsAymjk5huHDNl
NJXG5teNM7Xp+n8pC6vFIfjJ8GPRFV04JdjJyWg7U7KmnqNr5qxATAUDonPCcIPq
4X97i8vZXM9dfxao88fMXyDrdcSCaSxeIgt0kQdKgwUhiasHjfZKlCNw/lJ6NOSs
V4KFMtBKshPTIjSyeC+jxPkE8r0GmmdKlKGnL/GUdLzimnNNv4/nNVcbMCPvt+4R
hxiwrdQlX439ebqO8Nf2CD7/70IlcN1h7oG1PsVNa8WisomtqZWPa/dkua0ZJteX
nvoirEBxfHvqv5/BxCaHUUrdk77SLPCAG6RodzjfAkFnygku5UazS8+ymHHhjwg/
J/kNsN2vQ5pO18DNr3/nKXSUOwy0oSrEhVd/6zxPpZuW+Tum9dKDlGY9q/ufz+Tx
yF56EiCCBmESRxmw0tpguG6o199xiJLNWn1jFyHhxHdmB7vvqVo/S+uDEZ8vUJCT
c7fBAaxqumK4H2PUXxHFae9XvZhDzV1Au6mAi8GdeQ6/5r1/QV85cx4lnWG3Dl6+
sN0uyfTbh2/BoLqJvtcFDuAwf+SBIV9fdH4QIuEvWrKrDcvjFvkZimeBWgocBjZz
4P/tvsHYOjwdbelMYYFNTKtoR4/maFSfZV1x5RdHRoRZmsD1E+GX97ycnLoFrVgG
lSpGORawn4QUKvQDzW+IOX/X51J8jrvWz9V5Cg82Qkt1oDADkpSldc8HoZtF/c38
wEEY6ziFVpt8/3fkVB2RdyNK/yVy0L6UGa1dWTiydc9JuGND6IR6dja9asAc5480
z0kCtUTX2357+he+8mFYA2tdVT3UhY/eYvxmBrAZowoUPbjRZhAmL3rrkWmZsaL5
HoQt4EfuBbdMP5mquAmP3ZPUWa7mcx5p8IiyFqCfaUy0P5+m7bALEiqMnT3uIa7V
C4bERbG7Y5A/hZp7+qrrmvzM9M56vLAKgRFDZHxaSlZkJGwWUxMLVnUR6Sautn3/
MEAztDGW1A5i6QPVgFWXhDbW+4ZYxFACZ4Tve2GLHt+TVmyL7pH5GAYJvi0C6eLy
KFXS7aag1vik75VRHEoZj0jKwnAag1xIBpsX/7foHx+UVJmkUhiys5BcAAnowS7n
ICi6yUJshs5IKHtipzfB+qkwMYwIXGpDwWHOSyY+yNtfbPwUIs5suJGUBs9a9qe7
T6umNPayKbLsaDJvQRvNT1OLgAZB9utasjLWM3PK87MFH2j5WK7aLP8l3rNTYuWY
242QQYOLIyyef0Ow6qOWkP42N3V2y2A/ja75XxpPwTAekdO54Vxqu6a8gfULObXT
ygo61Iw1iDzF5A8rvrXZ3oZv5ZZmlLE3ls3XXSAxHvXVCI3xsSS0EDVC/sjuvKT+
kO9ocButr5BjSxUs/EjDdnG0UE5tJgaWZ1/9ReIeX3JGgrTC7HRK+ghutJvqHUJ1
k78VUGVw096L2nrlc+BKVJAVEvDJI84f0qv1Ief/ZKtaxxT5MOTspJ958PvGskHe
i8/W5i7X1tbvHCyfeGvmtMjPMkGtD5pI4Jp3fRMTEl46tYUdRs5yRFUDMkmVYBTr
hXwu6f3bwRBRvcXEfhYZ6FCJHOxF+gCPBnJmmXfqJPtcX7OjbA8r9V1JBVocDVFQ
9p11Q17mz2YCG9CAurOySf/XcCtAByyP7JojxnOqTCuKO80O7hh1uuLhgmyxaOUk
soP4DtBVzCsfNW77WC7NtgA+7HnY4HanHlZnZVQ3HztQumUlCAs6ZkAA+kOgSQKm
W2aTe0HoZAGAsbBn0abLAI9oxqPR5EQC6ViUUoWtgDdCU6tWahhQxaw6jDSlcs/1
kIwO+yYabrIpNW75IqzIDZKsjunCHolF5BFGtlXopeLr+aE3+Go0JNx3y5VVRkya
lXeURf7DrKudTGR8OK2K/dCW9vusdE9If3EOjKL0hMeSNbEiJXFSYtM090dmrI9/
pLBD+AKkU8TrqNxc36KlDyw7xQq7YJDqYK/RsbjLSt+E8449Ce86PKBBPDCV6bE8
0sTVlqu++B1fM70f71WTJl+MoAHvmOeM4e0gAkxI8FSC2fTdloPtzwRK/5y/+efz
hbM/tpsXk9TuO7KAcfKQgcFdKf6R/naGDSQPU0ns6rBPpEJRd5ojhWMNhgznVMk+
epylx+YqMQCGtgnAfg0a6m0OQCKYuYp1UL5wowNTP2BORMaIPamsdB9o93gV/EdD
/RnrUdQZrUaipUxE2BN9+6Vyapd6gdE/JZWBmEVnQsYvvFzHkCEP/EkxWL2r4qOx
J5kKjUTYd4BLVn4lAqYUbAOII54zZ1/kHEWV8ai0WEq48rY5fhh/GdsQ2qT0EL48
jFWzSlzDrr7VzhvLY4AstrWsYaLN4fd0Sh8e5eoFQj73PzWAprwrOlp7WUtmH6r9
LDz9TZnfhbfFcszCADRe+JEXUng24lqxJ4BX4ZveCiRJCnVdc0rRk6RalSagqnDt
/WPRuoPMMs3Us+Qs14Gr77uYSWqlJNOsRGywPHJVF69Wgb2Grv3a4Rv430C3D+a+
0dMOJXmE2k28iz64dfW/2AwHkF4A2sK2euvpLbY8JQW8kdBMcgGJJJWAh8rgWtOR
e3LazFgvxkhnL8winvbgKsqIyvqqSmLYAePPfV9YYTw8kNKwz8QYENh8kvDpb1vm
J/UJuhMXGmhWBTBFUhBIaM4M3zzsNgmzjpKWo+eCC5kF6c/jLMkczcInV0iPdO0Z
kpEIqm6lGFbuYEjOzwdU9RyeRxOTXMPHEgHfkUq4XfCjYEpyTItI3WiaBtejaEMX
JMAHY/9k0zVoO7VTEqLfdZhv905qFg5ZTKcAIs89e6WTApvB4FDar8BSm418eaAR
f0R9oH0JwXv0FaqNLHMuE4dJoMHHJt8V/cZWR7b8XKtQZ1zCrUWtmzNioSb1z3x+
0pJ3KzaEhqRZ8qZhIiPznrCS+JSFL5GAftjCzBkzxi/7GLAE5lkTSr3tA0uVz2Uv
ShpTQEDFfuu7VR7d7X5NFM8pvw6AUD72MAGB7umYrH5BqsEUIFip8ZeVF+5DKQcw
AnGRDfwTAh6Z+SQ+UUNMkbvV1TRy+c6mifmpfL6ppT8E6P5uEWoTPpxdXPO1tudO
mH3N/fDOfIhdRYaAyCIwcfOcuxsVa5ZoFUBJOST+toinkYe0eepsJMq7GuYPVT85
GATRw/s7WUVgy9ThqnJa+1Puu09QL6KbTJzCFRhlSoqX/DgI1CNaR3gSFZbabKbg
feSb0WTXlg6vzjosbTHFBAt0vfIrSU7HEdQs1B//0aKEuciOAbKZKR4hXBQWvJgB
tsaazVY9zKTNBvm/yTmTBoMOOcGP3ewwVgV0csPWSpPBNmnGoZLerjjDm1FzG9uy
kG0tp7EFh9qCqMGn0WkOyZQt34qvT4gceG91hQ/pqu67KGX5kHUzxQgCK4/uThsg
ACDG0qUQb0Bxnau2Lsus5s87CKhKN31ElWmy2dmdl8dYGZ/SZ7Gmuv7oCNW2By+m
NMgML+yWe6FF7ENpYYRpmNtCznsYDreSCQz14L3psHYQJt+k5e93ltbJTVvWp78g
eBwGjt59hSZ/SOF4nIBGdbghIfVAFKDfxQ8YS4a+Lnv86oi0c93qjFxozqF7YlFS
q24+UoJRAa6YAKTmoa4Y+eGau9JvxCMb9n5u6NIWphkjCz3okP7fr+wZxsfl7EBY
EM9ZDYQ4N5hh3GU2WdZvZ5uhBepcK4kRy44ntlfUw7WfdjCrCmc2L8uXuw5rXFSj
H3wtACnUSM15wt0VBQt0KALOg8aV6c+6Ar2C/BjeomZwXLbG98n6w8lm0UwV+R6e
QdAOmzdMxy3J5WPgzQCmD1UmcSSf97eueig8cWBjCx/fmOWf8t9SeeibYYtyTD77
T2gUWDXGHmvodwnzP2m607C0+7rd20VS5+vchlteD7CkjZV32iux6Zqy7IpjnlHx
aSrBU7AThNGuRBzv2dwa0TZox6oHjGQwzo1Q0TPo5oj+D5o3T2yWM9wJQf8MP3cE
4usGgRo1YgOndPnFtghFXrNHzbJU0H8UBXn4zBE9cRm4qGct2n8JFiNqeojqk0ww
nmVW2X3vks4tekTKidycbZSi5UGcgy0h28fc1J2lHtV4CIeCyM9lfKl1eMUR3myl
NY2n1PJKTFgjDzg8bZssQXt0Y4cB9Bk5dzKQxIZzAj4ZlzQWambgGJjMy7NCtg/B
Tv2Idh7LhQchWCXG9ZwtbeHtC5O52BYGDCT/dxW1Uk41UHWPPWrSVw4krgtoTHdX
PH7CHcQPSePP/L3UixMaKoUlKg6Ee8dWyHabeeEjphWQIiO30W+ALkDRYZ4nVYNV
l0MZchB+zUM8DOoB478s/7aJySbBtc3rFiYclAS0Jk+Qe0ZmIl7cTWmmZrsFRSW0
CAQx7KN2mqraubha5MAl5a/z3p3rIpl7ww30NjmSfb7vSJ4d5ov+8hqxJOM6IFLy
FvAt4XM4MsHBAl6r7SJWiDK8iJYF39NH/HotxNGWjbg/kBiky3Zt5fcBzlQpmx2J
JjrMaXItO/aA2ftaToDA+TqZR5eqBQx8SZAgfNnN7knl+kcZbzx4dfGVB3BET6ZC
ljksgwZBKC2ClH7/+AdkjEx3cfbvGQew7GRLbSA/pYwfQMfk8ZQqB7A/ko2e2bCx
/ROiTm7zYbuTQZ1OpWpQLswI1gfvHyVjbk0gl3VOkdiGcohDGk8qNAZRaxz7Tuxe
O2PAm2WXT/wcvXL3CZLAcmcEd7R1gh0MBpueFWJakZ4RZNuzzfafhc1EPxXWcEFY
OYJ0cC84wJ08rYaquDDCfyIhU8Aevd6+s6woMpC3Z7nPKEgCk2dQXelph07+MhkP
b/jGwC7j/mkCCAOweWK4p8k3zB3zsuEhKPuLlUTQDOGCca7oR8CnoIFSGtTUQM/V
7ZYnsW7PrLw5htGV0I4m0jqIERAz93FjBHXUV2Fp2e74Ju96DNVg2C36Vt7edUC5
kDwftbHs3vuMNOHBXYQa+hrTlgg2OyGpnMzeqkxSjjPCzqtnG9MtC+ESWnJZglpO
45HOLWHSnVZUIQ0tzFnu25I6MaHsuTIq2NwDaTuvaqbfuobyA1rsU6H1xUzavYnW
Dl4SsXbmb42/ZBGeYAg3Ui8EGylAlnnijsQAmEWuMuM+OKvfKlghNToVyMGq4P3B
EOcoLRRB+C+5G+m3RlvD5FEXkGgl9ZBIrAS0bBBk1S2OZTpX1TDFPQFXSUijbd/d
mWVFwz0NEwluUguU5ECuy4i4DLhPYt1EHJHWYYXLTIqpJmmKDpAecK+3JVUDEbt9
RAsemU5eG73xOJAfdZMg+YIIKo18C63VTjqHfm6mA8e00VJYrzW6x0o2WOLRX9qf
HlOIT707Y5YCKioUcUPcyMUbTGMYOnlZvQObqFPKw+nFzXhC/vWcXJ7iPTRfLNvs
FJLUNo8Q2eJTo2Z4II7cRx3GbPIEIQ5FV2TkY7pgOnSTjYVxG1hPBmKq+7rFWPzr
2M2Fymz2dJl/tXOQ4LOBjFuBqhyjnkwitIs8uJ7OEdYhg+GXq5ou2pzHtI6C/qLE
D5L27TGTPr0FvGlT7eddaFsBMxMr/9tmRDSs5vnUnzNRy1+0QjGgWi4lWQI5gU4Y
FZUncK3pECVGBHDA5VViQ6tM5hjqy1b0yMMlXDCkGWEgPHVzdEl+m2+E9xRw+HnT
inK9BoGuAwqmwzGE/2G/fOeVwvIvty7F9Vi04A/1HDSZKKlRgqMiqGBxRhOFcxSe
sy8S4mRWkzIh6pyij7gtAVnhWKPglJ8UU+sz5xWFKnc7fNh/yJH1CxbPQ1zMMVrq
aQBrUx9Q8mAW56ghBQVH3n1uS9flz+qmbDU/pTWfFRlfVXqTKGOBmcS0NVF+BPCo
QM6m4nW2tJEy9sYhBL4k8QBZVYjs/DTxlGRCgbVg7uqTSYzrfnGC+w/urqIfi/kI
WfogYkXPnIt83LN0Y7Q56omNAyRGaNdMbNau5weEm6zF8DfU+lK+f1TKIKhzoI3z
4NTaOlVdUe7LrWy1muuBaY9QieygQrSNLptEngrIeA0KR0kI30PdBwlNyOsypLG7
pRiDQAgMUDQBXtawvTOuern+5psyrrS6ARsTxn/Xg0TYPl9L3wcFJ9J6g5QkstWc
VGUjfWsRxu/SB2GV9fJZcRySP13WlOEu47XdE08wHolT4/S2zuG+oU1JMs+YYUhM
Ry094+oHqxE4W6mUVTzd8v4W39hXEpnx5bSxJnaOWsQi2+J5vRF9J8UNFAEe2ZBx
lgpxbzylNLhiUULrMovxSweWbewib1CB3DTn8lBq5TrCHDbTEiwmA/zyGlr8koaw
Y8S4T3lXgUCPPSSLy+ktRiT1eI8ITV1A7TN7L2l1vqNoI/UPhUJb+mbpbTI8jvDW
XuYNFxN9V0vO4XbNyOuDYqn54fKxXAr0w0wiAmMbYuvYXOoceqBg7VCwizcny+pq
oEQ0zKX117K3qjTw0pJKgeiOHu7dgBeF/w3+vIn+sfwru4PC1yE9R7wZPR7itmrX
hp6ke4caxY7A05NfF/TjIErlvHLhq0msOjzHQzH/rhsPki5e/3Sa6IlJaa71B9l/
CrqaWE7FJwRm1Ngbzz0+9NSj5hBiY/2ijyojLJV/sP97PnHmZxCHzGAMfQHBjLDq
4SqiN4//U19fpmHKccAma+SNhVDOHJdas08FsvAQsUU+vUB8l6JRh/OHQlYbZ+on
AO35VMOy8CEMGfTQu9KGYMbAurWMP/8NwW8hKuhywWufMZ+SbA1ne9ORDLLk7El6
6nSOu0ri4MLocZoritxKihPC7WXZ+P1vmrw8PNe4Hz9x2LQupbL+deRh0h8QCxYn
lgImrU1o0P77vNn0TcX3gUIalTp/HybMnEsu/U6bzRI3kPa55IhE/QqpHKofZaIh
ubABjx/JjcXTZcJFrMVRUZa5i0Yx63Pe5bHnNpdPLtb5EOAKs/k5VCQ7mHbtCcun
L5nKL8HPyIyVo99pq3+RWFct21f55DWla4/+XYvzTpdHlNVyF5O89RsB1wwT1ynM
73+1koBFA2NzLoVWTysolHDfifQ553AMXkL8aviqSmYpO02yQx9jU6wxfv53pus/
40JanRCTqjvNWSzQLEbMdGaL4MzRL1eLu0t8jjDS54/dJOR/Rbcho2CwU5NiKqpL
9vRi2j0XQ4lGZXAYVlnyR1GVQoRcWlrP92gZV+Mc5kTPHG0r3rcqEPckrmJMPu1R
OaqxqdLmLVdwrCnyzUG6LlLXr3gO9Lt21tbc70qTr6ymXy2HSEnSIVBA7hrfrYo9
qjGCmuOYvKeOtmK+QPBd6Tq6PXvg1Cn3E2nb7+rZbtQMDTX1G3kEWu/P52QhKcFV
grD7Cvwu589kJTVls3+PXDuSvS8kl0igVglj+71pOP7DV4Qe2h+5av0LZQYNx9+u
3MNgfDUBuC8fzCxRo49C/wt2igjsZ1m/VltyvLj5q9b6fndW8vDIn7rMc3kNphiR
gLHSv0dDgatljmpDkDVzPv0VnwTEkK6cF41/8cWyr4/6VZNA7dyM8DiV5kEQQDWm
VXlqEMh23/AXIODBzO6y+WjqxjLHLjXMtXme6pewmb2qV1zV/BbmHv29kU+zxuDO
m/MOep8vN3CgJNhxSmUa4vTb9u/j+jfyf7e9+RTq8Oq4vwazCN/NP+hKe+ld+1jg
dWWFKpEscDVE9aUr6pt4InUXcRCBKmgggc2U2rBfHft8a7ptgD2v2g2g+nv/nXn7
PmzDAzY+WJsUCmgv+4JfM1jXvmICOZ0xjXIHBQ8o0kRE+L9Dg5/vsjwAMd2jE+Lb
pQrSD3Q7MQkN4VmGU4AULwj8WEE6zRs/Wod0WYFsxjs5vAyWaDKv5NhdEAwQil1k
zIZ9lpxjC7wiRHA3hDrKdgv+8X2PQJ69WSMCHydq3lRqMEOiMGqRaieT036sqrWv
/OvqAMjadA+c8jN48Rs7uFqzfS7inNUzy2U7oJy33wx2/N2t6BqU8hM4ZHm1eH8m
CfYJnKprG1RlPuxM13PudSlL4dootGcGtMil2q1FrIoXdIIH0X+D0I1KTES3ImyX
BEZeSpBKdNfN18VfvQTRz0ksJ3DJge5vgsA56PY4BSfe9y4Z/jaS2JVXATtmHYpC
3T4nsYZRjdrtFKxC78qwewiMu8I2CNHOOpP+Ho27keXt8DpFIlUCckEEyAX3i4vZ
A9w9+IVVcGdWDbK9lZsqLWF2fN7uOfqgMMzjdzIbyLdMLADNZdrk07ldBMY7Pp54
DxIPb+t66tqCNv0Y/yztYEvDxdwFwJs+RLzi/bbNKzfBkzxAzTF91Sgl7AOwyW2Q
NQ8V/QQ6/icd3S42teoqleATMrFUzQEEa9l8vvPMlDhaYoEvA3Q5xDv0wYmeKJ0y
cypwStPYif+2/oPN9GxxaXju5+3JGJlPX/dcDXdeu8BCFFsc32DuX2u9jC0NsKBg
rJWLHamAsRZ2FWAlldVA56kk7vt1hyAM7guYjiGSRJzEL5wnw2eiA6AodRzaFGw0
5r36SRMqoGKeGLQMSYmZRZ5Q5vbz5ZccHLrfpCxwdy+dFd3ysdps/c08yCLUJAjz
XtWe5vgqPJvf/qbKxhNoPItHn1D3lQ+GZPSe1zqzfPhSlHVpZwOGCCFbDy8w5xbt
+4QOYlR1e89Qk8vOMSbKNDRJlLcCx+8TrYsBc4VCyQn+Xc3aF7l/FawtkrH6oAxO
HRANiBvRczC6OXhVwVN7wtFtwq6ocZNsv3Jv1YSSDBr8q7mKCS8z0m75i+jmyK8o
y4ok97BPwQwqffUbtLz2loWG3GumtwqZ64npRmFHZ6hBOcA/j7jC02YPXIjrcATC
zFMZdFuB3W2WFyOPxG5U2Z350fG+vy7RVruEZ9F5WprOE5NNch3xPm0pWt6OGlsE
rVAXMKGZR+8Q6ZxAsZv+Rcm4UqsVxvoPDMgkOLtF9Vuxa9C7BC8ualrv1JYGZCoZ
PcBeDFTOTOIrS4x7+H/jWs6uha5uEXP/vP/iksm1HkAm0z3wcmIQ5DeU0YwaLsqh
NH2fdDAO4LzWvphUOOAlbAbYSGWWDKoFTAOwZGCoKMmjBm/jmf9neygSyX7Ac0WW
HoN6LKfRrS85pJrStGUDSJfnvFWVJWOVv+Wmo8RsSJRHr3mRKAjaDzS7cp2cIavE
uuboKZ+SVuFgytg9QZHot+AIaaqE3vwtKlPsMn0vaJHc3apBT7Nr9s85pri1hWp9
gCncKhSsf22zPoF04UI282SEoZTQf5kYPmV3HxEkoEMAftHlQokOTVkqo+51qU37
JBt34fXwd0pszP8VMuo//N6Ydz7ILOLb8965J94ZzBIAGSPQeGoYRWrCNrqENsF7
N8o/Eeulft44QRI15LHWGlWChhfV632LUfMURuy5/a/0zM36oL8IIpj9Ek0wTsMp
qyr7mS54U4O7wYRylCsw/tE09oHCwQInkoiG61EI6gFeSceukUDxg51Usgz3+AgR
fubfQxCttQwEIyiH7PKSeuXvJUU6N+shMxXM/HxPDjYMcszHnn+QlZ3COU/j90rv
xEkq/afmIZXxkDFEDqbwUJWxuuU9hoUZ5PAScvQ9iMY+zuzZqh7Yw4OPEIcGOwtH
UzpGhbegSn8evjPAOsPCgOjzUgwne6I4TiRNPv5S8g/j8h/qBCIdFC0d5D0dQK7A
37ese69SoiJdRANd0gGHJZLdMQFSlSsRnocvqg2Zan7ylfMDPSsYD/xIpixCCSJO
Ejoc1Yx8SApF/fFWDSttpR+kH+uZ9YQPJ4TojByIDwyNoK+Ekoi7rToK3gV/gwLe
pKVtFrLBSUrCceazozpOhBvrQyGW7PMBa9qjHbEnnwW8vXrLwyyRNfSGyGDH9x2L
pd2BwIw/glCMZV5G0cLGaB9Q3LYYhOQr2sJ1JiojKMiLcoXvGOVEtctrNQfJPc7J
Ubfw5xsy4Bc6igrmdoID+f8+qVOkonciRQzB7ZgxM7tBT5iFhJdhq0CfHdpNyewt
ChGi5yaSnS39M8CHE3CoMdj2jc43rYGS+6DF3Wbluk8DfBWcsjYpB5mhhM35jHvY
A9tW/hivnJVQ+Rls9LWuYs+GTOBlFoa3Zv2lrZOHIFjzpS3duscWuVMbCIUPNpkT
q8KlRx/sXNpMtTkyr28aIemsoLPJBMlYlqad0vwtecUqktgIn7pBGDuhR8J7rvYF
9txkpDzSq0wss+RtQUzDO/acx6M5g9P3/CWojd0WXO6UpvLueL83yaJm15T/VNpE
hoDx7rDUdq26H7DuLRX137bOEfV3+lyQ9mj7djtYBuxaA0G80HI18lfdOSgoRSX9
SHvCPDkYKsjF49TOVZ6XMth9QEHlISSzX+B7CqvwA8O4/Dl1grjGpCkaC1uxRkjC
F6Lf82UQXsi9pnb2bc40HS8yMQlzpOq2XUCMNTKhKkrXccftQ9iOFAUUeo1xk1Jy
ialkLT/iu5VGyteB9Z9KQK4X5ibIUM5WrbiiIS/4/nuPjrW0MqXPPNNEdcrE6xay
HQJWKWChMEOzG51UylcCu9A/ZKmdtnbMvMsmNDUYggOBXxTabxVk+MXHvC1c/8Qx
rS5ieVDSoTwvuyCRkgP9CGOP9UgFR0YYlzhPuQLxl9cCSjZtOiITf1bUzhspWW7V
3bi6mWPJHexav4KffVDX1GRPz6gx+2q/bSCPOb7fkNjMnC24fMuw5RGTu+GzyHfN
muSoaiQ31IwhevGO1dEHqz5ywVo+EMwgz5ZdHZLXNUdsDy1re6VLlQffPltzfb9Y
h3ONvOy3M2TOj618EUGvNOWiiZbz6qIUUWc3AYtyFiVBV2iL2WO3gDpmw8JjQTsB
5yE6bTqX6FkYl0oOI0ki/Bw0M5L459Ffem4in9SuvHLdeO2/5mDwgwj3pv8R/uGU
lXm8jgQ3Yf95BJEhoMzToU/ZmPrmkTYuXvCEgKDYyklQc7QXP45uX3zo4YHV3jIl
/1PJMXhCNjqOZSEco1k8b1zqy/b7akHq0QBVkAz2kcPp45uO7Bd8RWV8fC35HWmt
ZOXN6IGcv6CYKoilHbIw1BUifzcODdMoDrez26Ioa7VCU7/O9skG33r3ZlXz6A/V
ipaO2ORCTNpxe5JR4u/my7N0K5zNevvEW286vyzrviYaD9kXBJMKEM5FA3bTrliQ
IGv95tlH68JAKlNOoxnOST9vcP7aps+K0X+4bsC4KPMP33W/pY3oLgqdK8rT7gzH
zw1dGtJN5vjQoHzcP/lvDKyKcftA1odrCAwrKpPz2dsFlbxzdNi4wbm1+UALVIND
3FnX5RVAu1Nr8eYhQCbC/1SgtyPKY6BJADjZXh+aEGJ+8X30olMrLmpQMb7Lc6e/
inW+U9kevSnWh0F2tbuiAxYeHnL/TFY/YXnd/hg/DylvAhEFITy7sEzPPbM3sHsr
ZAaJ+dUL/ortfp5x4xNli0ow9mQN7CWIzK7jo4NM3st4mp6fXqQtkr/nJQvEaPpA
bbUl84rhQg71Jpqg/6VO33xR510LXsVhautJloQuKoQZN/Hp1N6YvUYXQjJ5nwbe
pBgOTphFBtESQxJK0nC13RvpMnHIvhYxLhqd6Pm5IxLty/TTxaGYJExruQdigxvC
tpltZh9xlc17hYyCkvfZ2jzm5vR2f854UtkAOqiNysXDdtfEO2lcx2v3TAHlmMjp
kVihZwgxWuQF2hbLAwREq4u3XDhalx4tOjX46oPLYoJkWmfCNIZUd7pXM060XRfJ
i7su4jHJuFHFLlZrLrBN0CYAs7CpUeZU3EJdsEoz7mQmOz68gH+nuM5+6LkZmtVv
5wAtZXnFK5TIJMK/ISfFz8q7AFuYSiu1z/a50yL5dOHCljahtCu8Au08ZocLh4PA
zD7J7IzLCLv/2SEcMyNwPMHaBvPnge9SWffV2T6yg//GAdcqbHN4Z73ONRSC4QJw
srOxr0kz/1Yh3NS8ruxtKIZRhw0luRrBKIF0twi43efr95A5UP5NuE/1F2lP8HrO
npgQ+JwcJRahvSslAL031lNHykJZ6/OrIH7CPFpEBHhCQ1ab1fupBIx/qWxIS/Qz
EksIpl9nGC91sDguTMgKSLTnnOvpIIqWNl3av7rEZJ3l/FGlsxsVUvNQ2h0Xd7LS
st4jFjkgGhhPO/uGg5cW7g+UKNwwxJwQzC7kh5Sczjn7qw5vV4hgPj1+YO+jGNJb
LrsYby01+zlLPqssrbQb5dLQ1gmQcG049vQZ5cNbT77Ktx3181y8t1n/zIXU2tNr
AHlCZ78jHemJAd8VMSgSe+lVooFiAqCURQ+URpBhd/9LBnCoHPqKxGZIXSdMUxCG
MQr7QaPup/ARo6lD9g22Ipz79auMzcNcBcdiwQVOJg47wbT9qJ92H1eHnDbGwKaE
IjUyFvhZomGeJSgebHrtG7tDpPPejuuIsh23t08uTmdUkINZXxLHzJEvqLvT0+Rt
xbCoesPilCz9uq+ijXJEbZncvJroiIs6Ax0NFfOuvw7cF3ornKWEjEee0PzqO/mc
JMuKPv0cm6e377f+ka4H2KgjKOsc5q253gYUepN5por9NLVwn0Mh5YyIv0W507SG
U74tVpvAdEBft32UqzxLG8uXvfBu3ypNErK21rxzvJABoUt61lhjrmNuGtzbYOkQ
UuR1AL903bwQ9K/QlBSVR2J3G/dbF0pRuyKdDi4ghYtWBwvFHqlSCGLMgdwMQoLx
Ytt8LRLX6DPVKLwXlXlei7NtN2hkDA0hfqZ59uVDbIPhbWWpGbmOsAWW6UbQjBl8
mhow+dXIUxxUA1exK+bit1vcKHqY2knVFfVhltQo9nHqwRxu6YacrnkCRgpbWALI
6SMxlhAZ3X/sEYW2BvZwXHTYb/xQctQLWih8QQK6UW/I5k1gT90KTSsc0/Pi0L6m
ICEm6qDpyzZaSUMAkLSM27cq1eoGZnzjUC6OB+tiQG2Dhvh3m4MFI6FFA8G6mIuz
qn8dTCROSkHA9VFZGOqEAVRsmB8TrmRaK6rKIpR6+oYkEQGIGxY/ss8DJ5suRMXM
ShK75IwhHyNbp1qaqzUzxJ+GObrQfyztWt7Xbxezy86BD5ZT/G0JHTfZHBnnUbDX
Ucm3Jg5RhOiR94CJLYX3S5WiCG9p7gqll1mavWgE+j3bXMPXG6wBZ8T8Fg0mD/bp
uxUdmXH3OW/s3obCb2aC1ojFzxYDvsQC449hNgWIq3POgdN5Lbv13Ak/xR1dUSfC
hQOtH1+z/DzkGTSepw7aHd6kPMZK3tGLvlL9CULrTiGXFQ+YvjTOAu83O3kqxiKD
tSZ0dcism3IMXqEOO4AptHXy4OJ6G9nMZRSnp541obcsphJ8bFqRDI84gJeLHE/X
PP7AxMU0H7mvmfehEXKqUGfW9euDMuPI96mnQWAJHkdjUZe/Xylhb4lWi0umDfuu
kSWAWegIogpFIDJ4yZ9q+jbO5IPEukI2fTTRtg4GPQnotY8lvl4A6OzbQHk4cQT3
ZEPpoEi2F+rL2S3pNt9FZBdHlpTRJ89FQGL6MJXH+qaKhQ5reUIt/wmZbX7h/Op8
xNN0kbt24RQU96zue2R+OwfvL04vCKK7ibKDC27DjyaC17wrNKy7BjOFpNU+Pcjz
RybaPjUlOA88ghDnAB/1914ZgUdf4dsWvrfkuTtM0Ng03kuU4pNYX045/sHsMHXp
1haf+5bMFZ7qRnOY/+8ypYYhPtIxx1/bvqab5YGf3FC7cTG0Msq1zJmG3haXhk1j
PKfklMw1K/885HFDIJ28NWF+vTnWAEYv8zowi5Sucs4OcVajCyGf/ng4CckUNT96
Sm9jdyTNXMw0fJScw6LfFXzQG0sT//YE6YvChBnU70LoYgN12GwZ35YyPf3kQmW2
U8MLvyhWBfZr1sgiD0PBpvEq0KXhVPUOPTpsr05SFpnWvRMTyTvVjewwxd+YsXtp
38ge/vj42oJFCmGSrjmvibD5iL5AuSoTFy6p3aaDlX5wmyU43QjbiO8YW3ZHuM4G
gK4JPifL4WN5o2bQXsaSkMAOdFwv6iVgpYlvQItuOsmP9lGNZLONcuynkAUNjDoS
6cMkiQHKOkYM9DLvG+0HzA2oyWpSrBkPxBV5/hUoVcukmG/p1CvPFYFyaVH/fa/J
GQiVMH+0xuVqbEbnUhq4RzFRGDJv+GuBH/pgVGf1X51dfWCDKKD3HZflGI2LTO95
uZ6cRqERO5RvXEUmXRgYwnOjf1D7OB3KOY/isVm0OZiDcXX0OeYf7zFugsbrun8l
k6sSmqRa4aLe1H3rKqG9Kq9AkBP/em2Daa0+HH+kuxKLT9aMbeu2VDt3r4jZxNqL
Ar3O3IVHJgpdpo/k/D1tmYAZgxJVVLwHlkeuDPDb2j6lfUtchcma0f5tQHmTOhRB
/oSiINWwBq8XA8fxcxNl39mY/mfaZXai02VhKpDvwmKWqXoe2g6WkcLaelCBnyzf
73dc/l6tzifHtDEGIkGN5MZe0qBghv2C+LVuurCDe3pTGETYKE+8/6IoYnb76788
WJU7Lkf9uP9SMruRm6wC8SZmEYR2M4Yd9kd7DbnaLBM7VXOUyMvVAZ3fHlK2VQc5
eu6bT62rkz6w78ZAfEaSeH9RTUXg0VncmPoqdNPbFkYHZGLK67oAb53cjugqB1G7
4V2W49ryGoNnH50Q35wzn4eoetgpFPdloyP5h2bA3SgQuDnYAvi5/gp5q8UGRCTF
9C9v7JfhcNUsp9cdBYAqTRkUiJbwRU+LKyZHq/A1Ft8RDPeewx1kXhPyrYpMjfWr
PyUd76F+CyMEEnx+Np+W5gokYDqBgzT86XLv/XOldoDJXOb9jGpMfvCKuQHGwp7D
ELRGg8i8dKDTWBapHkS1BqRFIFWznEkUDNWaU1Z/08wjikIsbw4Ve6IsNVZukLBj
PfKnb3YaYwpIQ6DhNIymeKymWQQYFJby/aZaf5o30vSFXU9UpApR9qZMk8m3Hyc/
Y2+wOskX28j0YT9K4//X+lKaIXnBI8peWa2kGFDD77g21TK9VamOdv+kAQSn7mT/
VccVWQ7gWYmBMqb6mdmncUhbvP2fliZDWRVq3oRzXFjffExSTIxVKyjl61Kh7DXl
elhYLC+SzUbC+9YArhrzpbPGm0qUatn+M2g8p4ogvUFwhb6DdbM9jaG+mxeR/LXe
gEtBeQ0g6X499ItzmICCYW4xAot8UE3eVXD2gVRSI/eSQ8TyJQjofIFBalyJX9dh
Z+CT1I8CjbgNAPeHVLkWGTRmUJ2pWh7OZIBuMw1PYDnW8FFl5+834kL3ksCy55d6
FoBZwCI2rRn4ZpJhEEG+rZWJiJGVyIZ2zeHXkaYoCbGSgAbaiNIJ9oW8anpJnLvC
GTpGgcQtUyPva/7wVZXDXcVQe0UN34M16wpHioeyOy4Idi3BpI4gxqR1vdOi1zGu
gxAF885vWQXVIW9NikM+0o8uCSNcdhS2CNnHMK7FlgmOlo//xRZVe0EJ0m4Zqf5r
inOzRxMP/mXebGm5TY0ZJs+tWiP1WcoAzE3AAcs6kfRCtHLuxFpM4K3LdlHiIgrl
Mt//Ttu8QzSR3N38e7mkQMjsg37mijVGnYKU0lg33wl8ApA+Gw63YVH0rEmD2yVz
NKASjrTfJTa/bJxpJPSHXWxxYGxZc+PeBm1f+aoQYzFbpHSYukxSUfF73AaoN3HU
kgFCcKjUKqbSbJ87dv097qgVGU86PjJ4U3QYwrzm9SvEhEi0tsEt3szNNKr0AzVq
pdrh4+cREHXbymDXVjuMAq/x3ramT73EE2WmzicZs2pCjCISeu+osCkGBQDFXHQ9
4G6VQh05oSfvxjn77Y062RQE+H0bAzSYle15YexBZ66jEfNmq/uq9NA4p9E2BMPG
FB/Ie6rclVfaLCT9BN+Otfm7vahN63DyUT1wvmq9VsGGpH7aoW6Ni3oklvgy96+e
xeYpRvglWzadjpOWgrpEaLivCClOPl33nUHcOmVBzCWT2HIHauQtfehsKpyjSBEn
oipwZTXF5UKkwMtldniLHRtZQJA3AiLo40yz/0zFziaxHVQh5E/0n0HAZQmBqw39
WYxkV1AIcyBsykKBAbVGSHAPEe4EjLCHjmEStwjOxItRdCZVtbNE1F4GRsT4DnME
keQ0o5nhgFBXVama4g0At0kE/x7oUBZxzxgTylht1BJOuq/AZdBSiCHy5KA39DVA
J6gAbaY8jFNo80WW+DtkENeSjxm84hMhupDvZA0genMbrZUehckx80s4lharpYOo
laAC3hL3BLVaegnL3LSp7xDjxgcqH6c7V2TdTfiNt7N7E891/UR/IYTLlDXeci/m
mwqETxAXpZ9hKu+Yhex39wpDSGVboOXDQB2RbqutYsKCtDkjhuJ+MGt4QgwztPA2
8l+0EV1LILd1Uo1To3GxL4C04lh76sqLFcazgwG+i9foZK2iJ6eCqVfxf4T48MN2
FfFNBQTG7QpwdkwKxAllXVP6n2dk+Bb9Ko7KKNzwtZMVEkeiV5F+zHym0f9MNbwx
qLdWyF/wyWXBjVTB6dMs64ToD3tZZUdj7rrZjDnANVZ/mnL2IcJ5XueHaFo94ja5
rQHADP0y4R2/DqEDPKGTjLmj2ZH80PY4GqxmAKjK5Rn2f5aYSh1V1yA+HIc5I1Xq
iI/qswiP9b1Ot7Q50kID7E9lzfHzalIuJN9Bwv+nwNOXGShDV0RB0CJyuo9z77V4
GK9heKGoxblPNIvxsy9cv2WHqfOlCf3IESlx9/dpZDLxuCmvrRvQ7lbcvfom0Jg/
Ey6teAn8UEAVeiRBXwopA1BpQLpYeWIVJL8/038tZsClZB0SSEMK786+8E10ef2r
z6latVpwgAkRtexoBr0nM/07b6SsMRz7xgPGGNhJiCnbDSogrAR8aTsdhgbrtp+X
D+oJSyxnnqT1idPklbFK7BovO/yzLsUkyD6rqsGNqO+NVbbI4bcpzzl4R/p8lXV6
/dQqNZH8zacKZFydgInCbVKEoT6rR1tyQByEHiPuY7DCW3A1vp9yJZwDapNwP9k6
IAUpnnH2WOS8zbYwZFAvw8G07JKCUblWN3F+3g59mFnrr1LQYOHSsuRwqd6iNkYj
iaBJIbd4kevHaTMl1NmcTvATV8m8apeAZg4PVp0Iu4lbqjerih3Fvi0ATHliqrKG
u54JMOPhoV6NfVh61pn+8pJuqXy73KxpGwt6Z52d0kb09jQe1+N5NDMW5GLqpMsa
zMU2fud/GsCglqUtbSHYZdiCJA6bn2DoWwzeckARv5fRnk2AbmcRwshHIG3cOcSj
Lp7DPgEbndQ1slwxC3cxPywHxbKfJHWOnKtYPdxsqkOQovXy/541EVFPFeRL4i3O
BuFzyfwdFj/VbAprJvj5IIyFpBBcTVmjoVPbtx9daOmIG6plMainIeKKOoMiH8kk
Szj1vfWPdDFSb20OSYlul7Ro5RHphGMdTC+p4a4FinDva4P7/g9ND8ITm6HM+twS
GIlJr+X+fAIvfRoygyMaj+tI/VfS/PVG+9elYhM+uIrM48zK8FY23iAIBd2WnIUv
FUGIcGif0QzeUE6jO/GQA8CCszdi/o2NWdmdy+j46lJ52XcUUrWnJ6DA859FXMDn
jVXE5kc3iOLALtpYqposIhsL+XuewWZl2kXmV8rsh2xf8a8wn6BTiKD3LED447q9
04nO0ELZgD+IdXoYZD9SwbH83+FZ2FpZSfgJL6/Hf2aem7vgaTTLIifMQ8OL55va
j1Vby9XyJ9VPOqzVdRzbUFNCgTIhlhITmqANqtXWYcy1QPkYMyftxId0HLrURv4j
FCNiULvWPRdX5LGyjHVlfkkgOazVulr1j/w2/wXNdG2oBCKto9yTJFWH2p1raYBx
vJUVwy8REZ0iQiPtFEaTRkRPBPE+l/PLHehBJPPumNVDEuGXJs7EsU2F3XOIGS6D
zMUuJv7YlnSADjGIf4Cs3CWi4cfa6Z9vaSnyd1SGQ7HO43GZN2X4JZqPXhiEORsi
qEyRCLDzrQm/h5Kdv6r0HFXutd5bqtdlEoaQsr5fwUm3LKynjx0PXZ38ywKs2hjX
pVvBXQy+YU1fVl4sa/XHagsE2pXH7CEK15YVPFpqnKBvhZxhLDikH/kvKKhD/mPR
hjOfI2MZWpDuYZzTpBtgltUraPhZ7K3Q5uTyxue8S7emCrHUwIn+Jzx+cbgbv84X
uvm/tkhk53M2FVtqlktOlLLotRtWXwW2ihU7KRytU5agDCLvVNJ9wwII2wslXWHM
5XGMmA7Yl7M3InCBXpRGz6xGTy0i0aqP6gEFK3xgztITtb+umOzUMn+Ib0MclSUE
u+10LnDhkz8qOdifwdLTVzvktRaa6sj1HMU50QBDj55BRpD+vTfhPDrpVR72Ylwk
4Eo8NiZA9nUrqAn307XWcLpS9yVjDu9wrfwpLiAeZpQ2X7Tv+uhdk6qhopIKBwlh
5knT1uGeh4ZOwZILIdnv0O1I8NnMEILXTRQ1SroNTz3EJahn5JgY/eenLt/0Y8UE
NgfHMMIiVnQuGHuFTHQ0Ya7e2AaeaEzk5IrMobRRLPtw4A/Csjmh6a1CHMHyS6BQ
2KEnGvR3FqwAHnqpS2kKk0omi3iv6D7Ee7xIxVC4fQ+mtfxICNsTrHpWnbn32Zmz
05hUqJ8KAHNg0vAkqMvDnEw30qmH5hvq89HfjaukISP8YSqkmPjkGkontpCalwg+
4KCntnNF53BdXlE3Z2W/4666yfGtbxylqgqRzor2SYJ4jHWM+03fBVoe8tIkbbpb
oS1ifLghb4cCmh0HnmaVgpWYIphDODVN7t+K63Ov6ppptiygRZgP1t1v00cZkH++
Ui1QWru/9ErSoMZndq22H3IJscvWg3Q0F4PvHCkZQ/B0vqtGxfiFaEXIx1YF9Pgb
A0HSv5MsEcQJlYdE6UJIZbn0g5L/Jt/3pJ+yYQTuwKFRod1fu3Jis6MGtWDkdo1I
lnAOiXXFYzmXNTWyhgcw8MGnYi6Q81UMoNYDexONjycf+KE3TMRx37uTaCsXa8eu
HTmuY8hWmEL3h7u+15+wGWzUzMo4nJOhVhTCbAA3UZ23B//3y1okXEA9LssLKGn8
Qszo6rGsiOkNOJSDZNE9vZFcRn8Czi4FvQS0sYLDtrDdd+hDpSIDgGrjkU3joK2x
+UHKXvO/V7UO5kPQJk6lIjIpSi5MmMfWCOoEHCIJ6cO6rDwc2T1R5Pv8i8SmGA9P
phmzG4FeIOSwgKazqkH5MepNMW/Mu5rrPva4rt3Rc6LedsXWj+60I8VQdw+hsmL0
/W79e4L/LsqMOTWpzGtHbhvEDfkhl0t6eRKxXpZh1JV2eeS9zxDFY3Zy+yaEcup7
ZwbXZ0lBJ7UwdnZhydvgp1LYBYJWNjaGA8jM2tuujIizaIdJ0OkPzy1T62A/oXEw
Vu9++fGVJIAzsMl6IA6DQjEt/ytCUIcQOXzHBcQXFNk8xd0W50VbWuMCyScrjoYV
PKu+iF09lS2n7DYiN1Fsk9KZlfxIulMhkLVcPQ7d5yvn9C4jPVT5uLfPI8nW+367
C18TlEaYz4WjXhcz63MBcMekoxL9XqyZPHrgsVBJK6jnRWkReybPbXx263RoHhL0
ABP7n2up+/RSOUywTxwyYVA6BsJEcjSf7/Q+XLxdRm3Nhj5OrDRwv5k03ZdHXIhN
1B5VDzQOW7KBVP2+1GGrz57y2OqhIBdDfmQdisCeFKKJOQLeFH+o/aTUxmG3hSoS
uW7JuWMRPmIk4lwYvsyN2AFWQHGHjPF3JlVXMDb15FyxNqqjazR8mOdBi6pahzlL
Nuehe9LRohL/PAMbWS8PWkorx7UUl9eMTFhQc8MrSZf4wJuaB+VDnO8rFKQIZtC8
gNfWxofZ+uZQ9G5hk76VVp/t44hG6TWKbkqfqeelbx2mAcvoRR1uvRVBKjiwONUM
xzf4mLjQ4Dxa7pXxofPHXOmqfYujG4Newaj6Yu4zrFVk5oKuRk6WEfFR213aElWu
/O3KrM8W8LDtS1QTQjjS32Fey3zgJVmt9IpLkjdawGYAA1phXvO1qdbNAVxQrbKp
zbvrdHoIPHTiO2PSZ4AS51MH8ioDqXlGCU+g4CTnXjmDzYGCiAVHvOZH+kMVLqp0
WmHlvhWU2eKIU9IAb2N3I/vz75fJR1e5Rzy7eHPKUGHaUM9lwabSoD1IoPg1UbXD
/+wzAeeQwAevg3f/7Vzf5Od38fyD5Hw+r88CcSFx1Drb3mAa0nTpU57dbmgbZFIs
bsU9cilp6XAs84gsg4NeV/hOEnvhFlhETPYckXJujdVIm0dEQBBflgJxOkl4cSPK
bdYq+dJ7Zdvd45EvqQmCleLkIhztz0VJOS2hFwCokAVnvYOoH+AsNgQHXAaxMTHv
ijRMV9oFWO1dYuJQXvH2utg8k0lfsaHzY5YAr6WE3y26H5jqAYTHrU2sdY79gvBc
zStS+ZOPxryZ774it8qOmeYBbUDfYwT3uQIoWl9eG3p+ntHZ3uvoR9MyEdsKBsdr
`pragma protect end_protected
