`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k1IpSgHUefUp2r9z4PhtWPjwY+/anm4DjQNgE06frKRm9117l2cNCNqvurbg4nj9
ciqL7/KaVcFrwLOJnu6LavauWSjV8vgYwYRRfDBxYu5aibEbEwhhf0PK600zP5ud
FV3Yl0E7S9/ay0J0MQiM5N2simkf04Kzb3uzSRxAwsY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
goYhK2anl/FulShC8063iLvoxAwgivEjc0sBcQfvvgEAMzn5hfwaPDOLe/x33Z+M
/2FeKKQo3N3O/5m3XwKD6ovTfDe9PRQEnAJhvmy5Sc8CPLzAYyoXSSt9MBF2T3S9
X2gp8tzrK2k5T1S8RJV6k2FKmBEAI+m0BnAKA5kn9kEWUvRn/YqKBxnb9hs/5tsL
YNvpTCKdThFP2nXHIEKoBynhdtZ3qWUIdjGmZCuQ7za+LZuwZCK/W2lRS/MlyaSK
cn6KK85IYOUd4NrvauM50u/VN9GBD0uw4UuT1Otn5vtRwlR23DhRnlMExXrEpnha
q63cH3EDn3CxpM25BtdsIKl1NJtnGkpKI83qHnEyBMKgOu3Uis72ryBv3m3hEVAF
CX+Y2e0q4TWftl60LGjdLusQpiZqvFryk7OrNNJgmUPOfXL2gziVomNCoL/AoWTK
QfnxzFoMk0ViY3UsTAW19AspoPhPurvYc6SY3/sydjDX2Jk0jn2pd75VkEs5ETPO
ETTKmkqieRLj6uCuyCmFARe2lpv9Hyw7EL+pT2/XEw+yKOlvIw5CwtiCBs/pGQO2
PrI/6vmDkGP144+0j7fP9FfdyKnqDO8XNQRJCZER4WB74UbLfVl9GDYeGuZjWOXA
pcJbZa1A3GSoH6YjlSyIeuQXdZdlf2cSmwCzUnUtWdnL+6WQbMM8NoxtzX2IKqX4
ZJVzJbRGIzhgH+Rl/XWcqET/ibuDy4Y4MVHBeSJgPwNmV+9AXVF2IHlXs2VKMVrg
yyZQIY3N2edofh1pp3YMHbhtfu9toAOWoW/03cjDmUumyvNQmIGc1wDF1jdUZuHQ
FHPLUQLc+5S7UnugYH5N1n3eBTakL5VWX7YtfVkjZRp2wyfzvF2HXgJ8qxEv9pkK
PTMtw59LHEjv6wqVlssw+c18KUrBmb5dnG0LPwMR1LXHarg698CLMERuNHQgfCqU
Zi1l9QraSS8KcuBOUlJZNldnyUhb20JThxu4KDOPFxUM4rL6UcU0qFQUzcgeUa6r
qsnmuPbHD00cWN5n1R9Ml9bqM1q+4MTOqwHJbJ1yHxGN7o2pb8a7vjO5aOroJGiZ
+9vwAOCsOVHq06Dg+1u4e2PsZMp1gvd85EUh35J/oTwFESASOJZz6cZRTLvVy2mI
TEf12In6nZasTKfyltK/cmn652KZHaq/1fRQJMTITb7WESqimSIcO1Yp115rWNmD
XwK/hIZqk9U6w9r/dzGLqJo1S8cgKvaLCVjIhruojNbiei6ENRCi8OkXRAbT1Eu3
j0Grj+m3YwLp95Bre+Be43O1EzOyye+Bdx+mx11/qPB9LFqCWZXblZZ9uXXw4nlJ
uc5mq1pEKuab6fK/r3pe4rUxu6DUSITgVqw44dJzQWnP1K3zM5fqoiMc966gzg5Q
xzNOAAMD0ZncaKGf28/0gmFEMJkO3XsRgVOX9SM4EqV3oX4ksoN15Iazhjc/aknq
5lvxoG90gAL2FpC5oT3a/ITVz6hIl8snYidNEH+oELB+/KhiOxX14V0zXqIiRlhT
mUq0RHTFnAkUzAZdkkhNAd1WLqVQYVuPD0iO8kFqh/Rp45fl3eGn0GH6TUfCtIbA
5efLVxTIFzxASQmQQP+7dq+CiHdXWgUMIPPc+J4klnzM9kB+7Lk766B3J50IjCWe
LA1u6d8jYzptOEArKXPc9HMlClesaakgqXrTfssoYKlSmUTXmifl6vayK478oxlR
z1NmyRbaWgVmeO60QrMQ6IO4HdC+ObTf8RSjHPG5DHeMOr0fgtCXMLLMj3dk0NTZ
zxBsSb6ZlDASwxnLIgjeZC8Ep9fDl8ZM4/wUH+wdG2LqQjn6jEZAAAX/eXdYAG6N
e2DB/T+5JO80P4bR8smkeF+LoAh5myQM9iHQOZHiTlBxzvADlC3auDCrBj1sxwPg
mThU7aF8/34GBPkFtg9xAI6kuvbECqDkQLIwOb6Bp7Be7liTKke7MvEfYiAQev67
+t7NMl1+xY1jkHs+lrEdFd2/hDbnRiZLa3NyDYqimueBnQCRFY/27PR4it3YCpEU
4aNCCRCHQFIT1n9maeFYd8LeAMCTUNbdpDxsfnFHz/50msfBo0/a5fBdL9Vx80PO
ObU0EGAJEQL9yGVQ9HChxSxVosCnLZqCCTbRt75OAgue69y2CknZn0v7vOZcx9cd
HJtyr2Uvkbq86tZnqGFqQo3YaHTJMyNWA4IBcc5t/xfs4u7O71yZSZw25Z1lmVhk
lx4nSCeGj0iUy8976OIWdN0VhKaJKr6pmJv3r+mdTNUMTk1dzVEEFXbfbaiE2aMq
DIRLXZh+MRksPT0jk9L7BNcnSGqJZHYXP6Q+HGcNG4+rRIFFjruFsL4RgxbZCv/N
TL5csHmzndUpBJsRCzykJQqzHArsAR9f1G8/Xye4etat6HXcMdkpVz8pSpL4DckP
/k0ZZAXNfbvsjFkPubfuxXG104bwPdGBVGyr76oQ8iSOsnMG/8Ru5dZWSrRT3k2y
k7Szp1eG+DKHZzpX/2yxefnlgmxHhiU7xM/Np+vjZZ/vwmA+t3cCAlgIwKC5q7z5
eAWzwtcGo9tosVXLaDK5cj3+fyF9awOLLLNm3QYOSd+Z0LXoZLySH/B2b22y4nJ9
tiQ29hEGi3FErwbiWW+yLD29/PhYiCXu3EChDTYXl+3KEwOIUYVHOPENI4BrkDTl
EEed1DBk00AAchWn99jva3c/b2j0O6r7k12+T/qyTKV01YH/vQOUwx2Upb/d1S6t
jXSgant/18HhcvQYO61jOizdUnQdhcw5KSIJNJ+7lguAMMH06orxVhwn11e4LW1r
hN4XGQmczhpWo9EqQRzwc0QKMCCmZMP0N31RqGcGNZ24uYBsF5uUNavEqwQjQ2s0
N1b9kNM4vjFBBchftge9gLVR/5gN7rKkTBC+Ui+/s3vSlYAiC+M+jIjlxisjUD+S
olYH2PU+qk2HFuV6J5dX8hXj0PPYI56kbQGDMhNMT1uhBN4dXxqAZDMslyrBKw33
re7e3z+gpTkBt4/SbF+G0OJKBby7BQRYRO4vkWJ+4LeptImdF19U0VmTc6CDINQF
LFn4sNSEenaR4+stBUnMj9uVjprglGN81INzojUlmmlJfLmTg711eyIVxef81nv8
zBWhq+05oIQGKGNLsooqDhIenbe5j2jbEahX9C5TxIqbz8iw5d7xljZjI4ZeLwum
3mLNz8ZKVaSBrAIw41YtDDV/HGSNBghgMF+hjJSxCGZsrJ6U17OVopRz6tWL8WAw
UPD4bfG/VQAHwGwWZWafzsznvXldvzPj/vAlQW6iclWiJhjBs/uPu34SDzpiIeTU
qHBzO2N/7pemep2jodnT8jNg9lO5HKIpjrThSpp8XbidVz87oW4xQcoX6VYpKvP0
IrpYWeQctqaMcGkhboYSKwg0keIqWuBdB32Hh+/tVNjw7hIBD0+l4FyigLKTZpnW
ALMZQMIW2rTcJnWyLf97ZHmluRizMn+jbV4/HCjIR7qe8KoHd/bMqJi2FyvVCSow
siWVm0cvCx0wCcWzoYrOzaEoOrgkMhC+tBZGUq7QkDmOHd+IIN54qJL3T5mI8+T2
wAX7dofJl5tQC1nvfMtFzly3JT+z4MP92A0t/ORXqaY5Y93F/fmsjLZO7sK95FbJ
xRp9RaHbVixAyAotnpVjHTdYsL5DMQaax7/lkkO1zk0jd2CRc0gM2jMYbEb75nIX
czl2C0JkE4w1hlAauBn0uU+uYmdTRkj/qJ1OsqU1A5jtdOM8+j9+wSPuiR4u7Kpg
NCXGEAjyIC/k5p6o3Qh+51mO/t6e5Qh3imlUoBRsFg5X75EbB05O2fQqnMGcHW6R
UAoAwAccrl1iyjby9Zgrzwzm1XqQye3Bg0KHStsQFFP9PpYTjy8N5yHd1Y7nQrIc
n3EZeOAACVq+nI1KPYnPDYN6uLCVatp4DAct15KeXwkWkFNRFNYq9yXIH+Spbbnl
IKL0aQZmAWeRvfpKlnU4ZZ7N5tQEfFscpZpyRzEWVdTYcFmRDYgYsJSPDSRPXM+A
tPO7WM1t2lpYAaFSEvWnAAWK83euIHBdZ/FE93a52ht+6qvcxwJ5f/D4ok08ITSX
diBQs+Y1JdD3Z9B5xW7qzHHFw8aFYZXGVoVhLdSxK+uDCUyJYZktCl3J7Kt0iKJn
skI2ela6l6qoouMu9pCy1FNtgZn8NqMp7bkv3mVT+n6PNFfj98kMqxQWynLt60+0
WHTXkwD5sSkqSeK6s/qVsJovIeUxzKoNFu95Mk2nQUiJ/bm4W4jz8sjVrkGKFqWk
Ld5GRGdQvo+QIuDRedKHaMsKHs7v2t/1iyWqQaxLodAzOP5C3+obNcQ5/ZLohBEw
SGXACGxBxvQEE+ubKXzwkFgBkcne20B+lrE2PcPWw9GnyUagBzDqNWJGFUQxX07V
ONBWW1SXCgrP5j01WpmOiWgUdsUGmEnqQMlr3AW+WW6Rl9KgsGg5Gpo+mLvRa5AU
pX3anT6Wss0rI1VnBp0XuOb/SeriXhj7CftMZO/gff09MSMv1Fom+I6/oRnSnMdF
+PgyvQS7TqAIbUMlfT4OAF6JorLvcpSZyzYMcYJ9n1as1cJWQRKR3T9LsuVlJoqt
FDDD16vMDpGrSRYicwEx0XAsXdp0+QHW5dPR41aAThcj/MUqj9CiZoadKvLqCFJu
KgwGrtnPUNa3VwjhtNjtOpU486K0c1GR2XVU62JkXdBpLcQRKN6GZY83isLWBcwh
zCW+05ycOO2r4wUjQsyirmpcPUURwehQ4qgvzBTfRZmIE/8CkfSxiVoDnPuJu/i3
5T+Eh+TW+N45ftp7RCnLrrJXtrIRlliAo1e6uNrwSmAkhGg1yovBPVdl2b5ZidpO
UGstGuCqQeAWWk10VU4VEO/rZtR8pKoilWCp2zvVFJD/3DzSYByhQbAm21eqXLC/
IhPq601jD/9cHKFgTBPkO3NdEDzOZnCY0aIU2nZWucGnlf27E/VK5aNF7SDl9yob
m4fEa6AoHk2Vkj+fsSoI18GgNHlMVH5UHbZSUBhl2/j9zGtRhFQSkKWeypeEELXy
YGJDFzaEwVMvJVjjmosdCbiYpqAfWhMPG9gSswOYY/Zs9bc0gWGs30W/sRqSJZk+
Be0fbdYCDWNq/+pIYsnmRmR7s92Aqe54O2H81tSKjFo7RuWC5FDW7FAHmAEflTyq
jhtxlgPH2IzozhaPmWCBvsGbj7eK5UdtWqb5kVMWy0TLT1pDafiYTapPpSyOmhcM
9NBrZCBHEK6LE1CZlZTaewSW+HCQZFDlP/WJC88Rin8klZBCVbn4An0tDllDXlXK
Ww126kX/zEecNwUUy6Hv1AQ7utD+K7AjLh3q13puvIqF972HNu4i+2EDUR4o8ITq
lNw+DLP9NcirQjD0nIy7+CABaj++A1beULN/Ilf0uOO7k+XLTGW23daVYL+Onzv4
xx10dlPc7AABikGpOdp9fDfVnvNVdfQ35UFgoFs+qphOpGICczGEBJ4YAhMAGAAr
D5A2p1KMm0rTDmU7tYfiQWs4Qn0o4N+7wa4ZkW28l9ge6vg5j03uZWG5r75AiWXw
BUOJdBzELTQb3CnEvXkM3F94xUqmq8P7kLGYAvpkoOVkYhxCZELMn7vHfrKXgAIp
7i8vz7Z+rtwPBK3xzQY24Ui/M0grrZorXeY8oUsZToUpzyvnQKqxu3+l0y+Ab5an
Z0cZSBMGWxDTg/hqYGpmuw9v7hkFM1/NpISLeI81LEDLJrc5WkA5eWGqFUb6226y
8PtDgRnTMCZHZq4TN3Aq9ueB2ipoiC95/ruRjwkyV0SoNjJShpLQLTRc8xaZDZna
W6ECC7k0xrHDmFyYdCRxKwJEhpO4zcZnfHlNjzf+Ioo4EDJZAFmiEcxvdJDvTyXh
pVj9wQbf6zSe4FmwhFSf86zoDWyMC/8vSTt+vxItF8NCZ66hE/8OFqzuCLm/EFlh
GXY0xeBAREb61/BLrVJxubR3aM+G0JyJrPjrUdQxQzbHstcRN6C7MyTsAHkkvPZs
Yee7RD55X1LNAmfbhThCyij0knYW+xiMk5euiGAxbV/aGSngYnC6WXY5h/b9/pft
gWyXQq6yeIzHwpTGp8CrN8zee/AMACoXGi7EiKWSxkgvdxoHcg030NaGSBwRyy1A
RK8Ijo4qH+U8ISyMilKtaOPu7szWracYZyXnFaTH4yzZLVECBWTEIn0Vv1Fa6o63
9E7ArD9SK3fGacvNMdFbWLs6XXTukiKKWCBZDWCqCPwQpp3tF0TScFNyNfo/kmi7
8oCQ1h/eZhnIHTXX6333qmSO7VrWVCFl79ZXiIx5XyBJCk9wk47OSqNRCbQDoEbu
QVweW94ce2F0pMICXbXdnIOe4siMUPdfDNWiLzJd6llt5YZZbJucs/KPbihkzHrX
L9LNB1IsYNZOL2D5T3UhkCTzUJ+jhqC6WSXYaEGgs9HXkyGUZsStWU4SUiLZ9+k2
Tc5Uum8QDcrZ5bq+Y0+4b496qXZNx22C1cKsgz8sN5uzV6ipeXCzTxefJAeRDmIV
YdtPtcD/iAeAVes74YTkz05g5XPTvQkeYmWWWCHzY7vTN6zJPMfBS2t1mWOCUSW3
GD5Jci4BRz94uMS3UOAC1YbYtK6mkVFPF6mqZyCnrmNlI5xf4WStORl8dTG03BBt
LlEtgmzwS/ilgin26pQHHVLyp7duHI3Wr/KsuMu/ZO3AsU1C7L/CeV2D0PFWlTGu
2KABoDMzJt4R9k2SdyQP1LSo2VD9QzrHrEnHcsyq309i6L+y9G/YY5zl/wpjMAUp
uy53cGlD925Xoe564v6+F050yilqgY8JbiKI/nXxLVYmg+Fq1wGGYKRSclbNTtfq
CN1+4i5Z6QFBJnXhzoaVCCR0Bb/5r0vrR3j6t5Mpu8R5e9f8ornbetIOfWxYyw1Z
kd/1uXo7XYWgOzACEmXscecyGlsrIkLaz1tkCpoNGTDO00Nlu1BGIDarJcXNLFqM
ZCkm0iTNvFmruwGMcwsevLZcF07QnvfyKN3eHwWxQpdkw4yi98NhltWdd2ohuS+v
n4XsF5T/DRJdEU0Qk43nNNJeJJIrOf/Dz3PPqObIMme2CRqKQLX7lDmmXCxoVWG+
4GMP9ohytidzCqkqN4CL4XudrdiSd55DkjP9sV8mU9bkPGNQFpKZgUK6+THLBMRa
BV1A7B2zclTY5zQrNQnPsZI8mbMkXtaX3i3rXjZmyxI=
`pragma protect end_protected
