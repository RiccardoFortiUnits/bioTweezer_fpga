`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ka29r2C9P69fXZW8BORkRR4CPXr4PgQ7Fumf+kaosvmmx4Ihp1Z0sV1b+CvgGbJM
UuLodNfWImn6l10K1ooSsAgPp4CJtzEuxSK1yII9l0rZ38lusiiCLULMjPoM7bLC
h0CU541+3DgrotDS6WM1InIhikUHCbaduFCQt4wZ/rU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4848)
CbQgFcbWuVa2eOTABL1L7uGtRnbbD0Kl26FUdgFGKEa7mSzACmx2RD9YC6ME9IsI
wKjSlnG54rxqsYNb7F4MsD+ZmW8Yd3VQWiOfcDcbaiy58yE1jThgccaj0nd5eUtY
0/sq8weFWk97jMdxFTzNkPemumovMfYJ0rXSBUpnOXdROK7CCgsSJgXBW/l9TG9G
83j2y/Q+/EueYbBh5wyLGUm8f8NE05NNyi+opTrwu9XrGej0GVVdsUcKFTHrNW/S
3yvo2RoAGovsuUj+p07V4Ae+WS5uosxn4VF49f7Db0PmJ+P6ehnmftzpKl2No4DL
/exePGZnkaHQdNNoRmFv+unP7nd7EMb7vsllHJ6Z73bFgCX8oAEnuSEibu5kd+CN
mQHRA/BJWasLs4OKOvK91q8mvBa66WXywIipNK3V94u/3ckeUXVfNEe95XLa5T/I
1Q03i86TEq3/VuKC7M7zMSHeh5upyMiQOddQbyKT3jbc91K6wHw/GhcngThkUdMO
yVubltrwD8rY9Yqc1ERi1CGpMDzXgp4wjrmNTWCQCOTvYhAU31qv7kTOmcDQL2zb
Rqf3XehGgqKZypiatuua2BeXTICgL4EWEHRCzfakgN+b66SptlOYfZb3mI/1O7iy
Q9E61UvCNEm8mqqBEnAp4ADkazCh4V++Hnck2uMW86oqNKpIJ6zavoXxXOmahXgk
3uT0wQ/vcv0Ob47NXNUtX4Jub7Qae2G76W1plJhwwCgmVB7ld3YH4qq668wXwnvx
t/I6QWqxUY8UvrvBWPcHqnfGhFXv1XUXlKDg1r0MKIxH7+gD+HDYvEurPDT5DZB/
JThlc+JWazRjIIEhYQizsFdQTty2uLYhqt5JR74eLG07J1F/n1TT8+qMvOC/p+Gf
wOkVWgOH3fWk1dTaP5nstp3BMwYxhkwZZg+ZXPUVBwheJuWqy3Du+fJ9jzoTpRJ7
pVjxHWLC/EPBgl13bZZxfUt6aN4Ik7WCyKn79cGPuHaxEwiRFc9HzrtD1N9GANVe
IlgqszDIG2/gc4AMR2y1Gc89o89ZoFVolQcPdxfRoPyrdx5Mt0RyDnx8t9/DdHCy
Zmnb7prdgQtWVaS672zBFECHwTGh5kN4aeXXrcbSOLFmD+Ug47HI3etF8incW0gy
nzRH3rwKC4MyEN2F3G6YwfgMViPlbiuWUtOyshkQCPFXEdgXaZCdNdgHyMEw/lkc
LLBrwbtDyApnOe4kmmwk9sZLswja+Fwk766qtLPiLCQwzEBy7gqyStM8DFVlwgHF
GnNlalHCjJ06YU8PKDc8z0ITaN6yKUXkvsrVRBqIbm5ZV86IT9Eovkvk4T+0Ilha
WumK7eURtzmHMMdxP9XnJUFIeCKJ49xejbz3O4yYIwf3DnIVupCu6c+3cVLaWxrH
Z4QumP3OKpxZq+cIVD3+t1lBJF+p7YxaAJFIywxiNeOvMRUEvtB8qp7O73cK9n8a
jLwVm/jHNmIrQ3LUhX+gI90jPzGAFV9mjhkfY/Xn+fGWs4qKHYD2pv+2J4Aork8U
ab9ji2gK2d3kvWn/GowRnrvrAKTx4nzE6XVJDDd8x4yVbAX8cFdmQNjxwez2J5Mf
YkM9LVjjs4qHK3YoMMAk1ZyXqb89frVXZvUWtRPYq4w50Q1XCDG+FbsHshadLCQr
54WleRERH0i3azdiJZujBrnoy/syiWCBXE4Esg44ziLEXSzhK6xjvdpEOxVmciVT
qiuyIcEE6U44lEbJPRXHM54swePNaG9UKDFJ4ZaRt1WmME405OQlMI9s9llpe+7F
k+TiZJUCoGlSGQSZmaTSZjn3KlUZe9M9WD/8/JZTQVkosplaBLWivmMKC5miAmO3
g8qN0N5+3o1QNB37Lo8fJUiBk0wQPfu/dXESQez8n/LySTfauALXwxXV5XigA+YE
wST2R/ntfX2aTlebh9dNpqB4pTjLpnyp4x18+jvlxSpIcl6E4ue5V1ddXMSKMLzF
o1sE6n1NH8faS+LmNDOMS4ODRrGReYmYkYg+cBFCKa9BW80+fJfi2MIDyFRcn15k
c9LnpqULpccrNMuFipIFzYf9TaOF73NzrQy7XCTBjBttcXi0e/eXrNwul+2+T6mv
+icB8SuoNwtgdmHLJekpdgcAjQ0ptJzp8QmsmcnBNrdn/KEKiAiH4oTva+qCAoEY
lPLZv614cX1goo/jW7fZjAZxNRND1adZNCjiXhYQ5kRb7sfktMH4fQOJdUNYklyU
E86ROysQ6oV3Ow+X1CLXsEXyw2sXi2Q0u2u0SFD8vAb8Ir4zg0B+GN6IQVMOQRyO
jdQqnWGv1h5y7S7yGoRhW/E7ZRg7QY5IL6rV41+skej1Y2l5e3PMCePVJyvCa9nz
RAp+N4OLGHLXBMYrbGlKzrTuy5u97SPkebSGNwWHRhSd2E/xD+tPFF7CuHfDPO/W
WLj+M/xxolIr8Ij/7wqBCTL0WMpqQKy1jmyHvVtcHhbybAHXyoZlfQ+xzDk48O1c
MtVlPyf4gY96zg+ZHPKkbUIKSr9XNjnpH6RwU8QHz8feRtIRFOud/WrNen2hXP5E
VBUBzO8zTJtbm2zUATJWoFqByxkseQOAsDEsCeqhOxKqHomGreKS4bwmS4T5vVlR
GwICtsWI/f6JIOggXr23YAs/kWTn7TWxOngl9bwpqFzpRiQ82ltum4CwKnvsOic3
gmUfVYAr9ZKFAdkDVgg/YTu/3WsjgqJQP2dzk+TakZcZNi64NnTO6sklILEPN5aB
5xHWJQ97aGOyI264cT+YgsISYKNDEETEZ5AqiaJ/71S2qDV2tr1tq/5uh19g4rOb
9Nlzr5joxC5R4rlA0/S7TEuSVYMVnNsIQMR16wS0FyKzNxdo+8vu2gx0cjgRiyMJ
gZVXszDgyJK3iwLD8xEel/84ZMh4xrb2BdFIP0uq1jZa0AWrWRv6HITeHwUaYc8Q
45Bo1KuH9h45/N5repyEN+ASFgXJ2ZU1lEwmvGT5sL/3qriqVXEyUA63T/o+eWoX
pUo3vtCW/p/GJaRLeisWX581CpOf2nb+tzSvPJ9X70rJmvZX72AcNYbMLw374xGd
8fCQwimXQdhhWoK0j26XGi6g7Wc3eBJ/sDn2oPvJMjT+NPTJ4ZjwKeGwIQrIqQhl
bTdHMPfBnY3ToPP67tuJpimbs/7YOBY/099t0xIiPewUEciIZFs24YHGQTJnh1Zp
LwMl44B9zMPk3Fkk0UzwQomGn708ocMzfWIKDnHqP5fQ+OMDsxy8cLAJHB4z1Ew7
OuRfmiiHRrJL6ZLKSNhPrWL35WJINuEoXBz55nSzqEtzU1UaBUfhyIRXUA3WZ5sg
sqATnECnCuKtfRdf2smnLdfyT1M9qhvM3n1HIGo6nl0WQZyy052h8VSpMam7F4Y7
WeJP9Itm0SsJFssoNHrCt6Z81B0chrTYHv8N+6LqrOyL1qh98OcC4x8PWPgp5pD7
AOzoZ5SxH2z6S7vkYg9t84Z9KfJ+S4dPPod49PBKnUC9DEu6aMvmW2FkWWuXHWGL
EzEuZOD2sUNakV7/IxyMzdjsvqQ6lt/B13z+jbNVEAd4yVkDzvoaDNunodAKM/Ax
b/iq558xF4vZoG6iQz2JTgf2dzwrmPnSECr0xcarDsCTgq3DBL+UoxfGiHmyx4jL
tTQ88EoF2wVm+1hleOEk1fEYdqYDVlQLStia4rToH+ZnXOe1HBPWqEjgYNqISxnA
aBqsZJRWgzSkMNlmLdVXDsSMBtAMVcboK8wIi5IGz5Y6jpBnzCy+yilpC27Nz6FH
0GX8ItZnB+sLHwGDrgvmcZ8gS0SVyZly9kl/WnukbNgWAj5NO8OQjX+t5wV+FXf8
wWMTOVVRgo0XPASz9tvRkP/cn2eNAn2VJISpOld19cSjwSVQtEkStJZO4uA17eKq
1UQ9gWqea9ocIAjRoNuAmOKf9FtM2WrOYWdvuec4+PYXfvAPoWHRM4Bs8wUqtTHR
fU3G6Dc34H8nQBqnCOQAa6OoihBjgvgh7heOoPE8VeQddKF80UUTkRI8CtU3bB3d
yqfgB7LW9QOjEh+uFquzmyiLrWkoKmrNYLaawdLRNDeCteNxkfYIcY5T9RYg4gQw
+0+iv+91V9V/W6U5sdUoQ0sq5fy56Txz72qSJ6tWTAMXeG/LqfGwrdSmLGXxkax3
7Zbke5R9eIhNmzW17LIhj6zVWNokSLVttnRowbXKvjzKWUAaVEEy3/KBCahEzWVe
quU9KqyhguNNzvb3R4PsQA5OFw7Wq6W10ODrTqs01NNXG4pf7/WnJZAro3fc1ami
IwrNgfRHNXSfQq++6z0UCKWT5OidLHzhVSe1V6BOa7xaoxmGwKeyf8KWwAhSnkOo
YH/y7RvAtSS+M3bs77hMOJGASptS+9C0tn888VcsCioJoNvAZ6jU0cs+kpWGglNj
XbM+N/B1yncwKRXwiHmp3XQz/2BHSVPp7ZpOs1HQJpqHFBW8AzgrfyuMz+Cfou9K
QdJCRRJ0wB9uIuR7pIDdK1AkWqa2A/LrKyQBycERyJRK2K2oUW69t2QS9m6lNAzR
KOvjxNPBhB2wQdVOH0Uiu8AsSCk6yif2ajJ+P+m/4OVcTQj3bvZzdKRhl94YcxyJ
6v1qecLwW7jQtVDGt66rwMRzAe/iIUVWTyhOGqIGpV9TQHCdIf7UifQJAmCwo3vX
DqPDTPYtLX/84YXw9VzN0cgC07rDxyix3f1uVtZnQNbm95kiqVVkLIfh4C/kyn+4
wL2wci4rPbYN4Vr17nOGrpSPXH/JWHZdo5PwtS2+VK7436jKL1AnJc3r4Ug4hEP/
VqmM4kIm53b66oPHEn26qcdFtvWrPdZaRMA4P5203UVHS9iHjNirAczFXm3QPAWY
PTQjETuyYVdHwLzcONuouRlCdtPRSZNLLnXD7nbncy986qrq5vzzhTWJkJKAJC6x
BpvUJ9xk1k0fNOX6L9EAgJJb9vMMJDrJC4JDrQ5GFaX6zyVLJYBFeA7ORfQchmN/
QP6T5880tcksgKQgJnJ4wB5btTF1jgxG2D4IC6/4wcjS1RENxprAzAy3Aog3SgGh
21yaxRQ5nypNU0KFCtE4r0VfSBIFp44JHjU+XH01DxGmA3EeP+oYrNzS4bhYp4eg
QrKD93oALqFgvulGCQR3BNP4p8BC+QL0pO75JwCAXcAGe+FEF4x9WxtvHZ3gx3Ug
GMydxKhefl5x3nofj3ZYM0PFy5jcNUKLHxgq3YMsKPE+LOD9OG7qPRNf4AKy9w0t
28O7nafwbNr6M27Ss5a557KUqxlju0I/1TAFHkJAQaE/HG/Gv15e1gx/JzXd7XHJ
xdPQvOlLLNimQuc3L/5ISmloOgm4BANQ1vsc5X8WdZCl8vQexSSMuRneHRA74bth
G9PAsEWqRfkfebh+7nNFsogt926XYZQzqZQzJ5FErBaDnoC1gKfCyX1kOyCmLyg5
Gi0TwGXOXAhnuyqnA3aMeU91yYNR+UUQYsCV9Aq2KFw5McnDieZB8nmZpkqv4t/D
Mr2fWbKn4KEk/rSmpDCjxAOkonIAyAOULBFTVV1SPZY55fIjvMx+luH0LmWda6TA
joO7Yrwk/Yq6UH+8btaZGAA2oGtXIwXtQjeXgwyvAaXMAzhHpK6TaKWvz9O22Hup
kQjcf3O93ixL3L/mZKlbsb+WYWq6AT31LDlgeuw9Wv+rBvkBB1xOM33zquAQYK0E
z1SHOnA1u+1nla5jZFY0GEL/LT0e+zd1W0ONH4kmwzQi+XtjHc++xAcpoYD44m5F
FmhLHn+HdwxE/fF6IhYfyoGbF3mypRqT6MHit4Ua73ox7mpdOJy6A6no4YMaHcMA
xkvprBbPwqOF7NcRgm6/iVoMz6UkFq8d7qsemhSLA9SUFrs/1yGchBPzYxuV0Pjp
RzJ0ipVmJIDi5EEbNDtyInznPzGxY/kxKBJX6mZPB+gVs6jASME4REh8eOy77ik2
tL2FcdKCE6TxD9RaPOJLEQlFoSV38QHNXbEeFLIQO9ITvimw6qwjPO5GaXYNuYj7
Kfe4gMZPHQaKWwj0AHuYaHsf3k41DkoUvyctFB7LjfpHyMSXZ+L+twB/lbsdcPcE
eG+dPWzvbBFXGydY+4W9imR0gkks2CtRScdZXtdUl9LLwBSKb6Ub98N090EROpeL
PdI0TZaw04nEwj5pq+BYZKm/1REEtveb1VcijvhEduRN16CpbcD2kI+QYD2dIi5K
auMU7+phYV8iJ4X28GChvSxwAhpC7c9TmIc+BZPl1Y+JWboKDqQjI8mwvamZvYPH
rr/yuRgiclAR2j1xsw6KQlcZFR8h51q6hrObIylGyoI3msYNXnjlDnccOMHf/RH6
reWt50sP6PGys8Ca9qud5fFA8tL4qklnFAYVD3rL/rCLebLcHfcFEIyatyHcsteL
p9Ufmcs/+JJl1VfB6tid7giZ3k1IFYdEiSOCsxSPqXnQKbKTOY/AAQr5PBwrAY/D
`pragma protect end_protected
