// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
smD1/z4FhfLgi80HOvQC/yFbLCCf4kc3N0y3IAlTMFn3daEjeQJMc/clwrbAgzMWMta0GL2c1pwU
Ixx5/yPA13HTi2QhYMh7p/8qtGzxAeDhanWiBw9JcpzxeQNTo+Rt2thQSb66Qy5vyP+GdIkU/5Yf
byJjI4+khloUhBybdQtSlrEj+DOrYsjkDJIoK78VLwxW+Qpbm1m30PeVE7Hkw5iOeKzz1Zs4mreP
Q0xq6zD8iSwQwEK2+KBb5fxWsS50E1PWOgTWEq3SnIagpQ2cfyCpnp4YaQ731aP8SE5ufzgQsTLQ
ouHh0KHUUBHob5TpWR3lhMX48GM0Fvolc+XpdA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5760)
xC7youErk9EyXtBYBFSgVFuF96LsJY6JdVtMFlZcqSpSPt2yLXom4OxFdEKWIxBI72u9SO3uCVNy
xYKZa+DEdf9/qMAIcJRODOzNP6BcoNRGePfOqSs7VIrNg3Df0FC1aI4I1/Qa69F5EhmT6kMYFOlT
NC7m49KCuGXlihVjYJvD6FpchTcP6lU8uWRjyr7tXd9UZhXYLE6ZWd7Hh2ShgHkL0Pdv7W+wV2pV
PqYxgpxPgUgah8Ird7IRRsg+4pGw+Aidt1UhS1wt823OXKE+EzRGjrncJYGbJUpTgEkay5VPrZAN
1HrLTO2JytJCT45woMT7Ss5/8oCU9KDti90Wu6SBXywaTS2xWtEp4s28kpeVGDHh2vR0vhg2Qmi5
qolCav4d8svJ4A/cJUI6ex9ZK34qygYwql6BRXk6SgqLA6BaoqGdV0AKXIiog8tfIONWjSLoyNtI
JL44B95p+wTwI3OlkmirHwciLGKaytMBeYquOhbGUy7ivGP5VopSRUEEYO5f5Nye9Vrxn0/536Nd
No3NdtOYJSpjqzmVf21jGhU6BzaQ79oqpN+3JkCV556LSgqOC7RalzLhvCq4vFdTrHSNwDUJUFsJ
OXhDiTYydz2zJJdkGIz1TiPA5rhpiHpe2Za3guLOOoxyf526DDQy7c30977/+TCi5X77sMwqvXsD
mxmziNEgvPfY4Jpyn1ryZLOfARicIxZddLD6WaWgXYk9OTkUHA4OQLQQB6Qumvlg6R6I1E3W+wjf
IGdoIjYNDF//JlCeyh74gwwfIjXWuWPlLW49WFH0n5AbDuiI7ecKI971ECs7NTwFuAGKuiuCrKJ2
jGzgXmEVkBs57C7WeAYpLe6+D4P0EsBfauax3hnTzOoad3nah1ckSH1WRWm/gXH0F3+A8qM0q9iX
Wk1W91Lem9uA2H3BLA353rWPaalvlaoFoG+S3BttbE2t97SzieYBQb+8RCBo9BimmSXQ385NOaDB
VAbjyAurXTWwP1LynQpZ8vs1A9/lYBQU91q4heN5xPGyJ52i5IxBQK/cyhOKiO+WHJpc7GZxD+MP
sUAKMfXxDQAKkYjVxPkGM8gOtjIk9HdKsYfSSPtuNRDYx7d8vvKpku3zlfRZ66O7JVVz93YX6a2p
KFOBrXitvXyT9Dv+dEN2fgiaHF9EQiRbC7mQCXot4iLbR6+qD2hkqe5fV7Gg9Z5Nzcem+UBajaeK
aK7nygMsWBY9BijrNav6ppKf7ma6Y2vytP+iXFLWgJ/aF8mXZNAZxGcUaGA071PQZQrRQs5RrrjV
g4o/K17biGkkCxG4r8grTlG7gcYEbYIVkR8T0JRZbrlD1bAOLhuo4rAg5pK0zKKUeEb6Dnr9Mwc4
6XABpSn6fPbY5eBkhbW6CmRO0pqRWwAr7N7OR1HeoYxYfo+Sl0SU6MmWJryFLg9e7SJfC4kz9a1M
qQKW0xP8MEIdvUbm+fEwvc49YRit6ioXA1DUXozpWjh02NYyxuUlUs41GGJmNafnFCHrEnhvnhym
AALXNNxYrqMviGvg7q0s3UIRbNjhCnYzTaskpu+GDtJ9IyrDcXkmxLQ647r7US8qcDmnOdUbvHFb
9J976ZNjQh6cpEUqj1Wgbko9pignwigYTJDuV2mhzznl1Yy7MWAiKqRPvIywRi2o/1VKrgpXR2Yn
/AOtoVYrvVQjpi0gYmM5RVg/7dYhgAqxrxR5XQVpIs0+9uQsbb7nP7t6bFa8hxpshHEKSVS/GPNu
3CHxTNTJSTzwZmf0lG5ZUgTKDIK/qC/PUDqu+MgmEtTDOdQLFH0E2S4DwYlACGAIqTq5PyDf6nSG
4gIlH8o7TMp917D6QhYcrgD36hHGvxByeuD35GbPMR6ye/TLR/urc3eXT62NjY0YxuSs6kYPD5wk
/RVnWLCccORSWsIT9mrGQS2DZ8o/G9VFOajSA4BZxt7a+DKH8cXh1qrI1Z1iZAakv45JyUJFSU0e
SVvyCqHLSZhf/uvRv8pZQ8aKVE9xT+HGHO15/Vv9aBJsON/yP4GzXK0DLdueE1Q8kDnETG0yLqA4
b+Ct6xIdTdYSJTuU9si+my/SxfcZv/AWMk6eF6e0h4WNL4xYOePzUvPlljYeR42ZHzBb3GSVpuk7
X741lnDsEx0RfuyXZF9ok5n+PT27cUoE2hFr6AoeV+WB6zrM3wb6HP5CVRAlwMA8/td0EtJLfTvj
h5fogRPpidSJrSbYgzg5gHS8adcB+VksdSUA2O2eBOa3keMVF/KU+zBaKTOoCyuhStyZJjfgDN2Y
mAx888LknUPXyqu/NqWpp8dd+RQlktbwsqZ2wk2Wjn5Gm4gKlnA0K1vys90yNupmNEXPJmYyHPze
QCz2HGQKh2nL0KiGkZ+KgpkNUQz4lXcG57p5UUP1o1mjXpTa9FRUTgmSS/22RUpdzHN0BwF8pJSy
2XitZXZb9lNM9P8xhtXTHO/Y0ZpFWMg3eTZJQh2iVTW1Aa79jrgGt/YPM71NCZM6+zjaS9inerSw
b2Z8PJeNLYjo8YCNf2d+ldpPwg2y6KqiPrZCvIIGBrbuidfU1CLg4F7XInimkBfRVqouiRm9/L2J
5Co/XWpau225juxmvif2jsnMvuG2zIvZmmOwSJXMWdDjwz/eBDIsERsiINB5APkZ22l3zabqY/2/
zJmGjFetRjUkfKvY4eP7ajPKunofiy80Es6ftNBd8DuN/NBNTz9hzfFKJwCBgkT8Fgqj87CTu97n
kIWTTrETfhMZcNBx5sEERvR1twh80P8eKwVyal9b32GbXUuPASrQWYAJQv9tY75DzGVMbuZ8oa0P
8y3QvkCES1r5v8NKZkSfpYNoc2MHzVk14nksUnPvgHvW+ENlyM/KqHZKoUcJ0gdAuq1Qu6agtziO
5xLbr8uhYW91akOT4UsS4mow9X6oJEPiVfndgPEXjmrYW5Poq8A5OtjIXcPDXtTVGFKVLGyV7LMm
pDfVbg2wY/Dm7LYLgy/SQyoAG1Ziie6+vXZimLmZr08WXSGnmkW7aFifxtIqMSWNsoJi42Z+5xcv
iW8m+0TwbmLNyrBlDuEf+bXpT/VtIUFRdHoMVNp5C57hYMsywpC6It0mEy6yhOO7/nETJthJ3Gwx
AIGMGHbIyHBv2GN0NXsWFbZ1FMziF9zqM/1pZjLTsnqXCJOfoM3y5fWs/4/4j05yBXlvsda4a3Jv
pS+WEYnssmiwGACyLrqJT4FyaVmXrQAksTNT9skeEilG8WeFi7SMWPCfFdBxCoIcMGtNdXZff1ls
twlYbYHEBIHnaXdc0+02BuCqeJrdIURMSAywGnU7euLLOvmGn7cLN+4JXiX0fDTyQdUnfh1aGvpC
frd2qxUPoSjPI5dvahZHJLRurs3I8PBkKUlkuP6VG+XO6ZWZ5loBgJ1D9fCK54cGEPN5i9JSGCNt
4ik4RBkGKPlOMpblctvFT00Ml4B1fHIN7m++GJ9roZQE2JJyXnGF/gurro+2S7FscH9jwCW6ZLSo
Qk5DBUZC7a8ULZF+KdgP9GPuwfVZdv+zRd3MV0jKdwdKzvgjv/Ubn94E45bVMaRYlh1Q0Vi11IOY
1fWM8hhaVCIrDm9DTW5Nl9kRFZO1kXyvZtXXas0egepKGjJnYQby3/PqHpqJGy64DbXPRPmzilpa
ObYe3LgD8JWklQIITOjDXRieqJeFyk0mqYFT7yCbYcDbOJt0ZaFMjAsxz/urbttJhIpmI0SNEg1P
4WYKsjAKJAj4iYknvoEuy8os644dBKakNgpsKfwsk3YegNWQEfCliTxZHtzEA6VcIqTX0KH4B9dr
hNgj8i+cRhSBC1VZ8rQ0S7rcJ/HRG/3AFvcYNI3+7Esi662GL87kTq4Hhpzs41l4ZaJUQBEBlmRM
iJ1EqfiG3URrLZuuE+kZ27i8kD/aCFrMLdnD5uRP5718a7C6UVZQId9KH9jW8N1acCDc6FDqG+5n
7J3hBc04z5TRIhna0MZI4sNYBEMm7CEDmMf4/8U617HSnfXejyHu/CNVp2ryw6tROBck4GxDhk5n
f0enpXZCDTUKBe1jhb2/3e5+IvQAqSEr7R8I2zeY+LrS42E9UIVB0hqazwvSvphOgj+mcghMA5Fq
yJ7KtWU3KKBIi+4nGywWfoGw0zCsdF4B+1bko/COy6wZIgiU44O6qhhtPl6LUDgfSUxdYVCoNbNj
FYqBd54k7g9FT+P/vq90PgGSBr54S6R0ueWyFNbgzRZWnAbRBeyt2VxkUkAgkrIUEL0QcJZUop8y
4/72wXR1/UoQFHMqTc9jnBb7xPCObBQoJmFbHhYJyEGz7XrD02j7hjSpyz6Mq0p7RHt8+aDSVw1X
Ha1iYOySezFVR/HNYCC8Nr+n6RTiXGGWt1Oi2ZVOQFEueYg7AjVS0BN/dDiyKoMrUd/exN1QDbRy
zq8+lgV03UtrsqmlzhNbZ5hVa2B7tpge1GWsl+/xmNJJ+D25JqM2i+CstfwaU4iXibgJrjFavDCe
2ELs0w8xJjJ8yriGMahHBAnNExMikCksQ9k0AqCAXH2uVJmTnmMYw/8LkRyodA+GxmrkwP65z5iV
eOVHYIrOVp+ud5C3gAFoyK6uAUtY0zMu3CgVhYqmCqcQIeHJ+3AyNka/3ZwXH2SAZG1DthtG5VH+
btdVfia18n40qSom8ZBO2VqLJjbqzWrQ9BeQEKhCa5yA3PI7aCcUGDylBaSRKApX0OwxxRexs4eT
CZBQQfzcqze2t7rvp0iabcc6A++N16QfLxv0lUwl8EH8ZDtuux2VCrxunDKsoUcrbxTrMKFnFyeY
6CVdG8n4i6uZgY70/6GGEJJmPugHG+cpzno+jhXphnL3Eux2XhpwtoajRlHzF/U5hT2N1YrlkK02
vRbwFzum3ccPJ3Vmyf1nNqRZSPvqRljVIPy2OPLfHMgvmQ2US9MqrkN5qWHH/Xic+KKQQkWrGhYh
ab4iPXPEy6f5vqMNoT+mWFmSKEmE5UMtquhC+Kpj8msJfapD7MhUR4kHJrfTTg5N/XQnWDOmQlt0
7VLAYxFWgB3mKs18SRXDUy4r6xadNP5tnY44xMaTh/gdi0BQ8Li2RnO/hGzAolvJpQPcpqqOnY5l
Ji2ciiCg53aHqQIMLooQZkdgOrXAaCUIbKD5BM8NtkE3pI5ILhFSFRFfeR/fTzy7nbEW6+kixNGq
stRT5qZMk/HABFU84zN/rfGJDmlpBFga4ua8Gp0EFE84CEqkQ08ZBo9OlyG/qwlfsP7yo55ASCuy
dk1VFZlRsrrbGe4YyV05o1jM0bR7XVCXhMmSGWtDJScsfIzzysLBFJ/t3lncuvbppNMX+9gjz3va
S/fEpldG52Ph/7L48YGHgki0+Axpxo/u+7OQcnpJYEympvGXSTUTKQWEVvfAwiSTM3ftQ9uiUWeT
jQRtSaIeIjGw/N9BgRhCKmnSE9EFEuKXKIS8Ga2tIknIyEsbnuP+QvrN8OJDlUwUyMYvLmdyPEDT
fmnl+NLyJaDSCf2SvsPT9hJrU24fWGqOkagFddvxHphHQqZbVj2SHsrx8tBsVR4L6V0Rmecz46dt
/LiknX1QHZNMQZ0zkrh0adP3FH7aiZqreUpU0x+fTrLDQ4JI55aXlKGTNQLGd0WaBHUdpR9kahnr
NiDqq0Wv4uiQl9F7ztkn0aD6N1i7hbXSbjgJ+JOXMqY4T1O3rvj8CTEHPxDId6IAV/1El6LcHJ30
KoofAGnqU4EiFUxnRWkbOPIGEtPts7O3UuuyPsdoEco32zzX5t45iMVrGgiUV/xc2YhG3p85Ln7b
jeSJNZY12Rfz6LlnF1bQktOWCdO6r3tM8K+BXppaTfqcKn2VlZE3RdHCSCMDhVHgdY02W/vYKbmN
/pVqaZ90M8peoeGMjNrqynEWA7ZhYZGWFMvY3TeCzcbk1cY8LDeSd+y3oZ0MhfvzutSM2T31u2Qu
Mb0iHbUdQdsNR83DNx+Nk1huA9UIQHib1HfsvNchw3hDHbj2adnCx5xXVD5+o0GbriQAxryXAYA4
JQPL99ygDTckcDFIdKRIPH4TkP6q+1HQu2RKepeplN6I/UloVPLOE7AG018KV+UqYekr5XOpBSRj
xrr4BvK+9MO5RGO5paBmi6PYui0xRXlpmIAtNQbAQ7OsiRVgFJvsBn+4IlAdIo2ipTWBWlsvuuPn
zPOyQ7hYpMVaocpkKZLW01K8lyVF9j2sRl4CZ5YghFCZQ2eoDZR12eeQoWJ+mtOkd+b6Dzq9Cckk
10ageKmJ/40FBBO50W4506aiJi0fm4LER81dKIUB4q8JtRNDWD9yl9fmXDK7qtwgcDfPpYp/WyAi
siO/fPhopmTS8juMqonXCpS47Wf0l/ioO8nwanuQ8A2BGkj0Kxt4s/bpyrLpJlum3i+TNOs1LPOh
+tlivucfR1xCMphIOIFlJwv+wa2/RjoW1VkEj05+Ch54GU8bGgdf8XIy1sEv677PUwwo4Gyjyf+2
mkTUYoqO8DzZSz/yetBq0uSGQQxE0hcvKTyPXLCqOsYbyh+SXDUzvrQvIMqUHK3b9qZHc2F/ruNN
XwQtl86To5oKOJ5MqIEX3ftS8eJwVWd6cadBsSUsZXNIE9zRfak8hnJ2O6Cck8/SXtevdjminX8+
QA+75Pt4wiUGq2+ie7xLupgkLdkFze4DbcPFw1oqJgeo40sNYWy4hCsvBhhvtZh7swbc0AFhAOMv
6lvGuNmEoFgzNpIKreQfJQfloSK4zSVwQPUebj5LmaL4fBIypmTColnhvusOBI6Ot6Ce62uPTj16
YLbclS2wmHoRAmw2j0Z9pzkVcXnLENbeJNwPfMu4VHcD9KshLisfCU14RBY2QI1Nohzwq5yeBJ4T
cpynR8/pkjqQsIWzl04qfpPFYwkoujfy57gNrAt/5KMka/wx6u/6pqugAwk4UtO40920/+fhNY1L
f1Asedxd56Ty1d8xrKuZymjUwY1gUFjBmsivKrCntwAeGQWtuC/JQlHll9paA0nA6Ko2WBZFpjzz
qT16aRIBYzmYFhq2YncKRLLgK/hV7XBcEh2SVEULXzAnmCYVRiqePSZeEp8ooJ/uepuviNVaTUwV
o9AkRtgQWODtf0KD3kRh2zdDWd/GmzROuG2o+hycvEB5RItgpgeaaCOcKdjHmwVwoM1aFyt2rmwz
GVvQxgQ59tBZZE3dfD66CNoTAXMSlqOmJDguvPfeZGvZi14KYdM20wEeob65D4kZE7Kf57BN4D8W
SF7jNirMJLnERnf1NiGQGXdeJajGc8PKTYd4pZSy5PGAFJ+4sTIqRTZSZ9TXBYxXejBhmr2MYQOg
jzl66aZ5c4T5qLu2jzQtgn9Zq8X6vtxwzv01WZbaGMAuUTJqudpR+jCwHsYzIc4yZ32jNoTIqXg3
WY4T1jaejCApx1S/+lD3RdxKv5niZnQygH6l7lELfzAK6jW1UywT55YSMU9aL+X0wlyAKiz0s9Y/
cnTUWFWYLCAyBmZVcGx2JRfCmny63VMXqxq9F24geg2BCEQgesJ1v2uuvze2rWmBMjG7Z2oyK9BO
ADjxIwGqS8piI09Ci5SBJ/0FAzgeLx2CHQmKkYFgTYGpDjf/Kw/snzkECiDMeOmooj6IPiwQ2PVW
wggHJ/VVumHhXLvv2+d/kOuRAgk//r2WGO4FCn5ly/vJpKd/0OBdcwhf9htv79CXcIpf3d/2uFlA
ihW4
`pragma protect end_protected
