-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
N1zX7uj936VQwm/m1lQSJSri3DxCxWKun9m1KPK7dNg+eHRYv/mlP5Ye7HATGcAtYlLNt1i/ag4O
CRLPe/lCtMxURxXhSO2x/eOBaFYOdUYqwebfQHGKhd+3hqj0oxE/Od+ZkwphawD6Hi9Remi6n0CG
kfvTdNt+ZifQE/pdvbKJiFr+v/DC7GU43W1nfsugqDElVJWXWKIUQW/lm3MCwEDhI3Zu3mbOss6Z
hd5kIvFu3hs8wtollEFAKyiM7fYjTTVu4JYD7nW6ELsQBU0ztrU/qdIH7fa5sfC1oqI3yXJTxhXi
V5HKij0QB5QpliYNiOZFcRLAG2gDP9tT42aPUQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2640)
`protect data_block
rym5l1TLJOYdgBADwhApnEi8FtBLrlvfHiAZVt9xxTPDHDSs/YvVK5cFvDOUkyAHqs+78ebvc8OS
/lLRPapqNb1LNI4UfLIzvRul9CjSM3Kd1a6HWA/KK43ORZd4FhmeojHx/1gGFA9MnkRLSgPu1MIX
Lwbv0KPvSAwKmMSK57bvx+xeVM7JDjNhIS1HySWw9cVjWJHxixnrRJWq0iqmbCTHYzRQ6sMDD5BQ
D8PIKCJWnL/hArT6ugaFKaSIMxSVq03PucQaJmIypEG10vAFeiWC81PpLK+bomejikoXsoo5n7k4
cSG6JsAv9BznFH03ecfPbj/Yi/u0gxebvbgWH+GqmcQvRZDKctZM/p2z4Ie4OBsFEzrA7Sa6Tbtu
99OxvM9TlD4a5RoOWO2D2mjBfr2gr6nxj9aokZwUtjjLswkuP3La3VjIBPynrHlxrEQpCEBVHrUx
wWAKb4RG3ZoA6wX3jIFLkMQhub9G9f5+hyESuBN2Z+seB4TKvFAd3IY47ldEKI/U+BufaqF63iCv
W3OLUQGXaIY4GVCA/a0nKukkYPN81Bd0Hif3qvrl12S2cORgd0a8hszIqGliY7Mqm4avPiC/kxR+
aRMtl9P0wjLzp/nlq4/yK7WTodlIVwOo4MVjk8DfCIetCwC+Ld0TttuJo/W/AalntLYRYu7mAhjh
dovANmmQaGUPVdXe+UnbgQg0lQ0O8IsRVfk/iE3z6fU+uUXBXx4C4AMKz/zYueZmkWPlZnV1Qt7N
N4p0lGYKyafI512ibzfkuQGR9f9LyBONa522drJxkoapYOXZhZGk3EocC9QkL7S8wr3JLlMDn29m
X99ifapbufIMsL5oZ9NA+F5iujoIy4ztbnhX7IA9fELciSbkeVpYt/ZSM/U7mE8oS8X17rIxcpiK
cIaKJUm1haKyoy8p+KJLGZzQcKU7pOKlYPJ/7gJLOteYR5JPk0DGGeBcDRgFKZE1bZFk1DdSeLfP
yjrGkjYj1LJHYkdnwVwAHxj9R0HvoJdO7aT4mUkE/ceOjG1ZOtPlvVccCexJU8TK4uDfIBzjdcH+
pvdMFKHttGPz8hBXP4q38ES1al+39i2r6aZBIsaHCnHz1HBitDi5P8qJbnV5McMLAGpQpZqdZ1y0
XlstOlVVoQamNB118FCHpJ83/YDCNlJs53R4UX81Q5iDky+w/y1YJJYpXpFfjAkJ8FtXBCL3Jwco
OSEi1onlqHXzexfhlxsCOhdn3Lbg/fXDQUftcG+Cng1x+viMONrrA1E6xLiFjofC8vGZnBa6XzJo
RliRkaLQb3wl3nlmGhNige0U69ibCVIs7yXoPtcucfOrhFrd9uAoclQ4ECvwjbZogmObyZjSiFcc
KHni+G2+O3oZoA606/aZSOHEwPtLah+OXFXWyFAdu5KMP0iImFd3gRnwN5y3DwZz6X10/kT9zEfL
SDtVgt/zZE5A6fYw+zh++1prq3hl1XSPUvA8eiyy3Eom3cVoP/pi+VjI0uRF+UdFab72ePBPBJvB
cG+SVoFk9sk3NuEP4curKt4I9rPxJn8AdfPya9FrFsG01FmU6BCSno46FUKFzxWLwvGn0euonuyf
eLZciV8GZQGe/7j5rm72EyX+BSjHeXwTVDJMApa1TvPyXHX270xHk0lfbeUrwCVBEGko8noG9+pu
Yr2Y2Et0NXc9ojximGWhmGSBKq7zJlEHe4QwCWO0Nd6+IQSfBqIld52lxQvUpvWwJNexCintIAw1
Ca8n1RGDDFqOogSKmRYSeNR+l5SQ9KlAbsZH9rU45Z6L3fNpOdBxxpbGf8oYC+Nb1jW5oxBrSHpS
xCIvnYomrvqUMMc6tjy9H6X8LCJD7NlsgyMvBPwpEbmim3hdX1nHd09fjcfyzoffSdU927z/J6IP
OMEF4XcPs0/2vakiL+b7mNAnWJnPs/6JorXxuVUDBHfB2TmTxwhNhFiL6Dpl0yOH863pIgoafuLY
d4vMe3qeOt8qz9JkSLw4LgYc/j9x3DPy95ge/IuFIOGBBwjuXXio6svAQb+xBV7dx7tzjaKlsZc+
qquvyOJQehNY6Z59AljVFWXO237salCEUXpe8ofFRs9ldMk3h6b39+AHJRXHzeLIu/7B8rNZxp9H
K+3bS7lxIrroMBNek9LC4mMwdndTBw8Ry8GLNp+qL/mSnpNnVJzGyfP1ez/JQUFOD90cWHRufpE2
xqNnOSwzbccfVbeDnF3MghcESESt+1MsEuk/mF/fjMpmwKvFLsayLrnC4UpBrpjc0r8RFqBhzwTP
ybs3zhIdaTjKx5DIkSfF6pe2YFJ/3lnT34GjN96tWyPF8hbYnEeK7O3R+aGN/GlwsZJY/MGFoUzE
I2INB0dMFitsA2f0jnkwystMcTRFGhdnSSMd+bX5yOOULib0vB2S1d5PI70y59t1O75eg95jzyFd
nPlP0TGrhuQlk8KS1pxWtocSAg6FMqoo2hDrSC7YJgMpAg1YsRpcoj8RX6Cd7gChNpelkXO4/UJF
gYaxky8y+hTu71IWVckG2nqMhzjetR3BF4d0QEko2dFtPp9JglCAvX/DuK+Fg6tGaCvKLQhwrdQP
DCWYHHA8XrZ3VnloZrhM9eMVz1tgayz2jmJrtBMNLmS3cTkGy5vz6qdes+zLps/bUsVB6i4MAU/e
/IHi9ks63Jm3gQyJoHdUNWc1TxbSbMrBetaOGKQZHJ1OS673FoSHfu+bUXYYE/JA+UY5XGL3trrV
nvDSqWoSnJW1XsM4yYRc8uQly5KYUf1Ru3lVE3n2csqCyPLGtlAcSXZoI+UaS3b5Q8kwzNzaC6gW
DUvHYdDhibup2QBXs4Mp9u4XF2hOvePk6T70D7fV9cOfZTzxsPh8Tdunlo4CcjlnixgQkqb02sQK
b0m+w6GvEezMuTIIE6M66y6GksnGnWkGgT3++f04CS/qx1f91gRfoU0ZTBSsV9RdyDXD+27lGESV
qFPoQn2kZPDiLHK7XnLe3f0xf7fKmIYw386EF1JkxEuYtnaEpl6CZ2C+4SLBHKXQc+qmFyFIhtUi
iCqFSc2SHGJVSVetJaXnfhl/YkZJ3OSZhlCiM22Ag9uvAZW4CF9yqna+KsJ1brPz+zEwT8ZX9cpV
M3iFd3aPCxcRGcUtX6Pmq952VlYtJurgIyEwQ8aCxd/RnQ1DhOEeWaOiAAASZr1YQltBe8K+lo/S
Z17zypSY6w2pUF0Dg+98lNS8jhYMb4FeFWXvFWJmZALH11F98gxgpzgGcaT9iu6dnalyrjtzKflR
M9I6qk6ZvvRAVB+6GPuiiDoJs6WIjYXNd/9EfWlLrakMFl5kfGxfufWLzkoXkKUC6dfKYrrB/B74
goF1K2Q8knsM9pfpj04tG/xXJJ4RbHTWm1VBiBoHofdrKD87MhA+/DpzLc0nKxt3fUGoJG8PJFIu
16RCB9ICfwdcuUcugP7XQzMouDo2Nh01skSNnr9DIknRR9SML2c1aRHvRjjpvzgRHK5uHVkQ1tBD
z0nUIWSnh4nIr1zCcmQ+Co6e
`protect end_protected
