`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i0ZpP/xXmpJasyu2W953RWP3LFwrKuzZrzvaKLeoGnX2OV+UgxqZuJMCMrv0wRtb
aL7DOrwh+o9JYcb5gnHR0idA4JdzKDHTM9ln0lFgvtF4jxpnU/KmQTXDUXAj12G1
IJ+JvLBZwX7hm2t7NCpc9Xbz4kDL8WJcMrQe1hTW2pI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19936)
gzfYclH9J8hW6vzpj1bQc3Prr7FHBtVaZ0uZjbMVYLQjV/UqDwgTu5a4kW4C8a76
g6xJ2wCWJFxjDKbAw0NUZOyI8cgJtCXZzBFbePO3BG5B8VcHZykqMu/WcTOcg+dj
yU5SRovbe4RH0oYlQI8yXA/PLVJo9QJYh4Ur6ALmtqiv5tuJku/aLGRHkaufMgN3
hprIN+6oL/Fc/MngHq96VldZp5whfL/hzyVcjwpDYaN8gQ9rObIylS4mZZdmhgkk
TRxfbv+cYGMzkOVlziv0bd/SAgULUnZa4WuhPRprId5AmfXuYTcue2fPW89jOq45
A2uO+D8VpPDWlXv6pt2D9iJxUgl3WQKdkmron2YOFq2nq77dy76AWvllZ9Ne+SDf
G2+Z71S8/iOqrXu2CB4sKaXXbvwH37PISt5kugLB+2GlwRUpIQ9fCLNEGe2FJzRQ
IsWZbIpGzaSGLhSE9KOiW3+hc71/UKT7t/dUotFeYB/a7vhrZZKwiQV7u/qSJpDM
/Nz6xvfkmTo9mvCdAlrysqwvz0eN05DgHvKiihxun84NtxFQWJEJt2kn9kbg5au2
KALtK9Or1kYfwVLpL6xNkf6WPTD6cCeXkwh7d6i6/ml87VhJytnSsBcxKVn6QAAH
3SYXkkHm8qm8MroGBupcKfWunqM+vnADr5JYWiJKaOEtqxOzgtIU4omLMLi0X6nk
gCDro4dVgA4bllgq2rC58+NRWv6oZM9r0c+9PAXrU/c68f3fka77AfK83SvQunma
RgRvKXM4hDmp3p+zbxbY0RZMNZjbLOI5DMznZVNcaUFXfVZeUeiIt4V0irnTkmv0
hEtGo/g5mbVrOfWM5Mdk/tE1SWlZf24T2IK6RM/ujOfxCmLO0rZU3oVb8EcuqHQQ
yhXCuB2U9Rods7+uHjMWX1+MfEQfpp00IqajmfdGZ1avkD1a0wYkOALOhPRmOYHe
tHmIRgXI2soS2RWhpGyKowDSLKPnFWumojcR44omQ/sXYsWKvsQZh0Lyc8sHwBFY
TW3jfo+FEyZ03QLjzUbEhnpT6Qres3Zi6BRAoIFwayab5C9T35RCL21BWunb+7iJ
e5+tQaNmQLcexlZouwcQrAh/gMQ6HTxpvwC1unlJbDBfxJx4BOye6UTJvRYxdtWw
SOUaTxPxeyE8Rg0Wpxk1J6c5RE5UdEwfkuRMunFbMMuQlTrwX5syxIQy/J4ICga5
BFTfSXq/qPRLEllPEhvrPHlA84pMdYgf5UVMEbBYPh4TxEYvE7xxFmV1Wxafb2ce
okuMtj113vUduKm75PAm3FaZPrnzl8WAfnBwhGc/Hy1E60Gh3qFEZC95tFciLCoY
UbeE7xU3F1WQO031lXBKTzDIYpWsB2Detw6RBUcbz2Gt6yHMx2lHy6GjcRWbvePh
NS9xEzBiDedxJ9atAuMZfO2YLKxI5camKiN1bkllhJN7Rwt6w9BSOb/dI+DFKb3b
eGBR8fDqAzQJH1QKff1JKTsORd7YYdnGlzdUtV39fypFIV3HK4G7lkBmr1YA1O/O
v4e4a1JKnXRhdn2DazuNPVbaxFZrFly9isOx0U1SXhGQA2w8zd4J72tgBJBlvToN
i4zhx1Aor5htEzfu/FpTiAkVLN8EgF34HEFJKA7VpmLUrRai8if/q1zjHOU0Cfw5
BL95yBwYdH1vc8o8XywgFix5x8J1p+f8anAP3mE7uMV+M/qYiZw547PL7LiFaBur
T+9uZyEUN8Jl5WbEi2/WI+XuSBFTbUcI9FtGsjuwBYZc9q152r/agEAFI5d8+4cE
7lQgdzvWNEl6P0XOfWy3tEqdP3+lmFaXYdSDV1rRb1LKup18wqSzTOatd5aOPknf
GAonO1tLmBH+ewX6ChwGIw8QwdWfZ7laf+c6lnaKgNbyg2NgtXBOSlr15FcbrV+B
wRIEfnTrURWOLAMW/Rmcso4Xe8HKyS33xjzLN8zILPkQ7mad6aZdidaNLcvevOZZ
lEQ8AxGHT469ilUWJWMH6PO/g3MwskaIgCXIUnRjbbsidqPKKF/r7CMkOzwDYG9F
2sRlwXVaeWM/2ojQ+qMPExJVCTkXad5hl0JDvzZ36bTUgUPiKs4JXDQLkhnUYJ03
xLu730U+dZxCjkDtCEWU/fyGi3ZzsN14xn0UGQCniLQhZc7d5RbOJ74nBvzg+pqU
Tw5SzL2tqekEneAvxVcS3tGUKR90gbjNVA043rAx5UZlF2OKN8AmgmnliNog9s//
nX2Th/KP+WiVXJ9OO6Xuu7/TgczMjObx3JE/nv4U1Wp5iYDKtljSHpvky9XWBrgr
UfxUyKqvRdjgg5Nk4z+zi0I+7iyT40ZZZB0u86zD9NkaS8ApGlyJPbcFHIMGSHZb
eWTIRXcghGIclDy04EgzyvDHPOZ6alhTQ65hM9AdNhQf6jybJGhfvMOR+nUm8MS5
0wdPKLpeX1CpJmzzEDfEKpkRAM4CQWfCbzdrx6eb4QmJEl6c9OuS+1QHr8LTFzZ6
6m8kR0fi/Qgcft23pHjLr49vXDWNcG3vVDRfJms3wAdK4Hg/NTMC8CSvTqroCUtp
dqje500IobN/s4+MaZIVWG24VbPnAedvCI5vLbGmk1tfyd9D2A1XLq60ZjhcWGmV
aBT+5PL/NCj2sBG+yAc7ffDp/Xh5xQdYoh2l4k0qTPp/xmYlrFbkyKsO5kT2t2dF
4sRGPw87FMitQesQ6uQbWNPbhddfxViZdDsXuGlA6vF8ou5viC8TtCq3y2ckMTGR
Xy2QFk2kn7g0n5WxbhFvb200B0DW+aRshO6pDQFACmtRNQCORtdYGv9kRmjAmKib
m4boPeeOsWljvZmLaWX1w18qtvNDeJSnKsCWISU0LSFaaQTfPay0IE3Oh2YkYt7f
gKcwmAwmyRM0Ih7BEULZ7p03XRMvHPBFg/voPW3u46rv6Vox1hZLqfyVFO2J7Yw8
rN+YUo4enIqiOFOhouvNU+LnlSJjHJS138XHyOjlWmKGy1668Vl52xvz6B295RAO
DRGDPK41RZPMlclD+RsmFpku/eBYepuM9g98z8sbSlHZ+9tKb431GxaSlU5kcias
0o6iAgXe6al1hi07eq0EMjUaEgVCtL7U0VJ3x8+os6M+orhe14RHioGUpkHkSZrM
Yo0IKZnTdNlJoN2iGJDpUXuTGzwK6err6m06kecloyj0v6Y1m0a666MaBGYvjA74
27TLpPkVErbnVi5bC2acl7+Cs975p2XR8lSFaVrdx8hsqEceTz4JR3EzhEB+icfY
gyLtC7fsaiTKKdt+B3mMx2lt57dqX3vbpA+97WOwC8CekmnzOwtMKp5c/LP9R1VW
x/2nJiw1r2ICeZ5lQStYyNoHslsZtcIEIxVgFUKmScb0Peo6s+FHIAoqKIJM5pmQ
Zb0wbX2mEUUUND7fLlr//P6+q5kKUYPB7jgzKJR6e7to8ejC8DHBW/z1XTxi+CWQ
g34y/YUW8GgrP+g5pGSol9INevETOoTEfRgP+68UYUSYxhtSp+89hnVqDOq60xUJ
StZ8Oqmbo4RbIf/zT/bwobzLtf0E3wRF/jFAHjE1dx6VEWZvBHRI/p4wR2X2RhNi
8jCW/EGeKHj37rZdOTFg+a8h7xFXFQ5CrViuARDpLnWnKHzmHTEQdXyHYSLlRfk2
0t+uVIKg6gmEtnEdP2mGqyfZg4DjVmmVU8wFkxTW5c5Wy77ZtOcANM2b/64lfQJb
YDGV1MCrhiGphNlWyuZ1kf+pt5kGuuKLNpwrgLriMsHSRJA4FW181LxPkVvai28b
m4o7NsydTe65IY0DqlwZL4BWDobkKMzr9wZEgAHWNh3JhuH053scZBbSBPK3AJUQ
aIQNn8YR4Ly0KUSVnTPB5Wjej+LaX7Z4fw7rja8TwgOOjno3rEdp/baKtj9UOm2i
iRT4v+jGMLk1ZbMqXv74XoD486Sk5o+gmk7RIq9+bPx8kD+yNByBYZKeNUhdFpaI
LaIGhWT1SBbppXXkhzMy1bcM11BpMuON5yA1zrxhcDAqs1HbFAtbmlg8f5T6kbG9
JhOjsodZDBYifXy8yInjM0wr6UbgSW8Z5WUxB983VrHVDAVqCV8zSMWWi76QwlrW
xrchk/c2hePq15z42M72WmxhIb+O4mB0i4zHYuiOm840yqLDxtagcsH3+h3eIAnn
sQRYQqY0AJf7ksOuUhWszcRdqIdKp6Q+d4hrKyO3k1roLQ3zrjsvc/Ks0sVxw19U
+JPL6BFdKSjW2wNEPftoUdH76p3l1wdOaTMmRkua50ALlqo7Q5jv07JVF655JfsI
rIvAeJsgo8mWCPJ0G7E+2krO2eKu0qdy7VBbhMS6BW+xW3sW3B4O3ATSG6w6K53M
W07Z0h4IJMezGsHnpiGliBnnS9nHsbmnKJ1QZ5g1r7NlmWCg0peB3WhGWyqev2VY
YX1MqyYtqEoib8FHOjEj0Ct8yV4AcW/YrZKdTbrfOeUGFfGOSJCISfGglplsPG+X
+m2LsoeWz/e1o8K986Hha12+WNAcvI+fegsdrCoTl97ViSznbk7ppurZHb4aaCkM
dn6nNWVHtScZSWHLknVA7x2BXBSH1BOL/RAuYEUL+s1pC54J1RCswU+DJY3IqwZm
1GSUrKO0YjEvNdWgZdRzxxjesIk2udnePMZTXryB3EJnqeIzytp31KftGPCh6/MI
XFlAik3a7IPBKPKT4NTVlC37LegSk6VwPxzF09l30LCxd6+HkFe7qOQtGhHwBECO
r81MlHQpgPtF5LJJW7N2VoIE8war2Wtml47GC+cFCxy9a/zn2T3GQovTNt3yj7gV
62jyaMil/3J7U71D3cyF/AcqkbdX098VTQ46uflZXLqLWA9Dd+qMf9DtDR5Gio3r
hglbpE46M6OdJVb5bhmFemHXezDsOB2TEFiuQijbtLFK2W2u6RPKpmcX6fCf9xsp
2RIks29pVM+SfyP3etewlRbGVgUgExu14Q1nX6TNR5nLbeRM7Eyytv30oxDvk6+G
VeRqRfpzbKnhOTWaZU5cuTB0xi+VuOGCg7oatO99mCk9zr/7zC8sl1W2BrkAyupv
3y+IZC8KGwL3Edsm9Ic09P92mxZPm2jRA3WhnTbwpQ++wxcu+wpsBTD8Evd8Ad+W
YAwCbBqmh55ywMycl61hhse0lmmp9Mxk9cj2uwnDBshCuThl6JYU3+qKLZ03Ym95
9r5o+3BGB7iT4rk14ZZPf8p/BIP4+Xf1ACj5dc1fDrcdjPUGNHyZdruv/ookUJ6m
tuO1ZgyZP8C5JmoE1O8R7d0B8TqnzdhztnExyW/ruFvqmX7Fn2+dAQh9zYsq72mm
kP8jVDnGR3QfUfGs/eClLZFWFlEnNu0g+ztcgY8UBDtsvJu3dYNVK0Q6WLj6cyXJ
gTwelKnyuA3wYartvljCHJPiasImSdHgH7xj8uDTm333OWwcxyATuMM6lzCfAaOL
TS6TNLDpc3wP1XT8KFv81j+X91ag4UlANMYPtFRvVZKkTJi4sQFOZHq/5C2CAcES
lHNQ+iOvikiUsZDNxYwdojuE4WZZYQyf2N8qBqWA5cZ49L9MBZGV6FugfZ7ypOhz
kqLMP00gk1tE1vU/ZlNXQ//4DUCDRuNu4jQzVzmdVMSVEm5w1wvndIUfvxlXxZ+/
N4yGVxgReBUcgsa9bvqq4eucFSearBFSVCWTEIU7uiEjUvf9Rgx21lbbAghcEqbS
JTF7WP5inwNyoJSKvlk+MIMjb6yDlAGP7qqLXZAuSwg4JvBVHDCb1v6qw6yt18Yr
8vTV9/Yez/qqkzy2xP9KomV0RsCuoUgO8VsJzBMBUdKNz0nLXooIp9237IXo+9nP
/Vzx8hk6RkwBK7dmib760Pfh4xZPTiAfKrvbeM9MXbsIQ8jVwt5dIpPAhZDiP3e5
G/PUpnZrbkXLhiVYAIUH0oVyg3tVXn4iIkSCkcgc9GOJDCRIcNyE7HEziHr2Cies
8R8WS2k0NmfghXu+7gnV0vY09R9VLqbdshL0UALXDzxuSNLKI2J30ulcMhjRxIvI
ajOvfIjCfP1OwcByapA37sIn9t+z13uj0zYnozfHZNNKkLKJQN1ypb53VDy/n2BU
EnEE/ejg926yDuPafRWnmy/i221GQJfeEt4MuNm4KZK/riCVbRFN0fXbYHXugyP3
uDEVgRb1URKnFKeSjPB3cKs/ZF+ljrdIIEK1ashBhMx2omb6Ug7MXNu5rT2cDf4l
KVLLelBrSjHysfNSj/skzjNy8CdFjVck7fbHAmeRGKfM6PiZl4406VbuNwqPronQ
qb3xSxLWLiv4gkjeWpSwpGpC4pKK2NAaB9BN/1Qol1G4GF+ZDutq1N+YoYWgndK1
fUqVPGQrf43LtEpkP1QpqESzNenk/DbNgeMDC2s5cdIWN+fvxImE5QFe8kEj4Aj8
c6dUNp/CyYEY3QugQKkvvQuVXaXiGmhQEvx6Ls3MgHeA6OJRq99wTZu7zjLnd6UW
5uklzuGpWszI1Gt1GzWbO68zBfSNIW97mY/jSM5LoBpfo5zF5Y7VKmgaldjCZlRh
pRkOG2GkJ+uD+B+86DXollvLvEddHnMf9ETjc2gNU0AGhWHqpeilAkxVyP3xieBb
t25Al/sOTnlmpTfk3xfqhew2ncSvNupGGzKUJkiMSXRZgPyrSI8coYpD29TEGkwQ
pw39qOpg7w91lL4IChX9AsLImOrwHBGyQf8HWGMCWojNO9PWSIGtjXVo3ZyhopPL
njw0A84yolxTr354oOHgPlLfGpvPReQsc3SEHuU1Q9xSq0y6I3/VCpb62a20rsRr
OnxZ1RWvNr9gqsn0M+M5ZArImfRWECkBCd8LSGNNRtSN+jbz3b1lYO0p8h1TwFwX
Z9351NcUSF1/nKHhQP+oJi0C0CBItEl2aFX3Jp8Z3ud4OH/1d/kWUzijiPsejz+b
JuDontx2ZAX61MOQnW7pWAFzYRLBkdQyqFhKJCL/zhCMEYGNVXJ563GQQaHYORo7
Ml61i5CdQJ+GAZM3t1+vFztBwoaOt+brY7XUYhj52AYBb9cMikE1I0CTGi0my4R3
vju8uQ5GpqIQ3ggUHIxlECE6kbXwJrJTvlb8KvY2qwNTKxeP/NJ6oITe9I3OHw3w
Bhg/CwXTurE5JXfIfyCroXwaOKPEo6KlMgHWJG5ifGUC+JCSAlEE+iChBpcZB/h9
TgzNlWon5pIuoWMiZTZdMLHD7zmjR0kFESkyp3Ct9T0lxP1MeLMFN7w1vZ2WINX7
DEjromSypOTqtQXygVangow/HFKswvXwp5BD/MdS+Phxm0SGx6dDPeCo0C+mjpK8
xJcrhxA16ioOBrdPSN0teOjG8gVNBWztg4IZtVYWRtLw4E4B+e62XHO61ozIud/P
xGJ5wBscP1Lh44JGI+MAKhOOa/DwyoRwXqdsweyYAfgEOx/5WVJn4ae2tYnsguPR
W+hxnvF6D3jXNFAQ8uBSN2Z179jjPhD0SWy8T//Q7R9+827DxcduQEsrQthrWSa+
sjeMQczYlKkHwnZEvHldJFlUpwCbl6jxeglsLZkoGBbwLDvXzX09NPwS/kmshokG
cIFzt0DsdjjCn/Gy+6xa6gONuVtz4ogj/9H4dIpv2/SZ0Cash8uFxuKZqRCW7xwp
iu6HRbaYHCy/HgMJjYacOAV3A0hngP3JkSuY1q2vtrAMvnNZT51kFovL6I8ZHROu
sC3fAQVjI/Q6zCTULTZQ6fUAbMjUmYBLl1YUx9yBPuv/G6MCrNREPFGrhd4+Yzm2
AsCcu41ZvtNzjDFBCx9NhFJ3t4r/kXXVcOM51onVXPsMojjig5mI8U5Z6zDbz4pD
TD3IOItY/cZm/6ocmKQT+jnuX1Hl4HZWSn50m51lOQ/p5foOqAPLhJ6US75BBPox
7TD8hOW6JGroSZiI0/2o6d+ZhDQddB5+CvqGbfryxeoY9cnfvXJofYYab/RapBEH
cvaaaMgFERH/OttCVFnzSCv5vrvks2zzYVfKCxuyH8EDLQ7EklzvQqH0KPgeLDE+
ZdzoOJGYnMYiH3EBDpHNoTyU5m56ewDibGMleamiuDvX/sMvqJcLyUB+PY65fQjg
OhXKDs22pIGjFo5WW46J3fGK6JPRfg4WAJYGGtq4RMhXHGBSFtHKHkHbFAwedDsO
iETu8BoEW5ntqpnCNRSm/32lNZYZJYk0k+YbqeCMwMLJg6i73ryGXEwVizdi0Z4j
rYzLCz38i98q9pVM09Yfc02+G1kke986pjPq4h4/PKohpehshMed6pYlWHuJdvKf
du7+OjzipR65ENgsahkSk5Faa2MBhTNOivTKYyFqRsDEvdN3F4XwLUwjP3tBs72H
NHHjZD21+fE1kEbPI3MSCf1xzt5DZfAMlrYeye9lYhOsefsRZPyo2boMHxPZ9m2I
lIBZI+DY1dQCY7pDO69W9yGKKNF+NHYYWyZJI1504SGUj5DZUi6u9CCYuCf5SM+x
PLfuN5J6VobHBj3BF7T0Ive56IvMeJa35WNGwTp47Y9aff9v0lqGlkksg0Ln9rYL
9tJPg3+1qK1sgSDFoU4dC7PLEmQRLk5rPHZjsiOsn2sMTPeqsIpwMXgsG2N4X4yH
OGBi8pA+GaekHGNk5+5qjBMSWtdIIrnIflL2smkUFqM+QSCp868JMf9Z1lK5r45n
5/IJ8VlkWUkdtdhVAbGvI7jSbvRM3CoTatpq/Ew775FA4Un0G2gvCQD6euI77L5l
jZH9n/AjAIPe6FKZmZWlphzzj/YRFJWjUVTiefP/98G+f/Iu6KV/5elKbI7yHR6b
FOPUV6/D8y7wmzAafT4ObhzIX2Ku2UKoSVHGz8Pex74swzO2mzpAnWsromRHVMyC
9EcHhvHr0w5XJ6aWHohJ1KQBsPp8aWg8dzB95toJllDpOwma6wltWrnT3YdB7/rK
bW54aHTitw9UWduONnpiAs0sH97tCjsRekphBJO5xRyoh3VoaHubWJThmXQ9mRUH
GDWCa19grlNv8JtXmImnShhNN+U5mKq8E1th7O1roA2iHcjIYEqiOjJYb3QGdbWp
PjrU0kO0Cu0zzTIxw+VYGqua/DBG2fzpugsMFYE/z6K1GWjCDL9g7QhYM230kuMg
xgnunVHuuOjlq9zcIeOkwsRiPR3/Ph1TgFAIPs8sLbiRQvF8rms3tEE9e4GMBHyy
SLiUnQbiehJ1FEzElbERp56T3XG+UFRy2i3EXrizTILKj3D+HbxSvAJPqTYQzwq0
heQP+pTj6sbWFLsOuC39HehfgkPOpKVNsM8oPbipUcoPybzBN+vnlQFBYKeEdVZK
eJBEm9QF0JdGkNFmlgqEuhFqauKL6y61dy1z961tUN3T9G6taO9i+QHPuzbUcDbs
9p5Tg8P+DrA8L5t536G0g72GynONfjqrvw4AOaUFbJmwSHsAdDqa12cI/vdev5UK
/s+4zcc4CgVg5jNKJDvJiKsbOxWktp8xnPcuqQGW+NT4XOhahvNLsMylLsDPgHAy
jVITUcMiSAgSHXs6UcfZv9ucz8BkajO7QYO1mw0mxvlTrSbKyMaeFzKRNtlwPc9v
IA6k/RIdJvz0r+x1oVY3fNeh9FTf1enIrHgTrwge6MvgB715CQmXLGBwhS7d529u
FnrzZMhaOfD1rj04xvFLs38BiPxwGINCWoV2CnDlqbMkHElw0L9TC9t1hltiKgw1
fYrlaJ1yaMHY2zcmJZsXPTVLlHdtbwCyI79JQ6S7201koONdXLiEwkNCrCwdKX17
jEnUm1ceXeDZXKNUO0JJvfBiXyoHIdQtES3a0QklXwJZ3KfAvi4O/0swNIQa9Ctp
OhQHvuCpqCrw0g+C+Dkqo5uoubw/CgwIZZweDEviwrCoERvj1ckDBd/FpncKE9x7
ASlOXBBW5LgLKyuE75ABhOP16GeSw8HlQG7YIe0HR13+12/5x44ImO7WY1zl0aib
EGzrG0iOj+nYVyKg8Omo/SUnv9ydUL4F9bA/W549/7kVewuF5LbKC0jrqupGggP9
hNTulEwk5osBXL9boHOTD8sFIS5RuuGAtsVlRJv45WeXykmKzTywILb+ZgnrkhF1
eJpzFQU6HYDFTjvxhveA+iNrdnHgNE4jKv+bWfenmzGaexR6JhEAfMqHU8y8ZEJv
Gkc4j2ExENorSKFA3FPaIrDs7HVhe/9c/Zbo+0z1B4o0ZTr/ADdpPUYjM50khDTx
mnw2BT3y3dbX6qXMlvIl3mD94WdGXWg4U3frrFgAy3jA0rvN5lszEqY1gOpoWu0S
21WMiSxDktd3YCZ7fkgmVZ+W9doH2wGaDNNOKQqTi5DRN7CzHL1s7bOn23MVWFI/
CxJMLlPlV7yI9CRynzU8vxtTLGFlVF/rlUv02kJlWdMWoq8volK2NWai63LZJ9mS
nKDfh0beqBOQ4ncesi9j6ZLtk9P0GFwi8WcORDYpMndX4rUJzJ3KMA9BHYQO/+T6
8fTTsti1vsuq4YGshB4sb3f05bKPPnzocVk4V9PuI6jSTEMnKAHbUr6rjq9vw0Ld
jrAxSC/gmR5JB7iT7XsPvqhUYMBntVVR+aE/1khv1+z3phj25Z8C3sFDsaR0W5Zy
HGy+kNR/dntcGm4NaHYfDw6b7iHvEA9LkOAJ69f+yoI6F2WBp2l5F4C6DshIPzoH
ZKtXpL+EmXvm8nSZdwAZ/zXPNt+LZbo3ixQgg0mKG4y3Jcq5c5FMbFlNs5zTrlNa
PNxdpJ2tSGWWpDynKBwdSuM04Ofre0I5rfVeSccLF0WfXe2sB/5eSl+0pnFmx2ad
rhCRELP40qSiLWo3+vAt47bmIV07r+TrST0yvTl6sticWzYbBPHzgt2hCefSPYX/
O5kgqsyTlQapzeBKRT+kDXShYhcCr7x9Yk9Y2B6CVT5JH+fue6o2YSbDQlZ+E+UI
hvgGntrEQugTAfUzpAbM8egP8jlZlefxR6EDEBs1RKmRc322ulRzgbnprawsCiff
BEvNNR2lBnRP0qVp+cfYJ3tM4zW+spR3ziUUDrwfaqH4V/9WT+kf12N2PfGmEzmA
l4xhLOxxsiIBqOxQwQzOQy6AfD7RBfJV+WZNiI6Ej9PLntqaO8HE5DTJ3ZqopbuF
/XFywSSmzZpt50097RkZTUx1MV0jUVrqpkpT1j5LKjUK7StJg7NP7E76dTCJ0dMf
1zZ5pUbGyqdpGPr3RpWHwWM7nAx0BIEKhy8CSq/VJG2i5IjWwMUjvdgfRUWMeUEZ
Xv9R9gpWH0PylfYYE89xYa+4SE3oGfmUhLthJp/1qIl7zEoPmumlCha3qDbmNgcK
85CkmtHQRsCPyXZOF8ZbnJPib+sxLgMSJdS7UZBVAxc56tEWEJ4Wh5rm+YdYvBu/
Wg+wiByyzhVZgk1r85YNsivJ0Zwy3cy/E1ooEPctHUdPbvb7F7w492jfYXSbzDY3
+LKc5lc0AJ5+tcLgLyEptNXL8dtdwdLDYC+P7bXYnG7KRRkiy1C94WuHgfE79FZA
tklJzg2wQ4jK+ocKluTkYUmMahnb4UZEREWW2yonyMnso3kAgLBeGWGfE63lJmdw
cTC+KdVMWIbilqx7p1ugif6WmS7SYjhsqf6pWIO3BoGCjQW4Yvl1MuNAxqK5HnH2
3yaLMEh8uLxQ720823ndNFcY72+tn3K1EAQqAwrQZyBJZf2oWUSH9BoYxRX5t7Vj
sCxqZodm/hxbrQFycdgN0yVXTs3lxcmXcQ1SFpJu9yeHrRR+oZ0t0F3x/RgioyyU
zL/iXmEzspuraoxGUAQuN2OPDoBO//trr2xswIRlHDg4qL1pfG+Rw+lLpYe4As+8
jTQ1n4xpzI5fLrOlYEJ4w5UlGyqx4jimjuMqiYW6ZuyC4XK2RPZNZ3iXOpk+T0qt
D/Yig4nVv1KJQacJhxbJKMiF2CeS1cTWmH51keIOmurm4dkGUBQRSz18Kg5dMJ4f
/jyeU3yq4YRjv4PK+/BE2F0ZDCWvdEP0Mq8eHAyITjrd/BIUL43THrpGkEbNThiV
RbYN+0hpGoBmTnVA4eTjY/tZnDa8EKLe+HD+Iw72I+HfO34rUQFBobFsFpVs7xfp
pmObuIXP5I9+oRE45gzbi3N/u2DwbES5NjBIF5P+hoBm+m7UzGXJg3UJ537gfv/P
RzhdS/rEk5ZU2hYnca1ndBfEPuz/sqbKhZbjBOyEEO5F1JowczsAheJnawOdTiYj
VnXvMGYiY/MOX0bhV2pfv8q0ZPdIYFDbYBK4YReThYLS1itLdpRQWgVLhxn4K/U8
pcci9qwaONaL/t5XIgxtvQYiIzMMguKY6Q9zjKfFPXpJ78ucL5LL7HQkwzujSANq
OkOOkDHJflh0tdSXBNI7jtn1nbs6oj8290hCA8oYP6Mp7YfIxeRu4ozk+z/lhPv7
8LST8NNPF2A8S+Q6Q49j+SwkgSXaz11KWfYIX76zbYuSBHXiO5u18q6uTtE2F9at
myM7OoE9Y4lHNp5U5tpbBfKFi4DTp9QOfpcHpp75dy6o3RgRfXGtUKRfYTTdOZ00
+BfBqEGU8+sbEKKaT6/ccDWufyh4IpyzlaWqlyzalPbN/5fLNV77FAc0x2Mk3HGG
cH4WjNCkPq6qP0jdO+xCeGWWdZyeAZT0xQZLoe/4aMV/oNWevIE1Hv/iuTVgtSYU
kbDkSlXPnOvnLc/6o6zFdGlhkgFEbUOZQe9nrNy2WnD2JbDiLT0GM9dAAdKLo2gi
9K4Lj5g57m3Eyr+SYnfzcCUT/q4NK+Jp2Kni7Zhd+djZd8nCo88EddBUcvQJcdWo
Dp+h2n9CUaFN3Z5qbEOMghly737ceCWpP8rVPxPWPwhKCdygl+PrYIklqXUy9pk8
5F+KBmZd3NHGEFmIsD+UQromMKP/nL6o6qCQwfmidfq49ajQUMVGol70QnV4KLxT
kyc2hs1VmxkvyWHncDQHcA5VWi7SLMJR2fVdusEpR9XHYH9ye6QUAmpDt2pkmSag
Z5OxNDOzHDUb35x8vHyCCJMUwJue5CXuq2uo3mz2WJoGz+hnBom7QHX4Qf8QxHks
4ciVq5vFLuRtu+l5olhlqmIH9wzVMZCzHfAstYgJ9mGlUDs7ugzMUzzpn5nZPMfz
ir5Ji04koJLs/Jgq3rx+qIRDdLcJjicv0Kyyh4QPxSQZdHCfhpnUaBg2vhWCGipZ
ZNU5U+5/7crsFkzIQAIENgY6chJBp/tiVaVTC4AqEYhg+Y3Gyh28r2RoDpGmSvMQ
Csi/NClXJd1L3IWEiEkdv/kE6quk5Dtd1FJVZHNJJ7lOA+33U+yStqkLq+gVEeY1
DVRcSW3AAntwGXm54UEXXqke/9wgx0glQf5r/yJqtkUbQhtbpzjAHcXAOcQWvNae
LH1Kw+Fcl1kQDwXUbKZd2W/OYqIUtyPbR/Ikbg5QL+IUVZyQ7IeHMzOmILK1NGf8
5kbGljesHVMcH7b8ISaOUFwiHQm3xQA2+H+TEdsRkoFUDyIJNZRBR7YXggFTaGHA
3oUEy5nsuvvvKDyOqAJGm3l4DW+ZbL8DD2n6Bi7Ay7VAGVxUlPZGqV1/iaMn1Rln
33imkOBy6WiU47Gm9VXl3/5LGYJ8+EoNfTq22YMQzRLyfuqQEi6JNpVdpZ5EjwcU
thV/IEZ9IMYkmr4RHXGPDDaq3svJndbeIFCIhL4DgvsEo7K5KbJwsKQ5kncLIuC4
jT6PEiuezrtBr8PPR3Dlf9XvwjjNWPZ/zckLw1pNESfbIgpHsGUEbdGqtDn30Eyt
CuK6WHsSFP0Igo2YH3DjCb0Gz6u2yuVbKAUQX/3pRgAtJTJ0s4nW5zFOwHyleMb9
7WeCYLwT1STDaldS/5iQnBKP1vScwyf6boi5wBHOqY9wBjt7pkf8AuPkvycgGDMl
64mhREhBrohC0Y4Ai2PsyS7o8k0T0ZL8IqeE4COaal2EIVxzavxkoR5lTjXoUofE
uV6wHpypqVItVpuY8DfvA9EimDed8izW6cjhCC68HCSHzMZEx/HBrq+SiOtyG9XW
xAQ268eMaeY6k6VGyy799/vjqPI7ZqW5vXjIcdJ565e03ZN251kmwouqKLHp2RmG
+zwtysx4EhcfLzikomy/y7ANZFaqx74Su4b26KtG5iTQ/o1KDm7TJYdN12nPOwTr
K8p1/Ql9EwWsu0wA+O7EeK4wQllRKVlKAZjvwAKGMQeVLat1rQxnEHYKgnQQyRCO
Ko9f0U4MrQEkdGuGQX5FSx/3nB0yzMyKQqtaz94KEZ6h5ChqOI7vadYbjRHJF6zW
Sgbt3rWzJw1bZ6O32LFWpyLGoTUolP5kaTOh+g0WsdEQUcOQI1AmIK9e3MS7Zd84
sgloKkYf5S5TOiDkn74djhzQfX/W+eb860x8LbtWNChwht8HPlRjKamUZ7P27cz4
A1gCDJLt/NA6dL168P99krzInrygqNJURqu95k6au+T1BtEqhAxWDUNQaYh067eI
qnCca0JbLx5yad/s+F3tVFsxMBjvfzCn3Q6eOh3w7TwduSgeWJwPNDpFC9CqIKyR
Dz1eblMubVjXVQATgkvXRmoBYvu4qJlMwOpQI68H6aIhzaWMXXdNAu1M6WzX6dGg
io2rnwZIy0SF1dkz6vq6v69oApKB7wRCcSKApRDKwgcQTMhej4bVX1cDxZ3BHvQs
R/riCg6quuJVWcblsVtASfc1Y/IAC5sUE91uV+Fz6AJUsMTzr9fgEqLL7HgTsyMf
Gi4cXXR4iy3vM66JvM120E0IplurdD8DJHiHws7+cl8vOcUXyJNtkc0ymOISJ9SB
ONWGK0GqA8NkcekEZmr1cXMnronpaRS5yCwPaMhqUHXvteWxQ+vsomXPBK0rfGKG
BsckhlBrbR4b70ysuXbobxCVxs/RXuA93R/JbfhDQSRDl0V4RF05hwgrlalfQse0
YmZLHYB/wDbgyHa2tMf4yEpl135mhrKboO3o/tIac43E0gC/H+PjCWJF+xfE+9ED
ptVdtftUY2XV10G2XTEvHPa+uIRH1+dkQZsd2uNN6fpE25Aaeink2BoOAT60bu3r
9eddrfYfDejxlkkdxijCI+K092xVHhhT6TyWDTH7N51JyZv3yxR8xJBlzktbyudl
Rhkmz3nIpTSWTX86/thtbq3IyHF0740//27YZfue+M6ml1L0EREr2fVyLIYVVEOx
FhoilAlYpyDWIS+9VDyrKMpONANP4vj5LGYxnQDecV1WdBhXWhmPFxf74feW+iLi
zqmatwrLxTvN0EAB/gYg6N+WuOnM+rM1QAFo377a+cM+1K1+7pBe9kfMis6N3d3c
D422DVRq1ow77CSTSN0v/xf08U71xD1rjK/62hrHzpMDJ4NYrw7pWYv6E7nBUzc1
Va2/FkdX0fc+aUCoccN7NnkP8hjDqgQd6N0chtSiGDktHX6vH+HRg0stRDvXqEl7
lGVWT7Pbvr6tPs1ds83/tqQ4bcPnqxhhrzNbE7bJq2/Ti1vYJHU6UNDlUUL6sBof
6O6aZLxVtzhRR3qkMxrCzQalNoFf0PS7a5ItlVsK3QllD6/5lQPp9JGH1guHzIpd
p0AJXAMI4iTYilDOvX+BmJ7ze55nlmFkPG7YsckvOPavjP/1whe2BnXaMhrcdxLf
OcjMR8gDiw4T86TQ4WQAHkKd8l20oPx/6SE0mMlFtMAYy0QHqyTotd9ocB0FknEk
+xeJYgWEkfcM1VDXx3SdBI1INOh3UX8ubLzqhfpwgs6rncTPqHUuTY52dp77ey9k
yN3n86MkuYmVrR+/1FIgkv5ydHL34ZXbj2SJurtKJcGKZG/Li59X1eI7eRlK+5xb
J/9XmBxqUvNZk8O9MblLmbKQJCVtOwoRhhc1dagak9rjqKfRhAbxfoXhRFJaNs1Z
wFjTxLjDu33kslclYK9x3GBMbjqImp+9eUygTTHGKnx1FbvSKRjtuwdl/C4VWRDq
49nha0YvNmR2e0F3RhSD9yqTy0OUBShl4bDbHsfj0Ee0dDSAc4gkU6Iyd9z5STMJ
FlNrPoIBawcdQpxoIQjzqEah5kIdYhyBRpYsuvA2DIOTEvGE1rgwVJUoq2DSdDqe
z/bzr5tsx2RDnUwSutSvUWNp3CAakjT76Mi6o9vICBDZkmeC9szEfYV7TCznK6Vw
qfrJw3CuVNRv5xdVLBEb6eWZYtIwCFI/faydd5ze2hwaITVsgLvnFMBftfL2msUO
NUibgVO2wXkj6DzI/oVS3D0OOo3OiIRfijSdyBg6SrCUeYqVSxHD8TnEqOdaMel8
C5qwKeOGy8DDMUovDl/9CK2giIR1KBcBQ14VkwPXoNnk8I50e8CZ7k/2InD1Mz2v
dJoEfosZ545z1rx7/S6DEOGxixzEpv8IS1fnLg3QdIRUcfBav9XY/Yan+4y+FnIw
nZtdfRjuGSmxGbIeEkpTGiIECmNEt84b3tFyaJksv2w9oyhiEX7erQDxySWmTq/r
tMFRUkuVOI+0URqhjgxaW5FUkuGwkWEHP+yJ1q+pDgm6sqV4ARuT2R/5jnAFeLck
PK9GojE2f3vh4Y7Vap8XPUsN8lhwNi6ipl25ia/juSyvETjSf0eL/fxIQQq/Lc7b
ny5tkdlbCV8ErjtBm5zizNjaza6Y4EJlssYXvRGBa+/Fp6M4frUWwOTi1/6fx+Wn
M2ZfUK4yQNpIEOowsoRwicLc6CIUPfEzXlidHV0QbfJHYDAwl6UjYm4R4JUoMjkX
jsjpKzjY6sI5+osRz0u9Fhwg/Mufo2LeC2hNScHdpLNl1ZsFXiIxuQeNLOUfpQwc
1Vj5kRXyNTbWZdiSP0fkUMig1j4Zyvz4D7TlgQ8gXvZla8lgf3kMkiW/rq/VwWSd
oCGAGja6sdYhSkR/CnlsfG0v8GPkQKODmkDEnVz/qRlEDiO93YaYf9I2aPvBDrv0
ifhgXLug7dcLGr4TUEUSL1/BB0B3Dda+p6P6S9b3xqGT3BUU33whf87mfhIeefhe
uhuuy6Tb0qYgwJoLCWhnB+DyBX6Z6fKY5s1cGZwXYESa0LokDh7uDccdRar3uzQb
gVUFNNY+FcSlrJtLdZn1RWTjOSuO8sSDKQ70o5xhv0AMwruzeWat7G+xs7d1RHtE
WbPM7g2vx7U2clAoMRsr7scaWdDm0GhHzNLN1rPNC8zYl9CdgGk+TQISSQKsAGNn
QU+fBipQRGSnvxC25Al+3oaLzbFqNG7NOO8lsMzy9Yff4QWi76lOQveHeofOe/QA
i9hhrvCO4N5MVA20Esz5G7kZXge3GrLA263H4LxLJdioEDn/DOaEu40KsIlzgxEZ
fXfYBsbEiG9rRY6SzmddgsweleOHYMbn+dTpMViReM08chlzL2H+578s2I2KZqHE
j+P6u1R7sXuwYeNGPBLU6a1eCXLyQBzmw84IYaEEBvzUQRBJZSRg79Rvu6d68DdZ
JYexVDw53atS5Hq61k1a8FP6V+gRItZrl1yWX7fLFdtGBCOX+VtnDcDFCr6TSLD1
6veJJW17AbC/oX10aBAzfE71c/+gaiWhEUUsYMNEVUXgINMG6fmH6ifN9NKIP/FT
VVJV9O3xd/mbLkqRxro0+G4tiYJ2hjXI8oUahgDPpGnxTz7wae3LTzRpgVE2x9Eo
0kByYdjfSd+SWh8FLl1b8cEzO+cahmEVot+vL+K9rzIMjjJphbGstoo4yVHhcP3e
UBx3nwtCjAQoE9flJPGhMJyeqCnEB7jA+7VI0XazNf9bQwDtHq62DHoY7Eq5RJqs
DSU4bfElK9Eob0t3KpLyfB2h/oQfPN9+xo46ziMZkaTyn+kjnrEOLP8jzEu7b72+
yTHEEM09wJudnF9pXDmJv1wkP1WqDni2/LzKLXf6G6pu9vi/dZUZkshhXjbCGLoe
2o6Uz5jmbYdZJzr5itwr7j0DK13rqmG4skcH+lWlhzWf2FS8Ninz2xIe+vbNpTXP
AlFlAhiSQdFMI6D5rf//rhcraXh46IhKdVOo68xX6p4+vJlWKy7M5tRBMwS4EFwo
m1MV0errXLbUbLTzShNJrAQQKvrF3x28xYL0mu+YNo5GWXf7lZ/bXyUFmC12u9Yk
XJWfiU2sg4OYWaC/b+pX4C9vrlEJ9tvD6Z6jN0AbtAp0QXuoEhPQjJZgx63TZOrA
3WR8QgN5YF13MfSgeuC/w+fzYuTIVoklc9GMtZmz9XyaIOkAKjgXDSO4D7kih7Vr
88vuk2Gye5ElHDRP0LvSbyiWx0EuU/2S8lzxRK9HUQzlvRw6h6aDZIOEVqvCj6lN
p8ci58weicd4KN4EfaQ2ugtM311JEaVXgG6Emq4rvO9hu1ugcTXbs7cFDZUdCsyd
/a/ty/CnxG5vC3zaYnN4bnnX/yYzfj/Q6kiQWgfnzExcpLHyvHT++Y1ad+oAvmGV
9P/i4LYwFOk63Y+IHXonhaRlUCnLVTtCvlUMCrnkPSY9yDLEiXBd717EOM7AJGwi
3VBNZTcwqo8gEfe0Z/lNGp/oTqAGSpzzxEusbqEs2HgwZDsfjHze3Uf1HZ+Z6X7J
+KGfKI3liPIEMDubcrRVlGPgaiKg8MU0UTZ02NNna1aALC+XssRozzpHYx0sq+VM
YNuemOxrNmdFTkQZhR/jIiPGDaALjhLlC6MOTCQj9LnFWiakpmNH0oUvT/3cY/tc
ToYpQ8oytg882B8D7vs9dhCZ/6Ut3I9AKn2IHnVyFcgNyHLk8Wvz4l4IKtP46f2z
42+5zLDbYhvpnf84elDNI6Ej4DxxnRUIIsd4YSvXvaGemIQEd2GZvmwfjpaitZSZ
RKjSPXoxfKByVXlz1br/cHWbKJq+0kNA/qbHbF99OfBTLP1QVauCDCvWA6Qj/Vtc
xur05c5wNxksZb4i/513UK2m1zdT1BEMuZybAmI8OhO67PfjBSpA3aolq5iD/vRR
dNv3LQBD4UnwVE5l7e9qg6reVDLVaLXY9lmt0LkAVQbaZ1wCnwTX2GAqWQ3+Hydv
5oc5NJTqiyTdoNXJ8yCROqcBIO76rHj5EuY0enPmGwZjR2PFdgnryL0xztFJOgOb
YW0iJKB10bKEOs7gqqCZu3WDft0+CRdlKT5W+MyXmEidEN0vpTHdaCAs3hxOompK
ieaK2uu7XQulweV19ulEjPzWcHFxpHDoKxYJNn9n8TBNrkMGZ3cCfA9Un3pGcHRa
i9ZyAi66uLobvEUmBfE2YXqZPpQiBvBfanxARj4NmrCSRe80LfGDSsrbcnLioZw6
RzkGteWywS+HEO4zCI/X7Bj15XLdM1YvdScl3tpu22WH+gxp4sf9WyKs92RYz4+d
8kePJDT/f1hDYaLdkxWC3/kc21veLjSdsUSeLnyWfSBxrJb/zS7RjV4OuMqKIuY4
kwqQMJ7gKbRjY4ZNXhM713VVOJtY+KbgjtVIUsiCwec8ZTgd+aaG28xecYrcH6XE
MUPtly5HVkuFi8T9B+Q0Qtb4FZvXYyz9PaecCE9q5BYYyZZUT7BPj6yv3DfTFVie
HpAbXYKserIEYb/mepPQuuiuyrU0GuKYI6PdLfPSVOJh4KZhNBZiz/qKoLAii0t/
6g0SQ/6qS2vh3Sn6YvV4ZqJl1yoPARbtDuANsAyZqh6Tsqk6cbacV6AjkDok8Tb4
nMjCtd4RkNpMp4v/ApvEDQLobapi2FYYVXz0Eh4tHJ0rjd726L8A2Vizo7+LsmxW
WWLIpBPo7+mb+VmGvlQzUljcjt5z3KdrjV3EE5ZDjBesT+BsbPyopTLAmAKoIBmc
DAD1PcaHvZEZyrwc1ue4T6B6UmOCaeW4x+EWOmvH4nVC0mwWDOvtu9LdgCSvr2hu
xrBCujcDvdR7pmxnvJr3AIKWw695IGE/AP/U9Tt7VxifRqwLUjYwAKvRqs2Ne07U
yatSAkEBejq5CLlkt/3SlqRfzOhHut175rBtC3WmiJ6mxL75CsnLw3Db06q9hTFA
EwdF/1hqFF47i3Gk/xagkZcSDg/Sq5nWi0RdwWI9wcYCIbOgZpX05u7LpCEqjeJx
C8cSm+T951MWBNh9dPrZUqJRyiDE0ow/HK76XSjg2EDNQRbksdLHkVnh3yhfEZjW
1OIkwlykY+eTqR+GU+w/TII1Q2twUXOEr+xXGHrX0lzSi6zrxB0ZFzZ1ojQ/Yl46
bCwNf/qml2QIQdPBB3/CfsLeUEs+9PUKYRVdd8sVjTVuC6nv6WaYukHm51fqPqjd
ipPDvYf3eUoxPnsLziNHP9ELZX1MyluhtQAI4la/enBdc/MS6D499tred/QC11cd
xdKoQ10tFRDP+P2vr8kN5iGWVQ3O2psvBsxS8W7aHa6ZrYaYfeAC8uebuHVlgSZD
4cYO10vxWjZ17RHyRVSg7iu+++p6e3k2J0AZDCY+JFUhdAPH3BWEWldGMIRJzJPu
dbwJKm0iqOrbXaXdWB0dVxqVDbgQ0/oWCWMnI5eoP9dLOUCbZ7Unp8NtFLqo/JYK
gplwOF9dsZ4FBBbMjdWNj4HSD/KTl1ulw9Y71xpNURMUTOGKciZU6dcl0Wm4SvqD
9Y/5YAip45OSZ0LgD00bUOGiiMdk/5ZyUO+fSiZX/dsEqqgiH7YHuwHUvXI1RfaH
aytb95zgIijvnf0JjMQbKSTp9f3mQgxxfAe/tWkwzZi4nXnGbWYm6Pt40evl7X7Z
u+w3XfoIICQnNw+/QwgNzYVZb4R+p2+XJ7+UQS+KoJLZf+bFp/ClRrhNWoIykNDo
4NMrHdREoMUEBKPdc6rfcC6eQSCHFoLIduRM6qjKOHFUbxRkHM4EocRIHj+iFEuI
X0YDG/iXjxHaVv0e9UU2edVY6/kve8r4czgG6YvQhaeDYyMft3UrjW2ey6gk42yj
RKe8F+fpyPI6laiQbuu4RvcPPWEc23Vk1yE2yE7IzbgbbJF2Src1yF7jhXum+tg+
X4RJ0+D5Lyd4LvnrS/WeE/EE0gWueus0KrxrCaFL1QAZg5JIB86FUyO3ZVCA0nXI
OCdR6vSS3hvqpSilCDkc/zIM9m0cS9yTDWLziloGLiyRcHjE8ZRoHcWVZGhiGPhG
UjMUW9YWyJeOXCJyxDoZkrQZG5A/oqH2RRe2Sw6HitVBZ5xgaoZUWcZhYkIlLldI
T7Sfi9MIeiLRu3FuBNHvy7mmb1JPGVn4owuo6vbYgOXBSoDcBx1TbMCK1Ybr1C0+
mdU5b+GzpymzJqouOq0ZrUvBLe9/LmCBFmeg3kCeWyAE+6vq+5b0aT+hqvuSlplX
utoJmpZJIq4MbPPWHcphp1nO4WFMCYA00mzGhtSHNvAXGEkRwCJrCkKfzcQmWLGh
bQ0FSel9Jg9I0xRTrFZ0izQjaqrROcxYYBEjs5hFsMvBltU/U/1x9ZDFXoQxZMft
wLpU41shdXqxHr2pGtJWqH4Sotn6ukN/lEEH//VofEf7friF+V+CVV3u9ThHhzZI
uG4x+R2YYBckiJGdFedMaKWmlwiDs+xkcSMqmXT9la7Yo0rNt2utkEWIms7eD+K0
lNzRuhOJFFoCUjn7KRtwj3roGVKDCGlqJcDFSlnUwarpi3OTPJjXeBJitb2A2lt9
7jcKVp3MseDd+kxZrCJzfEcA0/AYq2gpyzXZFtRXSaTbgxsFyW6Ir/BvNiagEB9y
i27Faq+XjLpA6EsmAWw2vsK1dSO0hVnqzURZ7bBEjRom9fPYuF30QEZnhF/CKH3K
ZrSDUxU7O2jq78rVAyLHqipfQfK2f1yydGeXTY/ldxohTBCdf5z3JIcAZaNGuCCX
HSdZo6fdsFQSMTmBr+c6djPujfTRCGUber3jKNIz2+YJl9LKzJS+XD66T0yT8+l1
RJgK2lJfohk5znN/noYY/WgDIkBuEVY81kEn5uJs0s2J02CfV15SZQaAt8BFqlCY
+tYKFgL3ZzCNbXttEcEGMpgPFuGd67sjRrvYpQ8yFyHqyDkKiVDIruech+8DLOe2
FVd1t2/j8IixqGDOA9LWVvtXMcxtcps91t42PykMbmCUKCD+l0Kj/p9d7ChyCuIl
EKDgAMi6V1UjLr4evs3LHjkNWxpNOV+EapTeARnKleQSjC8vgG8/8g4qvyN1TapE
HldJu975DZxoeUC0c5iUJr6QCEwHxHSlwXrx48w398I9+ilsffvNrujrYpMrytPl
yHB4gjlvJMhVBP0L/sn2GbLHc9q8spk0yJoJWbFx0ks2N/lavOVTteZDoaUKZqjF
Qyepoyq9B9jyXJxSRGGCvuueIz64sdCJOueK4+94t5/EfYQxMBPsWQE/9s8GlLzD
QJjjJxjTTvQxe44hODn5Kn3C/Xo+/iOhD8A6fGWekNwmKuBzC2RDgPbUpQ7DNsaE
iBdonfHZ1ZyVXqYjLGy/zCd6HsiLeG9MWTpScSfHKnTG8hzB2qBWMlbD65bhcShQ
v95EDyZjWs7gAKDQ2Au8rUTztRw6/1niTXkeDtBg7OqGOvvt4DM2SwXKAQi0Ky2e
qHASwSBwbfmKEDENbYPtuOgeyPwyDwUbPJgF3Sg0K/l8VNtv8sxTEcSP2wKINGtA
4bjkw/s84V+3lvoEmljXZ7aVdu5SltwNUWOldIEPxaHt2hoZz0w6uq1W+HKHIg2o
au8X0SbAbiE9ehs4varvdyu9ttyd8I+ESQduM0ECLbMAmN7yPI5xtcTXf4nKXsAM
lu2Xl3iB0ylc8fqP8JOTgyNalfbtMvsBlqvnaZ1kvxos/OJvYMiCwBIzV/cTGVz6
B6lfDEJQ/EhjYzsCmb9yiUFX8W+1XpFin0DFb8ASYS5zofDRqs1L39pdoN3dvkCE
LM/4uLZ1uySlzrAzAP4aSSM2YCuOObEIkkjXiz1JkGJX52pcRIBvZBrymV0cQnPZ
gpLKzYTZHbep6g6vNaWWlA8BatUJihuIbkvt/DoI5KhntOluX37MSMGe8lSz2aR6
B5FELNqghb7RzJj54s0p8VhzG7ZND2Jbzz3zyklzqASH9JAPmJMc8/7TVfDWmNlo
7cvfPTYe41frtR3cd0W7XscXBhHWx4IzGRL0iP5JF6kRqKZcY6BWliVd45XZmnye
WVEMpYDpYqnry2tbPrUHoY6HCW5hSUNUFZvTXCR9TfIh9mQipUazxsaR9lDfMsol
IlI00zAxK7gt6jp17c65LnU94bHG4DTYRzOqBImQLxQtxD1KMzabrqaAWMmVUr3y
Eixul508xe0abNmv5HoYZk12ON6XCBstYOKsiE9qdowkyR7Hc4s1MsBlErc3Xb4F
nAT7Q8YayD/P6wLlZq4O1XiKGjV4sS8UYpyfg7kMBubWa0suq9KImANRsR7MY1Zn
oDtQlwr7dIECm4mMp7kt6yqG6Fbvb0DAHmYGSX7+1KYdFHWTBGsvYf71cJN/OXtC
Cy5aGZep9WPEHT5esEOglBGj7B1Lqg4YZ2D/O5C7uVvdcJil3jWk0SrUFUGoVucX
O6cDWl/CK17ls2jVqpq7jWoy9ixgeHYEcQ9zt3JpS+QBn75Bx1MFQqqaQfAiu32u
V6i1cRusWRbwqqfzmnoRPT1K3lvyUR7iBXwQzMIgfAGWyqpG407QDjYtp2m8yP3Y
0wUN+XdOWMX0w0DQM8aKC90cxxDSHFc9mpOCNxVhjEF4vp3untBzuxCZSwh8zLhS
CXMunkC9CvIO01oaKD3cxx39umk39tBDbqpsCHIjNhf8R+Ny3wsZZcbLuO4IwE5b
F3A0P/jjxF4HplXwvNGUlv7TZ/V8ypgznoHDpB/yqLxAg6UwTAX+wmwlRvGvtRFK
KCCdPJPBgiYRI5rbomfUaT2NQjpvAfC/tFnJQMY+eRlRHRJBk7jO/kw7WX2Pov4I
KvYdkhdrkI09EMHMXHKO8g8Tz7cmDU+Qk7WTsuK3JyYfhUR5FxzcRDWBdasI83zS
XWEQUzCU2MPXxyGwhR3WhHMVIJHB/ryFaVTKyrVWQIjs9SJ/9dFh2xggfEOYgeca
yH9bZlhSi0umHmn+cOtxviMMzQHdViKuaTaUFKw0aQPCaXet4sT7cyw/axtQKkUo
07mit8W8mPjJxuZMSHTFiyfDOwZQcwt4zfsSKMY+5BbYUrNrxhWYMgf1HG2+l8ke
/yhs2FeKlnd/bu5dv2QSlsHw4CKGf4vqOoBVhGALxIaygbAGd1JRjn8O1eY7KBum
hZU07eDlbJS+6q5EBlc8jcw3F+0e5iR10DelegVKwzDguLTqJfX7+k1jRkEZkUGa
LSgJ90Te0VoF7InWxWeSTxUORKIAZczUITqrzCm7Jd1OpHFPpmjog8AAdHai1x9a
cSr4d/tQJab2NuENyfLUczecZsOMsYyc93WQ/sbh9ovM5vNdTEAmSOrld0LS+5A7
Iqs/NiK2yVIZtqaQ0DdUZDN3yNYuAOYlk/3a7lV4oTnPCg9KvqhioZ5107up3ebc
qjCd4Q6T85k1jogZB4AUbZDYemTwkowKKR9R5/0DgojvmS+XspLN9c02bnP2LPQZ
GXABbkYzoCxReTkM4VCcTLTdL1HCYnqrvbX5WyNzx9YH8MaLv+VWMYCeKZMHoiFL
qGvG+fwfcrXszyANBSCgJ1+V5ggliKYoFK40lcBKeP3pFv4IaA06F1K6Vgpm2Lzl
P41/eN33Nl12H2asES5pE02ImRHnXXrPqz0y7/Y5A6/W9eMDSoh5/MvnF5prMad+
yhNoq3ntF5uJBcG960vGfMaiDBTSK6WC2mDJwHYsVGQdZf0i/EKzs+MSun/wj+9T
RKdIwXzpU3Vq+L8zdRm2YZ0aoItwsa3Mok/eY+BuYcVmtPOil5fHRde1o7z7w8Gw
WJgQSCrG3t+ga0ABIVMiwjGGFqY2Qu0zUAfUEqHTK5WkTKTLl5zr/DNWETIbaXC6
LgvZoCdS2dA+afUQYG5OKJw/jKoEkm2TMeruFCJbdXTjTeGol+OTM6qZd6t3+KPA
l5UUXVyeuXhHfoZu1JYuI9Zs3GKLpTKc30VpSIq65nMa3U0bGmmYIm2PreSIJAUB
aPDtTv9t/2w2iVt7p1lI6PYZiIitBCp2oOcIsuLSBEllgWO3vxYXLKtuk+b15ZcE
Efdebtj9xViVW46/glWpMdfBUT2bJMK1hIcR1cc1gAoBKT6IG1pGrzrPotjlBsyZ
nH4uE3jnfHV24g6y/qzw4EXrcCweefp1dyYsynBsl4FNW9FC7SPWMr5Vt0bpnWPj
ngR2IWfx5w9nMqB1l5MDz/rvImDT7GivI2zfBiBWgDAxfUXN1b4doR8NG4N7hY9q
Rfkyd7t4ZN7DyonMWmw0B8CiyWXPO39pbC2MrzbgVJZzFZ57NkYRqf6EqWXCRfj9
upH15NQmpf8AK224KftWJWLU2kyg7ft/4dLs/IULp/FBCqlzf7oEepA25B9vc+du
sdrZUORHEVfQWg6eu0CSmg7SRF0wY8UvvGDOuGMYx9Fc/TAZaq78M9SPiUpSIcsJ
wDvIS+UtFUykhd/utbZnBd2x7oggz5A6VZpoH83bRcWZGeWdf3nK4jJLhD4Mt+xe
G+zfSJ1Wiuq538iC3epzOqYOKPfQaQfznY0saashqVUe4actS+F6gxaal9VC0g9L
LvnqegdW9qLrPBK1M7dec8xAvbLk4LDqz7gq6hZf+Yqx4s17NPnMeQaN94brI6YJ
XRnl/7EmToE0NNZZgwKTT0VUTnan7bsuQrPAQ8rdFVMTYJ44Z3xU01TBzusfOFCQ
3AULHEU48k5YAEWwKiIB0rvPa60xJ1GFaoPojcEMabv3JajAitT+33/wEZoKC6Mg
zOhSEi2U8cSKksyxy5skxg8SnzO88/lYSZisFs2AwhxS+cK0htUt9nlVMMo5qCNO
5atHSFpHn7Vl+f4epE3J8ws+Yf7xqBVXWc+2Z57d1/ivWVG4eKK5tx6hipE4z9dJ
zhqHQ7Y/OEpJVqWWiQFpS7D3cvXI4I/r4kPPLikVpVKn/IxdPQVR8p5ABsX2l9j3
F3W7vcHbuqaU0v63Fz+jt78WpCmsCCtqRJ4x2CPDoKBNx6nZVvC1mYAk2DKyiXPb
67/HN9PvWUA50ZwLYxAADa0Usa+wezSa7fxA3RgXWaUV8eFxRcFTQISiwfUr/Kmd
WjZm+pyRBdZYzk67LmUiH7QOLTobeYRalSrJR7cJfWZupNwNPklQLhY4gDT6FnKT
qyuaoqgeVt1vKtgRhwIQr+M3GjRM0s0vU3XXp4EEh2K4f0zikQLn25PjBk4whyMa
dtQdubwK7HfLu1/2qZjQghGkRIIghhWvpNMrixT7imlQwavhR2PGF3WT3aFJzfIr
UoTTyfVywyLjwrToUJqS4Ka2wKebuWebvMoXkO8FwZz4h+b7J28YMm5Nt59euZpg
R6J3UM3gixwxlxdxEBnluQCcGyz+c3q4+Wn8erv3Dkz1hajq+Mj7hE7JAoQ7huYV
VazfMkFDcXEI3gWcBzI0mKaAwRTgEwHAnjbUNbHaz23uCKhHDT4+QyBCzUPMcjWd
R7OrhCN6tkNL0N8w12llDlYKuhFsGu4HczHMdkTfBTG3YSaROzs7/eykvtmEHRFG
2NE81XSwNZvY0Lhu+YldBtb2A/XzD6AlUm7ZoEV/s8inY/QluNIxB6PYLqmFcDTz
ss+5PULW5VnLPM/P7qbaHxfqwhaqkCHTDMs6kEx3IAeJZ1XbQk3z2Z5lkV4N3bEQ
M57ObN29XKSS12K4yeomc/7xp+1eXJBtQC+AFUV4WZzAWH6TSaQGqupwJJMHQjxz
7fsKuAE6Pbe9F9lnh8Dppw==
`pragma protect end_protected
