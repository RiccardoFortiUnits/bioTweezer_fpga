`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XGmR29X3PqjXHdXZjz6Vsv7HRqLeODhME8lBAUN0Yz95XJf4NbhofVlVN/9O+85z
DQwNXY4PZytgOhsSRFnhhM6nio/SeUmYnVvvyTcTzBmyS6v1VYEf+h03HJowLqmT
qmiPe51CiRxMP1xQXmogujgyGvBK49eslhJOOw4y9mg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28016)
ks+AcXazZOfR/g68hfmyhCEyXigTIMainD9o6U8tS/RSSelrNqP0raMsgcf7CRSm
U1dutOhADd6OHeRo4kvHS6lyQQvrIwGVulNAjA+M5/Jn26jplLcrqlepjOn+hPgY
WmUf9pq+hEdsWx1Vzu6XehP6/43V3s9GTUOSygdPj1sBT4uUooJR9Pm9V8QgnULo
C6xLxkeRlOcMYP4Yzl/tfrb5NCCtPxp5Sm0cLETIEt0mfVhnHji36SwQy++V3ncF
Ohmoq00ryY+0D9vH03UHR86bKaY98avDjQPzZeB70vmOV6b2R+BDNEjUnDdKtLo9
Rqcbys5/d4Iax8VUoxdYc8RgA6Sfi+C9Iol831LmGHLOe6r+p1ytBQ6DYH0Ruj5D
6XvqwcNlDYKplBAReRxyay7/NGpO6mhwqKUqJ6ilUfZ7Hv/wGmgDQVF9+ylgIhHU
UhIxcpgDCBO27+mt7/6oWg2miL2tDNXDcCxPS6O0JzkQoElnCUJnl1IO+e01NIaP
zd5kpwp9BvwqzU6q7ftB4ZZnJvadUVYg1l8sQykx8+SuRXNK/3q8LJChMbSt8ysA
V3M2rBe8nJkt2bg/3nN1t8YPRbO0+rXpKfH9C7yG/wPzkBFBGM9lExxxKvKK3g+W
dSlp/EqbfiLLY2+IZebN+8vqDfQIzoHGmehC18Q4O9f7AUAMWg2FYeSoc1M8y4jI
YdGeaYDW2J2Hk8F2K3KnnnRZ5E3kiBI8vAFdd+wFhN1xsgwx7QGu3LlyVhDEMHAe
4Rp9i+aLVzuGrGCBPkwV9Fa3ygtxNSUz952xbldEXXmWJA0/Wsve5bsOV1jUJ4u6
kx0AZXyx8uJIdw/ostwXksileOqFEclCEOK6Os5hkwUcYK8pNCsSkXD9eHFQp/gm
sCcvBBJ/rcFhKuczdLJojyjPVudJhmP3O1S2jo5zDoG/+8Xg/C8EcsYFBwvnR1SH
jfwA5nT7LDMHTGXpv7TqpbWCYWf5c5cIrhRWeaEqdWs5oLcv1Bi9H/IeA29VOBGR
a3TUInLwj4K4cGdwAtarz5136kpgjYABl5+e+BGHQJL35iy7/EHGCfpCGrC+ePK2
vjMz26HXgt3/lKoQNgzDsJEmVsA8gmK33Kko6MpxoQ/arMYGqv6Gy20Cq6Gmsv09
Nd5+FTensa78lT2PNIltiGQf+bp7LSSrmvjZyRasf1a9xXxtziKKqGxHdShskwJc
cZ/jUkRZC+uO6gfceGimr6wkZtU0M6xOvKsaThCRPUCg6JgavyOQNdkCcWDEg26S
KRwOsZyky8jPu4/ghmurd0XuX/JMF+EXIcTuSxgC1S7Qbl7SXUxOdfgP3k58z3aP
SbOT47GObv90g4BH71x9tq1KX7PW4nOZSrxZgZ8XAo7Ly8jQy25oeoxgLQbFoKro
MLVlz0NX5/1GIS/DQAoq/Syt80ONvNoZj0J0B8KrIakDW81X+GVGu+Ud2y4xMVag
3TrHqPzo/hPT1gbI6TOFnPOPpfS2RQ9Lo/OXwJOYgXlJQgMX6k9c9RWZKrUHGvNb
GTCRMDzzu4Nmri0oxGu537NzdPWwode1K9A8szBFjKwn0m6d1L1P4lPi4GguZZYd
xWjwgrGcOHr5uWy1VFMZTZRJJHdJzN65PwooTsOSIX1zG7BcamQj+19aBl7oX7OO
RHUm/v+77t3bwvnMMi/NiZ9YQjCGKQNY4KdiJlvEh+DyL6D9zQLCzhL8U72Qjlnu
Z59MwQKzQQVZaEW3+zU8DUc1r+ZzeBmdWCTW3SdM2DS72fHcOniG3NktUZVh81Um
OZmghmhJCqJQiH2ZjzLwdPgnrs+zfOZ0uTU3g8SGWPiGaM94OhZc8UPeQ/DsYiYV
VzDZrjvQMCXvs4AR50ptZvIGQh6U5GU5g8GM2naBEWrQVwusHEyPYkacHWGwRDRk
9JQ6PAlMYvr5rx01yTlCNlVHtRh91mDmXsyr7Ka2VCUDXhhWUjosPwzheXKyhb9j
dj1tqIBN+JcOpn4WatN4DkuKHzZpnOgJzJAm1begYxLjp/msKrro44pQB1uTQdfj
4eISIBh1NwVkPaNRUoh2tdNbe7Ijb70w2lm2Or85oesf6bv5b4Dm8u/8El0qIr13
/PbBlctP9omIKOjMSqTZXOzNsEVqenV7poay4W4D/ntjJglru+FWCBisKLgctMKV
pG86l0NUWXhVV/IsmtXFOlllS/aVP82DbuBpPknWjNPiK85Fp6tJjgC/c9emvLI5
b50CiMtW0xJzU8wGbaW7WQ0xuqsFQVE0Td+dIdJoglZBKVfsXisLK28v4frrrnig
08vgZAJ4FYcDBnRkMF2CtZws2LfTBR4mI+O/pM+i9K9hEjhUcazwGp9XMJ4sHJjm
z3sx5vBE6PbEEisy9udCeyoftJNVpbsA6di0rxv/1OX0/+PflnZW7gEUtfvjiWwk
5N3E9uQ3hbuKsV4ECm4h03C7gxWMaIA8zPHdsjViEDYA45qBBS/AFbjvmQuhTqu4
5A7QfIAduQLfZeAK85IGSgaJWqXZJroevDRLflx7kC8jrc0uSvRBj3jk14fYYzSL
15kV9dPOXInkNkjTyoNsU36i79dn37eIHgyjyW4SVP1sCoLYeM7DciPSAJlOPdAx
9C2WKidbMM/soJeKMYa1tw+Rh2VhOfN9ptd2F2VzZzV9dxjJup3lOJlA9f7cjTTi
sw+dKZB+Oc+lhqtsee4Abt/+x5elE5A6Phj3qbuQrVHb2UyN1GZg33fwkvRjpNuQ
TEBilab7T2oLiqoRyJsF1UxMFKy0tV5qU10Wn/OjXg6fxfimo8TDn1tuqGQ9hwaF
/9EF70uIkr/chtaPRovr8XNhBNwJl8X+mHfD3ev9xfEJ552XLl4G9jUpm7xZnWBe
T3vkblWTs57gpHOSrxbju5V1H+8e8K2rfs4C8n87fKQ3mtjV++ewowL8Ei4mYnUQ
P0VjLyFUPU+duduZZf3chVCMjNfD+N85ibBfU4EoczN39K5DH9LobiHKNyZIckxD
ERzDiXqH/BbglBia/XltwvihDLUQUlmmlMk2pvcnpbIWAacHIwEprASHAm5c+AeG
vV7iCxPG8JfVwZvtTO9sz3LUb7iwUd00+QB+sWbJIq8gZDw2IxDQRIUU5fLGgPBu
mEBCHbWT6//eid8Vx94FJmSr8MxyJAA8yLXbKn+L0XJE4wlFLiyrLFKZekugv4wK
8nr4C0Fy3/PWYt3JUpvir7urrMEsSisw3e1ioq5nPSjeSFHDWqUYyYs4Fmmpfd3f
GhCsHCjsmUQcQUtpMpK0DstW2Cv3dCEJq6YL7wK4CSjMK0TLgelkrdqcue6Jnkr7
HrGwCwHQi8f0TSUYvibgxCKj1C/704S0QPOJBI+EZJYnX63ENTSL5yMTgkNqQa0y
RyVv5SqKN1pXXM2TN50VHWzV1r53MZsBwtquiDVKCK3OkfVFlI7nAk/GE71QreAZ
fYR3bN/khR+MtGRtdbyX6n9qxfyQIjNsazaRe2IJGLAcg7YQPZ3doegfWaYBSpSx
NK44MjLdR3fHBNflkDPgoZB+wARm5WF34BRAqhd1iXy6ndstJ/IPBgtbcLvn4Hzw
ynFFAjZFR/2paW7odbPrSI7WPVHy3g33m60UUc6vwKkOmOJ5ImNdYXVg3VVwsd5H
MjKauaaQjmZItsYXvUU4SrCGFyCjIUWx5SIaA65NcC9/xbL9cLeCLT0JD5CbANdK
lct6n/v+UguD6Yj63B1UXb1PxMV4tlRlfAhcX5aMn+Zl0pazsJ1A8TtlDkRTHyPF
HiNKZK6PD37fsLk/afdzohjiXuQNzKuZaqr6/1zsJ43TQzdK2cZU9KPW9LWpNrMY
K/HrTkmBFm7+kavIUEp/89LbMsgjJ/blsRqmTPRw+RiA1AqXsW46mhg+feyKyfZl
IbOknZ7hXnm9C2cyRz/Llc1jiUyUYmVc0gAQ3qWMH/9cEDfrni9WcsxLAoWLmHPz
N4NfjNyFGwbgYxsmVlMblhojAVPfeOUiZBzhaH0ozkkGTsPg98CFLj3CE/rJcOnr
3LNxqES/+y8K2GFoV/LkmK0QkEmNgVNBtdrhZirnedBBhDiMzGXlWUvVUEKTXg98
hrS3gxECMUvY2LPsRDfAtwaRc8jm6MzHbCA8mwKQ9MisK10V03cfJiPQRG1WifXo
YzonfVLLATubTQPHuyz5c3upq4B2AgLlr9Ftu/LXyqZe5Qtqw2kldepL0rH44DlI
ol8IpaLLULmp6NgMO19m9x9kNB0YPkhSMNE4JSF5ZudnGKAJMzleWBwEe+bzcwU/
fnt8K/UNXueAVD74BvAgROzEWtEptrFQjn8rVu7BcDkEXYaZpqx0tv/BltjsqlBc
Z/pPSqqALNZpjj8hZ2pLakqkSG3Vl4OiyD9h3kwz07kWWpE6doCWyIOlzRNlkFMF
AZaoAM7cvEjjO7ymE5n0jaf4ajbntLxYPT9bC4XFUc2iirZ7ISPZESKw6jc+Tfey
juGw5KtY1EuVFVFN93GW8nYntf72VTId05h5Ss9G3VgCgyW/ZEkYcalJhpA0Up6N
limH4lQVIaet1Vzn5sD3y9Q2vqZG85JmcIfvRCvMrSP5Hh4OTDqY/lhnS6TrVHtB
t5xChzzAXFqrrTx8KbmbHcOGhqmrc9ofXfqhZIRghLWfTPAGIgb+sScQnnHfBdyZ
tGasiUm6sf0me1XiUF1Kr3MKZBbjzuMH59zNXUcbetpD08IrDM1U9gYZ9aANyJ27
HebzD4k+USecpqtlxy9ecYGv9v31+eWpWzj7bCJLYn0GlPgtGUtpvfZXsdxVzEwD
QFc51HxwrMYuMkvPcByD0kPRSGIKLMmAdrSmMx5ds0gNUS/V8dQ8FzYZ9u/3lufE
KoSTHMz0TXIEyUzSPlqeGsMnNSD0FIFl2YPxO+u3YnI41y0LyU5ZiDtbF8opwwXL
z7U+9GYcoL2EBlElNRH8hgoH7Ixp+R+XSxZdAyPZ3r5rPFqLj9Vd8x44CLCpUcH0
BCFzotNO9JelDTsbLYa9sDbubNxb3XEUe94Pw+N7XCGHeGd/djPeg0NBeuUrr621
iaqXFg23XnBOxia/RX/TJa8ZjYB6AB2O69pv7PaGAU3XZCiPGzUuvCp5EnIIB62z
VAObtgdHMy8kBL4r52EqjXoXe8a9ULHnBhDFEa4pcpBOt5teHX3g5vrVISa2uEsy
rB3mvkrPiap27MiMPXjMv0ZlwjEDnCbgaopGEX7fEue7rbx3QzigUqsobscZRmdZ
L/sg2gwZbYntQ/dLV7v1dKbfEdWz/6HnUluS4V/sPF9D5e+nFU0F3U6Y+ivt49kn
airdRYxC4hSwW9zxHFId0lzHc0NB+qlWddE6/mHXnYu9N+woX9OouqHHDPZwmGKn
89gWj1SqmyaEtrgbLnhJOp0CNA63hcbtBYv9jCSFQC0gq8agOC75l2o/SQohcv70
fTVbIM7WU6bdWjefKG4GYwIhbfIDEKYg8vNBHa8FDBiuDRxvquCg4/JeBGn89EDe
v7yhUb0a/bKz/UFJE37CiIMtfd/OeRk3ylwnn4z+hbWpXeZrh/HM67X4Wm9poR4j
W+JCgnNTfCjPF8D4GDU9TCWWHmmBCeP+9fWQ35XUIDJ8PPuZvoyvtVcidh337cIm
4rBA89kDYW8eRNSzLKMpbHila6fDjVkuSSB50a8wc3V3Bj/2DfdYe1iiGTM6I7iE
ZOqoUaTB6R+uDESMp4cC0ap7x95xSTkvB243b9YerQYAwOoebjsUupEuhhE/zVaN
XVV4deVsbZCXfbJoRUe/OQrfg+XtZwK8mQJ/Dyi1A+F9agvBJMOjPJzttEwSfg5J
+zVs3dn7RCokKKfI1O4SbXQ/vOcRGnlZk85F/6ITuJ1lGOsVG6F3kmMxAK/Lbzqy
K6p4Ui3gSZcyUG+blz9orH8zT9mJzFAn6/+fgoWas32RzkE6/6fv9rhSJTKlJ3wP
z7Etrct/NHuv+9x7FZb6q3l+b/y5WiTcdOnsE3JEtMQsNyOzkH2VZOe2ubRVVDBn
H+UzqI38I+Z+OJi/MxSC9a7jIQaKQmYlEnRzOoqJS4W93kloKoe/Olys596d+eqk
ImtgEpmD/Wwjfg4L/nHIizP1wRiXENucodszysMpQZwGINgcVuQNZ27ZtEjczSvT
Ms1Z3xgOxunA7SrHoW6b3eSVfhhRcXmMvY2IUxwvp9D9LXL8DXM9U6DC76cgXTDo
K0S2s4/vTmsGZCnADHcALsEiyz19OhcMrp/io+2mr2fKbdERBbFqlyH6ZaFf6pJA
wcNRLJ75qsQaKp3b613KtC2QzzSDJcaJxNee1tq5djVO/xb9xRhO1RRa8/3KCi15
Ovbbg1qXe1toLpVY2GBDf5r1xKGw9Z5CsBLVV7EmBAp42hqM/TpYxEKc0Hh7SJCH
sXDXrgir0BqstBp5zsHQn7OwxFTPvKLkVArCQck/w1HGMM68avHUl3UQSJ4lwO/B
UsUfOyzD8lG1wussAb+eCLI+2uk5rHK97QOV8XXKv6kaoMm21xLY48G0czBGtmji
5Bivg7ZU5cRZe9UULiHYUWaFh/iVZDkkIOt/Ph28s7wey/gmFDBQ4CJ0ZnX9q3WO
JrRqhIZNVq2O5/yFQh2TpqKxAbANCPkFdhQp4qCjycX1X4wlMihwK0c8Q3zjPpiy
9rlogRLMZfC7GYWvT4BKAre2i8UWKnbxr44LxQaXv4MvnRKBzPD5OcqSKYqK5+FS
IRWEHPIV2t6HqNxUC01Oe9D6GbeP0FD7ylRtScDAdDptsgitfRTrb6x2KF+fCvaA
Qo4br2liMJz9qWrbpEJdZAdHDg2MpzD3bs7KXfVbkCSj/jtVcyv9R99YsE30A7Mb
8Xn8BNdXHc9J5SHuTXLuHZXMVEgH4K6TB9iIStQxKJI3kO05CPI4Z6WFeS+hu7lW
MzL/z4Wj2Ax/LvekNJJWqpuwSq5EgWB3rm+cp9BbgYrIJxkXTIHTAfg2HJz97GsX
OvjX6UIC9nQ99KJ8KPEVmVy5bSEVKJHz0bWDakvD6dN2VarTVeXHC1ulOzjyeRdZ
B5DkuIcmhkO03Z4YBGXARqfo6b+z4WnwvqyjsicPSwq02tARJVDoDilQz02037QG
HQ7qmgOzg05D/+TFDpXi978I4SoRP/VqbeF/7SC+1NHRrKGMNRsu7GfaInsaZftY
uwTslOTyuXdTPxg4M7zvl7KKsYCO9mvrlltzmUavjvYGKpeFRCa6MYXxi9HEiEBZ
8PZG2FWmgZ09qUZexGV53cwrDciR7ftRjWfdBTfHg7Qx4X6Cpd8XTwrzNt7varEl
muWHgP2olsrUoYWxyLArne3pBlEaPQSzpRIOl2YsKlT8H9D/ZWLEDzaw2R8zxaMp
PHrF1FG/samQioBY1jaSjUN32y5Sms9V194xRGTZ3hKH91zwC0bMjvb550zSiwo6
PCJaQBrV1F5KUvX9F2a3Uo4i/OOW293ai9KzjPKe1ehnwJUIwP4Z7r7Zlcg4nLdD
L3IgrmfLwY3NP0iLFKGlWxHPTWNpP6WGNujVfJxa7wB0WlttoC0aglYJp/d2EUrE
6C+KPaE+w2GrKpEg51wcbMYka1IQdn1rBXO1xbT9L57VoP7yz19TjcQJD+nRUPnW
xs5yjyCivF5XxMVnRb8RLD4ANeOckm5eKl1qSg15TclAmEbkM9MSBKPLa6jQCx2M
HIV+2FEm0XOmIx6RliJXUWykjnPJzjrtHvuSrxSqD9c29e63S0BAtdq+PKkphq6y
eSCe/ralYD1Y70hdBGrTmpUIBwNHYRgV2e7TU27esINTmcjFncLqDdCzLO92OWUn
616kKFV6Ff2IMEMopLbjiwReebmGeNGyEOlQJYgNSN6bdUTiAyhEqzOB/lbkW0FE
kQEs4tRr0+BXb6tCKbhZAzTfqdSCF2VRxZSgWzYYYWhEi4qBR/mClXI5Q9PMXWJz
QmQf0eDrVg/oVqbm1rt7KiHqrPrlhKO60Q2j9bmQvzXYYLlgeP5F8PM8xVm32G1C
tk/U/7Uijjt16BjbNGpg5X3KJVzuHvQwWShmhkkSbTQ9PFg62cjCt+W1SP8iDh7A
takYJMtlERjHG3CvfXeu7Zl//iUkEOhXTvB7vm/dijM/DY2CdDIIMxUuR47HzfbR
2dP2smYwLAu/RPlr2oOnlVJASoQiuJgiR0/zKb42Hxkwq8PpckpZCNtwteOCCFzz
MaLXpHKXUYNXmd2XM5evuT0//vQAjTuG2x6kCkBdrwKntNZaF2Z8fnSDbPtXLwnJ
XpXqdJocvlBepTwWx5s5La+zv0vQKluugHnub0xguY+54aN0MwHFWAR64+Brbfe1
Tw7uawWda5ikFvM3amZ+q5unw31CUQGje5UCrZVdkoZvvVZCSTVWASlxf/9fWrGQ
ZP0/W9C5SNePuJR9YtqUcDPoHkJzo/KWtt7qo9fhShCa/zz0cyrfxq2uSVNioGmB
do3PJqrtcT6yWYqRs1GNPA+pJ0CFiXyR3l5pggXBrZ6P6JEqweaHUENC9xr5PHrW
kJuyXFn+jfgNm6VLyUPzWX9RWqaMW7nD7yGAxHFoDj6EcaJV65n/WRNE5tqg+O49
Ejvrh5RK3phi63R/xA+2nRqW3MilED9UokeS0UcZ6iaU3eAfeulc9RR9EVZ4wO5s
G7oNQVrsM51ItCI+NutmrK2+aOjnF5uXRMW8chfnkIP4VoyKz5MAYLMSjltk5kR7
OXl1UMUySrmoZejN4mnjBsoJTDolsThG1tnzJx8v3r1hTp7FMbEOD9LOOsZYl+dt
8QVvtUxCGdYWKdU50+sVA/0OxBHS6P7X0PdDfP/YRvHWF3kwUDA2kJDCcGbayj4I
vCw8DuWpxPShSZ97BTdtMN5dlmcI4DPLAtlbEiWaHFwDzwk1SI5n0WzrG9C6FcdO
jnZsmzsT7Cfr4lRKFnZatdEMyrO2hHCzX/uLTI+ay/Fwfqpaxg/wWS4R43/O86Gp
OoPUY09x1s8SPKi98aiCxaJwGb2sQDrNYF5ic/oyALaO/JZQmmc/z53uzH9fnqTb
ocZpPTUBmKJCe1fxSXwBbvEsSEqo0k+9vFg2X2xUJewmGejIJEIMrARmlcgH+78I
WASyJvsy10N3c9Fmx88qwfaDKq8G/mYOaYRy4VTugOsujpM1jGznrUkry/8sOSxD
Bnw0H1Jea1nI1giGMiIDdDxpJ0Gi8S2I9cRlwg7ZHt+QtHh1HSkOcYelz6xvl9+U
KGMe0EtcuL7iwyvfyxMrGen5No3K7PQUyd0UnJA1YuLTMkXl19zyNCL1meELd2NZ
izMmkxga7bSKc7IR3W6+GfjnB+fvuSdgbbB77CEDMMIltvaYaOuZLGDA8oqKj0Er
bA1U/GseqZ3CH6ayRKe/HtUQYFvJSC6EyAmTx0XCUlb83xCEQnJayY3dZXSxL9TI
aKGkpbt9/5YZXbWA9TkNk5VZB1tOhol/UKrZhI6elHgpUtdf8bunoEWsiQXlLji+
W6RcbL70dynyyySYwQHsmqGkFyVWdjE0Jrc/n+F1WVJSFOdX32orTrhjCCUxeIvq
YmXfVdj/ebP5YZPbCx/OI6JFLaN1Fekw42ZTHqpmDiwreR1J2eXVYn6DQlXmWGW0
QNvHBN5VfFrYXvDb6BLsnPIG/5BUfTMRQroPrlRH3P23PkAsxHJ1QCRBDIqsXCwy
2JyG0iDwvJTK2WIq26luq2UjdwgstJY2LnoDlXiH5Ar4l5nzmI+6eJHGFRI5lDuU
PnFFXXm3Wtsz6RZTFrxQ11qdzyVx39Xsg3egsHVH02hsUnI4O/DNXJ0PLG0OhJcD
EwTkCYoQA9U5enNCNTe85y/kjrWnu3opIYs3iD30f3F70o/SSiNGTjUK77UHve9z
k4je2q9TwZdoQQygLHMYJXjSp8jCVoe/WhMiEDM0nO4piksZB99yNJ+Uwtv4sVEE
25gIxtLvsXQ5d1daIm0bzrrjNL+rrV+x/qGSq9NXJcojwmC7UwsIUmN44pdb/Laa
2tGARW8pyP3+ceG1hY7kR5P+8MyrJiVGohc3koco8MxT2vt5282TWdxd1/dybYaq
l5JMczOJ1p5RhRkSb3hL6W0TFm+mLsrSsrimad/CveuJqID0BV2LTvs7Vbh19wHc
LaXBE5omLX7CaZin+LyQWrCWhk4sR0sjJRNMkpZyI+Bnhv51U23Lrp3kLuG+OdGr
8LwPmozSMUnuxUwA58Bn6hi1Sxdj1Fy0BDUhYi9H9sgk+4RQBQcFSDDa/PLWT8rr
OWuUsGM9rYqVoas4/Gvq72Y71EqqrdcL8atH+GrCXqBYpzFAIC09wUXqE/a//c2j
UbwBX0VCt5AhwT1RKQxJsI0ToiHbeSVG+panErlJXsAHQCuU0MCBO7CtZrDTQsdf
/ZSFE74kzl3e3iLebuykjxVMCP+g/qLB/DYAtWZkpWYl5Skk5HPsIhlPPp/IYIuz
iCmQQDw37T79rGWgF4Sne8Br96hALcLDqdaiV98PUDzPcSRCcbsS+Y5Cjb7z9gbN
U3lNqwJWaLtGV9oxGr3hwDISUabLSKLMoTrkksTBfwXcu2y4MQT6oSNpIYjtrvYy
aMuibLbu3KoDGM0N+kUK7VZCe+YwGc5gxKxvDA1p7HstTdhPxrC50nqp5u6V/fGN
536qnOLI3TxiSP4HvI0w9HK6hpiZ/PIZE5gdeZYFQlYUu7B1ihTRrcZdd7JXlCaC
BosR0mcMOUqzwMue2p00cw9GOz2Bne4JhVa4z5Xz/33PeLAT9W7abXNlTMEIRra+
prPf0c1qoIZWhHZJtp/wzDHPixKZkHAdhJEq1gVaGUVGvXQsMNoW7O7FYVAJYItq
n0GcavGfD2saAmW44OFyeNR5+bDdu1Ple9R7BqiiBQzp9pAuF2i6tOLpJD2WD2YG
apLRHuYdM0L6wVNJiGovS3qOtcA7Fpf8xP7cckdoyI8qSRgLNvQKjhhYbETZGQZF
CnOqsa29z9oWg9/zMsda2W4iul4oZKlth2FHL0hzfBN5JuJ5zHlUSkD0f5l2Hfj1
LrY9nk1N14DB61uhRHXWWdHdk/muNquxR3pZ6I5Wk+Hf1ZlIHlD621yq9gFmqlEr
0bpv6GIyV+8liNQrVV8QpL0NMLDNxTnfd6LZ+mjJn00hKn7ImHGduPe8oHtPeJX/
JfWZRrpA/BEdLkgqCsUnsTgfqpxzkFwat0Jfk+wr4HXaM0ugtRqtyon7gx3l/pTG
43PQ/7F4+9ZzGNMM6jaXmTFWJR6zmNnzUTUeBOJ/Z3osZD7/9PiPJWweEDoxdcw5
MqouIwZs2y7K1kAJe1T9CUWB43/ZgkGqR7fv4kVzXh4H2brgV0LpXIui1mNrw9bn
XSCkivjgIx1jA3St2c+E+qZgZVmWWddh4xX4SvqwZlHB8FbsnM+lG5yAjyHpuce9
Xy+vCD5qKBapxbfiPg+nYe4SxqRfpfeqHhrVhjN1w4fM7Fh/ZubT0NwvXI1Nl4r/
hnxFsl0lvyvja2RLC9yfB0v4uauo92We2pqtv/XhbFj/8ZRKdytKqY5U/+OUgAjN
Xwx8mEoIJulCnZpL5lOLzQnwveGbmi2sctLSmIpmvYoblL7zMP+mvHPyMrkHPrbn
Ap7q7hPPMrqfnanoWeispOw3YUKMtjaR6Uqv0YnqKqDycZdNs/Q1k5vdNANgW91z
4XwclTDeqk61qr7ivmmUzkBWy+YYcn4lQl6S0NTdzpW0JErDsRc9wR9bxefw1Ea3
7SRvixAAmrl04TxdJBRmmh+EiSCuPZu/LIDLm+W6E0wR3gP8n7l/IQOqggaaG77G
kd/C9o1WRGB4u9jYwh8d0Soz5HdF/SvK9Ou85gyqFizYy5yIedRRhjTAtAj+4e/x
LYX3Ree2AIkyPApHleeOXxJHBx6sRLgtrtSHEUuQUbGoU8RDAHSI5XbRAL1ygfV5
evOGfXthBM4Aps3WpnDU3PkhvtAYMEmv+wJAonBRbf9vpBrhPxuzZIm7O8Vkjddl
DacO+dyiaXz9JXbXy6aSpbavBZniDrv8uDQriM+UK+oomT7wG1/vtQzhYxPoIMgV
0bIALZOnTlxvZICnKCng3+1qoxAZp1pPlnsW8rwI7dGQxAm9MWwltqhwyapvqUwj
a6UYWedl68lU33BD8zTELXD0D1w6vutp23mIB2ArnphXlIWvSc9VBwaghbtpUAOW
ga6rBYmlwRAwrmQZAQySlMv0Y2o4EXSO2C7FeNpoLEyQXs/duEgbWeFgBmC05OiI
Lr9b/ubJ69gyxtenyjASLrELZMH/jV2M56kn83TyAGtPfz6xEUEQKyJOdix1XOLv
y93OHqTUzPC1ARFnm2r5+YF5iZkZg2O9AtGN1q2aYcZ/L0zwAKuwacGA1E6/G85X
eQpScWWNi+cshcTe64NqniWO29MinalE/O+jM8ahBno59NXORIlhEF/MG3Yj8VXF
65ApSdMXb4ZSrmYodpQH0oDhF7j3pxm5pZmOtHaj3jVoVwDiyLipD7/X5hZAnHr9
Mx50bkO5B7gTtAX4QhhATGU4GNt7+oUNJLI28Oyi70wFq1TXvgTcLXIL4LWfZSWG
sp+0mdhCJ7Y3YsARtraoke56LkxqslT7GxDtY35dGffyLi7kBdugUx+q6zKvg2Xh
0Mtpr79JKKRsIFFWyXhJlBFTb5a+agnDxCa0eBcsj9LEdF7IelKPrpID22A3ZLn4
1eziV3sdLCTV8gHJt+weHJdCoC0mDFqO79TlVMtfTqqBbqnUVqQ1P6OnRf/2JxJd
kArVk8j2jNn92/Q1T3rm89/0QBzlMPEc5wafqIZxv9MoVj48dn3D1bb4w/73amfV
IFcPqKR0rBVPOBirvBXPh7WxrNvrIt0XwAPK5F7nKZPdDYSVfWJHvGPx9JluaSRs
QhhQlF3SW4+dMGqLtzOPI+NV26cGh3gFvDGBJCIzStvHBpBipDLnfyR2hEjO3kpa
o2uo0jDdm8HPLLj8nX3WuT81p8DBbJdU+q+13wghW91YDJ/2BDisYvqQPfsa129X
aGR1pqZiPkiGPQg2V7gr/Q77cgFg4+ordnd/GiwgufOXR2U7YTcaZMwk4Q62dIOe
Djvj4TRHLYyFZmzz1DBw+5aEYfzOYXci1WEgSF0PEOdNUoiIgwXI+Rl1ZFPNXpmO
inlPZHSsp/V1IQH7EuhNyCQfn9fcC/CEq1t92sspKgFKduifxQc5Kejjltp3EcZL
IAyNRytitS8gsbQX3oz+1o2TZob2z21kSO/I8NNVYRQ3pAyzDP2mYDtOY1SFgD1Y
EU9hpofb1cW8SSM6sYDBpaD+HWj2KQaa6+tatM/5eub11lcNZKX8dqKhXCazmKWw
G0jmXC+zphtFSFS2mGY2vX8M+blNGh7uuEFhUPogU8p/jTK1IaMZ3Z0AlNEKQBiy
6ysir6lkk+ZhvkLsKFXFCXLW3BtWDxEs22NNngd4fWmfsmy0AEyMLazqLaAdPPbz
gh9sXSqXVbWZRqClhNRnCpd0NgiU67exlQkHV/hLL8CRXdZGUeDI1vLLvV/ZcPqj
BgIHrrXMi94VNLNn/YcOvoirOb7kdr59AMkC4E1rHESJrG7IKCzzJNqPOhHRPWX2
jYucsPSlJ8R9YaZ/pnc1dHFJSdVYvwRs73lJroS+yZ8eFKNFtXxYa0o8Mnnj8ABm
21XepaQ7WDKnI6ROPinmwCOQFEZUg+oHvqUkFfmLv57+RXNloqphXqGhg3aFqloP
nM+niLOJJvRUC7bzM9fefzZhxlUmLM+NRT7LLf+G+t9furyH3zqQTgvFlC/Kx+Lc
XLcRNwUP6BTtIH+WiTVi5+FShirOIue4kIFvBVlL5siM0oy2y/ojEa0Gf03AJEaH
hE8Qu+7Bm6HXbuc8ajaJqkA5IuJ6dN2+3iXxu3N1PWC+zd5h4neuzhZobswc1geS
2vhLDethYQBinZ/TNjhZxHpNX932kYtNHrzMPJXwN2ZJjPX4WYcrF2nINuuq0xSA
PeLZ5gckzo7sgrNkGT9CDFxTFHtTXO6zVPCARvcZRtEO0TxDH+nSHcCkiaYf3tqV
58s5lU1pRs9axiB2jw0K7UN9keR2j9vFauhQuYZINP7Z4Y4YidkFyJLyT2FLUWk7
Bu5IBGBPmCVw3CEHHLkPIXjXjQy25xkqWQEJEsZBTexnVlz64Gajeh82IsQZavyA
FvrSJSrueDm545RjKQqn1ImiCCxW04F3hVaUKxKIzoOn2yhSiDfLmqxvH9tQKIRC
GtBMcockA0IuviMJkXHcBLdneebklA/rxy31yU+M93uh9190oJ8QBjT1zvf7rzyn
QY1RRp8iW27jBvmgh4rPkSjFbP/XNNUUbmFoFFIHkYj66fBazE6EwBx8wClKZI3y
c3cOi42Nzz4B3rULkJMkaxwzoviDDp49GDxDJg10NSlyKlZE6EyP/3SbOcINGpdO
wP5LmGx5vXPa1jpfhx6WvAlecL1IErN0cHADoqP3kNJ17BjG1PxRI7NLe+efmIjY
AI8mW55HSui0GC+1qZVsW17H47D1NbUmW5uwfA5w9xLUjli7gzTZwFDm7UZbWocu
hJeKR/7djROd61Ng4QSwVgLjb25mliHbxP/hWDmozx1ESyRX9VmwgwZcbTCBqsXq
axKVTlIkq5+/Se21RANN5z2oTl/wBv1NJrr6FMchLlizZxqrwuwDzZ/jMImXVx8b
LLt8FVFSPlOSl6X3NWaI5+SuBqYusDuiekpI/Efy7vMI5pCffklvhRtR1EL8prtj
9HXF0aFYiIORSZTGVGa20BS61m7lJGFc0v+SD5n5B9vbE7rV8qOAmUIg1dYUmWO/
HteEyCPpRMN+olUjxeCdLRcKUOsQHQ3LwzIH3lfBEDdkJDW2f2S8utB/KJhb6aBR
NayvxtqR2p8z6duJtpB1jSfUBAR/sFFOcW7f5gKyE4zg8w6TQBP2nn2ekNCOAwPh
VaWVn0tMpqbk3G46SqCm8sgyIAn2PVGcB5Rtn3xAPJBqaQ678O4t4jC9+v9Reimp
10EZ23BT3CmhpQTEaeGvAn2fcCpltQxMga82NPFxj/n5RTQptS6mCdXYPxlmjMM8
vAoOqkt599KwPZTBKn6qh9H/TPCyX7wbKljef/ppIG99bqCrzHM/GkQVLJHLyG+O
cCkqg/6H9RGB9s5SDORYqcR6iQnu4LbCOn6vR0YxkQk/+Faj+zclZCr8bYBuh74s
DSirC9OBcfU6KkR7asFZZjPTa4ds6L5C8jBmrCRjWPkIqUzxWY7xA275Z8uWut7F
DFymfuPFiZYZoVjlDVpfTlq+V8wf7FSxzloF0sK3eKS9hjCslboUfYPlJ3g5PbDB
OHhHAhpUaFzql67/RJ9Aw7DoExgKueNyZgIIzwAUmKpEz3L9RKkWq7x0eGREpiD4
4OmIbW2SQNGhti3xgRBdvkwnVHlbZ6twn6CdyjHNiBFvD5HsavQum/R2PI0StzDm
Xn0CU+ib8FhfUJy25dIs3TC1o3htETFrddYrnKTa0gmWJmrku0QOO7giSc0+BDkj
J8hXWeUPzRP33PajaWGuzF81TJpOhOdRPpqoawsSRtjdl9zBv9tQAZLVfpCj6X8z
GCoveRUcJtqLRFLrIeRjAIzrOlz2vVi9u0HfjIKoa/xVMAR7aEePWLHnCNEbRVrK
BS3m4PeY9ahwSuJjo87z6TmjGpan+i888IPgjmeRclgXZVNo8+RzIfJFTGM1xUWF
Qq7FSOlYAJCnd/J8MBrbs9d+o84+wi90nVqlL7X0Q/003zG/5ZY1FXcCYNE172Er
NafJP7qCMYpln7TFQufoiaYbhabYc5Wgr89RT+oXtr6oi0WYgv+17lHgyAhlQWWn
B1ryHW0pURAkInDy6yl5PkOIvHVRbnBFAwXT5wVKMXC74a+2kxoRjxDTEQFiUkrq
uErevjpysk1o3YRlf+uzDtPvWLPE4gOfkqM5lbMguw08HY5pbMqCoFaL2mlVV8Ci
NiY9PGMU/1FnGBEeqMxio8Pby1dJVGKryS37eqBS+MA4L1lUyiALqehrBdVcQgpt
/3W65TREri0wJYh2EZMiMu4vzs5cxe/ubyDqrkDjwHmW+U0OPwFSrAoE4F+sYweJ
B5FIwj7Iu8j5S29P0jxMCKBxCIiKi4vLyAl8k80zUq3KmFXMaedhtMeP0Br+H1XS
8UuapWE86cC0nrrSTWrmh6DRShCs/3sacbz89KBUQNknZpiFSRqMdNsmkJH6bdM2
LF/j7kefZiFxddgpa+TJ5WwVsoltiMioGWVKi2hj9Zx8QxrmzLThaK83ZiATuJNW
U6MRq2mHBy7/vx7u2uIcH5PdzheY+WG6tjG1Uy4ghvZz1ZnqhNf5mZ+I+KKHYK+j
nrlyxsilqM/YCc/k8eSLQEFSF/qM/+ZwTKzXEc38RZEG8HA6KfHsWaxP4SSSgEZC
Zq8hdATQW5lGRwgK36BAO15d7DrP6AB2m6iDwct3qjLySsPtMNWR7OoxUSVprUTN
t4oEp7BTlJ1MYs5e696vbaJwrZ9MaL4h+T/4NNL9EwEX6PAtQnKq+M3S1lsy0VHA
uqqzUtwGvZlCOs0lHUe8DI9a2dHf8mWgT8U2LJRmYlAFATbi65fg0veoJSDIMK3g
7hTMUqjYjV3k/TMbet92248JMNOw0KAg3zAGKd14zsdoYkHwZzB7+HvV1qkZtA7i
tCzanhe8Yd7zambUk0bAPuay0MkcllRDCwU8+am+STTk+DQviKzkilwtFidx1ECa
teDh7LPrE04PTBfZGE1npTLZHJohYCLjERb+gBivjJipumLxk1FYVpX4PTU+9NaI
w+IyAsxXvSFKWSd80ouYozy18Vi30fOv0fh+MZzVnK0k0UXkWoKjXLJNCe7P9vZj
nwaWVyMSAMryRmZ9ubar8R+KYioZvnFtdfdjzvN0xagsTasocOsCS2+y0pf+aiyL
V7x90bp6wZ19mAEmfoAVTuiZCW0n61vG1SfDmcoh1sKsuyTYpZkGDqnDYRStSVdy
fjMT+HpA1KfgpGVTG4IF/S8GTQ3y+6AhOXZLzECr0H4G90gHTKxOHCzz2TM3kKFo
XotnVpYa4+7xVy6+Nj9YQ7JDnmrGlSIRKdRKXgWcoTMWTo7jqjPU7tB89vaQvE3n
d2T4vWYtHm1CMvbZ4uHrfGdvZSZ50qONsUMeIyiav1AdJbxLhzT+9aSjYBstWOxU
7G17dQxrGNtDbqWW3Gqo98XVmAKGcG0fkI90Mt1UXoIzAe67ADw0ZMUWbZsLzFnB
xevz6eQsVSgcdF4yEnemVbDK0KBE4uPDNf0BnxtjvaVusvPj5ZPx7ENaEKDgxPZM
M6FAXp+f/MdbH2vUDV7mW/+hDiyItPw0kXqdScDFDw9yka/ITEVRctG4EHh5AD51
AcBnwufKDA/zQi9PF2UAclisVf2nERVWvfp43Y7188wOGW7os4+jNmzOxEIoGIo2
ecBWXGpwrw3A5dyigzsqCrQvrMTfdNiGxnSekuCPovV38Ebt4aRYi4U7y0g9trEt
smo49G0GROaZMEai2gvU2hh749l2LRLkGEQDL4AXolkxUykSKMROP4VzB7xMx4G8
YMlOhSXzW+PUprNq/lJkEbjPRT8Hw3qB283A33FxjbGUbYw0et2t1Z740txM7VQ0
g/RzfUhFHwYzdFw1Zg/wXN3H6+zwbEPljiy4wWMgSVBIlRkM5FyRphPlebGiyi7Z
VpgtYv4naCz2XqdFY6qwY1igMiRNMn8vfZMknc2WnU06e5MvQq0YSJmQOru3R4Uk
9vJYX+No2ksIllac850g8K9KCApppMXvulAQv1nu7xyZd+ds3WxatYwILJx6Olr8
j0A8p1YL6XYzYFhKOtHlkUWwN6EB8LVsjn6u3DiPk6iEKiny33ulVnwCKcadv+4R
2uUElE/3CCU0skHNoqEG7A42CrGEmBNNNTIL+mi2ZEEDSzbTnEYVeGOyFSKx/qF6
WSfhUxY8oZuctewLuQaigpADCtnbH/GTTUdqBCit2p0VwAafdZX0LjAAlDuhvKFe
K0b4CQ6QAn0ZIXv8oQy3hfeU3ULTXqMXz25Nlkkaax7hzKieZqdl/w/rGcewN6JQ
GxilO3eWgS1b22oqOFdITZP6fIQSQmwmUxKoUamOMo2av8grLr+WBNAQqcrXwXCP
vk0dxPHG1txr/ZEGDNGX/h7tdkt1h7bBdlNxTrR6Jrk2CSzlTldHvM7SkfLkHXX0
76Gxb2Gt512eEd+mQ6kAfg7N4HhHUNv2J5z9Wacb36c4Jg/+tWOpfPZfQxQnnbiC
qwuo+Mq8IXik47BB1PZzKIeg/BwcrNo+89sgUQ85jt9Y8wJ4EXN4gH8/8YnrB31I
ESx67k+f4CKq1cDEyDQUZNSC/7/bTr2gewCyH+RVVQs0pvguTan41UFXpPIV17nZ
UYsBW4QgQkEg9A+68y/Ysfi9LI4yLZxl7UPHQLbW7SmRnK2kAWK71MFZgozGaCaG
XdvPvrauyZYn+T+Z5k3JU+B61Rumm9ldV/hvvIrS9TEAPCEEpuItIyeqA4fNknad
qZFKJqjojphXMcq5WYBGHPiWhKzJCO8wSlXZONrP889v2Em6+ifii1NZtbzBcePy
ZAFku+q/Plxe+5jkPN0KulKWqt7I2aQqaDeHUjzW3jjBXvU8H9Mi2RZJQnjOPJ5I
XRopHGis5YIefT8Fmea8i5LAIUN76CZ59Zt/Q7UVaQWwG6XaN48tGtdCV3VIJjma
cbCJqzN9GovbENuPnldPk3LdUywTKaE99B5EPj0t5jdaX46kX+uORK3jq+so9Xyx
kP9PswjbGj8s95Gd3yhmczE6ZADPPaQLbBJY6wLqnPJooqJBDHVWmvR+hXnQ0em/
czK4JtStSbjYzcFbIwKg0EaAbmy++lTcAWKUf9dEpat2LDr5HaYc6oNgCF7TncYj
4LmF88OrErqpQnmdpZWxF8nThT5zlzTIRLw6WmyaTx9mKcolICFrMZyBQFdw/Hcj
SAlILVyieNtwas6yZCalzZWcyXmU9vFMBC4gnU1/8NGxwr+G4p0mRFazwESjZd4w
Arxj5F9QybQ8VviC6CZbwXPDvzvK8s21bNIAXf0eIZHybZ8RbrVC8atbdVcbi51v
SuZYqJkjzZE9ivvONGMsQaeBx/Pr9N3Mc4brK+qd230xMhfQa4bR9tSu8A4uGyKN
eHynuMBpcjgwp7j8BsD5y9neJ6S5xiItbL30gXaGuKOdd0H7I6/esAZPgsoDYH5A
mOX2/qJPhEYLKt6A31APhRC2kpAsyqp54Gg6eRVnf7f4pQTMgh1kv8DvBcWmsmxG
sSHxXPUMKFhfjkFHU+A1Rnxze2aOLcDD8uLHAI6a3kDya7yoUs6XyvyJsZumeSCj
3utiooLt+i3bAJ/8tzK4g/U65IzrUIT7UXh8EyvALVGn1IxBCcMSTHIVf8LvTr1B
3Ur1zkeykT+5CJSHV0H1WgD+TVxkcDaydV9eEpysLY95mQbt9PYaeclGdqQQf5UM
cStcJdwQ8aB9TROHn6h3pQ+usk5Iy+xFSXVZRZNkcmVxS/7waG28/IYYTSCK8ZpQ
ULDk6ero1g0xfOfaTTXCgMLrV19JJg9QMdTgKraLalBxhbyuL8HmKyoXZ/hVwij9
zps6o5tA+nfXrdyfNx7wZeAxR1ZmowYkavrWC7iq88KYeK1dgB6RSe5V3ogdur2N
1q3bb9XgZkOW1/Rd+VFfk7zo371tvxi3+XvIMvI6XgqHCwdPQc6SbZ7IE81Z6WwC
YLoUioHjOJEdojW5AKXCXrakU3ahHblXJyCOH2uqJkozF33ikHpWCm+pnY52t1ow
wuvMqLxx5JZYEsidokW3R8nMsVDwICzWWE+/vHdPrasRmy/DG15NVZS7Zw4RVTf9
uNnJaI5I8zffodBrOAcvnSZw8D5Cq4bX/SPta1BHMwcY4OzwXA1UlitoWa4dMt59
I8Z4AIgebAB5yOd/aGkm/Jaa0bu/g1StO97TrAvbY1f7h5UujOfBf4r/OwGKZOon
Hnm/zGGpBlr0B/n+BVIEupTkuufAS+VdTz0dDSOxIGbmeAVFxf4A6jJnVg+SxAOm
p8YRP6q1yQv+BvwWN3VLIGI9iC1EpsfXSnsG30kRi1Ate0W0kgT2Pv7xh8g98JYS
NTlvElYWKNLjv+kLE7ubIdMSSwf604U0SvqYYz8Z16BwGj4HzDnjIxtN7UgXIZ0+
yW8bQeHRB3EH8Y3y0p0qQEzDgkSieAwQF84PHOPX8ZDHv9JFo6rhG8JOTZwyxBvL
u1Yskag7H7Hqn6K99wJobDT1cyXXRmj2ApWib1rcJOCHymPPlg6sfvWayclKEW3+
hWvwQJpNAyDCqQCVHwOtz9kd/GZGFpU1LOr19zA+V8wxDT3FnpyrFODQVXYFoJpD
t+3weuq9fUOAblJSh//g5OLCk9iAaEIpg5agquMRJA0Xw0N8+y9Q7l13BKjhIrQ2
n5qlwIpWrSA+OHuB5bi3xdKMRMK03oBD4tpr5wm29o4xkvj3gNxA8RZbfwCIIlRi
9dnnSOtyjKLIiW4V37VqjmAoPmNQFu6PFunbEtARa6GTrZjBE/fhUtX6Tvw6DhT/
LGtUxg8LspxE63LsOFuech2yizHOW0Dev6LMyrDIgvk6OB0fTWTdy64oTEijpSGP
0eP/RWLryBn/cIcJnAOu9c+2gD6TcYKieyYVMmBXenzD00jiL1dHFHnAfpQSBwCs
dUNqH3pOzVB64Ltg3nP5QG12+JkfjFidgTJi4lPpu6Jo/NCBSgvsiez0qQFzW3sS
rgCrmApRIiGwvRZj7aRceTqMXQOQwb5dQ2XLvHZOl5BdcNISLe5vw8XiIlumt+6H
hMmWCiaX/6JKjSzMIWEf4VwpnfJFjyteqxgO9pqT8DoTxBI+DNMnIyC+tb0wuHuN
KBSrRnWoZhEkAVI6mYzs/wIh13i8PVWf8441UDwnb++BrBzU10fqo6GnfXwDWAKz
yw/PhDajujaP0eiv0f/rLLt6eTIytr4+7fRurf1Tmrosln51GXYGloDkvpjk1wsM
Ca8l6Kbih4tKBdxcf+xVUYR4K6+Pvzl2QHbLT7rSwZDnMVTLjtA1QqLM5dSLVZwX
0MqPHCkrFH99qHsSTl8yI9Yeed5WhFiYVB4daG45dbRudrjr/SWZF3ykzV+1zheJ
UP3IlRiSuXEGVChoKLq1ryWTI6tN1PEqI/5Ke7sR+a/AgjNxzTASRQIYab6nFUYn
VdHdEdhsADRRBWFYkCB9Pu/E/9syhC2JJ9bDHbh7pAft1NQ3dCLs7LzvITXLMdDg
xj+4/xm2HiV2DOwlU3BbWOxBI1YXQ7TE7XXkp4orZzHwU+7AmrbKUX7e9trgPnGa
zOOMeyTEmloaagvcVmUJMMCQnVx0qgP4y4XaLbeLlOm21RUVF7Hd7i5eZu1dR5oT
I6B0+icCDuogyG5QudFKCA922TjST2sjIMOWK55gsjINjisISpZ7lDBCtT1iRU9o
WAeHz1VD4eobgTI1dvXuecA06q1DMFalbweED4+PHJoaqSDXb2tDJ4Fs3xZUSFoA
FPnnHI9T2BQ0X1+oSXdqYeEfDPYnSHp5Y4CPei/sHjAgaXWMupa69uBDbOaGeMqT
ptKP3A/Byv+EEnh+iWU/ZYej/x7z16gauaK6QKyNGRTbi+ZmhuhsCu50qxhsH2cj
02Io1TygLvx6JvrLHOnz+vquVFrroZ8QbSAAxGcOTGNEdv47NFtxC1RcJc5zhtGV
vOb50MZVMMVePFgambwkQGiIPbrV6IBG8rubi+qx6+HUtZD4IcQ9+JC6fCRDTjRY
jpAiq+RFv7FcK0aKDJQ+sZ1H+ADw2fVPyMKlxVDDzRCHipQPjGhKRrvgKf1Oool/
F/7kMfDJZvxRU9Ti/Jld6eWnAx2eX2v+GcAn1qol61NcqJl8sKyTNuj3UuFx8TKF
3JcN3UIcB38s4cOXYlAXAC9yZX50k0xFAuyjtpf2M/hXI1X/pqI2rNrnB7u63z0U
G4zKmriFZFFO5jCp4fymq78J3E/re3k+ZD96GTCKT0gmPVvwKeFmZLMrv3Miarpa
P+GjyBaCJ6NFRUMwNe/a2stjeN9gFZVRt7nLHLZeY6v4LEgU39uOA9f/N7qlDg7W
63aRnmghGyxUnK6DLGbxHyL/DjpVup/UyAbZ6/Yrp9a6fIJgFRkiZ/Xyu19GpdfB
lrQ46Iu7vLfP80+FCuUZdv0DXtCr8zReOL7OgpOotJBBOaZih+ozoYBp53dKaE0T
Q+A+Ae90Lvo5UOotcEtAH7tRPb/glKNsRZtrM3I6zNw6yVfca791rrV7/DWKCLsQ
wmKMt8lkeFV7eZK5TMZ7IVcZE8KYJ8dxU3CKBI5eYKdJcOxRy+dPMlw+iuxo5AtZ
+wRwgpcT14Tyfwg/Lkb2mC+/2IwiVY660KUFp+3HXeONi0XeAOjVZTmBRj6lN3Up
1siU32GcwQ6j4CqGgMY2gLlRgLnA7BLHgDzMgE40hNLdqfmZzTxD5wPwIFsstFG8
uPlz524UlOwDl5rha1g9pFyv9oDYTMt1oREfmJ0wwFNRNxNKYKUjxAaQ7Wk7CdHz
iCrkwgeajokYW2+vxiPlvWRQytSsf2jvmhMJXaVBaW1AmPlh2yZ9uVAhWb3i7n22
/fRZjpm35V1LNP7NeqiEAIaGkCnmW6JkmcqBS6Ta1CpdOl2LmpuzIU6fRa0d+aYf
/qki1vFPRmnXYz+7G52AiRU+Lt+QRdBxZvZoQ9KsoEYlQl0rAPzP/ZvNC1HJ4wMT
3ZmhJJge+6E0+trv7ZQRQDUCBuQNdSxFfpI9YJEoXxSdwprYgu+QfLS8j5Gu5BNW
uPxdGUOVRZk1ZGj68+/VCBrqBc/ULP0euGviYnKI9xLBXyor0JO6DnoIyyTbsoIJ
q6hLOZdceK2OKJ0Xsu6uEZ396hlpyNMoJ+RsSVyYmwveb7bqUbi75shIVOligPVX
/+Th6rcvJp5i4FUDTcGN8MB9CNq8HrZsHLW2Mtar+rSLus3BfgomAa/cc6OukYEC
eXSdK0tmgDnaiMvNxh/J+RvdR8+yJd8RvPVq5mutSiQF/j6TCOm8JdYiap5oTHIz
4zxN1TUnPckuAcByOLU9ZWSWeMlbwOXS7zYlopnqMKybEVtL3YjcWG2tDCJ1TZoZ
LQeHrIXsgh7DQDFXVFUAcZiCOI5ga4qgScXPCxwFWbdli+LKpzrk66Mq4usC+a4Z
6HLP1YKIefLwZkxAtiTOfP2q1pT/+HFDOmsdQUzmoJFAQHXMenqEm168SDcgzbKb
UIhQsfkhUS9JG8oSJ4giKjCGXyjkh9CerrA7WWNkZSP+v6s7W19FBr/ZgZPXxrnJ
QsR07/XOq0ZFDrZywApDHe0FrZqlMs5I2qSkqL57NAVciZ6hyDw7lw78QACVGSbN
yKvxTYx3yhdUMvXWA+WPfbwZBQDCKfxydvv9pdp3IMJsNLInSi6U8ZBMGgkTqdo2
e7J88r5ouXXMIFoAAjfpdM+pw2el4ui1ra3KXpRvalG0bbgKOQFNAUUUWr7XmqP+
CqSunPYguLOkI86Ezhzffki2/JWlGM7PZRijHgsOZ00xT6/tpIEvOWe3b3IQtCEP
kjHCql7XUylmwyJQUiy404l/z8cJpz0td6McZeBzu90DYKtH1QPqxiykgTSvw1sh
WlBAtMKjL7p7kNJiSkK/z7fNKBmmDPcacCv0ZwhEoG/BhDmiJP7tm70LrErbLWZJ
zN0IfrzDkddGOS5DOfOSiuNL4gleMortb7uV5/MOIaF4cRdLn+aOzQpwmyNSR4te
2ij3dNuNlbltbfpqCst1BK3BNVgA2rjdn41e/ViBg1AIhT1vrw6jBbeQ6TmEZyhF
HTUlIriHzCSTH8goBN2w3fTcEDnUswHRnkRrh+7LMSXzUaXayLWPkImmso/Xqre5
jTBBEdaxg5aEdxuannKPEorVSnIIsuozMgXh4I9aBLnOqwKgj4U0vvUj+Jul3BFW
68jBhYXb7kF0Ie8aa75987JNHwLMuIB4J9giZrnGOoOxeAZgLN7COUf5GhIi6TE3
3q7bz43DTavMv0/qEEFC2649ZXWsr8g8Mg9UngB3pQNRv/adqZFl1armzdWFbB3M
z9qgmPw72kawQ7KvbH5JulLhV3RH1rGHmIjXLD/dRxJ74zK9D5MpXk9BWeQ9+ey4
59xdkjMPN8C1bgeDWcMWeAQfve5JMYfNTtga0OR2CoMoeMGtOIMGfqca0WCIhhya
jDvupiJ72lgGzHvfSA6bbNzg31pyjFWfB6OgyDqt5HVg1fj2VzX78c0tZemlZnWU
wFLw/Ro6aZwILRx7kosXFxpRgJGHeDaH9DSFHA59Dh8oQpaTBqsVIkUdJ00HnP+q
gP9GErag+FHNq4lJ2ciD6DnTeDWNcGwfm5PQI0f81K4rzwSxEfoa/lBFqNSyQ9RR
1EWy4RVA8UjudP7jy0o1gzCX1b5D2y3qgcoPhC+SdlJN0j4EMiOmJMjTQtiMf8bX
SeO5Tha8JSZ95nGN0xH1FhfSGxctdUBM01vtFbZy1vyyR+opAiBEE0VzgUJ584Gr
TGXAh12EYWFNVxqHFiqLzTgmzM5o3cPvhhfxdWaE+cGKvgBhoxp29gzEeRyvSJuX
KV2yTA3btM4voC8QxPm90VeOmwuwxjMY0snP1aNyr38uPT1G73sc5jN//gkxFn52
emioScReKa82iyCEjyNoU2+tTCCbS5rhp+ma9R7HIPKZ8jMkkRvKRhpUf54ERyil
9J4pAhSJKvT3Pl2+/mqjjsjHIVH08emkIqtXyr6ipo3CjUoKRLN/au9PK3YbqJpe
/FwhLkWwKutSg97HXa2ExtATBWGwY7efmdMWJ+dTTQw9g5r57XEZOmo+gFz41h1O
C4qiElzS7Y8NZ0HwLDsfiKfkUMq4KoI67G5VPfpsoPpwpnMD091az6GBZv4sqyMB
gbIn1w+sFc733XLDJ+ZEKGtlWD1zWaWOAjs1Q6bO8RxnYcGrPmi3IZQpTxTCHCxO
X7uBa9XjaZv/3uUtwkdAMDcqxi2EWlzz30pLQGKk7fum8r0A6UYJWIJyI/+VtKMm
+V0AAkjP6aebbRwjlP7ErDwYRXeNjq2LXuEzqLoYvQKLnNNDpeZ4MKqAHxziuQDF
/bESnWnXXDpZuIo4ML2+Ao+zWzbbKLqPgY5p0dYa/6KgU7mK3AosAO9Esd1bI31Z
3nkQid3zRSZVoGIP0RrZGGw7tVZ6NOpqLkKk0l5pvN/3KOgSsRBdnim2DDVVNNAr
BRm9iyRRc/UlRNJYNuu7Et0uybIIHWlllARs6gj3eIMTujrS0/ZJPey9n9NVdHCh
eJSyDq3C9vE/XC28iIxfnXeSePNEccJH01yEDeZKEFbPxwYrbKaMUUiWyjoyc2/W
fVXCNEqrYr4h2yT7s84DGmGEgKcNoAs6p7870bRGLE5Bd4k6UIYF0oJhkEuEMTQn
yBy7cg7dUxHqZSHSmu3lVPNT8DRWmcijqYzqcHc1T0Ar3EYEwvE9c3Hihf5dliry
uzAJcQhnhlFm0uq6IjH/FmcEnmGIb0qN7aj9yX206zKM+1/zcN9KH8MjcncK7yGk
gxaCL98Xe/DP+LbtE/TfItKjNRrh/IVN9inV/JF07xtHRK9Pali+OQsYVYVMEUFI
VrzqkfOBuV08kuhcHS6wcXGlDJCCwn96QpQBcLuXExhN8lDr31S1bWHJH2YdJyAW
rVfEAinkE8bY4fsPtWBRDmbOHPlq4A8SjWyqdaHZI0Z5yjZ2TC3Fa0G2YowBK/Xg
TKJEXyGiR8yr3ri0hZJbE4KY7OXNB5hLPaycJrWjP7n1SLiwZW3ZSwkoFSRvDw+/
NjGmAwS5HzzBPYfn7Y8gh1SLsbDdGxm/unuhhwymv3CsxjgOgfsCRkPwKoFxiSE1
uBK/2nIJLaMxoUJ+p6KVXACi2e0OZ9JItOsc+ZOO6jhkuSV/W0WSoJD11MVX7ybR
umuYth85xDLekqs/sMmIPFWf9VeTrdB53VA0bcTqXKrqFKk0WHeFDRBS9xrMqIjA
pjMTXQp+Xk9Bd5F2YiE1DVEt/0/drU/bWTcyU1xYyzGQNfWgej89U+aCx49I+spR
eZJehIE3qJ5Iax6V/+ZKEX+dLOyA7tVpRbzvikVnAg2XogoysTX7j6xGKOSAJlKY
K3UmmZYc33uPYwzlKT6p85ME+oZ1jBSwTNoOZExLf/HDpE0yjWs1ih0E76TUfq0j
+RquOwaRh68D3afRl/poSmVvj2y8jrsHac+mVaw7Myb01JQvuE0pIn1wvfMeOHI7
xmk+D2TeQ4xqf1L2sUG0q2tmv3kZfm41AVpyiknwhuWmWmU3SWs50htIdzaMZOtG
PM3SiQDyDKJwLVdPqBI7qy37TFWjRYO0eTZd7G1wNndnGVKT7L1EDUniqaMJRX6N
TuUwMpY9zLEWsEB3Eis980K1GLlQ2YR/R2TWBh22yoL4IWckRnW+jbVzltG8uBJh
lrpnaUbRWWDinrONI+kuJZmU0q1vEhC7Vjtbc94JgD1OLCs4TtTe9iL7mFlyNLB3
JaOSBnm/cIVtfldJL6bpQYVb9JKRyqqHKunXQqFASyCkIBA0Q6hHOoRmNM0+oZ3V
kMo4h2KBb7DRzZ0OBDbX6GJipHRrNXu3UZt4XZs+elqjzERjYfHZ6u30Xsn3JTuS
aB27HZIOuxBF19JtO/2vkQS6R3v1WowDVLkZN8zyD29TOjkYDS5tXvYWgvchVf+V
gI8rPNSoXZNR1p9OZUVMuppaSOC2rrRTBPxoanJ3mWrKPmcuAea86Te4jRMG3t8F
kXEtv0WCPEcIpFFL5WiHU+x6HPTIgxBnxyCrWnjnLs2cTd1nH3Y/4fX3b5tMuI4q
IgG6zG3dJ9zkGRw5/fauEHK8vISoouYXC3IU5cs0NekYnyCSR/gYItkQJGKswRma
UBTr0OfwO+IWwAGlF59+VaoLypGB6hO5OBF8w3WazjZd0a2E9X7hHTqKW6mRZ7Yd
WoFz2FN5zGJDSyEgb5DM6gFoFZ76DgrwDkvWUKleug7HdmIi/RmkSFsnRQlzacfA
mDVG5CLPrgElZq7v3ku0/2imz0Ch/2UomzG/GIvVNOi0+la3lzh1nR8DURbB+bWd
igv2kDK2aJ2tvcEPSciF6KkIjtK9yujH26VYEk7sPhl4IxKA+RXqpVzQK6CnCUFY
nzDU3mJy8sl47pL0jtmgQnfMYkbJDtOnBgdndQX1/SJ1w5fDZyAO8Ofw/YJgZJYQ
Pq6CQTYGxtRFq6y2lUQEzD2cKVTt1onw0tDwtRVwiNFgs6LIkOsEPLa9p5b0u0ji
X2ckg+SjtRy0MznG5ppAHCjYK9fGgDoS+yOL6qvwJoYJK9+cHq9wx+X13DRDZKa6
oDQK9AX980kuKhXdCph1E94q0Lx/ejAeLvSwzhwvNEyN5YQsFkekGXg2fnhf+b/U
hv2ab79/PLfCCWvDT9hnfvn6D5XWsH8uAxCLhj+MBF9urJzJ2gRDul3OWp2a0PSi
JoPmEE83QDdkR2kYyLuwF1Efh/MQb3G5eNsi6UgqBzKAqHf/Y4F4pG2dPczHmYlO
tLaVPGrcbZd+hdLGxlWWIikJ+h4Mp9NvHk8Pss1iYxaCCPMqmGbu7iGkICBvVhv1
jiC5hENubtvM1bfmsxnyjK5Lzpos/8k78THM4/t6NjIOhftfGtAG7M07j2h/yq5J
kb3UG+TDUsTDaOGgDvLa/JvFtVXg68iiZBfDEyNSralK/rVvrUS+R9on2Yj/765/
lF38ugfil+KNYcVcnkUxekfOpYr+dNcl+rbLL/+KASk6sKR2HLgwnE2h1I/RpoKV
yvjUXJ6AlrV6+OWuLnBBIxLJDovP6UkXI3ZDKssnPX54E0V6SxNitaabdxIDK30O
FFDkgW3U6CfpYbx8VS/scj/aLl4BaDUQhAwlo5srMS4WTBcqM0cjN+BsaLcvltiJ
ufzQSN4YE0iCrVJAg3BoUcR+CJCYTHUvnQ1y+hYJRYF03rtlicah72Euh8sliHWm
kClUciEUOWJJ+rn1JHlwZxEiFrxNHahpDFX45I1WKACcK2CTfVU9AS967KDHzz8e
QEqnAomSMfwOmSpcZ8RLIdhlU8fzzYGqqnLrwUJa0JLpunU6J4/yJc+CqWlAEuzb
pOLh3uMXXB3n9jwNbEXBFqOgfKOM3jK9s8jbN4H8lSO1gboMgNANgQC4a7Q+6ThK
WJlPMC86gxSGCb1MEcjseRudz4Bobocao4VbM/L7ZvyAGtCUcEfCT4QU+Y7edXYS
L83ScFLGGqp2OSZYPuqMj050J6BBQxx7Hcy/vdvyFujr1JsY6BfXmy9yykFZ4ZAH
PqGGxo9HHP2H7pFWrvNRofiL2tJTfINzu/O6Nalchvk72B2WHBDZLywdc+knY+v2
NI/BolzvGQP4huSQ4CjtgTMnDNT4/iapqaUuaW0mYp33aItCDaafottOpfPwCAa7
UsD2Kdf+9D30Z/X1d6xy9CSYKPYa8GX/drGgUlbisPCsynO/CAyU3v3BbBTTa2Ms
Hr8jTN91qB6Ag8izOhYQg9m4n5gC1ONp4B7hh6lJ4Iv5IhjI3g2KvDr0UGNi/6HA
YlPDDB+WR/IWfEONp85Ib0vgOzHg2i5RbpF+hXPxT5thNhjEH8s6F52uTrnKYFdR
NuC3/3bTD3rmqfOcPPLQ+4yQoIt1Xkts1AS5K+HBblikP4yPNmpuxE3wYDkstpvb
Litn+fI4ea8lWd+hwAeSR9K95oSuxYqH8E5Jub5+UwBCo21DXgiqmpQ85kINpBxt
GaUNpAYsn8CSxCj5mU8g+WoXZZKnUwtBmgKiXPqjVozgTgpOmiUaDDpsVu4e/00j
IBgJqn5QLz+zKwN71rHS1wlHmH7qTZWTWEwJYg+74MT+8EcTdhlccJMEgaq+yh/s
fhhY+KVvzzBfV48A1V3/MUh2C3DGhK+WkO043Az1pVHAYStxR00Dk9QbT99SP9aK
K5h2o3/OFT08T8wgXIznsljR5/D6bFphtA9uG029gQkg/vlUB9XCsHoW8kU+nSgv
w+YRMctB5/8O2IReuwyLeJnCv9gjfrxJj5FvaaS3/L+eUAL10/8/Yn/ncsEreY1H
i4FGhfE/phKnvioxte680zisQ+m2RIF4pscp4UvTYzPtundH/xec3qKspjlJTPoG
Fyj+8plXu/a57vLnUSnY1gMXQ3Y+z4gmJeIPgZlo17Agkc1/qBFs7mULNdr67ZYC
DQl9ki5KQC/nSwSA1Du2OzVNqGUyfwtQHqt8CQO6gcuPoL56VKWGvXqeScxpQgBy
+nOEH78bCrTlFRu1ulx71Yq6qPAtE2k0r6KwjE8WRcvylflGJghvjZRlTrnRglwV
Qm0gssJM8Ht4WSQK2PClfgIU9Iby9JKO/Tpwy5d4d1mHOFQ2xfBWZIzU2ECOSKsi
IDBF3GtdiQOSK3fWQ6ociC4cWzbqBA01TCcQ8E7JrmNjbQQsSGF33M1FORhFbIL7
sTfBUZ2l64kNoSzHEgdHLobr0NRIaCCV50Mpkwrx0F8KPFN2NPr4KNgb/tvYRCV3
5x9Tbrjy67S2ywn6rkdNke9R3vsx0uDYucLU5g+oCxSyiXX0b8Ea4NsNd/fDV3RT
0oqXH3GWXJjyZA9/koj8wuHYdw76mHwJYmykPml0c2TOvIrADouRhq0dY67pdVQU
36THKFLcSwq04Ex1UUZHyFWr3OdKnaQy9PFvJO5Wr0ydSJToPLbjDs09c9LchcAR
6/kmWanpYotYZP6/RPGbyeytQyKqdK+otFf2eOzlMbTWemMf4L4kR+JDxTx4Neda
OuvaltrSka0HR+BX1xknrV0BtAxFoi0RDFDl2DL8FZze0ax5uTXiZrahjI+kMhpO
a9iiGDhdJyn2NNJ+578VH/3bc+ktiB0HKcAgvnrUmb5oVBX63GaRlfzQ6rukOtKv
mKcxI5NXMx9Y222siOJKWHVB7/HW1og89nQolAHWb4uW8oZtkx5ZK7e+1GqL9J0p
Bq1pHoOUZffFZised0hAc1GxmiI5XJmFEPwEVPbayetvH8jBNXCMvpNq4QFdjOM+
ZJuYC2rWEa7rY0xmrYdDBxVJh5mZz9cRMo0Ay+HAxHt0ZPkkgpyunRzspNJdBR4K
r34dCcickP66coNueioUlJ7AvECKUEUHb7konglMi9e0QXtSoYMRnWDRJeoVqoCn
gx3hFreuamCkgoJkyB1grMbTsC+t9pk6Yg0y4GYedxTpW8YaBRr8U3D1I6Btbiwk
Vjw/Xelvmh8hxWr7olSCf6eTeDQjUlc66c84xNtXUp9faHeb5v5GeR/yoCQketnD
kJgacoywoITK8/f4eaxzqoRcUqXeRXbg4fEI+Yhy1N6jQOLv35V738nzdZ4mMTBa
/DEhOUSIuFmQKFXkIgk9y1GsWHdv0I6HE+HSmF8cn85wDOosDc7L/4Ar+r+2vY6p
6PdObWac8HaMDf2qcmXsxz3XO1PPmwce2rwiWffISm81aX1e59cPyCqgb8y5v36O
P5lU5cM+zMl7BZB3eJqRRK6OVp4U7/YSWIW4Rz8EYSV6E9AJ1D75iH7qVAqS2X7l
KOH1iWenNSw0f1Re8mxCOZpEU7E5fyMBGC9r9+FHt7UUzqWJHtk17nO/JDrrqQ7O
Se1KY64UceK3bFhWbQ6G9JBaeAUXEClQ3dmj+IPhZyk2MUC5tPWKCjVUP6PRP38K
RFZWnYnnywwHPOEySkeXUbRpcedbzself+cGeOPULf76ESA8aO+U2E9phMAx+7b8
v8QYIMB0U6kMiWMgIkQWAR4YpSaymapHYLwR16U5tE8E3HZzsGOhJz21Qcl+B3Me
llYTR1loHvUkhp2GUZsY/DaokuTLC1+CnoaM002nU2YxIxdnC6+obJ1v7P3czf31
IRfP/6D8QmqrHr/VOWtVmO/eEZtuuT6NNd1SUbT5z/C24zp+y3MH6dF329mmW2KX
dptPR2dWnTALflqQBVzUCwdkeYQGfumc8jVz5hk52PdscoLfJbLkCUmV6nZK6Jv2
ucvrZEuXxKyZeKhpk1IoWKMdYjV7vj6XcM0o1LTaTZE7L0saL2HLnZxoFpCx7Fe9
0w26s1iMRKT59hsgT55D/V++K3HqvfSwtIK4u7ViItAw1BK4sO2ARiZCDjrdCt3R
ef1HNHPvQ+Ew2ZwOrgu96MQGWhXgT2W4v6Md9lzaP363dyEnwNEvc04K7xxDYIdp
vWNa23FaA6i0yIkMQVpBeQTkJ93TE9jxz5yW0e7inF5/tQDPKxoBH5G5Y0QDnJ53
DEeTdVIJfh7Jl0RwQ6rsY1vOYnbvRnZRqH5QDocKphziAGuyS5qLCzEbNxGpj61M
S14cpMSY7BXoPwWUKvPXGbwSJs8Df+WGP+fBaCHnXhRW5KWgV38utyryCtbqBDYk
DgK0bJeOuSn+AIHMR4m0aH0oqfKxjth0lI5ff86Zij2TL+2cHZtHmstS2ID7Zaez
Absk1d8UEmoTjpTPWJ9gKIvYSTN7AAh5XR6wAHJPBhrmfcC9/SfbmcPiz1+dhnE6
Fv0xwvKThdphrFkKiezRg4synfs/T3ZmcN5Hl8/GtYiN0DYSGvQ1xiVfwTP4A18o
KOTTw7Ck9rGoXf+kQyWz2nZ/wgXp9rOz4gZh+YrYi8jUU3nRFqhqUwJTXft7uPI0
fbkiGaOqVLVEbKz0rpUeX3KRP6HGTTsJWHVkpQyxDAR1xBKBsvPBqnMmy0NatUTp
hoyCBdCRiUCk9numy4/qpbYPoSC5WAlF8UGiL+13PaQOhPQmE/8P/StXVsBe9JZB
Js9d/zihAQrqscU+S37jpZ+D97p+5I0oHdxjfPY+mzV0ITfzdJvcMEFXT459uvHr
+sf6qpIvqGclrI6np3VlqITAqRmgkotfvQuK4CWjJDcJQlhx7jP/pUk1qy4uDtoK
X/LpjXaCBHfpZ7FkXpaL6kjcd6WvL3ENWu1o1EHC2Xj0ZjB8IGqDf7BaNwU2o+Jm
SoVZwvSibWFDJdRJJOmmziRSBYFWgx8t8/Altu/0nqYErd7OeI4aYPITUyM00HWi
a3YbmLw4ug8vXUPCr/CtBL9g0bvRLVZz8QFTbVMt3+hGFCo7AowkOAC0eFIGsvzi
Op9LYpfOSFsjZbAeDOkp7QcBjBJyS6uuglFTG3CdrY672JCaE2Q7r2dTxonEjEK+
a+Ap14RVH58ZLUXXxytca8Bpx8dakuB1BGum0erS7/v/eA1nRPxwLzgqyrhfQBRG
nlDm8g26D46AOabe15udrrmuTj/US2tAO0Wwi9B8VWpYs8UfRDObonMcznMAppVZ
1XechxfVu6mgfEmDVP1h/i/VfmAp+LFVTsnv+Esh+9ed7RhEY79vc8qVwPokIutx
QHd5kdHPtno7PXm3cYbfe9hTSzlAkoI21KRjjiZlWCbSINgkm72x6iHCnGSmyPyQ
SvO1Wo/BWjg/3HWATT7BVr962JTRdgQr+8ydU2Gc8nOiVVs+sX1wSv6iGwPvnF2f
i9W7hyRMIdKORIRFHqUoKofi52EiYW7LN9apeFV27/6C1UNjSZbZSorT8uDPdiDC
/ujWnhURJDAQSwzudxez+VBYY2Fvl0otrZXleieEojRbcq+ODtnpguIMkLG4rwko
3OveBMBcHSwQybWdFL9FgHijKT1k7V6gJdSmaRi8wTyGzV+vgz2wWHom7/bFJzv8
RNtOlFm+Ju0AG4TaKMYxMYP3AMmxquEYBHd3Qe4OmjDUX5Q0JtfE9zKe3ymL9tnr
PY8G0WtBRtRfKhN79WW+ZPC8p1Yfd+Y0vYwBjNDw+IfvdfCcFj9KPMfYnNMs+cJt
/6b9XDJV1ZZUx/VFhA1hYUMSo4VGXOAOl1yZCTwM3njy5AdEoFlaUZ3LZZLOjPL9
4vHts9JobKIeDQfhV8/gn1SM5NBz4sQ+zUz4JfrQVcIT5zEgAzX5mInUTghOu2up
/GI/N80lm7/QLqnoIbsUgbcbGQaLi1jDsk2aRz8aLuzBS6hfNCP8rXhEdmfNABRt
sPoPRgt7zrCYIFoCSVrxGpcOhtdKXBEm4Q9MB5GNBg59nLzQxf5R48itHtsB0Ogs
35HTVsXRaa7rMv/TnL7ka4+GRrkLWvH5HxcooSvbWYlzuoB740xxr5CItzBd2rOX
Cz6ESYrIJrj+xJDV6knHrGtMaM8RqyhXJ8KkRov6Vl9ouqjQ0diLJ5QQ5/mSrq3s
mWMXAG9fU9dWqW+dxQpQewBGQcX+KF0+IHcQ67r9T1lxZLvCqn755u2M9W6IleQh
X6ajlIw+6O+5DBmE9B8sVYb69b7rkf4wEcrilk4yg9C5L8CyCEsasxLvT0HZ6q+p
gq7vDWt4qu3DyI1QKUz7pCJ0iwN8nlx150Qtdl1h0bIaDBb2u3xqZn+SxWi0CfQh
WdZMEjgoJzfsiXPOTqs/prD1bl1HEF9IjSd05p2O5wlpMoL9uQn2xRkVdgrdIp+o
4g/EcLJJTcwT06d5VyoH3AQQsWmfgGz1le5u2XlrztPcTf5MjCk/fXaMbbeaPdeG
250cutkS+CRiahotAjKe/dgs6V+ywrVKv0PssqG5A5LHiXd+fTsXzyK7BysNmM+I
fPSt3cHPAv41MmohSge6OBruDPlPUEettjDxZwuaSKgaYHyeljjEeQxC5yc8cHkQ
dz2uvROWWQHh9LHaLD7ess8rw0NcGy6a7Q25JFCf3Yl1FUQkirzqwKYNmaPScgfs
2EZJGrsZroyfqab+Zt38GWdfJ45bfJWiaco0BXPGQeaLbPUAmpX14kHp/1LVmNpq
BbzRZS44uqxkgtLwZW0NpmkPa9Zb+avPzrI5ptwGFhYU0t2oqV4qzC0tHAUpNuXd
6bU6cbjfhDRcp8i1e/IJ/+hgFlKD6NG6lzpOfthT9EisSFlEuRzfLhoJKsDQ3cz+
aEBrDBPApJWe7GW5iNNsycrYsdLCpoKRtEZ5ixJUqVRybM2/UB6UgYsfeTT3LPIP
N7VbsXl0Vt2uoOnejW9vkqZ++Y7NDVmCHk8fyJSB5W5UJOevch4hE66aVefaFlF/
lwvtP6mbbhLfXCL4wnng2tQ9moK9XDNWVSGvSFNbOBPGbHKl4uqC1G1Ebcx+8JHD
tF5xAov3AIE30vSieKxxUuVsE4olihHCQzc1vTm3Ra4FcGcZiaB2hmFqzcxHfdW5
VLoPLZ6laOVWmgmq5kEmee/hrC8H29MBCm+q6FH27+F6iwSkLWbUo1zR3iIvProj
C0EhKt0QVFcHn0dFX59rqY9BVV/eUU5iE585c4gafU5rHyUAwXL/z1/9SQQxS3IN
H49Pza1SzPCuIFwNQkj3JVUKS1utJCsM1VMxF6fIYUT2rnmN1LqW0kiXKvoOAp9o
XCWOmj51iXHMeZduWPPNw/yUcSMBu68H7TqnIddFlhpKspW7x/jETBRXYsNqLVLf
38ZQ+lFLWmhvSxKHAQfoaUNDEcNpWC2jFCeuhJQ5YJ72hAy6py1VDi9zkPPV0GqX
goZmz0UIBlASAadm8CVmF4MZHYJAKC/zSHR872SBI74em6+teai5dPNkVeDzUOpO
4xNrU9+uaPXap9UvN4wL22Zh3TuH4jqTNy7Z1ASFKElUuBGn1inj7f5PJau6pydA
S0V6eMdyVqSQOSxwwOOaeygrN/KjsHlCYQzRZ6RKp7C/rRRscd2ewDi1FQq9yiuT
vUSGUMDEqJHEt2xtFsdIWdZfTPN42o6FxQFO77mR6Fw1sA7luV23tSackXKi6hfU
V+di8bUJJA6OoUfhLZtWpoLspkEd4chAFWJerD8U5jlcrspCe7xY5Fr85erEaIGh
yj/4oO6UM3NKWfm0ZLmP0ojpPX1uxNox5bPiq73XdLtChQegdqIWu/X7zXaC9HPa
OgzCSD3jUyEImIFRzTzYNLIBekGciXOaK9tKVzf2EvXMcbBmQlURUS8y2OZF4BIK
VaROPywq5ksrTjfkDp4mqXSTLxEUddQpgZ650fkbVmzXcRszLEk4QyvsZOPBSrXs
pZ6FoKd0ykwOTbJ4b4XaqukbOFR3EVCaPe+v4FwtsaxdM+AzkIvI982mni84xPn+
e2yl6eikJKgOuE8xjw8t9duxQnRzDbsc+A1ssF1+N7iGNDnuHWFWlr1iFhyyVqHW
FWxzm1N9zUIepFyJSBMUiu6WqMRBWfr9o0lgi0/J1BrYJ6toB5NpEwWiED0xJt1B
IyQGv6V0EfFPH2u585bteK2GN/Q6eUMIvalSZ5Gdw6jxJIhI+EbQYS/V1DKSxFcs
N2OH0P3gNxVJiNksOscVG2gg/GDr2g0LvyxiSNbHgByqKKuCnG/ZUK5l1Ve//UJO
iyI75QQDmRMWJfhfchPLkNOSlwCVsHXuzc9NrWH5kCrAHfcqCcZzXx7qmwJNmUYQ
teUfVAAOW6uiQeYfjUqRnRtuMP99k4jdRSZONwKTKphDchMqiGQzL320MiWWRZcj
P3xrkyGb8CQsoFtOJ5MLDWHtxnc6sWz9krFRQTAnhwxm8VXy/qrJpNxpb93040pT
a5rh8atge1QILG7yLOVOYl0dE893eqk5OSnl+puAyb3qaTZfZhtFfjf9hXSFTePy
kggXAZSWPAMayjfAl7h6BaqxROpeKHbD1tyAK2q3esbmAQOAzPo3xXjV6WVtd5z7
zrxzQnvnYeEhGd2vP4Al73ovKhwWwvG4p4pAqnFKvYuslxy31JrUD6JpP4SsNjDE
kdnzmQV0kctUy38hEiUqkl5J47WeBdOFmz+4kitocRhCssoamWjcgo/giFGRPlPz
rg781mbmwcv+krhToAypX8c/vlnuwBwXA2rlt9gdmdY/jrA3NzGrRiK5hpu50DOJ
8g6pmTcsBeryNR8thAHL++ALhXBIedf63PNCgxv9esD/JnRt5TC1iQ0lTtAgA+mw
sgVEGxCH/UuI3unxGrc/ag8giw+0oMpvADzM8p/oRfp/D79XoKghGJke2/8iGcMs
VIX28mZMvDHWXgcxTeiwEbSfSjqkaUcdJ6HxSPzLJKSJHkTHE5xdmmhsoaKd68Wl
X5b/qgiNslXjNhpS+mtwYZZOFSMBtnepfW3RLTrTDcxl9jABXF2Q/jR1Fjernq75
r/ARoGAbB5/gd34KVrKmUhaCMLntDMbWS2aNA7h0mLuVAQdVzsIf6E+ramnoJRCL
s2iu8TAVqc5sOukyqAAwEPCSdiMqIl7+qr1zvTruQ3Ct4/W9kNa58MypcxREFlIv
dGG2vgjR+y0WrGm0BU3G/OSLq4O+Tcsvbny47GB4lV0TJFF67DU9a3FwS8ePT/ay
mPUZMtfACVokHNLgNAqpk1ZeGeEpE8IAIjfA+I9t209CtvnBFIcxOUPLtvYa4m4N
SBuhweG+CFoQ2gCYuQ1n+G4G0cMiSROdl/3aDem3rgESKVOUyFrNt/pFZAeo6IUw
r+dFXXrJ1u9jV87skpEkvjZX6Arld//dsM3QFm1/tpBFqoyd2dME6TEplUFYXYJB
ouGaNBiPmTkT5kM2wkzzPRpdguLLxeqUFUlRocmokSTE7EiKfQkVL/Uhwmw8l7E1
3wreFoB5hC8XvG89CpffMfpT1mDB7bn8lIcwNDPHjhSUgpjEKFLmDI+Yd11gDdwQ
2U1aK9Bds9lawCXnk1MzZPjbPQ14g0Gvl1gTB1+mxp3mgMOhgz6Y1G8OVxohefRx
8y/UuWxaN3JCqy7N8zEhWWSHSjb/D7rswlMDIAaBwpfmLp1Y1Jip332NH4UxZjoa
4FqAHCmRzuzdoUVXRHNRSBiOPXcScmZF3IaH1S81OLEfi3jUtuQ72ZXPMBPup9xs
SHRXcHlbikfvcS46uM0i0zx/7F5o63T8eEy+6OE0fcPKBTpprm8izQCmkNcZRaWG
pDovp1CdVROVLfMk46aA90c3bBKOMcO1aVlDDIJhPg0fQQQfoNW6cXu/c+JAdAW9
6DKaw9l6ybC5fhQ++zEETWmFRC2koaI/w45v1mJbPUQaoOStDa76M8qZExOic/Hm
EYekXSadUZva1Gy/8ZkmeHYdPlIx4t0dde3UGRBj7ijWa+noJ8rOUd0Q/kenpz5Q
erorzBXfgW0iKddpp69UPgUCJJvqqPlQmP+AhDLRv3vxTUL6nMpE0WEJfeWTjk4z
eiZkz+7Z8SwSREHtyctaRavHPwrxaWvUk5zH6Xyibk3a1KyTiMiQlAVl7iuDPyKY
dinpwiKFhaVCQViOAaBsPdfV5dK4tJqRx18cv2QyyQ81pX0lknhIxZ/hjxZleEwB
97QkV1Yp7zRcpCxmlcTQYh1yhr9oE6mT8sAh9drSlAagE7gvZFF5nlkUGiUeBuLO
WOiENIWljwlQFkym6/rHJbnquNzrdIbE6R8fB8EE6r2SklQlx2gDpArmDcIVgm8u
bUw2eOrV8kPyVZcdIa44MU0XYRSWaqjxofJOCIraGdw=
`pragma protect end_protected
