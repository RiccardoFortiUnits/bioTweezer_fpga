-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JA3pO6akK5qOFf4owxfgLypUXCUpIuzVfp0J9u/0wt2Vkt6I76d3XGj5Uxr5gAsLsqrmph83dvbn
ykb833xodPzf89Y4Nqhs0BTm97bn56Ygyee9Uz7PN7iNq7mY9jkJoThdN+VNez7JLPmtX/lXC8Tc
HtiSph7blov4FQ3uCvGRlKso5/TJyco/UEDyIljdWiOsm5TVic5XpJFhZg1qgZhJTlpPZLt2z7RK
mpuqS8u5Atc2FloBSi4FgkPrmaIiIKY0wKstC78J0pEAgmBIAGsAdhCoNGWJHD5wick3y8BIYc7e
B5teo72sWqqqPcYBRlK1ttkAIcAphEK7JnPcGQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8560)
`protect data_block
He/6z/OI8LpJLne2bnnKgEazGx36H0oI6qdypLglw8V6fgG5++dArQ1YBFwZTW3xewvrw5lC97ps
YDdJYkFLAJPdsb+J0jLi8BPWa7ufxzBkzPabsMzpbLcXHTFkgIH8IRseFF5JSLviW0FsTQgT2gVP
iggFhBUCBBcIvYAjiJAMl2wDo4uHt1DrOin8Iqucboq/BE0DN3abM33tEgxJDr3qfgZSMq2dfgjb
xi6mKKi6di5xcG3u6W0G/efxZSVMo1o7iAHgi1qWDixXpBvMwoG0gogD3eK7Nm7A3/GZbzj7OGUK
GL3KzJcZMTt9kY0E5PrpAfhRhTqkeY5cqUxx3181zdKAbYXFzFRwO/N+jmQQ6wYfK5/MyE2Zd1Cn
/abhna9vcVLuQj/IDVmZtUNhLzFu6Tt3E5YOWUlbO5L/2csi4sEYGBvC7XpDlfRIY8HhAU17AxIg
sQSGzeL5c1bMCnj5mpIypl2LAyx/ul+PZaBkTQvpP7O72haWNrntcqhUmxTfeEU2+jYqxORP1goE
YhjUARXdi2XupVDgVMiuPrqVI5UVGTszlNLC72AJwiW+LeFI6jd5JVHucVhIASx+Wdaa0nllgybf
x2pD6trWZR14368WNhZJ+P443Ri4ifgGTnxwxnRWcqcsQssQFTmCwQjUYgnxcw9eltWzsfWgrPe2
SOHVhA+6LwtbfNHLEBeL7QCfgH7w1fOAqBvcB1yQXpGaAEf4Rb2liuaC2xeGGd0RXUQrskL254TT
xuYehzoEMcXhkcfUmLpYFeQRfngyMA3pld1AyjMLil4eWqTxgXVgmegF6zJz1DkCsgeBXvUU5Xs/
495Q6Gjmt521q97H00oZfAGi8ovL3M23IdDYc7Q/a9t0UIclfTP4JI0DuHDiz5pVqrBzkia1pZI3
+SKDnKVtdz3HlsyXeV6cfOTs8gmQmN/WtGG9YigLT3CH6yovJOgGubWVRTDw2NNnec7qPL36urSi
shE8JiioxDKQG90k5y12wuVNFjek1AwFrJHfjOzmFqcshC6RaaU0n/A2lYzDzwnGOGfB1UJTzKbJ
IUbmaI3n946xUWKhdlSlF1sjVaodFkU4yfmjaN/RZWKf5ihGAAt/6dKiaCS4gtIAP2tkG0mUUhRV
ZqRB2f8tTlJxQib/g+AjoLGo0L3Y2xnWQixdJSbtGF+jkJZdnI0PsoMHL+KEWuHbPor5ODKxNntd
BeKSnH7s9fTIIsKVNiP2SQyAIQ6FNSrhGm9S9A4Kf2TnO2vJpmIantt7ina6PnNnCbQaX0of4I4X
78Ga1+E7FvH94OhdnFAmiy1VQTkRMftAFkmGkZRAIGBSYluuXCYEXMLYGmJOld+1LHxnlIpOyft+
D7pUi2CP+q6zqL7z3kso9l2MngnnfxIcAKD1FDF8caJIw0i6O7Dkog+FTlU2wAWKYJtTJrrlN8Uf
M+9NBtXA6/P3CDtQDpYaTZKm5yGRz6rKWLEsh59TbsCVAxkKbyZZdL5+ecdVzLrVZ/qyejBFU0Kc
NJ/BEQRjJc4ThH+7+2DKKcu88wX1I2JC2T9f8HcVpGwMMIIZ38S9lwj0Ppco8usUqnD+YwloGB0f
A5tJekULkapt7KspteZBTL3YAcv6kL3vR4dX0XXGUovsvFeSORhyLOgG4zBRh/s0k+4jWqUGFM2w
GT/BT7VfopzI4Ut6pH14JPC/XqDBj6qE9gETCpZrw2V+3kxZAsg+UQNndvuzjv+4pITNoALU8aIu
Z87MQ7HC1mkpPgykx68K/ZILmQ+tdFLpK22fehAzJz1uRFKg4ffvDdfymqqDPzuDeyazrngSjSTn
5tFPk3yNRdZfpJH1UQHUYu6jPZ2M7JFgmkMjZwwEYZGKYXo4B2fYZqCQFoRhn7JvG74k2abwciBg
7RwZx8BZBdU6U/EJqZ0k7vxLWDjYGZ0bJLAwpoiIVZoO+VKh9aaewBgSROK24biSpTKRYJLLc0If
DBVtsGZYVteQ5IpPUimxysw4FYSCYPQBmPg7yTmzpY6pPegv72w8si0LtIrg3rmoD+MT0ujixnOn
Ov7ZdOTAn8UeKADSNc8apED9MlUcAXAjiZ/XLczIKtV9JpIGPPM0LDMf/V8Ibwp3EF23O5bGYvl7
9Yr+VDablaeJPQGH+3NMppdeLm3TAJbidmtm/LZjR0K8fnZiHKA6k+Dk7y5RKwvHIiFmjKoCmFYJ
wW7q6VkYCvxVZ3DdjweXAni14rMywMYXjrlidyflkfl8wvyz/f8+KiKB6ChMEo4Q7tp9o/H8mTCq
pmGci8foaTYuv1tg2vFsdgesUbEAIYHwS4zv9hVFLaA5yI7Aa9cURaDTUQ4TFHOJjM1wnzuhu1Mp
5Y5WGbtj6Lkh6mOVzhNvZNZn9YQinnJD9L0ALhtAEgCvSD/yvF+sbTiW9zBXXPjWnklHcDbS/A7Q
BFMO/Yf6J3zib/G+AJwitLYusPfskcm1cM2qUjU8FJcb3tEWObkZwxwbubn4dFg52HoSEt5xmoeF
8MukaC8pyyQ5tnz8gUBZGfNqFnz1mnx6hotAJ7QBFCgGkevV+n+JfKs7tMV1smWRzu9CXGzamLGQ
uLHP2v5ML9C6NhUg6aruBOwRx8XxuK8KaBvO9rZS8SAqUPqrnmmuai9fxUPadXlnoHEZpuZxjKI8
5ks0S9H7fuO81k71KHT2/tcGbhRo7IiILkbvcXluZ9FVeF0RpV3sJDFEPt9K8wW6hA6cD7tBYvYG
YGUL6mCnNW0qp98ANYIoLzoU6HHMdMTNML0Xf/Zqf7mJW67VLnc7EqTE8C/fl3OUTxrzOGbTOB3Z
PDAFKCrKbKOWs3CWsdoe8hKn9JaiwaQUm+LaqJc9wPg+NK9wZO1GQziUi9SJBXPct99+aN/FMSUV
ETwFvYOI/AzyMdCoZkX85Bvw54GGz8C0dk4afURf8XrczQRLw1uMGhIRTb8Ly1wmU5FujgCRljV5
XzqPs1evC5ypFSeWmKZyAjiA6nzUpV/4OhXyfQgpKvTjSsi0O9ZhyqAj7QNZN5e5s6RmdwSp1tbj
mLbkOKMmFYfGr9DJ9rJzVaFtCFluFxJjOL9MQx1aKzFBZ0jkO6L1ldNG2LqOxknIemXIrKUJuQe2
Ks/yaxcJrIx08V0CvBwhjZa+guXYzHe48F0zoWlwxjjLfab6cnHYOW6WM311WMuIcxSk4su9oGkg
StFYF8eLMzpyKflNW6ufaOEdaY/v2T1exYdnoGgxg8zJh8BSLGD0ipeSKinqa/ctEK2i6sqV4du2
elYJo1Q+se/VxeB+0PnxE4sL+etyYndOPetG3RigSC0Bd8Gq/D+9qJyNuz713hI8kQncVjMTBKa4
ufgmj/Chzw95hD9dsbIzNphhX7p8eND+gfwYi2U8JKmHVaDdBS3E2UmvkW/YdrqYgg4bqlkl0qHt
QiwKtbJalTfaSHy9biFslD/fyhlI5q+JOgOXAkI8naY8nB+YxBLsDVy7eZ/BZVXwhXx3reSAdm/l
VPGzp9vUAIheeeNvEhzoUM3tEwbrxYPZGWlHfGWRXIpx1KAZMFtDYK1jxg1Fqwx62ag+Benxqw+F
Sz8r7QGxr0e0pZaivaH2OcFVhdraMRYNCGF9uBt6ilXh8iV25JDCq3V9ykta/S59KSY+TZ9/ypo8
WACOJArtpLC+16bq6M+cB3LEVVGpdNVumSE+ZYs0MEW+YDcw0FFh1Rwkkr5viZtIM6317J4cZwO5
3PolSra2yYXEdBdajTZ81zoLVyw+LS4gBHB7abouZK/TeacjL0nRnB4rzttamPoRBeIgXvifM2V3
Fb8RMjrRZOkhzKu4asPLg9/bAl103NgFqQ96+NWCRnm7ffO3ESapkAC10bKXgJBE5c5bkaQ2dIkv
01XitUbVfmXioMYF11ljkrrX2wBee5D1kFUDQ4+m4kJs33J1WoTlASeZlzl7ZAnRcolSKq4IdOlJ
EJqXbRqs6QbmN6CFJEiEmU/UFGmiJdh+8A/KFKk9rao77f1uJL1WJIzWukP0G5OUg6y7CD8Lh0pU
vJ49beWjB8OPkGuIpl4PyglP2FckRJxlfEKT5XNE70OcpjioI1GjAlT3RcQrnd8jSPGBHUHBXsCa
bJXOuNaV8Xw1brQ8yYEvVPx4cSemshXznQ7qpnRYxGJ7l2y4JDqenYimnRtUCpoAd/pSrmZBVbCe
2qNWCwywFHyIv6VcdzWaaSrf3F0/cYkSNgrnvTvkQYZ7PYaldxlqwb9U0LN6I1swDUnozpxxnJWi
ezcBgDG1S9aNenSStz2Zo/i5VdxDwTWYCq1qlK1XN5CtkwcZ0JEKQXYK2HL7nyznibI5UY6bvXyP
BzdeQ0Ckeu/v2wftBrlfKNhBvK2O3Dmf9BYYLzhByDHG4xdTTB/REhyn3YXouV2icFhx7pb5BamJ
GVAUR4YB7l/AYhPb6ynXhOXP3RXUFoNkACNlcZxz/CrCqToVYHSAcsgps6/xYBhoSRpoDaa46V9K
ajbolFp0DhjLEgpko41AlZhqSRC95VITRiCXhXPM2MxmHg7mttHXZN0zAzXyDg2w/IIP3dEMdzUr
eewEidxrhwRolrh4plsXZKKeL65RlN12DVP+5FnsIxjmVLZNB3VRRmIC/csNnLZjN/91dzUO1ky3
Ib8WYMOq/8N6SO+XNbWUj4b6oXgqFULEfsCVxSDn/BVgC63TE0diirkhXU+u4km0pqpCIHq5oZqT
sqrWteR0rTY0npoxn2AdIPbvo7AMO46fgqejySHuTYpAr6FJczIcsWjOD0IAmQZHWeWrh+soi6Sf
Oh/u3NGYF+U2aOKPsctnoCXhI9ksLcIMQJIoyPopffoBLGu9R8Y9nTm5s3NDfwMbz2tzjVnAYwDq
gN3nn+gEKLAwY2341ipahQsetL/a2/zpFNPsJ+Vc/TRDGzh7N/RqIU1Lydv5Wbla4lFLp7aB1Rmr
5Pe5uwkx0W/g4YWaVRlP817JBSw4CMo7kLwhYmXOvttOZ6cB7QjkoL+JSIcdGPecjk49CJRLcz2b
d8wwXJfzm3ZwQgVLOGmylPrCqxg1mlOKhxSsYLaXPghETfYEy169QBL9XTg7CSobbceUQeyTYzuY
gVLScUS3axmuaFnAzJ0wqg3YZGXn8bF7l6gZBm4630/yS2zEcW1f/Cw6U4t+RvMbA4fdBHTNXe/g
4EIffHo2MT+/dbNlkCewOCQLoDYl172RMEv2kS/YrHjGnr+k3RebyxiLpIcLfKYFIqDKb6eiCBiN
1dMTsmrNAsg6Uxg3VNuridiyXdGuKGZXa5ng0LtkkyMm0qzyalwPaxhBgpSpohkyWI36xcjSFAJO
HZoJhF7Q2c8hqJB9z+ikry/T9KkO66+d8l+/qVCDVeJ8Wbtn5lOp6Tnh2m4WukjRtrLFHXAMo+qu
noBL6y8EaAMHFWBYjBRF8W07rhMOpU8T5NDc8/Zbavp42zRSJUFdVgGWiw+t4G43pteqYBYvoirA
eoCgPN+ezMlQAaRRxDWVaAMTD6WBmMDpaf4zzJMus+Xpy0XEpNyAVw6HWGto00zI6VhcQ9cu7Vsa
fhFNGKuYIJ6dhb8WR4AQ4wHqsxfGnp8x5gKBCxr2v+NPx7TRSbgHnl8RW2cC0wvHrl27tTwB3ESd
nHO+SJCD5T804eGyfHeKnBKoatRNJfY7l9zKj7yMytkvUY6o3YjIQ/fBvOgD/r404DoolLhm5P11
+N2J3eDN0oYIG8ynD2/dapjwuZV7c5++j+TTxW8f2GBDdyWy+iwlQflxdXbyyyb6vKdCLdiL3DRl
MOusiad5znwgaaLoPBfO2ASFbiL+fpuqr3zvb91mNL/MMWqfRfwFyK+D+l/t7Gz/7j1jrBmKQWGt
u3CI6Oh0bS1orlZ4Iqil1DvT3S4K1I5Ktj/8F/yNaA6/n9uHQNrGYMYFZfkW0t3Ez3/vqd93Gf7D
zH2ZTyw8kqkY6nvFcgkl+kkkFdTIo87+c5VRrpO+NuNB6wjy4KhUWTjzd3SmdiH6rUdlnevOdFBg
3HTdcoPE2LdFyt19sSc0esBaw8WdSCMcPAANTFRwVEkWGbfgBGPe5DJXKOqnmtwtgi7S5vss61KW
AEUCYp8JB887FmbgHbA0KfwPLY1hZkxljFvoPYhfEifwz0KXPCuYLisWpQb3JSUAPXuZBHGT62IN
xoYuzNOVMwPE/SPlUvB7cWUFc8BTf1edbRJ/FdesPrSAs72iDr/iAvUEonAUG9FMEUGJtP22ssOe
sJvwFz7krqvHAGO3rQvmeTDcR2XgDrJGZTBT+RAcktCMv0TlISxN5a6J1EVLJkduEQhQE6N1IRhu
j/FgYMThONt+WNqRBFH7lPWZCjQuBQRbfVjAq8OVSfDoFGs2c4V0pdfnustMQsdzLAqj7Ng6bLXQ
KKpr2thYVY3Dd3tf9OILtvaGJpOm3otZoq/apd/fTDZ+iyb2QFXVJE2qj2hyrvAoE/f2EW9figag
7yONITgEhLjmD7t8pR8kUXgGRqein4nXkMlhxNo8/vTs9g2BQOQ/4APVv4HLEuttc4c/kxTcDZcJ
kssiqDtk57iXCuJNhaSiELzvWUhTpU9tK8zOFhpUpzPEabNQo7GbaLU6AkyxWGK+V31P3iaiSQFb
gmXso6QkCnJNns19nivdBHnmQX/ueHCtE5WZGqYobr20KQGV8YKku6zV+gg2XCqWIW1Gh8j8BByg
7ATssiS4GsPRR0obImu/j6pOwcADeT1W7MuUggnCyLGXzYyAnxxa5Hxwl7TwBC7StFovDbk7LjSM
KtCRL3P7vY+e2krzHI5Gzskj7y4i/lnPsbOGl5ISCtyYJytJo3Jqygjy3HjeoJ5jw/XNZ13lnvCE
dXtBlcR5UhKyo386CS2mRHMQQTx8061fKnZqvZN/p4UXX9OgDjBgiXYFqtFykNtwiZZuHYy9TR62
oOpeisknmiL8WnKDJxQ0KVCPJ0E+hDZYGBKnw07qSjtcBQiovMz815TQxPBmvSRPLJToczcu7dZ8
Mb4uORiMYrzI1aXYWXcTKvxTVG9Mqqet3MhA6i0+rynm6A2Et0rKCRGt7rNa0jxPyPNTI7AT/fXr
jQP7Hyls7fXhjCVLqiiKz0Gp3yiQpEJ0mhrSPkt9b6xdvJKl3uNqO4CmrhWe80AsVxay0W/h1zHr
eEg8YkdJRuLZqQfuF4PyEtiHQzfsgtx/thxe23BMATCe0gMyepssvI1YcvcycnWejhvIahQmnqJj
STRkpO34teC3AAg5Hcjl9eqUyFFpMoppdhlxlBBWk7gxQv4KouCRlqPotSlY9N6koCFkrvo7uWKC
/hM7ZkAGOwZZUwa5kujqum5gVrVOHoDwmY1ILkzmGHu/cj+8pj5GWZs99TkcenAijKC9b65qQW6V
+oYE9SmSnnEDQdLKN0v9HGVhNKbcan6JweR0lbXP0ySE9gzO8mVbLK83QthgOO5G2fOcfIZHLnNX
sh3pNfSVWNqHrX1nNAE1ztSUeVCEd51OdqKQlR4IakYQVlDkyQCf6mmJASC6ux1T8U2W0lI9i+5/
BXnZkxGVIn2tl+H7gO/7qG3bmfAISA7Jzus3rWLoRYg2Z1rlN/sBcsjD02FhBMSU3cVVMoY8yPb3
YjavU9FhGIMXzRO/crd9IeBS9Qet1I4DTzxPd3lgJbc9KQAeTaUN5u8ORUaA0vaAWe2hZh9fW0VH
VbLqO2jE5TW7F713Q+tHamDh7584mymypxaIATXN+b0/U1BaWAeTfVTTqVEs6JxhwNyln/qLob5H
p16o5mn37x0q5m4sFqyaKV14P7RmeBAgk2ly8QBtcWiEag6OHheeI58l7ZBkJ/VbrmtiaiDln1Dq
yB7ZcjAlt8ho/k2hrLA2IwTSBCtyqrXDWmwM19iDbRNg5DNjWk95MlVcq2w3gLvM0WBotOb5hiKr
K6tplqEeclNLvCXLtNfsAY1as5rb5CSgsTjaFkRlgWfQkkQledr8jH3kkl3f4jrROqg9WKMKMBPp
fTRHcRl6U632p6fcnGjK6RPmxGECYYH/HzFfpl30mPAw9/RkyglDPFKtXtLNspB4wvvbFlOq91DP
0jIs8uJ+cDLcFDi+yjYfZgdxsThbajnLYa0ODyShdj+Vq6XVBUlg6dijdU3xjvUXszK1WTYIpW4Q
AAj6c7P7Sbkz//SGqrx9W23LIAXoFevDnUpvfDBcku8OV2WAffq2l63Vydo46tIaxa/0ztCOnk45
z/Aa3eBuEb6KbEI7lze82zriC6aF7YthcoTUu5jaivK9ZqwaLSjbUwPUAWAcHY9/e8JB84u+x/fv
jEqLgM2vCIjBdgwdozCUS4xPOj15s6k0cZ2ND9Ff1Ogy7ROER3fyrFzvbIToz9ABrVNaxUceg+YC
xVOvym1SK4/rGnXCSnLYGWCM9yPa7oYQOt+zSnjAuImckdILuablQAGNNzUuf8M13R0anIuQXK77
FBUs1iOeJFQ5mHlivjKmEj+ALGzIHPULVJlFc8/nNkSKGjhTEFXu8HlJHxsv3E59cmWSWJFE2w7+
NKHJWQ/MtzZhIbNm9LBY/YWbX3l1BWPsnEhWZtwJMPln0qUjTKrKMPmdFEnuxlvl+RI3pd51cKDh
81vCd/FW84883Oog14fK+zrW/h4Ym4/7EEUYsfJteE90j4TJQqK/JN1WPpvxnYje35KHlCc1uJfl
hAN0xe/EofIwDXDJ5/eFBpITxsCplUg6x5+w/deqEdcx5p0kB1KQ8OYS7lF6kC/tNG0SUy8HuJCz
GXshhlWjh5JSp9YhKAgO20SDBTHOw3pl2Mf3WESN965ZxEUW3ZOhY0ENGszuhyWb03ytyFSy4uDL
+0TcI9wi072b0mt2ucKolRLWfwa/naEi4wYacFQrjnDLlxdU8BCR7Zudq5tF0wN3kVOEjO2tJLih
RbZfZoTI01mrthB+6EfdtSj4x4R6Gem0a/xcDuK6GCpper13pIExQKhbP5cCzm7E3db5ocES74ko
AnuI8cOqoOgqhY4UolkfCmyULZ/yHTEwpLDc5+UMug68JTVUBnUEa7Fw21EC5oQR/sI2BMTRkSLM
c6wEjLPBS5BYSvR7HAWYKz/D2N+CzNLqhumtq87xy86btjZ9E+s9LKzjQXq83xLeG1s31Futd+xR
weOLa6nRg846a2YFsxphAPDhz6JL5oRJf1qBsA7T9Xbdi/SghcmJpm5Z9P4QELlsdHuVEZ2eAcb7
yFrVkfVH1oEuNrEoQsYYPtZN/YEpvaN0165Y4tuIez3CQRVh79I5ubeOKlQwEMvMef0RFwjn8Zm2
Vs57VnZ/5xYHxhAtVAwXnvCb8/gOxwL5iymGSUb4HdAx/AwI0AJOupWXkOsTawQ/72cmfWf9PlAb
moNsW+B5Sg2641n+5LZBeyTa98YiRBIg6yciPUiKG1efTLkK3EUWJN2oUtwnAHuMMBopnjXNFAVF
D2AVo5EH6MnZKFY2RM4I6ka12rU3qvg/Y2nHtZMjzsbNhOXYWlkyZM27c+p2xrqZuzckscolI5Gn
643SPUtVczpQNoMy7Jtdovgin6IzAxrDIhCZpbxVosqVP6c00uPtGYBP5nyRz4BSYIicbuO8oF2t
9h5R4nzLCAXXcucDVK+kKILoT/wFHKwblONHS7oUenrlaTqseCcaf6fVRCeFZXT+9RWy92FBiobj
S3ZSU6kV+zaHCGJ27BI68m6bFAZ15cXjOnO6f8nKzfoUa3/nwluvaberpsay4/0YN4rHILuonwLH
MJMBpXOI3gkAn/rjL22sKEA0tcdC8dcOOs5VLxcGKbThM9q9TrvBLYL1l9rfVU0EVhCyAraYYVNN
KE45JqMWDgelwo2q39/vLeVQ/cFME5XSB/RdM2eGw65mMlkfmZq7bVIlJ55rEGzoAxBHovCokyep
AjUo5boFL8YgJ3SV4ZsxsNdvYjzf7FdIXdLkknbz8Gk48ynUp8Rz9kQCiRo4M1QXLEzr3ZMKdNzW
+qa9pVi/GBfLCawzMWACuALYQj9emMUrZstZGaXF31Znw2S4gvJ0yUfMr8hr3hxkiG8h/KK6ZnDt
bN41CkqwzsDXiz1EBLIIxOTB7cXY7qvAMEtEQxdsXilJ6Cb1jrO/+pCO4iYyyNFMhT1mMuu7l+Fa
zDzekXm6tw76B/geHHIzJjUgTiR/RRxK/IBosnr5MaoMudG1zvVFHvNnMaim6iSyP3GBWhTyr3zR
9FvEj41wxi+c0ptFgwlD3Ls6fS4sbGENMOT1h1JZ+WUTpjLaQO3TmJqINrdrbvpfk0BtO/MD4OLO
RN9b07nvgge2IkdY5N0cUFFe6Ra4gD+uMOnSiEVnIphKPjnmiKrgagG8Iu+4K0YASTOJLkO57S7f
gT95Rd434T/VUqhfJcgYtxBZIlLnU/mFSBJM43N/vMacJpA8U7zR/b/4RBF/Lf6D5Iy1IzFTT9us
q3i86e2FK0n14lliuP9bu0L20Xju6RaL6HvTJIhZNwk0j8742GsYx0S469hzrtvHTj7g67tAin99
aTo0Ma5uzQ/8Utfk0wSNvQfTctj+BE5/S/pRHoVde+anIqRL58HfIiDjfhRv0aiJu5nhEM6OQWD9
01V+Nvuixrj2Akff7mqS25dONjjs0SCXNDNGsLThr4K2VFXgp6n59k4H0YYmOmdAQBooQQ7X/MKK
LpQG6eBJyZGxNfgWef98HInwKkQtSR4rfz2sbd3Yd13nr7QRvbjaO4MJU3UYFxrEx/8xiXzLLfpr
9SMlFdh6Zc9fJReOSgnE6MTBwGy0vvN2dLkk47Rhqo0BbTXRbfCv9hzseIBgyt8BlLVZpw914hhG
5a4PlTGvTxhmRSc/m9izUnT31SVyJtG1z88YCFg5LX6KcszzyaDSkXCGiB2pp+SeICWDAOC6nvcm
3SuORuFOX04gnvIRHhduObNGYTtxg1YpbFye6UdFJR+QH4qKvSTpB4L6ImxhJHIT7lzEqdq5Ku/6
H8cS4GAQSw98G0/RDZFLJI5UVXUzm7NZ/p1pPUTPTjFZjdrN73cnEVOT5+iyCokt7jhSiIrkGcCR
lwyrHlu7JXJ/08DQtXretorz3YA51mwayykrBXm2AkMCrKDhapYoiNah8psQWQDNAKRaRvVVMSNS
qiW13Hh3lO44wbCIdxRXcgrL3lKsSGSIaIzpNPi5ZASQf6HtulLg5MO7mgYjLCE2JMdqUlr33iSg
XRDcyEDHxmdBv6YMGhttjBoSlBsfzw37Dpkilpf91FbIFcIWDlkBJ2Zwiu43xqZyFR4FthWjSYjz
MFYBhGE6svtqrzRycXatLwTPm5XJ6npPw2NxIjpZyr/L+5NHE3me5CZ2qkX2xXGnFqVOiWrAceZD
5/kDnb4srZPMTF/MF5HGUv6k6Mea/Um7HM7K7tbz2n9RT0sucz1gkl1JqTN8jrxsZJn8fsKwJFHM
rZ/MMOqKVvArVA==
`protect end_protected
