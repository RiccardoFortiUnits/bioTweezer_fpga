`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l/9iUJYNYSh3xReMbCiJ6ka/aBGe5fLfFqbQmU1i/0QdLvKD2kRJN2n9wyXzyVRo
nJxjuNWJx12B0RFOomI6vm0UthbIIzdpzaWhieBABei3ORHB7yA4/4YdMWsb2eJQ
HkhWUaKLEpZwtz5Gxy1KcvBGjiWJhp17m7hpI4mPF3Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
rodcLB0pxjMKi0QAVbDVdYshqN/2o6K05JhJz8SE6VqwrNP8g3Rz6+CihCPZB3FQ
0RqSGy2I12YuwnJjEmjf4+BqB9fy99LaUkm+0ZB7Ps1EgkT3/eTh9aXWsJVBXEj3
IWPtMfZvOA+bASC6aROLEqx0erN3l+K94A83Rt6wDWaZFSnvGUFiL+NoMJr1YG7I
Xag6ASIgz31/HX7r/WvNk7ICECZkliH4vGyJa/f0r2cVZCg25TfadWUvMWceoOY5
qRPy1U/KDvNWbu9gGtl2tfK3/xCeDnIIIYUbAF2sNdC9jUGicAL13x+c2LOAs+8E
3PENGRZwdoYTgsUbhqmQhjBYMvRmDBNSf4iZqRCWGjZ72GfWmrWV1jn45XQggzdn
S9XzoypJevHQS/Oh45oE8BaLCD+XzkbZsf9a2yQVVxwXSpP/ojAWnB4n/SDqzh7b
l8+qfQrbQPJiuFShw2jbAGTnUUKDWaqudHku+29+7ZtbwV6lRs04OW1k/T/0jDFc
VOhojOfV1otz/I84Eb8e5QxnafqWwJzsOTJxgWxsMV9BBdRqLMzW3S9HPd+Y81Jy
7uEyNnKAt7u5pjDVsfhJuZgi631BjX57golztOQxL3k6GN+eZJxUb6+6dkIXXupw
I82mi+DLACL8HYyFQLCjsrnQdnjMeMpa5Pg6Pv3ZgIhvCb7Ak4JmOuvZa+zcO4A4
BvuY90QUu9WE27XJWjKPPbF/YdzY7nYjlnSxURQlV7OlCeuXvPP8AcdUpAWHwsym
0mQEMt5czW4FitXFYmUmBgH9QYP8og0LfWQsnqTKM0+dwEn3/cELjMWKnw2uDHrL
M4u+aOBpy2sANsd+Q2zqMpISQH/JMKppkzXC6eDCjGC+bSw/Q7LV7+EDa3e4jbeT
e3aqY1mZw1gscI7BzkOUbgOh6INLbCWEX0z9YQjsAzJu4UXWt8VqIlju648iIYx1
bXGAtu7P/ZRHC01YHTNhfp9jmQWZlFTGL56ZLpnE0INm13e/OmUBHFq9vq4QG7/d
y7UZaRoiskcprd42LvNYB0LHQYCSKv50P0aklGY3MrTwH5D6llqL6LH6zhUS5RoA
SApbzTx43Ew8OxxEndfritvqQuqLDZB5qKAfbzudJoFua9ya54JXzTGrumdJdNOB
48rMsxZGCFyWTTT2rygMD/BK/4e12dWvZ5FiybfKHkwKLKiqeKQHdFVINbx2ku58
EHWTsLWS15+UfYOcEzil3v2ZYntzOLwVg9UACB2T9iNLP1dyn3ZU1UhW7P42GS6K
RRwRtpDoG+ftJQwN9BGearpA7z6PzATTb5bdGOo7WYygXJs/LX2HnRCe2rurVdFF
A9sfaQayzoLHLnLo02UpqBp8H5aZsWcZlDJPlB3IS4nG/zWEuks+EUG7cb9WEKHK
tcdpCJasUNFEBaIk/kFhTLyDalX/WHvwFcBNOaxwbehY6s6JxUytA7dXkr5ODb9m
YcphpMPLOUq0/1BSYSx+pVV1IwxwhtkZ0usuO5I3Q3i8IeVFKQHh1/wOywMt9kzO
p10EmTurPiGMB7TbPUFWWaWuEnymKITuGrQs5Ut8vVZxI+kU4CMgpGL740KYGZO+
UobKu1TXX5LWIOmvDqVHz57V8UTxwm+BBSRekCSOChG9gxRUMBD9EHXiVrjptC5M
tdFypYu92JSrWcIvn5LA8e7FQpvRwzlaTPfyCRbubyx4KU2hH/QntbMs8tDHsXBu
N5K8GhU3NrDwtWTUJC3D+DmhjoUKBr9Ch/Q1jntC9F5BAhEVxcfRRUpQg9SOj9Ay
NIff3Q0H0lERqwoKUhIpbANEw94rN2TPslRd5fwnlljuJRzi/upfBJxpLHsErG02
BmQV4e/XoNTos+60uMZI9faBFTyrV4Aa5hp4XVnxkp2G14iR4a9A9b3305wFwSkj
E83J47bApZwjnKTztswHk8m+02PZkF4Lof/RbBdx63s6888bGAV9D8MLhONBZdp0
AfX/yTe8O55mpzZCEGAfz1KFUjHULogOpgYcpI8W0HlLO+9VllQq7SATj8g23C4G
G1NkvLfbLmE6UbBkCcEk5PZ6gSvrw7nC91D9qKEb4W3zfOjUpicegGJGgr1zxWuh
MYQquN88e291s544Wcwm4Abws36FlPZL2H1UtxTQIvlNLhCYoSin9GM+4LYAddHz
JUsGY6DLC+hyAAuLrGv0j0ltkayJoG6guv8Q0EUr94MWUfoBoWSZMM6We/ceyjbk
ZQmMAr8jbYWIiHEYiGgLUoJZsIsFZDWK3Z414Q4JLDIa/OQL1IhxRPWtMzuLCLof
oSb7uai1/wn47r6iJ8JH+G6HGnMqQn0YQPOCoimAvp7i61ok+nKucZA1Ky+KTc+1
xGqMGl3hQilEsaEoGJxMygdouBagpFQyUvdbGiRAwkU/W0G/WgDu/HnNh0Bqnm3o
CrSKWYtFIRL9Qwo/mzvgdBjs3pacqhtHH5zGVO+/DKUr54MiG8n6tVP+YNAlQ+RS
PeKpW/Ao89kP6YekNoPr0k8YbkRyJDVtEJiEsMCVSVl0J3D7aMerSwYwyrnBQK7t
xl3CUUafENWebWLajAfxgUQyMA3JpZ8h6+nps31yYlYsnxLzHwpkGBx6HVrSic2j
dCIrbggch/DaQWjhVxwbP7RjgJbCwJpJMCE6AGAhiJjDvyq/IP1cLbNlQ/PAgKPF
BUAxhxRovkwlykRvmpQPs5yTllrkllkXX8cjzV4IdCethlBwGBGFK2Jk8vVFrUFF
5Oinwx9qmDyGXlp9JBwh76YFbKJvgmI0JmE80kqlWEAH3pBOwXnepOwax1AfsOvm
cg6xL5W3q0dZ8auhapfvAYhshY054o/jC0FVxJvhhmp/2I8y2B//IKG9d9nOPbHI
TR30mnABo3qnAI5JxD3AHouqZVtN83GUzGta9Mj58pw//faz2N4PQel1RHLmC3fu
Af02o/i8LEF9AmkxoY+4FW/vQ/wGE7EiQTdqkZ2h20WIn8khQ4Rosy+1snZCZWvi
V4F0RRK8p8X6J3coQXUVtbyCfqYhIN8cuJi4Kr1LulJwHvLVBmzPPZner/1oXfMS
u6GrQ8QKBcjrO33NQvmEoKzz4XDoBJTWY73sYFLuZ/hdSs/fcTu/w2ujDxat4jd+
eZjsUcau5Mnqk2l9hjeAyBAqX+w2UcaxvWzdyOLvNmsH5AlbAbq0MhUjEAVwP5A5
kJmxBpsCjxDkQQlfCOZfaH2vYKTdvN7Baqp5IMiFBzUmXmfGXWiQIJAax7dIme0j
vw3DSERe8/ToAj7eS/kCIX5U6tpSONfH5oBf8yoqNmcLL46gu6EjKfF1Sphlbytp
3Qj/MtOUB7yN22d+xxDQU+HOTvTM1//IXy+apiEu64zGAx5QsxbHFPa2MF7AikUB
toonKEDXp2wPrVJm5GavSQ+cX1U5WSaijxgaAV4JcMMaZQ2R1WmpufY7l59TdCSU
ONV8qtvdGYAyXHTKE0EftbgooOTVAzSaBInNcu45uPHCVjkDod/CuWA/9+Nazfyr
HpjBePmcGjswUPgV1e7zm3xLeqNP9dqrVe/7a/WN9JzZAW6temMV1X3TFAhY7RQi
oLhpyDb/jhI12kX0YKElL9SuOTSkR9Py1TDyd1xgTFXBrVAXbjbeF6EkpZgkQab2
Et72D2Wv1D3aOSUOHOtOu7eecNxyt8N+C7FAkEoe1Q3VOhZHL+Rl1NNoi2Og8Osn
Q6a0vHYUx8rYmOPTcbf9mBpp7SfVwEhUoTmRNmlJEshOX8Jnb8hqG3N2sz3j6baa
JbwfmG9qfIYq/345wUcW0YCa3PO9oADnyXlfPlreW8XGZzG3Y0bQ2z5i+CEaMXYk
33v8UIfhNP1w4gmea3if0roZ00SNM6GfEGTWsYb5mImZiqJao+hBkj5lRsmOt1Qr
3q7rS+du9LLVixOkkOqrH9QkcOCoRfupyXiDr7LOy97CivVz2jra0HaWb0G4WC6E
/RclBcP0544tPJgXGym7E2qBNiwQwC48bLTusokf/Uwh3cIPze3XmIzkFo2Z0h7P
7RZaVRCxS2HzS1W4EAqtGk3w2K6UNlRvwdqT1FTgDPy4+aRN9iVQU3V3ucRPxN0z
odxH5q5LEtYVLUy4INccFy0+6V6ccF1XpsEOklmukobuelrnlZwd00jzVzbHTRsJ
Q1HxOXnWTpeXwGLC5L1zdS7QJmzrS5b5euCwEACiFHLZyIjucvJ2GJRmJwteEhCi
2H7KjOaaAPaCrwIdhbJwHeg1X6Ke6oBpm4wVyH+MdlYudPITKYRKBGp5SdHoDyaj
rNaARieabOWkoVywIoZ6w8JC/xVdSvWw5J8QvOptO8lP/rzU0oIzMGuB9S4exUx1
BLSFAIVIhmHYiytgZE7CKlbL33N/D0Jq5BpqLWNLToFEHOVvIpdCw6m9yNnHILjl
jeDZBhsMNbFvMilEvDXhWsZVUvvjyWycIjCHC5PELPqjY4AsJpG69L5w6jy10vfm
Cyr8/d7WXZ/i1eGflvGv9RdcrLr1Xnp4S+WeqQ609OiNG/ScYwDY4WovjShyeCa3
nIWKuJ+tlPLtk9dwCuf7Fn69rw4O3HuM28urfPEzyZmEVC6xy7O4EW2e80AFeR2t
JbECI3nyDKSPZapAJmkXhEGti2v5rW2mnNnjzAegQSdS0gAImR+iKdJE6A0b8wK+
bq7UHseYNnFmkbXDqRu4C7jWQgdeZ7BrTtmLz76iXiyjrMxrKCbGzTn2TjBNZROx
v2FFqNXvhd3xTz9l4xozJngrOYGTTCEymBbyvoCyeeMpmCnHnqhTOPP1F+q2k4yb
mXP64+8RF66Tlj1JEU9A9AMZeN80DKGPsokYftIzhc706NfzN13gjE3DuawIr3Na
pCc2gJ6AxC/NORrV6q4LJaMHupRGzluYd0NKrGaP5T3wKJvzDg+cTJorOeyiEo7F
Nd+U9rphyHFlPpBXrEm5twPF09Vd3RI51qHTSbGQcK0joaKON0vzhrnDU5tZkNwm
4C6D5qxQum4NJOnXUbqCiU2dgRHNHz9Sp54Q0yh2oy4IF3PGIA85aOx6o/TGimmf
0oWe/hV4S9PXsKxTGR2HtgfhSjwLQ1TpP5G/v0FdCLFJTxBQiJeNIqSNYka905M+
vNfJI0skEMZbQAAsR6bWpP6pwh2M2oJ9ALdVyCGVVcRHjIIi38bo1wOb8apyOpxE
WjM574hNOLtK1xBg4+QPjdsizS7vXwzzNE41lwl+yAhm8lffGSyQ1qRy/7Ad2znb
cQLXgrCKFvDyrPN2jmgOzf0NKBShIO4giIHn1N6/iBUa5r2bp+hrlxOj+GZWd3++
9d3hgzOdCzuFcdYszOXKMEFwK5c6EPbfeznLcRvIqyx62PTNb7ec25a5zLLdqb8O
xhK8n3LDf3VRxM+QR1+CX3HvSyY5YfX1KOowylefdDCKSvSQ8HhsT1vlWS29UjvY
FoYR51+MXrYvvm5iYx8iQdWZoEEaYx36aANVJ8FacMUphSRnQM/hVZDxOlRv8Cs1
sw/okMUN8I1xfqih4Vfs6xsial8NYGnhAtGRi/qD2mBLpknvHuAy1CiPSvJoWuZ3
JCrtxs/ccImhNmVVJMvP1k29BgGrauyaQRyVExyvQ5s6s8EQlqqOWmus/jzPjC/I
MTU5F+SvRCJlWwSCJ1ZqiIrp/H0xxtVhnSpW5Yy4WZH5asyHx2G2DhE7QAPYh0Au
jdJUcCYRrx3j483neTU6K1vNS20NH0dLFHrE325WBGFSdHTkXsAex1E6lC2KOUmW
uGyhURujGugeLRC/vbKvVTGg6D5PDLYWxqAFDaQZ8YPEl/bdqW/W/TBhFDP5RnH3
5FtLFYS6K3aTle9iY93Wv2JbLJrCI6FJgdTVLsPvqsEzbXgVVfu2nb1L1T2/Vopa
NulAnPNAAabBhFy6Hxx1N699NK9rNaMI3RxI9JssV3LX48/vjx+lZfy2Eh/Agduy
nRD31BVnZBSpyzEAdHdonyVhkqIqvc/GSAdRS1XLVA/OcF238OLWSZJ1O7VUA/5K
fJKpzM4frN1BJql+qemU9OajE9k2lhKJtCNx7NwDVzFHBRlhqegYcKXG8YbAR+Qm
1vTQrZgCnAqoGOKsKgo9X2EPAks+lbBMIHMPql0t5SSyQRH4ty7Le51lqB++Zs4z
Se3w057aUTUQeFuomGHfBPutovALSjH92A6fBtYLfZR1FDB8elNdzkSwjfq7OUnl
LsUs2LJJAYd7WaCUyF5pEUIM2Z1We9ZhT9zPsoWtrx5DLAG+jLoEEgLjHuj7KqgF
3F3ooaONarJ0adsquvTYGv1XSirBe6FM5puiKcDjxdAtoXBDxo6oksKd96BFm9+V
v8zeLildGVMURzkyrpS6aj4vG2TVeGxxoBKSzxxJ3mwIYddzEcArtl7V6UbXONXq
pbRBDFRoxInvqoaZ3sZpnuLhe8uYuaEXlQawu+OI17pW3OWOl+4esqPp6rv6sRV0
T9r0yuNKeNZzWeZZrgnbUR+KTBu0+oAJH7QgVJKH7q2eOP+qZxdRO2YrqIOhibOZ
MkRZ4QDmuEm+AzRvo3WQRqyv9OB6vVx/40Ls4EPhVBEqMCFZfd73jj3Z0Z1s7bpE
+bjbzP1G21KtxP3DyUoP7wsCpU5miMUn6rzysMLBdiTH8j5/wrlF/DsJOelzW/YO
fcvhmGRUnaW9cunY1fjpV7sDiuRffy2/uLL5KzFXqjC75ECFh81JB7rmarefr5et
gb0wPwi6kBsK3Tbio9K4t8TdelV+Dax0g901yBAAdb0R+GIk7KDS2kErxHRzqclI
ASgaWftV9hCpnFFdJs7ViSv93Mc2wdFYF6SRm217sna5ZZmgCh7oNAymfZDUE/p7
+UA9h+xO4EO2o+Q4dXbAkN+tplSI7FAYic4HDeKvSjKz3tFDXdLXiep3HkIyvxuu
0VaIZrhiMeaOmWqcMfdgodrXZe46gLez9NyZ5QB3xKi2NKuM3VyeCRlJk+znWe0m
jJtPTImPBV0J1dSSYcbC1xYKdl6jRXb7/ZATGfaFHm+n8bebqiTLaInXJ09z2wk4
jYuWJ21HUhj//KWQ5A+TxrPBrq8Go2yiSEcjtkzMdEYUoTehnOrutUROxiBqcCpe
AeMjWaV6TGt38QHtJgsLbqDQDhsKf7qlbEh2jWpkPnjPq30dVcqTijydoe24NZhm
gLY69lIO3poiP52eVityMkhGIis2O9TkrAhRrOI3o6wbqZQBTD+7Y93w2IpNxpkw
qFDWBJWyY03MhTR5YvjLD+kikmclpjYVSZo+ynV1xZo+ZW97Ml6fpD7vFF0x3PAC
uqWqys+iEuSNmByjy9ZgzXWGEtd0zvwOBvnrk42MCFApW2ny2clrkmJ7r7gYwFG8
p2wXem1typuC7T0MdeykopwQxROh18zkUNHM4gRfKhqo0R4kbCT86vxtbigqS9cm
G5iHf2b9sgv9pFxf11lpqVGIZIiYveY441e2+i1XnP+1zd0UFAsSKP86iHvyNvb4
MbcQZznuIV9YiWecx9K8VMMR3qwYWkC3qXUwmr5Iejwjax9/nYx6jJemWWrEzUXd
ATUdalhDeGLmmMRxGTfCZo4dVMz6iwMKWZ5HCtpsmXJzp4pHqmyJcVhuEmYe0I1y
`pragma protect end_protected
