-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OoBxdGZfHg4Wb0ju9ro3MxwT12FIC6nb4evSE3zkmqi/GWDcH3L6vgPSmKmblgiOhpASpSGlFXmT
9v2r5EflHkbBjPb2su3Q/+fVPoXJVQcVvkbDh8nh4Xonf92eMf+eR3PAcJohj99gS7ffLwvP7Z1I
yq57kk64gvJBBCWuf+L0iodSrNFBXAMzOZvYLPKomakWdtgydVR3IGXxYP6ouupT3VkXBPtHiNxJ
IZJRK/exByg+fcaw6GmqDgPQ6SR36/LZFX4GDOSMQgSCan4G2gYJ5gXyfItF/0nHXNLi1hWlZYs8
EpG25p9GqYUOMZFTcxUeHzoAhfXZ/B13yAev3A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13456)
`protect data_block
9XqZx6KvkVeZ/6oiOxF+VhVcHB0b+gujw8FnnfEJXXOtwJOU7+RyX3OmADm/qrVXPCF6QLUFe+bQ
mlf3pF9KpyM8G8uKEYz0nKqw4dTh1056TSNSa+RC3o9zsjjN2JOoCdDbMq8Dsv5g5H8lrllbB4mY
0kgX/2XsgLxPAeKStx4wzPA6ALaZH4nno70Y5mHTkfH2vnERtlm24rhuK9W0T7pfyfcgsp16OoyZ
GZR2+v94oeeYrti225Z3vFkcL/kwl6cCgN7N/o01tfycjQBgPXERmSmlUME2QE/NF87AL/Es2R/j
kQ/4O+ZzKslasht5aukoujOH5acD0CwdRWfFaaE1xsJmjHPlv9XUscMBp4/hFaE7rAtYkOQD50es
J9wy59FxKJgeV7+K7JfZQ7EvD/l67A0fBPh8Dj/XOH79iTVJszTvdRDIjZsmRKjz59UJyDmo9YPH
HGa9w6djGoeKE49P6msn2tDzd54tzjxCu+N+mAMuL+RIo44z3G90byf3SGW6snAxUBXEuDUO2F+j
BpaLbtH8IXksp0YZNFmN071uq3Vu4NhLHVsgx6If3PzgWbZtcWgV4RyO0pJBZHC8BIlvNBdiOg1l
n9DKvodCqwIgv0ldro0BlcAVulYJuyynERDpKEHFL7QX8cZjxd8Y2u4qRGzUWx1OQJp7nMmsLbrC
YwcCYc1hzzXNafHNVk7BHKISMr3TlEo24NE299QzMwKfRA7A2HnvESRa4tnYE0mfD/Ss1ztdxZYh
XIvH8cJ1Tv970qKFAxJetLv5Ij1muJI3unQP70NGAe+VvRBa0t3iDr/9ysUPV86KNl8JouShHgSc
6LlZpYsZjFz03zJzpl+3IGQsZsMrlRPIQUOSqFc+dhbNwkgabsOsFiTbgT63kaI0GpvJdq5s2YFt
McIJTf8cB7MstaghYIMcGp4evpc3OsNfU8y0Ky12zFivgT1NBUL7YmpexTSiImUiYMVIHTSxkd13
zI0VuPmaN1gMSZZ56VYE8Qum/Z6tldGboBtdsCI+J3x9VaMoyoAllwXG7D+3C+MLSHkpfUAKwKuK
9azt5/wJl8sp4/pHqLFqjbiszzk0PuI2keBwtYUkxCFgIXX+9J5UdHiYipajd6z2NzCp624A77yt
rIq/h26jjjZsGHeUhM2bv11GkgubuJfVnlwcmgUTvU8+dGl06QIElXGnO4ql8+Or/N+kQKumkOIe
axM5MDyQXgwprhX5vxWL64ldFlWi6oBHjJveSZdjAAuAxspu4Q55m5cdDNqODmuZU3P4E9uDth6X
ge0jmNg+yp4YckSH+ENs+WrswlRfE8d1GTksacmBeqzQKjAq2dI1Ts7GUQBHGqULIXa5YA7bZ78+
DVsHWOXWutrzmkNrR0ozpcv+IG4TW55dWzyxy0v/ZJgjnXBtYmVBTBq6Sv2pdonJnVdiVpzAYVfD
ttoe9HfVmn6Ru9Pkwt6dYYLC7bLCBb7V1CU6Kz/2YFHeyAo9YROlE0GYEKKjYg1i4wyyZNFcfnD4
qoKRHQAXWhU17iRST8NBG7ihHwOFaFO+u0+v+EEea4+WFLQASZnhxTm/z/ek/rK+Bj8dlabNakXi
qsfJMApj7Hohvf+tOc0L1Ow5fxRRCO3RuDUCc9D7FL/d6ZQbQABmSxij5jeJzDsE4CmSFx4ay2co
r7F14t5Xfz27AEXmorDsr583nkJXaRm/pbKOb+j+ECSuyfp5xxtcpxbTBB0QoiZ1ugHCwB4cSasf
bIog0h8Vb6X/Gle7Kb7E/kwb/lUpGqit2DzumoI9XDLa+2e0Ct6E/bekKOjPeH+u/cgMWGEs1xHE
7oWyQTS6gZ1x4XDu45AxlXblCvZSD1rCegZ//9CV85tnRhBT2Z+Z/BfUHmvEG35EWXly1hyxuTIr
x0HI6o978KP+lDh6ScvVbQohU7qArxWUl2zHyvT3JvCo5mvmvOHSZD3Rm+C+PTQGgHFKBaP8WX/R
tJA5qSC7M2WAxcj7CcKwDL2m4KqF2LL/8Is0Nuq0asj+OHx4C0zhsfPL5lsxiRKd5PgaqGG3/KZC
hjLSF4UA8N5iFbgpRo7IyIGDPhdMA8cyhaUg7d5Rhs9Av/Uw7ZbI6e/xQvoPPvDguGALdg3jrh0Q
4xbMfDSMaXtKIt3vOZTeggMvK14Nf5y0B9vG+FBYDFQ/k2/bHv48G4CJqvQgav7pz3GS/uWLtR4R
2F35Hf+h0c94klVddFBOdCpT1dC90ieSzMtwzaigLsv4L69QbDjtyMdsE+9ycbnCijw5lKI4d3xl
mT2DWVWOKlqSIKmcMjulzIJIFmuinZFE/AUAdh7z013iAzOBlkS+f2PPt8hYzgxL2wFbFDS7ia4F
6kLQ/q1g63frcmsJ9N/xv885i5t9tuoWoh+XXjlhrTL37sdna0FbLGQpk+6L1c6Xn+h4LfFRx8ed
nZF9Gi8YveYo2V9kd/AO5eTzI9C96VVCXXQqno1dGKJz1c4jBoWgT2BFE/bnpzC8VyPkNeVioHIT
Ebyhn2MqDv2VW85bT6ipY6tl8HA0mc7yQuHe+1FKUMpa0eEzQ5LsLzHvrA3+b/1mUJxz4J3cInlY
oK72AY4ILcYJGMkvZYp7xEAdbNxkwJL30jA3P8SND6xB16weW6HhvrN/bHKRZ5ZkGPqgAc0aj3MP
QGU7cb/da6p+EyGWN48R/ecZVlgEMoVGsBURXcxuNKI9/8/D7N7y8Gyg1QrfkdRuR5GtLxQlyD89
y+MhU3T0930gr2kDY9JM1naIvJhfDKiYGvUe0CDO0Y/ATuhIDUYJSs7VzR4bjLLEFxmOmPgNgQ64
I0DYN+MXhv5M0eAb6qKV7pj8UTzcHqVkCWq8/Mbft+UTBHdgqau1WUT1ieOOAR0IlvfjdLcTkGij
2sRZCbyPput6HBJLOR/jW2OLrdgyTDmu2AuVCeCDsyWVxsQZUihTzRrnnTpCLhQswA0YIcYCo6Y3
Mb5TSXq30l6qFp1kR9YFU3C5KaveRy+jaibDaFFY1NHMynODSIaIElpfyta8/1xmwf5gVlniezw6
GiuR0FLb/eegywwN7tS2vBFzfT01mAjggexYfiyqL+8wUOGLuqdy9hll7ZN6htK/0vNBvctpsfhP
Z+pRlKYMPiikzejRUb2dHbMmO2qnPCgomrzDdFJK1/VdS5//IsZYrP+mihoc2FYSSHFHhL5G+icM
PObWE3cmbxHraUKV+zxFpBWTZScn477uaV862SYnHR8WMbvZHxJgikYN+hLU+sfNmeRhUitIu2/Y
oSM20GZvh6r5Ij4FW47w8UYrgExcuInZGjyLAIRqaKHMAOwquKFniSjzYgE2W4GujpIDTQRbBLTD
bwz7KNaJVaIKy87AFNQ2sTKhC2k+WIKd8vkqnhNtwcHe3e0zNURs2/tr83GMUxBZxvfKzhAtVOM7
szYeJ6jbcrdY/1xAgW1rE/ITu8wkCmMEJfKd/PRpn+lztdrS8vJFM7dEs2SfcKNsAIlMymRaGWkl
P4DDy/CcG9u8K6Kw08X4kOe/MrMLjCUdlR98X4MDC0Ai7zl/VPL7S3kxhKvlp1dCSW2wKkJNe7A6
/N+cyCvksgYjJ5BiV9cclu7WriB3Hz/9NgxazV/kktX5bod+JAN5KRQkQBiKMvX2xBIPl8Fj3D7g
yQJSV9VrwlbSqNycEnoX6bNGC/xvILf9A8fVuKdNKoHknlTqs6fFv7crGuPqLURHb67Jpsda2hyF
Jg6nAPA65pSVoPf5MZ5Eoh/cmgeUl1fGHlME+ZFN2t9EKXzjqtRMcDv6zWfhUSIvm9CRAHHwj6yL
7KNXPIX5TqP4htaXH5G4YtFDjkImC7OEFxGzkcYq/ak4soVn1cqClbdoF6SWv1M6sAHLXzsc6mnn
cG88Yp3OxuzI/hN7LvPqovncnPSK+AUUz3oBVsHkZ4QP3e6+FWJDbA0W+Y5SjlMHjrQ5J4l1uVz1
BkiRWeAdK+u71oGQG0pNiWg9Ps3cJ56nxBdzRNnSV8o3GZ98Vh028vzu1XFSgr+xVbJd+4hTOnM8
5LOtrth6Dp8hFzvaCARwYmxGev+8ZJD3yhkkXa2aZ2EpA1w+hJusRopRY3D6IpyaSt+UhZf3EWRg
03Ndli4eJWxalYHDZNicfmRTtxBj311zwLqGqxsc8bzUq+II+op3dJ1Yew6Pd+O0XIcuxD4I0J+m
TI0tIxNiJqnXn07PuL/077qhPHtvaGQPfqSXZGVDw8VA2lbCLjXVeUKQvgvePJ5A+Dnr+ASeyuvX
HZ8osf1Q8bdjXUj15jh3/M6aFhXcMUAQdICZHk4o/oYMRP+RyXnzNc4CKsNymJc/atIdrWbCgvJS
2xpW0fhSeFJ2F/zFcF9JwevQViwCjYlX9BY+VGtJWPYcuvKeyOl+WQe81KVMG76kMX1SywdIfhQM
bSEId5UO1GYTVm2qyBHIMk/fiYLEVHDm1+Hv6cttxsH2hmMM+qbQiNUJb0JTpvsWp4zjRwIwc/Zk
ouGBChbmMQihFs9gJL4M6qhpWrrNg0llPHDa8RXPWz5IUwdAITRbyKg+Q21/xFOUQPQvvgkLPPNK
RDF2MAOjgTKzdv5yG0jqewUJawRqgD63DQ5HI1gaoookf9uZoIgJUde7G3BPwA/McUN1igVFB80C
mltQOoxzzSeygA/7NtApcsXoJ7IlDxmkmo4rhYtW5pnMoERCCF+rOu8pC54JCY2d8fQ9OiY3RGnK
6wOxS0I3ttTbnj8vMqy4HIH+PYsPepC+f8IpjWzbHgYj9jjBcLvmDRD2iNHqnisoNC1OdzR4Ecr/
uOlf0n763e/BDeZ1Int1RvWUJnynlUydspkHnCMW41NbAsMeJPxZyONHI8orY9ZNkbJxmMTOUsF4
4oe8E7w3N3voISZFTkF2CRhC4ypa8WcAMF+0BtESLRY4xVZNeCRSMiqh3tMLNzxxb1dEp0w64tRo
v/EqTIv9zX/G3SAcmPEllk3oOLwwPMKLoaWlW4RHtSmGjKGRjMXEco8O2dn4iO8hulxzbC3wIOfb
i4EHbf6to9YZdg9cSyps14LFclobq6yB5TEeWyYDA5szrIbHBZ9VwPsEZMLxHipRXH41xHNhUGcS
de7shmzedjelLbgZ+BfC4TxZLqDw6me8UZflfEkZvbpGoL/+IXKXzoa5zemt030oPtmenLoJ4ASO
Xfdt4vT6YS9bOjGMbm4Mj/TnjGRq9m+7DgG4icLcjmFLWF9DDBt5JI6dTD1ePLW0xkA1w6KEos17
Tfdodja2P/EnywJULfPisI2pX/CKDmUwLZRIEMP31qtO212lh8YQKlp/UfMNVc14rWL1DPeLbXYK
Xnxl18hWhNIMpX7EDPsnB0fvIu5fKxI2Ty3t3SJ0TWVcUZtTuqV+ATe3HQEImi6O+dgEKrqeCQqv
ikC0AgWMCMw/0+7SgHC6UuIZEKtsqGOMIHoq43u1ST2rAbOgzLK/6OT7Swk14ED3L+fzN9t87KiN
jZybcx66Bnjbmer0RsdmReePZHgYvGWMhO6ZyhHIC4GXYESSSXIHHh9Wkq5ejGIi6gWFccIuEQRq
Q1dOoQbVTlGGX8//IIUKriomkDhN0wN0/o9joP0S9T6abc1MUL5sgNGspC7kxzLjQL+4ATKedeA1
MHF2dMbFF9+t4I4vuEQYh1cYynd15CU7jUamQruF+B8vGUBbmVKi7t6RegVyeZDxmzYj59gnbJBj
x4wytdx+L2UXiTPHGyyN4IqBwjdLCq38J98gZlzcnws3WwJLay33X7UCmP/9c0GR6TdD/iQJfFlm
oOx3cX0m0WG2G7rfuRukYNmebHbtJD30KgeC0Uv4LOJv70Ai2XvHkkJCM0wka1jlLiLFAck0UvDi
yTjH3vz4pXqNgITX1FjEGos44hpQUkMHVTu47CvFVQRgmiWjM0Y5W9ZejarJOIh2RIqNo6ZAeZ0Q
EaA4HwBJdDGp972688n3AsDgMTmj9GvtQlvef+42c5K+fWW6ILonUGbvroBzwQ69s/MQKIZDR+nb
8WbbTCvFjyA75815c01lrSPcyQmSn48KDXiEzReLumkq7YH8dopVm0ut7hyeTcIDCbe/HbAQ3Y3r
C3ejzCI3CLbBWSosOGqAlzKUnZIp90xjldnVYcANlGm71YyvP4R7wbyhj3ckEg76hQccrvGjUtn/
B2dDeimw2OqD2ybl1x8qP7ilTQcnCMEdRGwEjWEfW7QDu0G8UVajSvW6WYb5W04zfgxmRLDrjd5B
p28eK+vmaZ+9ia4FseIpzFc202saNJZoh+g7CVxZe6ws0kUXyBLvjlbQfj/NRApjr2hay7NUMR2s
V9oEcoqKN5tRAmfPU5OpoZHU45NnZlTPWCrYhnq8Pt50YHPDGTwtywZ4cRHwcy5T2xEEIYYZV3OV
u1Rr2C/xyn0onXkydGwzLwNzsdgH5fy0TAqdlZwBNVXBHBRt6Cmiu9tAaydNgV+1/2x8DTbfkUAi
XUaIpLxHCb9t0c72ZzJwGOn5BTK8Lc1548NCOnSRgkSqwSLYQEUw+g5B5oD/TSPhuqCxtNJQ7cSp
C3KU2zQDceDXfCM1idOBHcy784+gh+CVZiyxJO7p90FujLF/vVTWWIIB5qjKLEgHAAuwek07ZZ2W
K1PtPZkvU9k8VF8uKGc5U5f8ZcJsZSoYnVY8Iz/N65+0SVrhn8SnoC1C/Ayjf+PY2V/tscLH4PZJ
phKmE0wqbnWkLNA88tpagYV2AlvGwe71viTsVk0GiypHv1ZZL1KMIzzQimR8AE1I2Kh7lJiDtx/i
l2IXi2W5PnLYJpi1Gxng8xGM7l2xj65mdHyWCOKrgBOgq0Ja+aPLIobftZO/nB5jfjOF+5I6YBDS
ZabDBHTOgy2GP9j0hGxfh2iwsTjJJlsbmuRgdnwwvVUK1nNYIa6Xdg1zMsIzxtdwmtWo+4ZLbJi5
oXI7hj25pMP/JFQ5m/QmpG3VDdO2vnDRA+8zFBejsqxRYcg81L4idvelB+d840I85piYI0yE6XVD
zwLmkskSCprbpMgyONXn4FtMt2rkdbqj0bSwUh9aDjSXYSEXAS9dqjFnTbSYZzhMpL1gROwrXiF0
o/M7Ga6Veyemw34OThzWivxSLX7TJAET2ifJOCb3qwzNN0IK9irlGMe24+pOdaI9TyuqHqRhzJxl
fhi5incpVumSBWNPZChlkGQ/XHSy0xcxWYu5/sa65jD7x2fdIyihr8DVqivkxWZLGhWw7D1YVybQ
aEDLaw8OZ9j+OeF+BkGpVuvHNtEpCFyVgKUQUrKbE+05cPJJndbUxfplO+kUR0pN9tQiQW4hHJ+X
C5XgIEmsvlQJlfG1aYYeZkhOE3jwAzpgQUWyQWunh/ocp0PY1qdWkPSO3sKeUaFrH/Ol/FZ8FqOF
Tai06warUxpfa8Y1YPj87r8BJhpoo+IExjPdtxYNtqyd6+GD0P07PTsXkIU0OlGJG+RNL3UDVEBz
tMZdtIPYDpMqPXcikraTUD/vXmfVxH6dzrXpsI9R6HlooDlr/Xw7QaXl/bbs1slcUnwSt2sUDEeA
xm7KXzeREBCKr1DMSAiJtt80A02upBV6J+RlYil1TSVFAD1HNdBJx1dhjLXKTX1aZlyBYzYyYXqk
InevkwPQPV+qIOc6U8UAhLhV8JX6T4zslUddXLlu447//hDdQ3Ky9sT3mOvou67Jj8RBtnGIIxYj
nvhR4m4lR5N6J0SrvLgqNB7YkS8gBsEO+OMzBEMumgid3Ggb+riKawZufCMk/CI18m5xhlO2trQ5
Jv3Bdlk8Q04FKYy2VmHybJYSKb/PNOyC4Kz4oi+dTRO898DWq8Z6XO+AXTKpPqZz1cJWd9CcVyUq
mGhwRInLaj+mS3ucJaa9vpf+emEA9fQhEL05ojSZG8ESFZOyRlfAZF8b84hT6/YCQ0LqQ0cjwOEV
W6+afOyf3cu3aO+ENEbi8Qyf6ryTCBFoGgMg3KvpAAvLHtHkOb2l+HJc1/C4XzJLy6kzkQQodDzC
0mRUMqcktQza01NXIL2Vm7gd5/JlmM7P25iG3mGcB+MnzMsYuhfNvaLDRexK+S31m9MUrI2nwITg
4PjhBTa+QDoyAAM1bWtRFdxJ7udPdWtXXZ3lhZmWw1BbWohykhjmUlN/SfUFC1bDvrJ81M2z004N
y+b82ieoCpxHKnhiJrbXJMAoy0YbW4MweBI746ZpO4yp40lesgrBACjizHAAYu41ilXkhbqpPXT4
VX9KvrENXz4uv2efRZhsgh8Grth2xaWE5PBBd+GnBzBcFDd7Gm2Zyy3P/YD4ukBlywDrEFDj6uUx
7ff+7nVRg4Ku+Rorn9VSb3Vz3JZKbCF7ohUEn4GOzIS2MA4EdSXmA7Xj3z9u75ltO+4qJ/UbnogE
uqJ0qqnTYctU1TWx/tsGPxvTpwE3mdeYf+peNSd5xVWp8OjiFS7uGJW9DuxbDMLEbd7OtjQsxI7U
+zdBWcPIs0w+v129BJCYzQaCX0waMOXRO3O+AmarNl0eu99eGMatN8bfuBw8FXsQbA/29/2V/Frw
iX0xL6d3KUlKvJqYqsBhTAxDiQnINBn3kzi/z9iVN/VXq70apVfYyFEVftbtYR7apBhDqv4LziEP
yJF14mDYIP1bFGOVs5DkiHInV2sBgepb6QfDYUHONSp8plcv4lOmpF00EW6TQB83GRnWr2XE3N1h
XJGQbqR8DYYcAC5rt2bnJ9mDCHPOciwoICICwKKlGAc4CKv0lQUaIziGE76rv3XXON5Y+p0l7bZC
Ibsh37Vmn5VEuw5hI3zLzf0UFPQf7Eqi6P18VLaVBQ8q++r+elOfBEhJpBoWqpyM/Lw9KlL7gABz
yoX8G0OrOcEfrtw29M75moQo1dL7IjssORfLzHtqLSGVtq2jlxfjW771STaGEGHHKWOW4flhsmgy
xJSZqRjBOeQ82kaL0ru/gLtAEcjYgs7QZV4HMh6GUW+r07GmC661hS/wwe4vP3HokY9thctrOxOU
H48Ofr6+cet9NHkHSPLiDx03wqNpHJB02Ruant9L91numlWp7G2V3aaEFJaA8IMcDGFE7ZJaIgfB
OWFo6DZ5RdOPPSUl9Mg2urFX1Nr/aVG4aogTGBvJ7lfNTsILph5pdKHWh9YrJTshPYzT9Cn1pTX5
HiM81QAmARBNpfklsU2CT6GRx7k7I+dxp2viaZdCaLUY35L9o9PUUJ+YPcItkWTt629quuVhTrwZ
Dc8kTiMg25K2hflBKurVpRqLkc0acCL68eT+fqES6djYEhoz288P8inQIh0M3b9Bfve0rvlQ4DSi
iUoenAdIIFfx2KbouP/UMrG6WXYodL4I+mIsKQQL6XsDJFIAXhN1j+isq5sSdQtrSxXQ2vned9ju
skLFuqdURRnFs46MK7PcGUJB1KqyePINMtQnfX+FUu2wa8fnd2U3veQiC2gR0kdNbOj9Wp5Qjh4X
+eGoKeV5A2jCduLZ+OLioD/rxtbgDXawRJc/+hOvkRQ5wuBmNcsiexAxfUSigzsYLduv+Mg92DeG
EihHE43lWSbv5/M1z9cqCS5X8aiRbPpCPmQrW8XqDu9+8wQVN5K/Ef6IjYgvJW2Eh6tpxWbk6OK8
zjx2v9k40vwfKFfjrZNmltLmO87BACa1ZNxOs3iU3fYOql1ZsACjpqn/L1BVsB37gdQRsvPSWHr/
D4uZ06L3MQKshH1BczYj2WGrgUImOI0iHXlr0Ob4uGUkunIkIw3HKkWsx98NnYuUn20n6zuMfztB
cmahdBHK8U8jircJYVqPtF7ePsa/u9dOAAK60xIRy9cM1l0bVE2bCzqv8SZlM7iaM/sgOI8ZZlxU
XMsOlY9vRK6nEp4fAvbT+DzlcfNdx5oWyCmRNnjT4RlIVu0bAwlUXM1wxFaE159t1BCdLts+PuTv
Fx7RFTaeaW61JWaUCD/3LCkZDlggOfM9/Y64Fwgur2EifH0CIxf2h2igkWrHPtqknIIT0y0iouG+
VzkTryeNnJ5i/nuqIP6Q+kVuQ/zPqPQmn8Oc0SFmRkcRMvtdQF5JMk5FYOK31nPbfTeUsUfYEEV+
cklY7L+PDSD12i6Gv3i4HMuI2ol1O2lru9XACPa87clJU3oq3J8qvb1hc/yeln9L8xpNkOl+yyRm
Qg8c+kY9/ssFxVu8VwApRYBTKeun1+iUjxAafpaHYEF+YRCk7R8vZxhhC+/1aAf4OOFd143rSGWB
4WQk1FR/cwpaqF2QQuDdCMaj4PRhMl35tn4a61/xtHDE2LtTYdd+dmpvKfUpNFkWxdHOKWxQ5fxd
r3TZhYqpdDgHEb4GjR1fIw+1Et3KVQHcrjh77eatSwVnrUITEE2nhdz+G9qA6scZglb+heZfFe5D
nrcg36xzxdtU8oHDi6RFBLq5ah8oX3o90fZhSkh9d7ZWr4K34vcpfN/vUV2PW/OSiTEAqsapN+sn
BGwWrTKvpC5Zu8LI/jaZ1PYPjcX+yRoEeguspF4UCTuRkF6vs+JJTfMWTMQqEn9/co+zUSPQgJoI
fVZEj+sfDsxPrhJSWbxJXmlhO76xGnmtnzjRVx1q+9kzRH8z3xIXxzivhaMJsPSEF+SF2RVxp1DT
3G//a8QnfgYBe23QvWhZ6pfeNy9c2gtx8vwy/IJW9zbQdVgsF/OV9Au5Cn5O0bmRUOnma3sN7ZK3
1q5EH0jZQ+s9Wm3eYMb2H698/+OSxBZvsTjL4HRFBX65nbtBwGBaWJGM8CDVqkSf8eFBe8NKPeb5
0AiDvoD+YDTG6SQxeWVZ0b/U3CR2ZQP8ZRdd/sI9LKDprZRP6nEsRGuqeayawK0i1ovxBJn6V7DY
6smErL2v9L2ijOZT8f3AUVnRQbb1rmI+o0PvKrE7KKIBXATMGDLj2PWpv3cS3PQvk42VUlZmaStT
rxZXiSd6yg4qi/sm0qaJh2lX9c5Ib7bEGvDZ3N2Uzspk7mAH5eDPEijrrsQJRsrECTU2adUk4dYC
mNm8F3V51Yzz/aUU5aGwkx3AHEsTqfkzrW+LrX04nOJnJwjJP4NKx7H7SaRhBjyUC8adNPmfowe8
clAJ1r9v1fLuCWaG0SzES0/gERENY2OlSxVtARng2jH7MwPluHeDMyPYJrbWHrfrTx4DwEo7UbEp
oB1XOFKIE6wGYqWDcki5xGmjOeyHicCKaVF7WOv1vbhe9xtk7MS6RHAblwEsZCWLe+l9+tTRmuNr
tQ2vRwfK8V78azrvM9dt3A4dGPT37612r5yLIw8/eA/k6OaXLhmd5aKwx9gUxqQ+FgJeyw14b5O3
rLMvfjLn3/rCC3u/5Dltppx8+1LNmtJWTlw9/BJLnq6R6IoR1kSQE8kQCPpsSSrhvLAgBn41Sljc
bbdXaYywBWreoDJZ0FMV5QxVB+3ApEylZY/TkdeWxYRlaZ799zP2R+XU18oWoeu8hJ4UnsRqEmME
+65bt7X5mWdYCggqjXTUQNb2TMtsf+owrp7d6oILSkXFVomfjs0RTdrQ2XmEXX8JC9kl72gb3HLF
ZLYs+6OvCVyzy3hizK+L98bB7xJjUAXJUFL9zJtCF4iqtV0d7c9l6poWEQcCeDNhNIQb7cwN60hq
pm6AWphd4Xy8ntR7rlFwrWXlIBnM4dByLWDSahkgH7k4uM82ovCd22mCmBOxVTLLF8pZ1QmMaq8L
QL+OJK+K71PQ8p7FiLwAvUgTZGHaLbi458ysncMr4n6pl3PQo+pL9UOnw/Mc94buQF/HXHgu0afg
8z4nQbbWX7jiFZyVZvc1+zO2r6O7JGNEArkwcBWnmsvDsabPudY0BDRd3DgEGoRDTZZiO6z1Nnve
v6WojicSvnLPBuczrTH6tgThMdUr3NJ/kjV5kGkqm7v9NiYIKvQhuBhpZcDP4yMGb6xTP03lXoYl
Uf1w5+sHQb4j0CbB//CCYe6+bJ0IcC1TxhCKAZOs8571Myk0dd3DBlaVQJUQTmDXbbJBSYxbUDZA
X8Xy5VEUZp1g7vDy24xjYM2bL5/Bbii5K6JmjHKLFsUxAy5N9CZw/SVEy4BW8Orp26xDQ4Gb0gwV
YX790XydjWxA1lDdMZvFQ9Gd8CPumcyhp1nL8yYBtp6pHFVAQnKCqp/GWx9szdNmt1WvqhvbesJ7
3mqMqYpkdNmQ48tUZItPC2eN/V3d0s3Cjia0CN2uXGtN+IW2c1Ykh5ljtIKj+XskwfPoAvWVSXJH
DDh1QZxNXydzpxgz8Sys+I/ggRx/bL5XM0fi9lOSd9/LDRum4V/gvjTIzogHoBN1IDoKLRKNCj3t
uNn4kf4a6njbQ9yvytVs5njpfT5lauddpRU5yYCvdEkjjfj+E+5OJF1TZsRCMedCySu+6WKHqJWe
NzS8gJSDcOo+t3OD26NlU+jhOysy781oujOmPdy1BkHrpz7nfWZw6pfI5Jf5/wAkKm7Mapb9Rdjm
04NlCk2LUC4ktZqQCPPMdzu/9mwja53Yf5sCY3VXVoH3FiemmF+k8m2HekCHJt2+NH2E6sfbP8Nt
vI9XzQRSUyi1v0rlqaqfdGMPWXe+ueJrLD0Y0qtfKhvk8RPnoBwzSEj4Nj/2uhzCSNaLnCwpvPcp
ai4G5EHA1NjYoliaIRTh4uF2N7Naky7Go5zIBO4+kcyybZGNJPpJ2YIitS0km4fvX413FZRMtMLJ
YL3JpvicSrE1TatwfNFWZpePPy+bs3RD36m2l2sBGsyZdUiB7dfK8LxC/BGbnT/fO8TKw5f73pOn
F/NtTyekh7Vvv3F8/ekn4BvcBdzWaYkxuOfwNQMKx8HrqX2u8OJLFlF9vDgF8fAZ4eFTClvT8O44
AXtNEgL/p0OKFYhwzU4F+zbPv2lix1C5s3xrwaK53vpT15A0xCXuxuyQrCpJjr6VohUM+m2CVQqj
OLATZ+e5y+1QaLnffiVDkpwcttlMuWnYOF1o2UBLnSD9I4GbU3EYN5dbyKb6+4SSY71Jy2nEiPy5
GXDwJjJB+p2oVla9Qti6pvD7UbKkKvE2Xq80ll0N0ftw86K+GzWO5x56nIDBGUWH4sH3PpHL8cKm
3XchqcOs3UnI613syPA39CCLLXr/orj5aSllGNATvItSIM8CsNUXP8kKLhJRO0N9Gdh7TumiGrSB
6U2iz+I+Lm7cQ8FVoDYkPNcaB/cUgX89oBwUPG85ak+i7jWAyPYIB95fAsPdrtWcfS5wsrX5KLDt
yXptT3ih8/r9kOgVPztF+EZtfOvG9o5+J4LxqEsuSeqnnEGTvrDvgh0FNZFkS5rSMzoGzZrNEPDr
q5USDnNgiAvvjR7igLRajr2vS1fNjibS2J2L8rj9s3OIZUXpG5AFBR7ial0yFJ1civq70WWtTb10
cV11afGtEHChk3a1sQSCjej536JJ416hqsix8TMr8o3lijlEfjgMBz69pmMKHIh0jZc3g0FnSkde
64f2B0wgwGuQBq5mvQMROk4KVCGD03BVagiBHXOdf6wj0v24roWAPr4gRJ++Dmg08jc22chUIeHg
dq8dTYLqt6xv1y0DwVClhIfjp6wC6AE2IznFzdA+TgiZ6ouElX+SIRVb0QnJ/WcxDOEgAhcXjdmy
MWoI2AgufacWROtMD+nT9seXQy45z90gLx7Z+8rgEUHrP3CyiKPpQYVdfGla/waljMgK5pUabkMc
iw4uhIKQavSneERSTq05KBeAGNujR3uAreyFDUbLEUF1Mc5WOe872QKdznh6KmV2Y9fuV1rvjO3m
5xvZACAmJW71pyRTdJgUDCrsjswoTUaCUuSChdUap8KSwuJljbvTQbOfzds3nWkNcrscj6QORyVG
JU7/AVFtNrWFw1tmPoHfgG58C67C2oar97Nig2tfhJoGj1uIa5Wyk2kauBqTm33psdcogAGYGfGF
4+s71Kcl6puwFdmwp/mf+Q/D9lpN9xx4ur1gSOEflGTvEJtYiJVg3mbXfYkzjQAgR+mRfxQO5SfY
yjB9uQnC3Fg2pRcHo3yVu3mab5i7bsiyA9Gaq5ZyzFqqkjHb4ZxfRZVPUcowb9UJfphx5500KONE
lJsblDkXzjSHpFIaDmKdNWV2DfH3Xe44/uyWOQbR6hfexs/SXxmTwM5I5y1eDnCVuksJ+5Ld1m4k
HswhwUhd8225vNEZoxJjYlzgtVxlwOb3wa7Hegp/m/4asNOw0iMoKFJ3FwUiNP7Ny+cFu5aRcJFx
p9IfdFdICqXLS7Sy1NttAEyGPl8tUmZIsRlyHbH325CzuCBOblfxmWTiyJO8eU2E49S5+oargoHs
jvyGnTSavWrNLfV0by1Q/vs7XClH0n18YzmsMSsVcCyFxySLolz6t3tI+/r+LWeXum9jx+m50mFp
Ti28U1/KmZ19mZhwglWPb1Rq91c3EOPfQGW297fq2UgaANZj20mNWU2lN/QGhNtVpmtKityDDSEM
O68ELyDu7KDzQ23n/bQqjy1rx+zz4F7tReQaVFtUO00OgukNlsSwhSCH5MDqaZ4sFlo1VOc0diKF
tm1jKOPivSXTiGjEFnicAacLWY9GfzEPOybRoRE9wdxjfpBEXLA2KeGKGT8245PzSWA3hR3Ca5J5
3qoD5LPMoB0T4OHtxdgeYKPgFnysO5GwuchVQjMCFFRU2ruKnghz8H45ixViQIf7cRs8BazbwPgY
wnstaSGWrHhbcLB7xebbLKdr19UP9Itz5/s3rq/z3gbTW8YxJomss0ueyak9yzz3NYruVGppdHVB
2xEtb2e2eH+/Gu7HJOWYmgpNGgc6It1MrEkI/M2TpVR/YYNmLsYurxTznFheJvAISprlWYd/QmNT
Z8BDh7NcngpSiC50di3vfJl/Q9Src0C/9pS4f5v+hzOrkxbVwu6Q15V4mCH6Vn+IrzoACgB3OwRX
hG5NjScdS2T3wPmEx/hhRC5wavBVETe8jEXaBP+0ZdfzbGNIxA8xUCXQz7KypiKQ6HhPx92kwMU2
BT+wjlYSCM/kFnod8WJTgeeL/CJ8aSOz8Fu3E+8jPMvgIfYc40etRHy2pEsR+wCKD/keRybtZ3Q+
j/GA6f3WgpkB3g4C8IU7YQjWVklwcaGkNJzugPVL8PhpA4vStHTXBZwyYqne/dqy7wSwFt+PvJhW
lhe2fstm6j1X/mvpueDamHiiiUjPHzj4qfZgMbN/buZpr9l7T5hvpxzWtJfTSDD/E0rqrnOzMyhh
p2pIFaNtFSSMia1206RdsKedp1Q78UN1iy1mVaTv7et2YxyAE80S6WUaJya9ukT17Lob/lZfWw8D
gfUCBdhgYiUbV5epFLsEUTjkoRAmmEuRBCNnnWICuqTElPNGilp5E5faHaQEMpwiR708mUd8z9YE
60mAamCcWyi0KwrSJGJ58xDiQZivPcFocHuCxNeEIC0P5h0eRpUlumlsdPNtXhovcVNbYSu3dmMs
4NwwZv3IVUHoMkHZ/KVe+sp606kYV9abxLdO7NiM6UtgtMAromD1qEj22v7v01IZ26Otz3sct3bq
M6gnh4DD6KzcEoCQceirT0GwT9CbWhS9PbCVQ+E2WhRFWdJOJPcYgVq23MlOC1nZtt/bupyeeTwu
0GluqtE7e6XzIU9DxbKn+KPTMfQMOtejDPXvB5t+7LBizRR/Nc8HNd45cwlMpZkVeTSrwiQu4jab
ckWT5Il4UCIfKfo/BdLsYZ3rck2lZRQLfmQmhvAORxEyyVJctjvFkhKKs+NDqryymSou1P6dNDQ9
PcWEUlEGgML0XCjGjMFl/ZJ/VioBoV6GIXZzZerLcs1doERRANXGFUXH8O288EPbrqo/ZK0xQy+x
tMRTTnXzbIlKMmkM7DDjwJ7QPKOCoop7nKkGkijTNqdR5AZzH0s6y4IvMUwKu9EhPkmqsh0qW5PQ
P7xAakSfQc1ZTdf2oLXvKQqt8Z1YI1LkNm9nsyDcGjrlAQB3ji5x2eX5tQ1ENeaoi00XUXvzBoKh
KuBS9mOS+Lm96aFGjALaNlkrMrOoSgZHMLHsTxBpPbgQMUvNQTz/rnkTrryxCekSgQ9wOY9rUgxU
BCw0nO4DIG0gjhRFApTGPDNl54ehv6jkygGl9CxKIv5jBNhakj96+hPI03O0bNcYzznL/KzhsGbt
kgkgmTVMWCxL+StOW/6f5zGEB3+fQ2mdtz8RZbp+5LBxv5F/P0kvvrLbcuTTHjVUz7k7g+r0cZ1a
s2zV7c5pJBEKchKteAoAr7DEmEGwxfaqKdonNi6louWlpHPXT8iwbbk1b0r9y63BoPpyZwYo+M3s
seTqPEVMNG2KvblOJ+GeCv6VXFEn4ld7YNDPUUz8Rw65bZW1W0PLL3JeG1RAC5aAZxqezdpIkPJp
x07s7glH4fZFIx+nJmxg9MKzcMOvRCPcTRlUYFjrwJPR2Es3ZXK+yePpM8mza4m6QGlW2c5jz5Tn
30yiAHfNdteOhHtF8jfmHBmYY+0mNQ8WMbNZuH1anMxfKmR9DKFBw3PkiTLtRBskleL0hIkN+arF
bL70e63V8mucYNIeN3wIqkTutTgqKJnlGkYt6ax+fu9Ue3f9DtKANxiT491dxGye5LNTWYrZC8GO
9Ry3r/GekZXznVmpAphHOwH1zniyyvGn4eOqK0bTIMpiRqWCq9L/CnqSy+iREnBS6Dg0Wq989oWp
3GSBt8SG3V7mcRajoxheuYgoElJ/uvnbuQvwHoSwU3/BHxsVCrlWD23rqKPUaPhkJUGlPJgsgzGS
bphwqnkv9g0kv14a9FAfGjj1osKymVg59WDsSDUe25bOP7UT/TesNxsmJvXR5uBth55iZDuVwryE
6P66RsLEWfJg8iH7ZV04aae33Xz8sQQ1bRWKCE4Env3HBLS7LQF1KR4Y/b/445r15+315oYlrFtx
1SLBu1bQ/bfw19OtDCOtaDt9B/Sog4NDoGK612Jo8nJRy/s55tC6Tk5p+oR18aXkMoGigU8n7Nkd
nSNTB2b82gvMUJ1JuSUdaGXvWHBi/SmUTmyt45uhH/0DtDB3W5gxCW5FkFAQKYTFsVecH9CAssvB
KAby8BYlIOZnfOGDgzJSJ929qYug7rvP6etrDESEx98axnOAhfDirwtxm44sUFCMPy2Zs/rV7VsE
SA8009QsnCQ9AJTLJf+qWXxNpr0cgpoh3JrCHsoj4Tvf/ldCgUPc5qU5xKIARVPeX3914eXXyb//
1g5qZaf8N5bIe0q49FKgU5NSxpr+BhHpAvVFxEjB+7Imsds6zmu8Ax6T0XpMmaOCxIYH+0UVbLUB
9UnlJwAoRbw16sjSHSw54IWQu22TpT8s/1iCnTjfvReh5pdIXjyBnv/o1p//DQiclURfkzA7nzin
lfAzN7uZi77BTTZiLT1tBMR/GTFX0WD5HKmeXwHm5kGDjF12LkMmuKSXDuN89BNB44T0sQ547y+0
pqSC8KSWhw4WXZ7RihETEutxTuaHBMi88YH27qnpfQySP+iXWyFPpKcE58IveR6pd0NE1xUgJaLh
SuS+gN3dj3OmI6JMTlJ6mFyDWAn8CwMrCZnUTS4MU4bbyK6Q0rpQqgBTii3yCkl2NY0xIbDwq4kD
XDEGCqBnZKlbbtKcDPtTpss2jA6UjhJK91Cv6eShOohhVclpXDPTbpQgHggTsbpSZuGmETTT3C+J
sbo6pN6bVppdV1Y3KdU7cyq+WzbFhfu+y9WhJI8v5KVeDfOAZJS3kC5ooPdXnQ2c6i9fEU82sBj/
LvdGatlMY0iqGz5+6p2oE6+KOBrFCXZ960PcnZZLRWYtqUPJIecdOAzcRTDk8wzD/Qn3gH5TtPRV
6gre13A65nfSVQCOsByYvkAwrHWRkFs3H6pTdAWAkJgEJez+1BcDELhdPZ9TgQLLOzd7BnZun/ZS
v1TgByLptA0eUFmbOGe8LF8ADmYyk1La91zBesUPrwewHbDV3yphVSamJ3XZmkQYK6QVzGQXtdKu
ZHSx1jyWlU9PAyyp096AiWNvb06pxLn+UcuwBqpfk+LdYAUDl6t6yHZiWcjPmKE/JvqSPa8NuKJM
RV4uUA==
`protect end_protected
