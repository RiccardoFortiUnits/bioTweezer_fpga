-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
haYepEhP7DxBC4gGJxGeSNpnr5IOwU6wuwN8XTfRzkgENxJhY3vujujK3nujk9rV+aZxPg9v2VHE
mNYDufpWyo4cT8VsWUOqEUfC29cn7RNmsDD5dxC2h6gtRJuky77OmPdOdDRAWSHJ+CN5laqZKzXH
ZEVN/6FkcDP49HtM5eHq893Dz1Xn07+lTkZaBMz6valRjzjFqoJ296gwdDzHj3konxqdzbvFuul4
fOWslR+Sg1bdb3pHk82yrBZ7RthR5HP3gA7tNmnoVYtZ7EgA7Q0KMb/kNwbw4F2BRe4Of/pXLaQ0
K367Oew7LlULq+n0dlZ5mjN7ZApmKjMRivSbeA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7296)
`protect data_block
e8agpmkWv+6w7yT30ht1J5d5+GLrSnI3AghBz71mRp3Ve70vPfuRfSNNCt37GDlrlF18YCenotIa
4FZqAclkTZ4lioZNILXbwu0KETIMH3DoOnP8lNOpsUwTUhaiO0b7xv+TqKbTw6QG4+mNXVSG/bPd
3CU3b0k8QOUWLxEPXSJl0cRSxA9eEZ+S11BhVqE2GQpkka8d7Sg7ixEI1k45S6Yuf8m01iwnUWs/
R3hdlQoT29An7hMqhBCraI9MP0AV8Jp/t2DgofglMIJuciX01kVH32OU8HuUnNJJxgPZ6/Ug9PKn
eroK37UDdckvdR5tUlgVMhJdL8WdvYWbiNCRXJ1ew9L1VxidyLW4rRPfez+sw7nKMhfIxECVkwTe
VD/BJBPdccBZkPJEysdwxZtPCy4KFoGKjztfqNBojJfpmKkE/gqoKetukj5WdYpdzXLT+uf7DSKX
uzQrCzHTZG91Cg9267tPFzaWbb1dfswpl5g1br9n7/AE8DLgBAjB7P9o3ICHdytxIn3qw3WDZEEF
TNb+BK3YZelwqS0UhuLwKaM5Y3X6ask7dpoXL4dyl8eQRRQZBiTICHJVZj7naWqGTRTY6C4nB1Nl
Fg/YQAE62jDvIj05aewUJFACOI9JUt9YA8Lxod+3xHkUxDOFaM6CqINEkcTdyffWoYU8YGIRgZ1S
fEc2mhlze1jDS8ThL1gIzAoubhsjn2DqYLW3MbXCPNuWAxP9eJNdRa1u0nmRbUbGoPcsW39VTdty
p4NcMoxPEw20toBGs1mWqyUTYFVMH8GV8hKLcJg6obkQ2+gRBF+9uZJ7AioCm2AARB3+cbE/i0eh
g1lpCVN2QxGNDkPSZQA5c5eGSNForZ0uLK8fQiJCK+dKlb+dTY009Lv41jkF5NCwItgRur9Gwpif
TzBGxXYYiNJD/C75FluDRTK9WnKxoPm/cdyphZZymlowYRSBTQjjNYmBEUcr/flSxbDvKojLJd7I
zu5kTeTnotna1xNbPxj8NZ1FIE0P9CrOl8O61CWMFsdLCjq4b+exmrNycnTrG9iIjtJAURKzQY7X
/B490Q0QH6Be0KPssI2RaassNUZMC//fEYu26CeNzLD9sBAD/lKH5KsuT1Z/ybPE+9t0vpUdsnpY
xa1C5/nFjUdOokiP/llz03NDudja+osJo31GxTlwgN5PAxtsbrURsaotUKHzSo8+elwB85dxBZTT
L26/cUKlGYL3NzXnesZw/lv+7AaCt5RcuHpD1nkawSaP27flTKrtXDGFS5TD5JsQYyw6o/JrA5ct
NtjeMaagk+d/4lQFPz4sjbh/FxGji6wML7z1trK4TcR4f8Fb2LKqpno1LzW9QnpG0l5V5XL6lhvk
QBAslUccSYFJhXJweUvNGAejshY3VyPmHzbLTlkg8itxKv5Q2QIK1/KIBCbLXOkAxC33ds/QqF7l
z5rwFtWpsMw4QVKRgqzzE9RyHH3nRzXxaWXhXG8tTd8ZZqHgPemnU1aknHJSfc0oy+z+yCV8jaW3
1orJ1Dea7AnJuSdlIMwmxgQrjgQkjKfyCu+xvN1i4kuUdvmXVNwTwyNNOr6yHk0Hc5T46CUuOgzC
R0rY8xGtZt/5wvCeKoA+ua/JVFT9wIfJAMU9070V10xVCLuz3XTo3VCYzuqJo15eCopGsaOk9h8D
8lf+jGFd32v9tTW5li5ajlqF3+MFQhmBdoOclosbk2aDk9bmgjhSN0Gpd9oBxUIPF8yyAjuCojiA
PqtEs2r3YMshlzxfuUD3miEiPloxVNnUloE0cwE9Weh8kNbTSsE/ALPQjFBkvdcfVZ8zk3Z8ih1w
By63qPtXWOfYQQC9YMTOskjrzyZLvgfyWnyn6iivQ/bE2moWdB+LTlJ7qKiK2+RuBzjnbaMtpoKj
m6Q9tnN0r/4Sz+i6kTIjrns9ktQVuzrWsLoFXi7OvCqH9YGB5ub/XgbqNsLxzPs3WB6CYX+iHw9c
FjCNHI8rN/NdxzDKaM/ZYSrWiNesQYms/Kq/3cYjSSLj6jA3VcS1ZV1fFVQUaDs7q3psWztVAaRH
dfvu+rjhihv8BNvBi39j0tHMGAAJJG/X1YW4APYEgMugBm+GlCWJHKtoZuUUBNbZCuODK7EcSg/L
1+YE81dcFf3I7FILO1S0yBucC317D7bgeA46+B51fGKuAh5kEDbFENQorJqYo2HBRGlKcvsrYZ1l
a/zPf9qlNV5bwgE7rIKkWl1NlhMqg5JC2H7Fv3LKqYuiIhEp47rplwpMcccnMLYNXJyjElbyJr5+
BBuJTmeetB7NlpJtGZ/xcfBEy0ckUavt2qBLrLF74lV9TacDazpC3MVx+Jbqchss0aMl/R9uhXH6
8DFCbkEZFhqUejMz2xxSDv/MtUfE21Nh3Z/IKf0KWhEgdQG+4U41W130fuTjQTLMLw3rQ8hh5Lyg
No5l9Lca7hQ5inlVCXTKzlV0/7h1KVpVUrLW1j4MfzLdjmFfL6Yq6u1Kt7hrjbRFVwILzbms0QAi
6WKo7oVLQA1s04GWqOKpwCV99gvFvML0sZF1WbYDNyqhOE83wLXvgon8mU6XBCIzg8mei5HBh4ue
vife7EYqQppTYgUFnpmXjpm00f+liZyo+RXQKOXJeNImP9Q0kK3SM0vCO6gjU7eeCKWNiUIY6FrQ
k6zk03d1CxdhwlXJpp8HLROg9q44BdcHckGaqmK5NgcSH+fv6T22cMiMQEizr1l6LYZABcSK/xWb
BQHJWweEG8GMKWi2pEWYx9XvE3M4Wc5xGuR4MMZQouPP67rQQdd+EmkT2rfvlqjv1YnaI3BjtFDC
mCEvSszBk+xCSOXlZPahmkAZyAOZiuTz8m6K43K7BIHN55wUmTbZRvmOFPYFDSl+G6P1/GueiZsx
rIoDqiUKpy7MSxfI1Z+w1cl9vgvfbJzlvRsfW45ed11uimtIhsxa9k/Qr8EhEX9NE6nff8hEgEuM
mSq+CKcMuwEEZcIthKX3J7skeYchIGF+iaLA7WT7vev0dgOLLyWPN2mi6koxcoE7Wb5yCuV8rcZJ
/5rKH76CX7v8Wph3+Pn6pFiSXnwc9r7B6Wrp21DffNRDJBw2RXtwQqZl4I3iQYTr9COrgt0tplsI
YaVJb4iVYLFY1b5vRP755LRzk8v9LXcSa9MfV4TjINxE08Aa4IuaeUyyBCH4Pt7y2jkXOlMEJy28
/xMrcov7z7hboTyEX4sOM8Q0c2VorZWlFjWAXkK0mqUSkXjtzB4kdXjdnz/tg/wLsSKLoZGeVTXA
FMmyoFsb+CM0yZkG1gYU9C5xPocmx6PeswRKQrU+lN2YbwktIt/mZe9PR+Mj/YIyUVws2RjFMV8x
m8itpBkqaomZ4q5D6VieSeNV4eIyPxBlewbyABfmYh0r4cUJD+qN6EAwnPHnR/0+RSmeAROCREon
SXoFQD/w1NkENW0Mdb+vk1FBkwGnzY5T3zz6/g9h25GwulZ+osPfWsm2CqGG8kNRFPjh3n3G29V0
G/bckSueI8Zxcqhyrv243vez9Hk+V1vfHK6EYeXhpiQPJ1FlzARWdGVwqM6WSVlNKB1FkhniTs46
xYxCuARk3Daxadvr4Wsfbfm8MiIxKY0/ax1WvTJySgErgkYUpZyDS8q9jwF3UWALw0zntRxRvb3B
y/LCqCpKQ4Rlg5OhGCKkba7CM4v6BkBfGUmnqAa3n74BXuwiQw1AFTfLwRoNAYCDKaSvAImBle98
3G1anG/Za/PnPQz3cS6msocNuDYABJmtZfYhPvyS+jv347u2f8uNX85lv3q9yhhYiJlsO1LxnmfF
SHE1Jcmxz60ocfxB+edj7OK2yKNCr5bClzWxZYfL1yTWrsQ0aMbGujV1f0LHnLF1ygAvWi8UUFAN
WiHz6TKDAyZMhDKYgGM5lZg0/zaUtLFjsldrXRKHCgCVaJ85w6+9EJWUNYVU6bwMuf2aLqiIzF7Z
xG+v//HK3Q5j/i+fp4S+WgKib5H5zlfwaeHCVwNaxrmw39e/ELXI7I4+k9nhHi+Dox8zFndFGniu
xPbWSuwlHHXW1l2yRZXqTa1IJzbXWhPzKIrZnAm1xZb7Kdwnq+/RSDVYiHFOinImC/1FTNeM+BxQ
UoDrR9NDbIKeWLWScULA+mC3alm2HPA5A6XRDVc4+c2geQKduv4alD3JZjRpISCivhf8jGv2y+iE
V0Yub6pG7M1W/sJmCeGU5s587yubJt0R2det+satEYZONTv3AKifyFb1OmCSlWjxLAulQm/BUZMt
OAIbkCbi/k9CWuzNPZ+1Ev7fFqE4LVx49LaRXuVdjMLopKVA6eJEBlE6gEcKi3j9F5OQBeLEO02o
2aTfkYR0KXbCyum8HForB4SNcTs6jHzxwvcve0jHa6/MdOTKWbcjVbQkciZNQ+a8YJyfsWh6FejA
mBisY4WpsYMfoR3eESzGDI4Ls1QzI7H7bWMx3Nurmxrv2oMyibqd2VqWr0rZPRgq9QjgLmJfCAup
UuQ2TMSU69vV6edkn9Va2RSodXgKJWFlToVe06mSKooGKMTx2AF47KdHuyHfRJrD51csyvcT5OkC
gP9xoaS5qnZAfOHQnK9giiFG4HpkfIgv28b7stCYm71s2e45ap9/ndLG7ER0ipqxpnEWVBPnMyP0
2TqwZt1ToJEOIHhqMT+bSVyRN879fm4TWnZ/uJLDnHaCi0ak8VzhTdDnBuVKjPeTaXgTUmQmwDFc
EXE7RNNWB+h2R+bUibfRoW/uwrlCxaAZahYGhPNSpR4klsxLgqjSXWvsTmLkzoZkKv0GQWagFnbL
EqIVMe9FpN04OVD5jMdRjVVjt/WXfYjMWWBomG4vPwmjIxiEWgL0M6eaJ25SqZ7H8rMh05vhYvVo
0rb1+jyTu4RZ5u654q0Whs/oEKyR2K7YwDbxF/6KvV6rlqHSjn79HsBwZREsgENp6TFGIdJ29Xpx
uS5jmlQOIloJcaVwSrf27hnGiWUpM5l5O14lmCC3g3P9Jv08ReeE6MLtkxmdAT8y/7k2gbmapteE
Q3gbb9ZX9TxGJNOAja34t8WdaeSYymQJarBDBFMQWlg8tvsSqwYb/PfHrfLqQpTiMNlUOrltcvdm
4CIkm0zeYb/IMU/L2+g0UYAV93OIqks10odADUZJyJ1s9QRGDiwuHwhRFmyVTx0t/OjqG4wx/59K
Q2RLEqOa6q8YcSa0yfdPRII3o2uVlpKjnYiOjOLrRKTAZmI2Z77rPqa7VB1W5A29FNfayzXT+AhZ
LAm9BukJg7eQljBjTQ60+egCsu1sl0EuaN3DVZCcS2nUC32YSNyOh65bSWxywXOyKZEzIIpnzRcC
wWcfpT9OPA66RFhHCGrCeKup8mZcH8U0Pzcj7rilzCpIboPHTBSqAF/JkzsUzMYdgmxZ7kpzh9mx
ClqbYZryRfdUgPWcYsPPGF2RICuIOLGpMapNOIFpF3UENpsEIFCRB0I3UartPcoc2+S5of4CMkQW
Nly2o0Cnk6qJ8Zw9H63OjicFLVzdyofIOnDB8m9ZecerCZTUvz1VhIDCL9QwA6oSdsl2I5hmlyVp
AG7WBQaVTIeWlSHE1zGwDvHUsKjehx1f61UeeSVZMPiAfhI2KWtwNqN67sIVkEgpyPcuTrb/TbPD
qk8ihECedovAqQnosSYqC8x/7G338wcgfta2sEouQdUDS+4TLM+n5HmsuTu5HhNreijWkxHnqBlK
ErhvcI4cuboYId6/I2TwbgrG8MhIdbDTuCQM0yKwS5tWFbBj6kXyue7F78iXfMliq90UgN/q/Zzk
XjCGi3BAwtB85ab46Uc5k19sAkDC06SOqmUst3fRqEmvc1C8wqlqdXd0zKYntzwHu3PGK0sWEZuA
Ca6kiYbeg53fZnxiVM11wLJA/7mAlRwvhr1rYm7JjfGBpnYQnVyK95hGckNqlh1uv0VQIgE/+UIC
EvsvKm46XPD3BHLt3bEVZ/TtWGyMYh3rqy+Q3wfd0UvbjoUhmhH2U3oMB6Zhgnaeo9srotYi/TQO
RCnWgnEorqOCd/EGpdrPUqHMx/z0FhGjN0ACz54+SJZAkwLrpKFil2Rac5fjb5945JyIPXZd9Td7
iEiVi5b3HuSf1F66PJWmnQzbD67iGfJ9AvZ8X1RKL2rHo74pdTmI9H4vR/PRw7+A1tpnhBURWUPK
JLW6xkjLImNFocyYrFzollmkgK5STZlI2K4XdMzazf3fMK8mPRqZGiim3nd+1TXaxbnlDj8YH4ub
WrxI5xSLKD3uMmFv/5fTho61mabIes1vptPeHzVm8OsjIGmDVzkLHz6c0cKCqAewZYrCFwjJDsVf
CZkFNIRugT+HZPonpo7ZpMQ3Da967pAWdqdFP6Xm8uKOcryiWz7bPgKYuWWuiGUpuNGcB+0BIGjl
xg2BcZ4YKQV8k9mR/FOT46+mImQhbqLMWs7eQKzby7HgJFuZw3eAEUyuA5eLXtx4k54VpsA+IleK
0Ac+phj6sdcrXN4OfaE9YSCAka2o7naBlRLKeKv1Ym9GF/2khxZ4iRgLXBlPg+PNN1oqIkNZfqM0
8hN4Spw6F3tQDVn/VgWyqAP/FHzXj/eOLi5xC88/Sfx3TFQplmkOiq6YW8VeRaPqatwIBlp/D21t
OmlWZUvCUp8AXahMjJH7DubBk0p06dKOiX1uQ0hvuA6wfTLpuerlOK5PSNk0t9F0Az8xx3hP4Z/Q
WaoiiVgaIRAZzG+vR23LTF++JSUm/PL8RFGNBmaTottXXTTsA4vMwjDEKzI1qBTpbJVdddGRM08f
oND21GymCToUTQ1idRPMQneBOkB4uXatN/1Z4autRrR/9Tkdygf7LGpIPDF8gSJMRe7vCTzbPNZa
vxl4SSkWNhj1HvXNUVydhadd1BngSQVOxjoprDoJhtnLNHwUl93f1e4QWPM6juHJKga9sWFMAe1E
NvtYFaVQvVC42MgF3xuAq2WkHmaIbKjhFJv4Nj9k/qHvIsKUcoFqQRU7Q8OB7LyJW1kpKfVDExuz
2kC5iANiOTGJr3r1Czy5jSa/LQa8UcAtgj8uMwWJr0dALDkj/yG8vxWmaoW7IBVURFc6ULxeI+0n
X21Sw5gAnE3v0NOAUR0UMfJioEDho5YqUri2GUPdwBtF34cHvcPe3ce2LPRk8EtfrcPbpslI39BE
a9zwLN8aNOuK2p2Vb7vBPdhAwlP4f86QPjt895Hx10mVgg5YL+NV7rlvrmwhSn+XkOAC8cfrFtNf
ycJqbETJW+2nDb2xwb6CeohgG4xr+icxshIoTV5NcUeRt2K/cC04HbDbM61exptFRuii1CSdf42M
dapGB03upr9PBCTUgS0CGDwkaDAAa87/Us4BbGCFTH47pEP3jN1B9ly4aZ75+Uorxo9u3SmUnhQg
vk5+q55HIrYgXtnfSpLKdWpNKIHIz4wJ2t5qWsR9mx2ZdKDl5wrRfC0xqiElRnqCqOpelmCF/OsB
vmsV2CA2DkJSMiy2nFA/kHyqbzGjscYM8u4mV9ZTQYL6zIqe82GHx7MLBWKF6poi9W3fy2QDjTEw
hLWPw8YOaAPXdDFkQEYmyVJAN0Xe6/Z+yoYihwlwbHgDnbM1VvkmrHpWXmvCtObNXKpNTrNmexDl
YvJuQetdOE206JJp8guMYZVFcvBRsktuBNHc0z6v8MRPMzvDx2Gql6PopEcS/Yv0drgV7Um5Y471
O4NPx0s8cl3mi6rEDfS1/KkEFFuAwkhephXvqLVJjn6Max9ih8l4Y9bOXOOeIn1CA4ChKSev5WVm
7Nk+8QWXYUVrTY5Gx3yIJWC/hxSPVDbfVkXyWy0AkDHl31vUdkOnO9DxdIrNuBh7SykskJVJrU5e
TWLIoyp3tb4xClaaJfojtcuJ9qAwPfHSa72xeEStV3cyyUCnm8VsGNcKpwHtLy/z6oK+tZlPCwfA
xNRPgAnuaMhJe+HBeaEvZ01ue3GcOb0c+MeIbSTLB2eUHRJVChmRDn7tkg+bylAYbqSDDTp1fuX8
grpHxLvoK8OJZ8fTNN6zEQg7Olr2Lasjx8j6/TOLTesw4M02bMlLZUHRliXKfOfVdbre7+9Kjn0T
1qXNiCUbTfTgM/55D9e3wgONv230V2Cg+UpZC+CITmy1GysYPIVzwG3fOaHNo/O3QF2eGyt+Qdn1
7Osk2IAy09tVs8sdEUXwqnGYc9GpncvjHRpToP9043/1hOVeFKQQCVxoRY9hUSig3wGen1GCjki9
F9uzYD1I8FNTLSkxrz3b1VstEkpdmUZ+qDNM2ZTanSrqJA/F1nlBe3MicR8Q7qvvwikJdAcwIbeE
pfdoRPYmSfOZaY9IJ/F1cq5kyt/NSNwAJBfIO8bIa80YPD1E8Pa2lqa37Ob35VMlUqLUIbW2kNIw
uscYRQrDioLYRw6O7JQ+ihzvg2CFFRQDRbGHcDVCMLy83LXEHbo7T2Rc/fV/o+SHGrUEskcEMYes
063FNsWGaFBWG3G57Qz3dHO37+zO+tGXzWDbpy5T7yaG4rzEnT2ii5fMnYvYbAqdNrZ4wDkc/5vi
jLq9xNEdXVUjKxl6xnJ5FLgaA4Z0qvtPo1tqxC4DfaDQEsmgva2/Y4E3LW6rDojj5MtOzFVfqcCv
rCy6SXtGibmrD6XMVTPKrEbPOIowKTYRPux4J7SIor5o5aQd7gdKVRJ1p2c0NjeZeHtDnKczVKuw
Warc0xdzIuI9YT9dTUQ/C445KoFbzCwPOJAmN9EWbQZdm1h0ZBBRX9CLvksTYbE6TNlA2rJT7tPw
sq7lwbKjGCduGdJzPfcaKWAokh/j7bd1kRZJkeSgx2wAXvrLjBElfJeC/zTfePEN0UF2Do3gQsT6
Raa56fOosVWMM+efYhXsvRC2WaRIGQqVF4XxrEEupLzzJi5DwIa/9D6rmj6j7JONnKcOX6fYdqd1
GobHDxp86rlDBZyKjQ8Yjxlw2Cb858MEhD7Dv07XSsLQ1RTO6ZRMJabtpW6o59xMGjAUWI0hPT+B
+Fqfx//qDFzubdLdUpDAfgGHc+k/bcC820wEfYxm1vYHDnk43mVx2iLjvhxpPxFbPrxBPGCk73vB
BudH3lnNVSTcdVzIBG/Ae9//WfM0z4D4bQ0ZENPyFIUzZSQiivYgq25+rq3hTHsP4vVH87v63WSP
eia6XRyfNHFUzNaa1E+KrCr02DYkF0s2L9iEA32cK9bgiUJUDsVKv0xEn5DhIP0n8vkJ/SFyidoP
jNFr59NY3zFiaVVZOcjORGRo9UizABPNM+aA5U5fgSJwJEJ2CmVKQcAyfQI2sZDnesT5e4QMG5TF
AcEkuR9y2o62Mrae60MinwZ/OQVvYCLxmj3zsSzzVLaElvx8VqueQ5jUHa83xrHvRVAD1BR6YdPC
P7q3mh+GW3PnUkU2BNnFuKun+18Xzh4ApJ2cwHt9gVJUmkYcwOQQh/q4rerEBQr7T+v+CuU6SsrS
jK0QrUhOldTMjdgTCZWNA6Dk5nYIoqcPKE3nNju8yr7g0BB0uZsl18CDqecS71CLO3sJQu45X5P2
yAgzrh/gLxoTer/yDo5Zi+0O6Lu9cgB7fenQL3SxLu3vaaKXYF+0lYQwbKj6NuOL928Bspqsk3Ac
dP8gHipot3YXEytjwxkqdsBVvQ2qiyIY7q8n7ev+Hj2sWUI6eZo0eTJ84+wVG/JtzVGU1FcVtEbv
UL3G5ax26n51UGcsjxuwNI2m89gJhIkV1OADRE0NN97bYwzwTsZcSPe1OMPMC376nDyVnkrQ9kPX
`protect end_protected
