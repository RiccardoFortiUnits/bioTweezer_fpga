`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bt1veyn3NiNV9owIXgwVMOGaeLRXPx9wgStu7stggUw/OisF16sGahz7qhglfUsJ
QQoaxTSU42gYltgGqz8sBxy88dWEhZE89uCQalqzG8m1Sfzi7L9OjJ80Dnt8nhyY
L2+BGK8qZKXzLMR6e+G68HkJ3JLm28fC/nX3C2hCT/0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5648)
ybpimnhMjQyhEZJt75iQbzAI758ZZuE7H2ABR62DnDoiux+4qwgPF6IC/Bxj7iu6
hr/oZmDyykvJj37SzJldU793YVKmBAXPvhQblHdyAccjlujlM94m9nM5v5GE3ngc
F0UInNwI9fXXEykfp+2E/r0Wf9ZgBFwbl8RIBCXQbMAZQR73bFPFGtIFIkaLNixu
5dnmx+u61kPV7XNavVy5B8LCKlbFxb3QLMufCz3vfCsSubqFqY4gSJOglIYUwYBZ
Lv569MPOHpsR0UUbsYrzSDDZDZaKHqGS+0NkQpjHTOTzvEVTn2sPrwfj/wVu6akL
6zQdxpoKruguy+RRftrYAVyV5l9FBBSDRtBL5tfV6jWzJSejo+dEZLxf9cXIBYit
nwb75Ph5u9VK7p4eOPpUBYAwPjdqJEHlSvA23UfMrJ2rIXTHazJG5XaN2C+a0gWq
koj5grzeQQphUiTFl8E5U3bES9ah6CEz22Xi+tcwIX9UVWv/0QDwMiQmctfhM890
KD7rBJ3LLlL8UsBYoJMDIEb51nEe+mYN+Wh7EGNNZfSkF6AiilYnOpq79oWdhuE6
ZXctK9UeJNOW2iKq2HM4XPbqJva3stuD2AaF+m79i0TFMqwIBbY0/t7tFSRSM2nq
BCsKzcO9xqGcLEOXSjNGobOn0mq7uGgp1B5GMqiWA5utTVHlyfT5M6cS9CdYZXfk
DwufwnXtFf8PUIwSNm8lW0TX7Xwh43kewk80xCurK/+AWxg4Ft8JUgPOpoFmvD7f
08ZEBjvIcDPeagRO13XarDkakztfcwdDZ/hWPn1sakuAvne5ET0VBzAB6XMXbay4
47Ky90R9jacHT8WUP1Kj2P/BmOCeJQePghAt5EfZweJrRoyq+crNCQkrRZ0Spz1W
KKJJ3DRAhRB+V3c63ItLhdzwtU4oz/bgWuHjC77H0dbk5tdwU0qu/Sd89TiUxO1g
HyeZq3INVoxVfZqn0iw1nv7BTI8UcoZMcsU8Oi+vvmUyD4wWEH2RIpf2qKYBEHWI
Bqe+5aIif/A400+Iun/jvBqgk0eZSBuhzaFRgypLbp0p5OaQBs4r4OgdLB55bPLD
NtfyZa9hFIrqjJUrmwv/04hylJBxTJR0JVxznpysgsAG/F31+9+EX8bMVltja6NR
TrvshSNbV7GYigjh4DniF7ewVqGXmJXiSpg0CKaI1bNKK2cphXbDQ0LWGDPh1tqz
CLC7esRXJACHtfwhUzk9plYcFBvj9DGhXhpk/xysFp0MYSd0h/ly3hKwyYtFKsRw
G/ysKbRRTNmFRTSl6JesLPQb3VC7kxGzF54oVzZrBEnk9pNV4HFwVrLbee4FbXcJ
VI9nOsXRuhlJRB95gUm224Qw3xsQil+uFYSl/+3Aq1D8Dn2CJARBq8dlQ5T7pcmM
S8giTiBg03VCPg017TK56gisKRK23GjR/2c9DPtZxRZB1voZhoao58uVUTaQlLla
04nufEkCK5FJde1+EWIGYS38CTRp4ZN6fOpYguPaJh1d7Gmv09UFx8qPBYWUe7AE
h0RR6HU1o6/Ba1nyOcN7tgXblQRLUBPjg8ci26L77cOvhYjKrVBo1Jq8KSnvtjWQ
CtNyFHv0POYmvdwHDHF8k1dJ3PL+x8gmiEU7fDmIbe4CsLaRahBk4UPy8vudFHhz
E1mCpndc2RlFrPTJD/GD7nn40OTn6vMg9SMs78PHNgBzzEmphdx/4naDGYa8X6ta
eq0Qi3nB35tjwU+td57nojh3cVz205tvet1RxEu6MG+la39nzTftakLt31pqubgO
byeloRwMR7sCckql150EWo25/bKcRxrVC7qzZlsJ656oeuhkRFQpatYJeZ1iDrNB
tVhldm8RuRa8RLd/nMhuQ1ayXmCQKsWUGiEw7X7TuYruvk8lCsDpLnsJIkVhaRRw
v+IFLJ2zg3vtDcc8b8qknJEA+KkRb+gEqxvoTZFCLxXXrVJqp4RcAV3ZbwFpavpZ
Iwo7k1kY9SiaumTlxtj0Sqpgwj0Edt/NKuBVJv9hF4vnrFcP1vFUXLbxqu9EHddu
TRN4h5WBiLuNZCzvyhC2GxUlNCNaPYBcvh8KR3y1V6EDtHAgeDn7w3XYiJ3HES/X
YbyaYuX+zsWHQWfwJ/YhCNJ+EEPFqjtYgIyizFOn5sgPv7ajqfl8CtKbKDl+42wO
8YLfJY76lYZswUQ/ACQq97TOKgN8a8fERTGQEmLszhNy2cXODU27zZD79eCGkWXZ
sST+oCxDSNnPxkyq1UfbsdFR+xxsEaL/wc4g3HO51rybDgX16Hfcj3NMPlLgwZd5
4FBm8leYLSyGqDRJXhzzGxZTNnk00Bh2JDo9j5gkCpCMmeBx0pS72wl0fbCH0KKj
ZrcfGfu1pBvteZox1cLfUJ3a8HvJhMo7FNvU6lywS9SWHTTl+82TLCRNCzfthQCH
1ZUJzMZs/wfFUzRBJR4KCAiSh/VjCGwv+KvWZIM3tehvs6fLYE9e3GIBUE8h/wy8
hTpK6x5yvXtstJm8a1VzWdDN5Rhte69dXro5hyyi4avPn8c8VVfDml/xxGEkDbE8
3+6+ApmpWArW7jyIDhZ+cwG4dnp0QqC0e5pt8cjM/KMP39eEM4u1su027uSmV3vJ
6Ls9e2WKN9XETfk++u/E+Tf2vlW5Vz4qSmsWHWWKp4BqBax+HWDv94x5WND/k0mq
iR84YTdD2sPf6vRhCUHdYSapUOmKEwZn9hYp9TbM7UdYB8fX0YO79JMCA9z+sTnb
UbJt+hRJCUSYo5t8CN+XpNb6j7cQswKFAVjIf29pQDz1i4S1lrLccx/t/pAqpYzS
xpxbxEkVVavLzBfHXWzJ3NuPtYGBpNeBlP7PP4PG2L8WGA0iqljvEoB38BVy3vta
XjMJ11B2ew1pCy8L7Aw1CaGaUo7Fktt9sEX/No07dtrIlD0z0LsPbRL+vrCkk0r/
wrvduSLGUGXp+GvwnodpjGIEg3t/I35aQGbua8gxrgAlbq+6dKmqwStOUY1u0TAw
LONknpqUJBiAf4UBBECl4pkIPVMRlTgwx0yAZG+S0MbkBvuw1BoVKNOaILZAYwjP
rz5kUCgEG5uu2BZjf7FO7v2UXGhNh5Pr0WAHC4A6pFc3PqkSyFmSLukKaLocSA+N
ZUODAKyOfbZvIT87z7gQWgYyBIZAU0VILS+uWSboMOjzrNKQPALqlqgT3SkKyQ+9
D3+hqiiD5RLGWo7XlGpKFbMcdIWCh6MHUyy5fgzkSFQLAM/WC0XDfiLvHrYPINe3
D3q8ocHtXhJkfDrDDv5kqUWWoDedJaxZ/CWZnA7H/2gzGf6R6jhJIUqTWHr5N0D1
UkxX3MvivF7VyTUsnbHgY/BWjEWhg5lX3FnJSaq1aAbuDOHSyrrD73qMwE1UDCbn
x0Q9aH4VOsQAIfvdNnBCip46I2VTjArt4HuIaTdVjLtA7MC4CTKM7J9v8VGGisHZ
/Pl5z259CRmCBP7x5y549SYYrkm0FyCN1ab/faKfyT6sdVJUh9G8cibGSYXVyEuw
L8PUegMOsoldhpFewIcBx7fgwlemAMAcRwEm8bKN4o1nPjDtouCqw2IH0i31EFjy
xEdU13Elz9XcbtzpP4zLb1PsLRes3xH1SuOGNrNfCPEX9UzofhIxegT7quqG3lGq
lslKL3RZttw8idr1hZHf5qdsYfjeHA3b3zvF74OmclqTQpSh9vML1vKokj2mWPPe
cZcH3IhZ5MPtqJfKCk+XC+dODTWksEizEVmkvHuHFOPcpWOm7Bzz99YdRalkcKTV
OY8AvQjyU2Ck4bncTa5ke32CELY/CqQMJY0Rl4LrmR1s7hdJMlwlwkG/x+ARXev3
A8Ltd70BlKrAuehKyp+/JQHPnYxATmZ52bj5tu/ySwBcb1uYidUcZEfRVSH+eKEF
Daw4DKNkjXZo2lKOMrfcFwiX0SGtAkXKJKZRqGZgUYd0OUWJSH6MOnVQbgjuLx5P
g4UmGMjevPXAmuQ0KthrrU8i/VpcStlR0iYuBHO3GbzimlTFnnJysWqmoMmnSEcL
StGR7oWahLgWxWMfXAeYF4igZzoMZ5sXxXqiNUcC7i8ZkzKwFr1A6vvVcc3CBXHa
G+Y09wEzDcujYt1XWSTHhMrH+XvvHpzgbBpqbXMmuZMqLEFfR0a2G2AglHFO9ToU
J4w4KpjtCi9Mghejhxl69qq/HSfYCRl9SWVB6jn47owtTNujfOt2bULSaybSa+hX
4LEs1nCcOG6rVbBkGyxJtPqtd/uBJ4j/qj5cSJpiPnAaX/t4aq6Sb+S801TQkm6Y
xOIBK7bBJkKNeEFvFeIY0ceB5qUNvgjs7nTkSqytxSnEANUzHT7C4VjI2BIS40zE
oL3oiLSYVBd9OoTr2ohNbOeX4Mu8jWV8k9KvXqI3RRjfLzFAbAA4S2hV6rtUrmdB
Rw09Y0ffttZJpCZVQ/3uuiAMrBrYp8E13IfIRIfCaeQVFjucsghWWgbntOBnJKVb
ZnTtx5VgVMcbp+IO3xaKu3lOcHEgxfCrcvNiGgmfuTxo6NZsrFgjgGyXO6n26B1T
X5HuQPrY8e9wHyhhMgh9YhrsWbwd/rsQKVzABUXGngzo9IL4AHZC4U64weqdAmez
3WEF3Bx6eNTfyG/sWbNv6xY1nx+kZsz9y3KOZjvN6O1BO7tCfvVmhnpoy6ohbLho
Y+BrbDX//mRnWyr8qEBydrdm1IzsH5EE556Jqh9i07F2Kvj9f/1KKI12RDSKhuzK
3R6HWsXPfDsIu7q3YGj/o/S+H2NeP9cfNWGRna3SSbSTnUT3K6OE8BJ/4TIxb8it
3Xs2moRin47FDemheQYx/nHHC7qc3duWIEGf3/SO7lK+gycwgUROIaM+IUaYXe4E
wcc7RRIXmjpKFfT1ufkEKGQhWxi/eL/xHbit6K/J2gs9WlzuZRJsoC/QnlG8HcMH
W90zStuKeMhHVATaXSxH0UdXnaZj614GB/tsnqkuIe2WZBJXxovsGM0QUkdmzOmL
HpkB+AfrglmDvGGWq77koOISsTuNP4dsX9LVBNn6ju/cAOFZgRHNC6ZzOYsPH1/W
XT46onwUQEyN8b0TZ4VCQV/7YDAtZtGzff7BAGp63edIq9ou2oN7K/p7dGEU8o65
z2DBG0UssKlxhRvodu4Njb7q7QM6nrGOvTPx/RIouFYRbkFqwGYI8Xo5V62+1Pf/
VtVOE/NlRgOzkGfd7dDObc1or0rqIMdH2KcHI/1+ApfPcMgv6E4ycZs/BufAvdSc
TXxXOjtgt/D+1aVZkp9+Utkv3q6PmNk9mSbBhcw/Ev4VH0uJCB3FUUtcBSzcURv+
zxzfZVMs6hs/15d37P8zAG1mBm+PaMV1QhLmLj4ej/NI3BpnbfUemcqWRVtCuEL0
ftI4+Vj0r/kgOWi92eYNOPM+OJ8AUQolQzQeKN6en7NAb4aEdrMZyOK+x2/VB037
Qo7Cd64pmwoTADnXKdNbOyBQXbmO8kYS3zJZoEEgjJEOa3cd5emR8TLiOfq+MmRI
ELE73GBxpYZebt0h3Vz+Key7k9YI9OAWasj34JCEgonX1Ctl98UMvX0iWbhXzaJF
dVDNTCfuj8Eu250kNhGUqxGTYPrPSEME3NY8fEtLeIch4ykHjQ+nw6apeYON74kD
UljVO0AVozzkobYn1gKwbwAM6AEY0TA2/cVygLbSRAEmUAXKg+ZPt9h/tQbqgV2t
z0AalmzbpvoiJojraoTl1KSu3WzjqMFkC1nDpEaNvdmLJklcx9Vee1jLb1LLnvFC
isODiR1qitriCy44bmIYoSIIvVjwk5I677oPuQ7SPhc0PiYYKLI6+urfE3agoVA2
KaZCpGvSbhHr0wb0wxbQUdh5zlT4XFeIufIQDDJQMWQCYo/xoCBuR1Z+1Q5Np+Ub
a/oK0qAbOsZQveRme3Kepw+0c/YVLTjVVGEEwIX5JpX3p6j3Ip8WbjVTSpozWZGe
xCrqXo4C6/TB1JuTCTuzpRc1fQDBkImOd/fKQ0Bl7lkp8IGKwtXCgWAenjA+MEGC
fhmUV/V1MEN5hwN2ZMe16Mxo4cC3/R/ra0EhRx6n+iBaosVlu32p5t8Img2FX2zy
PSiQZ7E7YCvdJZ3xl6K2vMhQBeikBEWyrDYrKgEP9cfBU3fE9JdSj5YOEnEO+bIt
keJjbK1AUj3bCcCog8kKeGWsRycc0PBq176yVv/zj3lyE3K+accaaSiBrVIqdQfQ
pLlwcGhcieq8GLk1r2c7guiwu9OCwbP2eSgUvWZ5ERbYofK9v2DyKKOEr/oZFymU
2YAbWNPg4uP6mJtmIXq8U45Nzry/QlgrVjKKf9kGDQ3lgXOhLfPunweCeenzflE1
fjGCI2EavTUAAYcerf9KCQBg/wH/qD1j6RSDhv+VwsIRUxS2a7YgGq6f9jhGEP49
RV73LyGeOx6ZyupUKmZWXeHSIQ+P6aljshAC1KWjCthptN1aOUd+qmYd7uv15YGj
6OsIbcNSN1g8mhCzGAo/UTE5j+c7id/IiD09/c90CJrPHwRojT/6//DVBL4bJpJm
sSzylkPiocXTNVwtY7o7O1Fod9rycqukkRwFPxju3yrRzgPf7WsIGKFeh6/pE8Lj
0kfPb47QMnyn37XM7NReH+nCXskJHdezwzlJT6nxPh8LWcTAn5cTY5cGoIkYxJQp
AdGeeUJCPbHf2F9uXaNSpi8/kbTuM8ZfGDylKQ6T7m/RzJ7YXEhN0pjLrKv2Gthk
II5KxFbjBBjAUYpv42i6FeS3Xrxnr+Zn9XvyKsyHCx1io9pd03aZZBRWMkZtYvX9
/x6Tbkoy2ZIDg37MUbMzhePZTKSr84QiGKh6vlYF9mXLG4cAJH3DqFdjRr3LYCc1
dL8sySfUbrDZoXCGOfyU68t1FED/zYO0Ib0D9d7hgyPgk/dbJrazwYzOwe4ZJC3A
+70fkJwtk9qtS0atnzkkCsnvf6ud1EbJH5VlqYHtnr/oP4hB77zDFdD5FdQmzaFH
9uN8Wi9oUd8pQ/kuRCNsRpXZmarisSjdy06B1jiX6vQ6zmK8vlMVekGK+9WYqtzs
eCQigshxHMyuwFr3YbA07MwAZkRPlh10cvJiU5upVNHu/D0gKl6coJqZCE/0I2xD
/Jqj6p+5hT0khPX8it8Loorv4MAL2JeP68IelU3J1ZK0/RZfBp4ifulzD+tzT4u1
Qk0Q6EaHfm0T8zgWTvzU0o1SYPRZlbOFZN0kSCWK6CeBVh3XR1ELH0zDX2If16bw
MBPeIG7HVtxE2R4YvQf+D0mIptq2LyKXjaMjQDG4QM6X71/DiOINW07xev/0UevI
p/CdnykjvwTKjn6pEieElFhHEMVCwgiB9sXlzMmZyyBIX+8sjb/fvpRHGDXzyYXe
dCjQSntt/WDHgKmqmlR5xXR+AJyC3BDLBxvRFJxkA05CAUdt6w1VPqoUknRh+xGj
WD2eRyZG+SheYkSfvR1ZdhSlDrutq38RH7fXRJwOmqZCG2ScvZMD6zYYdI79ySx2
iWe3hr8R+AF7AfVzqRbGBESj6ZjDw0HpZUgBEqrmskU=
`pragma protect end_protected
