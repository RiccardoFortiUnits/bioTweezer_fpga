`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WAKwnW7XGBoxsLYzLmCTIe6+aPxUPoW5gvN7abBOA3hdbVgjj3me16IqNN1cQF61
bvRX59JB6k1C5n8ozwDwwnR9vIQQEQPvd9weMtpps8Jish/hp0X3BtelCO/fNmoI
XSLI0YkQ7alv/BvOvOXskM5vPd2EPkknnP2l8Yzkbrg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11632)
Gy+b5Q21pFtal0pBlfLBiT5Guq1n9dHNcneg+doaModF+6L95vnL1nAj/Sc16mQF
vSWfL4/rmn02PTjz+Yy1EmIWbHD91oqzKi78otU/8ivV0GbyqNF6rd5ykWgHEfyQ
sUfduk6i46iu3tTrZtTIFh2ojmz+2GV5KelnDLA2GwvJ8dhPds0LfUNe4I4igvDJ
ScQSzlYudAY3YngfTPDXQqnk2qi9qDUeKKNGuNxDr2jnypEQtw9P3bqIB2ihKFkc
cbj8LAKrMLh+4yWrokuLSt++6H4L0BQCPjVHcG/AGtWCnLnDQlIZP8QlfOVHI/mT
0VCib+ZE8i7XPcEBGHv6B5l2VjkPBEGeJGneLfYvMMXtpwOmf/Ut8JroaPgcAIIB
L9gtfk7EdTP3qqb698niiLgUmVxXFs/84nUfGjT192gIQhRe/NlgpxO2VHROej0S
R/0/PNASHyAMG97gmxrS5BUhrIfEReWyQPRPmq9Jv0VZj3pFS0SvvkEw8hG6ns6f
dMr23jcv/xFolirHQjD7MptnIgNghkdOqMSPs3MOHi7pF8QmQRr6FruFoevOXvqS
KkhJ7JUfUtkl7mn0jcp+V34cbwwP8YYG8CciSzVAxb4pVty7MRdLz0THjNRZ64ts
yxEyUcVqUz+0QYN9Zknzi6ABY3zGSGCuWbwhFy17GFBuFdMaHbdnj5scE2hTF5t0
CXutQaXFlDAKEZ4txTyfAUVmsNMv/DHBE9i6OqYxA0nqhbyqaGmDx9cm+fIAJMee
lR+dcd9d6xMkNYS3EYfhI/kGNkvO2MNgVuhu9NGG6y6OwSIG2T87BUeLorAmQbWl
6jRs/zOTXUL0GPRKsyQVYfTgd4RTEotqFrb1RqexcWEE7JKIL2f1kQd13ZZpOOGD
UIQ3z+Our/lfoJCiavHgDzCZPPlNazlhCclyiOaFcQufLwuc/s0PXcbL9XcuNtn6
TaxdhKvATXU0LZyXTHmuyhYPvjPWNcRiY8wjnAziaWuamJgSVjRQE0PUlWpCvMlC
nvoxLE3QIkMn6CXrWOtDeBFDnkSpf788H7OSw80vKve0ydpI/XbPKtcwa5FwnO6d
RS3kAQEGcltotAMV/9EFkIgzwRr2ACZ5fexllvFcKqX9MTNz6bsKfLgX+TnadMZ9
b4alSC6uiD8DfRlcVeejWPi8QCY9XCVged4JmI8w9R4l66Ao9d85j7fondX/R/W3
rOElq36a8UjsXsiOM3iX5pi09FcA/qxghLjtnihbkAo6baNyh6PJoKBzjHY3xaZU
/McgO89X1tMQ6Bk2r1BtRH0Zn8c/9nQt38h//6G/KNt14TziClNwvoi/5A06Lyry
cQfH3bRCV43cJ4ETKxhXo84iWhWdqEIb2X0h3dtyr2Y7RTzSUpSf43GQ0dxhimev
QniBDVSmHw+cKewPbD+/ByVLdkJUksEmRdz5CCO98lEZCzrgwsT1SMCvYJzSu7Dg
BgqIKYK7dxqIF+JIs56mUs4jrsJB/nyPqg1laQZ2ASYWVK63AeKAEO46WR5KCJts
9PhPrUx6TQv9O08swjT3R4HSOv+wqc7cbQCCHocTRAe3C1DTxKndw/b4qbvGJjfl
74sA3OB/m0Rgn+ceWYN7h6Jb8b2FaOzepoWSxtr9njQGe6raZnZ8Wp6bTRWpWr5a
9DcT7X+mIongOscR8hUcaVNRJoPcvKSQdAQ+8p5dSCMZAMc/UNwg/ml6erO16ziI
kJRcFUyC05kDiT3yPGDebZGdyml7XdfWBGuBNjJ79YboZ1AOAgXfyrB7Yq5YVFls
iL7LCm/crm/gUApUoBQfkaaJopH4zOmMyWOxp2BNAhTyagg9bKnoHrnPDBg6rZUk
wQZ1hf0uDxmHqilpzB6d0741G7gWF2wi7sEKf/hYWmvcWrHP8SXW0a1WlbRiCs3/
EplzN3OubiCyfZcTI1TVFYoKWX6qx9YH1bRIZEUz/Q7tCy/qAz8MviDVIbeKOcDm
6iEqHWZaJyqvzshH93cR4Sn4NpZRGPDX/bTOWs9r+3SymJsCMEe3/gtUdTlX4B3b
XK7RkGqKWKUll2PkPeFy2twJTonGE4fzczTrtkMUROvJ2q+I4114HDwSLOZ7cwyM
X+YTdpfCkDQTchiCaApkhnpS9egrN3AbDdNfLPW/Ua9x3K6nkT+opYgiG1X1wt3g
gS/c1s+eyPR31UxUKkCD/QuP36/gYnYobHEOJ7XDJgJYN1TlxxoIypcc4InQ9zyI
ccUYWcudiS2ylIfxGIcWtmGYp/rxWODho3uypGirxxTh6w/8/okXn4o96bNTOzPy
cy3JCLZS5YoCnyUwDAjsmwDkU1ZdzoLRu7F8reYv/eZbG3or4/PzU5ovI3feDbIt
yFmmieRTqXxtvl0JrHlOGba4PRNjZAaY4IUFQDuRfFOSo1wWKCmMlAhEDVcWkFWx
BGx6VLMmMku6ylOXC6pHjSQtfrNuojwyd1GzPuH0TCOUolV67oz3MWWoTdfIRg5j
DAJb+NhPO+KDugEu1tOzu8HiM5iTTb6GdsAqg66kvfw7H8zRUjKMfRu7x1DbT2Z+
3SQ+AWkgdVPBedzPxQsb3Xtmfs0/F5WFJzskqxWz8XbnwUs0Ox4Qj+67YqOXEYRc
AdkdC6L2sXfbd2X7vwqnALtgKnNneWmlApL1dXyrG77kBU01NK+Yn6DKRHNX9bUh
8fjpIpwueKKwef7QY+TiBep6+x+6oE1DvLScwgFrkDQEtZFPbHMw6PxX7oJO1EPK
hqU+8h5zCSrecd2wlEMmbDdYAWVYeeGUtYbbJtuaJ5FczS87/IHrbNLOx+vk4JGn
FCV0l+x+piMdCYNucIm7a2rAeAEw4C6PTGVpn+fP3t/+5++6zJmzsTti1NN98JA7
euOUUhA6PLPvOL+uvEWxaUusrpPIyHjDOL5la93uTFOdIt3/9JHO1ecP7IMkmiEs
yI31q+WXeMRq8XzpVmJN1KN+S1q8ow0MwKEocdUmYMftlfAcJ+30fuzJ480zPRYJ
CF1kSVJUt3In2LDmC15mbeK3XXWS2Ee8zCPZ6eUBvRu8IU3UEiiBNc2Vgy9+wGJZ
gObqynpkMTMyGUo2BCqvAMbfamEg2qZWJdz4BdOrODCuQc5I85+pfbyI4IUji4wz
tYlviOyx5ddPBcDrZxz6eohHFfBPgwFkztjGqiFpY9kmRpOwpEc6OACHAbuKtfNQ
+yb+DaAPBSntzHU+R3spzlUbCFlRWkT3TbVq/w2qfmc5UWEam41ErEz/B0v3Io4K
LOvThdZofiwTgW4xe9nmVmL7lJsyU7Zdi2w0hVqkoY/ij/ywN0MnyK5Hu/2EE3gu
9vf2b92a0lfzHyKBXPRU+fHEiEwGqFS5I3sVGoScKbFJBA1nQO+nG1/EEpAXyFMC
wOlgHx4aEV7jmBNxRHqgbZIprIRYUNa5r9fFwp6bJ4kxTIKRpWZH9MV82b+2c4sv
PmvA0fcvX+8SkXy5wPgVO0yPhXEYV+wOHMGnp7NITNqJ3EfrbHxDA2tT9WvL8vr9
R5ju13QtxWhBmuZD/gHSRALFXp+Mj094PmjLlxgIU5NOEZomr/GDwIJ71N0t4fN0
6CrRgYdvQ7UzmUBxuFgmr/V8+uadpqi+i/X4tw+u7f0cqmF44yMUF/Dq8dp8nqs0
jmerlh7BlZw/WSoRntzWLI1uszXv8U1Zur7puzKcPtILDoysaTmdWkN4qVYFsTGY
bmX7Dq3rrpQg+Nhb7iOq3VMdJPOR6eELM77gkZSVRRuJeRQXeAtoshwI2cdJRBEo
N1C21ow76YPp6Euy9edVUwpaV3URy8ZqvEbK7hrBxUC8YpgNS7LGgdUAB8ZuHBjp
PYsatzMj1j0UosTjQsZNALBRkWF734ecLcKVLzelTjAg2xyxgO5ZDCuzp4fdPKOV
O8o5j43F+gwGtbEUonwdd26AiJStZA4wnxjelpXyFYI4OeuTeJSWG+UWc1RbiUzQ
0GwFF4gxwp1y1jOdECPwb/6iDWBUUlS/YZdWeh8xIYeqsixKw2Ga5cBXGeZHh45l
P17p5/Ocb9r0a3P7XrRxGizje7SedIyJ7dhoxOwWbg4OK/p+dKDir2Onxxpu7odM
ZIqI3+vQb64oRzz5AzgF0klzTnhJnPgZKcOLaVoyhVnUT1C2X2a18VYHdzqW2acX
v5BJ8KOzvzIiqU7Fe8N2bvxd/tEdrrZ+MAlguT8WEb24njheo+ops/62hPh7oHQl
AYJAxCgjSKGE5dbUT8x0yyeNUT994fH3bjKOBVdao7KaM5pquw3ArGDw5JLLTIKz
ZVkSY/+reAJtLf6VmW9y0ERAH3idW/vDU2arIqBrq0lCIM5oPfZfWDvBy8oDDtZs
tN60yhmtU4vaGgIxYJVe4cjQ8v+rI0xAx7EebBFVkBqKHTZIqW3odBtAdK9GVRBF
QdKWNnWBulSTkvp8/PhWfhBHkVI4ntX6m4/LZqVDRSOUtJ4rfMVoNEazszrRjvyH
JaW5p9fTELXLdAGevOfyPdR9PDnqV6v8QRc1lpI9ixFOFi1NYD0WwblQmsnUDnLr
1GCHrTc95NPD36pKZcGXK5+95MN5F2UCe0XD3iDngugusE1S+6tU8+sFzZKoOFan
3Bh+07AbyBZ6ZGEq8nEVs41OF4qv3iuPGBad79TQ6eWMf5Abb5L9nPZ3HgGGR1iP
ZhG7zPkoXSeMJevD/EZspowqZpPbGgO+sdo5A1E+3P5C6Apjd0LIaknksljsuREx
kXrXBkuBIHIFWID5tqvtucRcUC5s9Cy2KjAKeI8bfb/i/3BOciIAlzfTbAnrusGL
lwB5Gyr0vSPATlyEmhrTBA3JFOGA8M64x/M6sBrFXdiGVDrh7BBoOjGPphtlh2Hm
FSSMP8fGb2l/869qQcYmfbeG+n7ec9f3oRhZU+J30aggtvKwOWx5ntQz80vXfzKV
1KLOYC3U8TbfOllQ52HeK0jyJtz+q9NA9DKrPygALq09uBEB0qZD/n39Dxr6wZ4A
BHCltwfKMngxBJQWwHtugJYBRDS3NIvMCLaUpxlfX22sc7iy0K+oHoZZZPBX9XYk
ZTtxCADFh0FdVJui3yR50yMlaNUB5yd1KmgvspOIaA6CsDpIrxbGb4DeacBeuDz9
2q29Y02gI2H3mDf3G2janZYtc7fBZAWsjWbSwtJ5TSKI+qBaNP4RNQ7pSbukZFZF
yp1cC22+ZkivTJvlF7sDOb3igyrUPnZfp+iOzPlrnmSdgYZx/N4GufF7ttwvWxpn
gia+PnTHGOWOSUNC/gLFSBATStlcC+/zEN6L1oMya4k+ZDcqca1rYGp7Jq1+sRif
IU1uer73MNh20XpjhqkRlxt/hEsDfIyweawW70HHqvwtKm9HhA0AedADcyNPa9n0
0I5hzayi4f1fIQ0hzoyl8sL0vwNLDkWm19ua548jEEAGNzF9sRKk430Z31SXBq3v
o4+udaDlb7dPpYakIhDA7+dmhu1/dt9DL84o89gqNqmeTRbxBGnuGK3n0hznUuGx
1FDiQT5nALY46Od7j5N6dREpx8UZOYhnPdIkIlDYonnuaH+/tmcCM2jvxSXG5e+D
ybH/5l7RqL6Bxog0+cV+sXfEAkDoHqKgZR2zQujXvhdw/UX9xnukGr+DRlm+npvk
5QIS6DcK4UCfXLqp6I5CTSGaqxWFsBYcJtg6viNS4fnYdZp8hwGIgU2QOk0zsAUl
/x148xoxmYjhHFtcmoe2ehXHf1TfD1UcbsMoy3P20a3m+xe6f9FTb9Krtm4R+3DD
+UShhjQCvKf8aMrQC/1LWeSgnPil9YVH6oFxH1RTKP5sPcFKzhLrIFUSXwtEuFsQ
Lc6WuRF7ElT6IQ3uagFxIbYE/oUc8G52Moc3RWxjj9X/0Cs+rLj9pEvyuvGdfp23
jYpjFm6yfUTaT4AEmBbNUWRAGcQ/IZJHttdlWNuheycDpwnGNLFs+I/UyMVf6Dbo
GkcPHiPGt3tn4xMWJubBsj34fs45Kvg3nyv4xGgFt/+Y/FE9ZSiu1Lw/2Cy0BMHL
/O1INO1BrB6rEq/Rc5HNcjIlGCm/cEZbnWvpXyN2E4A/Q7xADffTkVNx3AdNKXVQ
AGgkyCequojFSRq6LXRRR5vj+KaN4th/oFkKzXGCB0AjOzuNU6e7nRsezouIWBo1
tfey7vkD1PU5P7oMpOhAWifETWoNK5yo/yI+hisGUQu4t85kNez0zHk+8XFWiIKE
GpdNIdr7LQlrx7RvjRt5Ok2Aj7RKlzRlQT0izzL0bDqKk20cuPy5ae+bYMSREqJx
Rt09fnied5jl6PEw/eWXce8l9D+vBMxN8rRlaO5xj+QCNwxXygiEsngn0VDr2DC8
IPctB9LR/Oss79rht4inl7eFLlWPyzwe5yakQRw0eTubUW6PlKk2X8UiSLf0Xg+7
co/1lwI8RjvWTH02y1xyLvRXY/u6dk3u9yuR+un4OI4ufJWP8/CVVhqllURW5EBO
P86MtOV/oJNTmiACccjQWHmVmNJahlHQgSGq26+n3E8wZvuhMs7POJJd3/6mBI2v
bHSzPMUOCFrMhj5b69l9YGQsxYto0RcfeEGUSm5zyCD07UMmkqrGS4K2zVb6rnUA
EzCMoveYPanRM24h8jCJN/AHLliQDsjgrGoctqtbCHiYEWqiXN0TiWPcuw2WidCp
kN+cLPikdevFbr9iEme20uB1qwptkfk36OtLe2rMm1xgYcld/AqrzPDcbjjM8mYH
6fPGeGPgicWSZLFOdGgoNm1XuqZyMgsapLxO4vq2iU7NAx5JQ89mtyXvKVdVHhFo
8dEUfJHycIj7HFThNPPTXbqrgzSE2xaq3WD6drT7sVtYlrtJqbB1jWdUH3iWWAMJ
czaogxQUPi8nGZMloNeM3+XOzyM59QqUhyzZQMTCwAeZoVOiD+m2lAFxDqGGN86G
rEgLxsVX/Dzl1ReAGap8Y02xKaSQYUv3GaLXUwovFN7ODpvQLQFdwp89xsPgkU9T
1YXZTcSaVq7OUoNfXS7OiYPkGW30HZ6tnwVsBA+4C8j4JAXfAVuWexPNOqPaEgTm
XtcAsSqkPpNbZgCjwj67P3G+rTsMERkM04Q02zcvR4RpupTsbF982OsQRQmcohUH
na7OCoNxmD2G5Y6/maU+a/0S8T0o1GTd8jPaGEgZd4JqGS1iEK5feyzm3+FnR5tc
3IsCL4L/bRytfqz3lbSOaIHjyd3coRtbRaJ9T2fLf4iLuIQXDnrAA4+U+bmMUYfh
+192wKUhraqSOd6+T6a5oqLG1E0Fy4AqweT4rYHwxV92y4lFXLWSI3wwlCg+rDH6
stRT61MyYVUgPMkbEy5JyZpkB1TJ+/vS595BZTrIqhWpIiPGW3HWypIiQMLmEduY
9O7tuUiH1E52EEAYFyW0oS/AQPd2u7brGLd3DdrEciye0vcENZYAI0J82j8+QPE+
txCovteIai28Wb0eq11BJRFZlMnChQM5lcYbTLaCb5fIauITKQyGY2rJ4sK75E1d
W8zoEIysX2duX78rPCQBvqtMJLIYHmr9+gCUxENsOCkzHsLcNWa93OZQKzkAq+N1
cew8YZ9KYsZ97O+0vFQBiqnc59zmT/HUZN/IWABRI7Fawx1mbpAGpU1F9gQC9JLC
aiQtPj5tqXdDhFKwWpW5lfZlq5dp/yNL6NTgQRYSNMwKkgHA+qpjdJxy74Qje6fs
dF3IZqpdisXOxzL2sslfI4GOwICHG66RfC2OE0FUMPezjcbYPFh97+T7STHyZ7uz
gIOplCunOMUPBpkaIZ6hSIqEj85mAKRrR7cB4k0nRNvQIcWfDWsWNFXIr40E4aH8
hGJHXWNuCeV/ZjrwiaSRxC61lxI2aSt02uNxEpWEK4d+leGzSRGda9QyZXWv3y4M
quOJW1irxt7wMapUccKbFGW0oZ8X4AsCNt8vfBcUWReMO4c71HcwRX+A3WhUkJSy
NpxCtEuysjFvIchcpN2vdC5eDtY7JQXQlpOIMKpFJHWV13pmkweLea13NZjaD7ij
vNcBMD7jHf++DvfIaEYpQbCYXFfzOLOvdssmQWKZMfaatTzYk0TfUpx8h7dkGNjv
Y+jjQuSA8tPYl1O7u0Q6B8UFMzDR++dsQUp0uQ7HroebzSDV1IZWJWhtT987lSY9
qm1ECAACYyjVNjn3LiixNLREV4Ca+bNKroWb9xJM9EuD6CImWxCKC2u/mvPXV3Cm
UXPJPcCvcV0EhDpHnSFvigwmEyleCjR7y5c+iXpCYasUGNE5O+uwl22CAaARdu8U
bNcGdGseWh+rYN9tHmXpP/E+G/l6vLMEQEwXYLWMndIkTWDgLnZTeKyFmWSvBmgW
z66QQyATK+n8CQWy8yvqbhMfX1/RlqPSMzAbRdMBubAbqko7bebM4ysn9/dWQ3p+
vR4yIpoAESG8HNXMFRBF7ouxdjzfEtOG2qMDQBsA+ahHwlWB3KTA8Uo62GIZCmPc
NEBKAuxKaMM/Wutnz5zrN9W3g1ZCl2en3yqF5l9aJtTbGcw6CeUfEZQn+IZIVomI
oG5Rqza/Y7Qc64bk5+HHcE2QfvG4asdwgtPcp0iKBDqZr5Q01ab2DDNBDtneGDm/
T+9Xdr9++n4Dz3WDIc8EDf/50jzHnDhCW8C+1LBH/koE+5Y6QRL1v0b9oCClngbM
ErFmxpdIWa0/fDuPpfeY5bRrqcEatKvoLPog5dvPmq8Op6rv+PF9dIz283vCgvIM
92Ls09QMWK8rPCaQNWJ616uyfp+V+wzeJANeJr6VNKSR3tVhBZxq+iIuHYzl5i/J
gEkpp+IsWHCyzhN0HP8bk8oTePDD+m0q4fk3ABsavp7yxIBhwnh8+nztgh/WXMfV
qkzPK1XMNPie6zg0/Kmw28ADUj1HwqQqdk5C0iEFQyca5/wIYWQy0QhKsfPyw03+
77pVel61Il3ojXJf1GyDCW6dewbN6DsGe54uXeglFOZ7SSInkTIvy/HE6N5eSF1I
2zcGxq/xCvSX6Ob19ETxEnhOyPbn9vCVRV9t2UjJzYyG1SV5AOvaSEAS1m0TZkKp
15k10XbxTBmOc8HfqRfdjT3mrVWKZRhBM4oLtSblbhhAqKGECQ12tSLmVRRcx6aW
MlApTnQxSxAxoJ+vZXnfsIIvR0Ub3Sf61NyK/Re9nkK+QCY+2JnAWKmlVIY78qHO
keUELjNdhRqF9UzUm6GufYS7SRzOUXmSTtsnCM82OVIWTN6bqVVamcuJzTuUQfr4
ZlawFLq86A83YRYCn6b4O6c0Phhkl1YMnNSp54QqNFGA/Dr6WqJzzrLwQn07bHfK
OsUG2CBLZVgYwmEnCdqTKv+Fj71+leQUGXNUkg5/ychQA4P2edXLM1By4yd5E17q
VGNf3KcEIYKNwoG5swpwc1Cmap3QJQPun0gZJXO8hdNUvxMeQaP308hpH5fgaGgw
Zg4qPRCbAbcDJiNKSWlwf8hF8ZecKURWzNC4tuiOiHj3NvH/IwDUNWPDEb1A3fjv
9PKNPQUTnAO7HE9toCNqMRoC/zIpgY9im/wbyL4DIpVkX0wR7hH2N8dG8kaeg3Kt
JZg8Pu/UZcI1SfJRV9kDHc5r+PMnanM/kNRCMB8YySLzLNt90+E/tTzG1/Xb4ydb
Ij5otOhhvlUgxCtyfaEtrusZKQVX85VX/fMTFv7thCj54h5XEmD4Wa6alC4AeMO8
PkLNGvwicEncM4O2lkB6RgWkxJKvcXWrTpgcXPi57Fh0mazcNFYzcM6aAMFwD6rf
HWhoZAhsKKsPwLXw1dzQ6dai8l0oqHFXwF6NlQasTDCtRRRkgGSMKpmJALBr+4Ls
2Ilx7VZ4JjwmaJei2JFbMddwiEC51WKwFoeqfN7wzikBT9tvRNk63eGT5KV59kgv
gsCv7d0j7E3d75+Ku+EyAAqCOs4ZSqKkSWJ8ri1zAxNHzQKv4ly5ACBhqlgyc2qX
+VAOzSuAzoBW/gqy9xVhc0hDsYcv+lMJPYSA1JN34NA6JSZk5JlduUCg4Gl5fU6k
aYRzaFiXo7pCnRA012+Zbp+tQFd7eM94flRCNfeTs3bcxK7uADDkLWerDN99H2MR
mp1Bw4/JLikCAacnnt07CY4rsWitmWl0Qu81kfwWtbptPMuxve/W2QaIkiwQeCJy
JNbGT9Q1mzLiL4icbfRnncpPGsFvrbVbR2Tq7FhGCobi59tXy6aLn/Q7G5ML5AZR
MzGsGs1Gcx5g64Ty/gShZ1+eRaNRVBkunZ83X3BNkB5i8v87sn6GDkuxVhsgXI7u
AmbxMHeZ8T39yBFKCs8htKKjGs7K1g+i7G0xmn8ukXUfDfFHWGyuUrCYdBh8Wn4l
76AB97EMZDL+ZqpaNWlemFR+PolDMBTLGpLczEcsq/getFNcz+rRzTXEWJu625cw
XWlmTEHGZwMSu58Mj/FrOcslJ1hT6GrlP3/KY3pHpYKl2dI1EdMM7Wq/5hkl856K
nHeOqzmDm+fYHNxRph9eW5MO3fNwxFlu544oqo1kFjyNq9BHnQG6uDQ82UtDviYl
vpV6IL168XQIEi8cGDyUUGAp4P+i/o9reNMhZm9D4QCwN2OdLXGPgox0GSjOdk6/
esu6VaDNaVMFbPG04qlRUyfmN96Ii3hRW84mNozn+NoDFvzhwqgBOsZESvIMsQD4
H5kNg2PxcJWe845rcqN0UYHnU1Sc4Hl603SWsoikH+smdBix4HD/PSHIVt5yWBva
b85ij3OhiqoCfRTL32BRjjpNIlMbzHyO+vYufimQJFcGS/DpgJguHzvVpOJhvFkw
swXfjdnwaLBx+JugNdyQ0hB//rU7/CuMtMtFHTmdpoNCavxhdaxtexGqPxvAV6q4
LjPn6D1j9hbin3bYye1Sl1fGaLyG7PdwA4p41CEw3/kBNa05KiGCGC1g2AJqBHLf
q//6gYXI6qzbG2Vsj6SgIs7Y19GofHctHGYycGF6XOeLZ74jfKfv1vU2YfKE1zRM
P7+LwECaLvqF65htRoFTFuRCZIURrrxglGAqTRmhLHNq2h3oe5eOpUGP8OZi0VXL
IM1K9u/OF3trfaUaUuJLmOtmiVwlSV1AG1H97ahGSxJmF33jjml/fAshg4Ab98Pr
G6urEc1ihGWYReH8h9yy/1iXfaq8TyzJEZ2rD6pMjm+8yxPzfuhRoIqk9WULDrSD
MrHNrEnK0bq49AkHhfu2Uz6an/b2nNExCyA9k4DqPtBkEUexPpCt04LWrQTFSosj
Zbl94nwRUGdgeSkO5FGxTVbY28UApMQt2TTUccFIO4C9dsqFaz+yq/7IL6sbu8U4
lWqYeBWKP2KLnV4nlXhRIZU8NGs0hv480ttoq0BnCR3lDc+oIRxneHb9dU0cG9fC
Bh0clRQwQtKoxZZzVVNGKVL128SD3+kxlBrTtdwNx5TtznhC46AajzKzXJgHO5xu
n154PNtbmYfPpcCMqfjIa7lTKXsRoR7YFn8wMhVFaVp+y3qaLr4sGUkmDYYw8rvu
oFEGhPepd1nh0o5cXgLfUr2XYUYJkNbr+MIL892BzYHVOO9vpCfAqTAOfMo3zrHq
H/+r8hWXlfJsBwMWRwGRMjWbJrNvpmUazjUiQnB8578Kvoi3Xpb4JtbkeQHbl2D5
dGLDuRwG7dl6mKvt4H8i3qREQdQww3jK0qmxsXSnkebKZAItkr7l8Dr0RIesT6Iw
LfR8ikobYxiNVVb/3uAfHVxO7N30TaRpPh8Fm760AwNxdjsShztudE/zfu4V9PrO
Cf1wXSEWaH7k+qufsRE6ERc3E/4Q9WNZLUUpMZE350UOrNU57O6r3no75pFABFj8
Ll1SFoX94ZElfbM5+Ub1B4eLzc5vt9j2blsaggwRQh0kcez4fNQCr+t/87DnHmqI
ieN0A1PQ4rlJNidRKtUiRFkKSxm8YhmoxGRjGyWmx7ivONFdG6XLYpUMEAnZnuIq
pMmzWRYGZckQbC1tgiaNzEXTH08duf6dIceeNRXdeG3kCaiPFCXcwSkkBQLZArCl
F6mimcYPoCQ3OHIvuMiJA7+/lhNz+7ZsitIigaQ5JoG9AilOfNclD/eJZ/KnzI/r
7WuzClwRrKCrZuZ92axppOLQ3sB0aziN7DwJuJrZ5ziQSUpx4GR2Yq2+g2ZgYK2S
JvbjsDgL9Xhzy4P3kT/62MbEhwe6AkFLk6hlbyZ55SibW1uY8KLj9UsjJRZfnP/G
cwvfjMPN19kmkuhgT0keSCkdG9zA50VMIwwEADquPSEshHV7AfuE6SvvlZFL7vjE
JufDeSs9UQMIJIjX90ODtqM0qIyqRWhQ1O0F5p5qtsFwJpmCMgJ/dghsDHOVpmJu
mm7d39YCasLhctJhGV/k1A3dQFffn9IxtlNCQJO1g5gX7kjo0jGYUL71+X1vTkWA
hbmRoaLsze4OK5ep8kLHMHpPQU+slv44tHZkH/IiMryYAYy1S87mZ7Nm+BXjKFgD
0SoxTxxF+NeQRf6QCd4BbIrcMessBgghJAWcBIQcH7hzcbou47Z67JgO6yp6HfVx
4oQnSF4kwMnMjVqx2J2qzxGXJM43aBDHLw2OJlxHN4hL1/YZ6VvP50dSA5t0eB9I
Ag8gqSkKVK/DxTLgSmhP1Yhk2sH3pG41zjsesoqVbdCmEHvB5khU+Uikh17AZ71u
TNA26YXgpBubv9tdz/KQJq+63hjSixuZwU+wn6oTgHhwTM37+zAGyc+j/zOJR5IT
Y8TDJxO62IA++WO/qnjYC+eD7Vwki1t8BCO3WNfSPkD4wUVb/xpRvUs7zhaO/McH
rtOCqW/yyPjjfzok+YCpEwuG0lPm0W7xHYi6U+UP8W30iDxvXlkfe29ELFwJxWrk
JHub9iXOo/wgQkUpgVhCbag1mu7HnMK+vI2XGFdAaReO+elbh+7litTExa7X0Xrq
obUeDE1Mod9HrBZaj2K1v1HzP3ZNFuIJTHwq/KzNtejNFXmQ2vyiVRGI2ZknnOng
w/LIF0G8SQYLN0eB3uQzQVLwFSC/M9QAbfTf02FZ06166XSrDtJnKQ6SYsGY+l9u
EcqKyReM88uSNoYaMqLnbmT+b9Jjg5dCXx3lErU6viu1Sbixn8xQChDUf03vx0/I
48hWq3fJVjn1QNSimw0TKcd7TAt8PSjnc+pA8iASqGv9Yh/PFTnIkdKcChD2I0Md
yyVCvdqYnTprGIHOnE8VsMDTBZn7G1j7yiKHWXre7+xpx+3fzLXVDKB6f9Tn6KLC
BXv2xO5qzLyQT/CyIaU9hg8uQsG0T1UUGQRts68MqXqAdmctfFergffShkBL1D7u
a+MMRNFPI5lvE/oX/+s95RoR6Ep9hdrixih1pnS5ewmCPgRNaeJkxldWJ+l/YKHA
1U4B8h+/PRHjOfuQ4l5sxcf6cjLM7c3GHcnYLBnN2Wjsnh+dPIzpmSuvu1481etV
zgFUYa8ivOHMdCAv7mSCdZZGcWEAFwjwECNj16S/sJXVkGlAFw2dxp21djbJNTlY
7qe8rJztH0kivL0nreptN1lt0J+kiymOhGhQ1yVfuZvghQLWNxRvKCJWZmQfETy1
xFB4NC6Z1pD4fcxT3wk+VSlTkpoE2J8x6XTTZ7pVtBn+39duO7MucLpYlndHA+D/
LC7DLDCkG+Db+DmpsbI1gHql37H50FKpnkgVXHQI88HcZqytBcK17A395394gm6o
rJcJRIzN3isPXU+HOh3NCfwq8TuN+Uy8JeKPA56SMSkorL4qQA2tkGR6ynmY2Xkf
KkH8uUpeV/mgdJ0LHAoNKz0NqSpN8Soqi01Sh2uzIUwmjI/Td28iGYqD7iMvQaCH
+t/ROzTXKsyTbxS7km8pCLEGULngofyCEHudRyKLiLnklRuiLtwcU3PoqMU9uxC1
Znpp4jJOv2ze5V1IPiGY+qCc4upUVPKqj8eWqWrXmE69OGufZ1F9wOZbZw9K40Uo
S7vjjpAyTTP8jHphGtGQkS4etTTQk86nkFIu1ayR/H+P4dy6DxW4hdK2x1svz+0k
K8bHnODOO4EhO7v84OH+5iLQYCMKNRAYAhWU+pBj1W98MlcC7JQ9OwJhZRSCjvmw
5TTjHQGH/G6fu+a30dE3Gd+4bKt9Yrf0CvMXbdU8AvYT8QpxZTxVBOICx8TKUVAW
81F0S/wrzGzVHwHk11eSGGL1XbhFM87sBE6+o7euG+SJlKbIcxDPrQLBqLwe3nu9
d4KclGNrf2GsAKeUfSj0ul29tl2PXruazkR/JCIn+3hKheKq+wkGjAGCeddfsdlv
MQI6U/Sempoc42P13C+XDHwB3MKIylCVdUI1IXqMJZ95mLdI3BeJ2lcX5nchM67Q
qKBvG1pZxUWLOoe1UObcd2zEzTy7MHjzjAz0KobJUfGexEwVJcHBewjoVzBFFu2i
eo7l7vfAjVeWHPjH9PoKNbWV+k6oA47ODLYWhwWJ21/Q6O96Hcwlq85SFHsdM/Px
MsSI/Cwpglz4vcnU0Prtgp+xWI+ZKcZ+luYlPTf6yGx1mv1r9z5Jycc3F9RXXs4i
fEb0YcCg/3QAorlfhyCMHuGRjNjOc3rZ2hub0FMHQIDUvn1e2+rWZZTMBem2ZfU6
GjZgPILI4BBN7RPCQ7/T1Zql6z3tGY2E6AFTlBY5/ytP59hRGc3Hr5VUnY4Amwad
T+HpjZ7OhPvXvObwCyHRSTB6FalMGfKWAkOEtvROQW6FEx0chIPZfpyyn8sWFHjO
wau0nrmyoTp/QA+Uzh7ZPl7GQLA94bBU4fxI5WO6zjt5nL5VR2EXIF75iHUcrYlf
HnHYogKb/xhcdnXlp37BbQPPXaY308ZLN2mnZnXXin2R9OG2gXO5o+Vg293I+gwE
GrmHubBTtfs8sqcLvH6ylTiV7GlPsIRLIGCmTqPuev2KTCs+LFfPB7WNpEqenbDI
G1QD8II63tFPa1f+M6usyrzZvA/foBuN0UxOunK/jxTvoraF/1TEKh1td/FHWWVB
BkyMxfRC8LV08Me3TFIFiYpIRmB4FIxA3C+epR9oOg7VOYFKJxEaNAf8JGwanTGn
wek55K1tGVxLItbBLDn+oVBbwLkUONDjCk2xcgJDzbtxbz7nsEJGyuFVwyRsfolu
bHGiGk5rARQz8gGipEJd1hKAbL5ONf2Op/4xgkmmazqX/0otG7lYq3bQxLv7nJq6
Gueecf97xRgCfJBtCtW61c1AcvRqQffhhnC71pIXyBo4uMj18LbJyAcGmY+uTS3R
DTBoOzzzsjN58pEIuSFj/WVZc7oUxAudU9G0fk8/FDU+YaZjT1V+8WhcBNnxmMXr
HrkF3zIK32IxBsorX8jtKHozNUE+pm0/oK0/pgTizEda1TWLY2O3IsbMl2DFNthG
1gwXtDVDVCcql2wpHwEfDO+DmuCvDOS8lF6aohXjmsCcXna5jzO4aIr43yGlGiQX
+JUUXyf4vTqI+Vb1iBJSWAyACS02gtFE3pcnMmwOjp8H+Ccz2YQ92IZ1+2oM3q23
o3arSe1nE9xUmRj8xlEk1qmUDcG1z5SM1ivIaGdjBwtdDfrEFr4msnOW1vAfecls
VjJkewm+yPLDd0MbEaMfGQ==
`pragma protect end_protected
