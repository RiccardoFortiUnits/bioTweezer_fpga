`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AhG4RIJ0yC11OW4J/WpBpK0UVpC5ipnqf03FgwQCswPqHhlVRvQDPv5KtgGxEuN3
MZBrubml9yACL9zlyqt7ccwuyjAg/zjfyHSKFrnRxx5FxT/pqwzdeTQGMS2wp+RZ
NdEzA7EaH45Dt33sil6eXIPDptfC3b/150N4NxArjMM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12432)
42WaeGLaLpY4hgHPl+I14pcgBQRK2gCjvINNbVu+nQFLyWeaLRqvRX70aJMhJHPd
ufxVqSaZh1zoGn5IuzsBizYd2cGjjkP3ZprT2iGwYs3t7N+VUpQqw9OQKLBlKqjk
NYJ2f1hgaxbEZ7hBBiK/ZI+rBoH/QsrT4yYxTflOImmUA7B3iMYfY7nR0adKAjEs
Czte66+QZWRgyPWLoIMhLIUh8hH8+eCNzCiwbZs5Qxx87RM1Fw2xnNXiAoxIRLkC
T3Vb3XUlAUTd7fwbWNwNBMRQWTWuaA8oB/SkhPqJfR+imYwUo3ZLdeVOuO+XUv5U
12tSQA48GlTvS2Z7ahO3C4QcBODJt8gwUp5xr5XX+C3w1dQIdMLdkV6pXvOxQ7yg
OfS7ry2vu6NU09xjpFn0pd2qvxA74Dap5JbwDiIzQKXhTYWgKt+qjpfAjvMvjZTo
eW+uRg4WPL8YZHnfU/8GB4wxdSzSmgvyLLk/Mljvs89oh38liWqFVM775zfn/Pj2
Gd/xsswCu9CVMxCrujzgxqDEmxV/LmUAcLdGcWjB7BG0BysJZzTG9IhCwqgDIq0y
6bjJe/rduJxgoSi0Sf9jikZfNtGl8ybbNvMHUXO+B5ZqMi3elma8E1DVWlR3EIxv
R+q2ebIVby0OWhciObadkC5nx4jTN4ZDW0Owv25390iAJ7myzqomtFki2Z1QUwlF
cBb37pvoulxetCv7xTASRrA++wdq8L8NQ2aaPnohDB03fy9WFvAtB5FRHVi1OzGv
UMZOHbfkvE7Xo3uOKNBLze3XQL7lY8DOqKRGAMI4shD2MB0iiTg6wyg/G/s5kpZ6
EW1kLZSROxDgifyqbIVQ3n7uTkqHzO8BZJI5fpKTqIFZ3GPI9fA3XV6q4llUdLXs
h0RxRWq5JcQmWVV9NRkQAakg1RDNb3X1Cox/vKqOpx5b15vPGryrFyM5ZPcGSMm2
if6ZkrrqEPTcX7MXL7La4pKRodWqPNP/8ZbxrmqO8RiL7bBU9SC01W2QH4HNO2YI
SWbLEtO9Qm7N1GxggO1AIeEm2m39eO+SMadcWP4nN2SypZQQSUDD7KUacXwB2ze2
vP63mTznqX9NUvycAWI7rMaikFXbOhSfUBlvzz77a2v4Ftrdy417vHao5Zl7RKiU
FyV94qgxCl7fqNiBiTRG3bgTkgbmj9LBec+kwMNgaRbI06w3aslSbleSSpBFFoW5
u7N0ofYl4GbdAJikOM1uviFe3wlder5WII6E/Q0JwB+z5e5vO6BBXyqTe3/+5WFC
8xPfz7JB7TSTrFyyaH5aHWkZ1mALH/NvPIFNRjcLg+pLgJIEzJeV4aEeYjNALfVq
2uhn4axxve6ieqt3JhR0RhNa0Ng3TdfkNrCiMZHx0XT45mM6MOP0xXlshqLrVQiZ
bCLN+6FlwXehKJamS50E0Eg8jpxz0DW1HqQwnbmCgNvyueVC06VuotG7QVjYAR/C
NUnoVyMPXK7tN3Y8OK4bopUv0AqA5J5J3hV5+PtmKLMLYaL1BLehVD2tSxTQHcTc
ki6kBlJyrOtLTT33tYUwLHgGAx+FwAoBQ49ZRMaBOFc8wwHooGkvIas3rGhtqr7j
svBljBGXC3asBGQf5hXCrvGxjuyr1imSpLhpN/pm9WqlFaaHMJlbpEhKjhRuonFd
SBamPQFykGLSmgmp9WlIBT3ND2MG7ei4JQPZAWd8ZFjJ1WCd1aeSRXp3ZC8SDIry
GxEEelGHjemQ/SUDgol77q0zQD1s6ZbdwslHh42W0pQLvzk7QSv1t6t1xmf9gW/r
rhm+avX4yPKJGoGw4s7h5ujcJQR0f50g5eKq6tQDFKM3aMv0dZjROHXXFRxXNMl8
b5KF7TKPscWyWBstWbIRjTf5MnDbinPGQcej5EnG4ig6a2h7cYHMZMiNnkDqxszY
7GsgeIlmLId3XkdWItwtl0LShhV/Vn++EQxwRCe1YWEMV6V/2mZ9wHogYaFPO94T
2KdfiWNjp3OfDx6b5JnhcFDSvtG4tWxyEAi+g0a0PCitiojS04bOOTtFIwmJPtOj
z9hJygudf7+gICCvfEt20ZcQxvkL9MIKmf6kT9RI6w0E8cX2xc2JGEStEIYZsffv
xDnyQznWYLdOlVGCzq/HeRcBoDWV7IbkRQLz1nXhTzlgLbfvJ8Oa1orleL+9QwnW
ISFLvAMKv47rdKdI1WRxy85rkLv0P4E8F+xxwmR86AYa6w87AaRs5al3gDguCAS/
79uzceiEOQj7Cfz8ico3HojdwdssN90loXdzTnoL0fgFUezQX8pijZFKMcXD32/6
5/hQ/cd6s+XHg58Fu1HL+6rtmOeJGi4Maz9XPmVIlxYIkJ+Or8eMZoFX1VM51tyO
9yFK/6E3fIEQD3fMZGUciB4rFXZeVcsZ98pCkeap0u1QPOXKY46oHVRZHbIkdJ1v
eQ4J1qHgwAbwHMl4NpPXMr+7mkudDF7mYMXamGqAkar3Vl757qJDSwMrY2zIffA7
SDSdk8qsa/yZU1aV8OFgwR+/2PWX8FGw9ad43RjXScJAqPqmu/V4XSk5nGkmn+Ix
guJvEKBVDAS+4gMiYpSY+nabL561mlb6bTxZ8Ty1f1euxPjWMQZAIflIiBfvu5Do
3kmGYAHCzB/dy7TrcjUyro7GfGSGtGBQ7A25UCXRHBuzf5D8PsAcsLqaFNXaKluj
hDaG8EBFo618WBmrhGBjh95VmE88VyRWiOjXPNGe3+SLMjB+MufuqRe6l//CJE7R
Zj3alrTq3YEYTiLFmoTh8EN4bGsgzZshzWuI/KFKSV3o2URzc8ocgyZ7D6dLJB4J
VQpqJ4VSd5E3jvOqD2Xkn1cvzd+mkHHG/BRAopRuw2+2W/C/Rycg41DKRVqR6VeM
NdrXCFNM+eFgGDg41qZ6BvrnBYlewiEnJ+D3KGu2QqXe35pMAJ5PC3oissEvn1QJ
89dh7BdE6OwpIStUxvdnmlIION/oS3C7E0YmJZeE+6K5nB16vt7xdvPgUQ+UjC5t
LikQczBi69ksl1pwruBityeOvcAmta9RW4p6B1DdA/RwFkXz1w4fovZ/TXVleEc5
K6edbue5Z6/7nFY/qvRSnqqtZdcGiTSg/R28sDbSO5A5IO6Xuh50Q+CWWnhAPBx1
aGyQkx1pq99Imlh2/VSF7kVsR/eYCEEksO64Nzsj2k10RZFVmQMDgOu2cLtvJBB8
4S8WyvxSbljy0W00MtZKFZpJPad281EveijDI+0MCFg4ZiS4cwHIPwa9Gl2nZ61a
FmemIGM0+dgX968JMN+4fX182LUDXR8BroRoPVka9RSqqP26fWDmcy/7OEE1eVNn
vi+eNxYwEQhAWgSKbgDwVQgl2v1awCh467nUMfAIQ6f14YhRUJ6N+Mhaxf6CZFen
/lmGD09iI7NVjGUWiSksNDZOuqKXN8HWW118/xU2lMN3vEDuPYCuDa4ZttbjslBU
aG8xR9jKpL1FfP69Ta/6vvDyEfckfFRJTbNRYmCcAN7Y0j1LrTfffF517DQoD24k
IXQ1Xz3LS/jvrvEAwNlHsqm+p7y1+lzNd+zLXtvDSxKGPd42jub3hvVF94Ncbcok
VR8JLgGnYokSX60Krod5SGnVKi/WBkAjpK7Pe53dBb2dRxfGDNFFa6idn8onY7hC
qTmq5hddVJAKrfoo7pVn861sJ6av9gtrdPzzCiQWo6N4pWbt3pn6PtjdcT/VY0D9
VWWSWNKR9v/EBdj7QqPFlIXXGTzf2/SDhrQwi/U1x2IjExgfXhWIsMw3SP3cD/li
IumvpXm8QuHD4RY484LOskv7QEzX8CPYzZPlq9KX3Li7zFqxoEXJnSBN1vefgGb1
y13nEeIqKtk4jGZ7gF0Z5rKI3fgMRTTyMaftg/5yui7apiPomY+Qnp1zydQIULmh
mg+K7SWOUsZA3TdCYm3MFFVFSWpZ3dF+lzpenmAr4RGe2PjCx+BCW96bzG7sC5te
ZTd9zgjqSMZNKtsxmtLStFq+H7kjf3qYhLQvUF8BgiH9CAnfhORnwK8tyjOBR/UJ
ISAF6IN3buuQWzb2GM2GbdjILz+G4rP0i3XOhv/CrwdFhxMbAyZpNU8xpwdxKEss
x9qKLeEmlnXdstZedhdixPboGzvCLlMsCrTGhossSvo94A1emS2jy1lNw6HMJWZy
7s3YMS+vqFeDTCQShqCoKcGmvOxsk8cI5Z0tnsNv9Ql8SyAT2ioA0JnP+D1VPj5T
4A9eh+kbOaVR/5QiKdumYo7P2hR3t5GEHB02pUt8tVug0JJQBQpDpQh9nbAFLMAN
7h34On9e7eoq5m1XWNrqv2o29jUNnj0RU1S1Xe1JJFcOECXsFqjZeh1iHF5S3FQ+
oElQME08bmtttKYbGmPD5KAgcG4X9d2TXt25fEduZkIWoiNGM1eK93ot6uOvlyjW
pTF4VAMYokXbCV9xqjy+6PoC6cYSBxs6ad4FVEB4TgZMBgO5azfO1xht83mRcz0d
PQKWGnOnyVV6puJBHrIJr0lZSjjP9KPFcKEBtAfWT0QuqTQ5lWj4/xyPyaF8+ros
fihXZjPhUreNFH3ZuxZPt3sNM7BoBaecZtHz8zs3aINDgGx4ebLWv+WlfVhk1KMe
AJQtO1EHRDwtY4msxNAEScvHU1pK0nTNqfh5ixdusLDS28VRZJj/e09iwDIFnCg5
XpeNmwHMkZ/ovt/LpaC88AlkxSVQD7XONhIzhD0gftMN/HdGF62ML0y5Fkb+/qeh
k8eQWZk8Jn/8L3+TquW87P7gcPcAN2a568sN/UZOd1bv3+G6pVKzSNFS4XBsPf4W
J5qz5k8O3uEkF3jbviYJcxTH6Q1pOvyQJhcsiReRrSE9GVxbZoifOrUcVD3XMe1M
B3t0tlFmUgykp++NeXTvNRSvrUHOMelFuVCEmBe6pk9gLTy0pwy0w+of6ao4BXGs
A4mVuJDUqQ5OBeLJYlcMyXHap77PLqtBDHTvj2Ftg/gvwh0gz8RdfUHvJMV6Sgg9
7fLqnjsh3bldC1XnuMFwdySZvMTXLY2pefyrLk5DoNIBlv25IVlEhSb8RWQgK0a2
eAcZtYGGEaEnc4dca6JpzmIt0h2FnznF3pCoR1TB7QwWjcXC00Am0x4sbvFEMa26
4KXlmiRtRneFEzeuuTglQS+6qGvays7ZZI6Pa+vTZicPML72LvkuFwT1eUYvQKlC
+CkGZcrBe7S4teZ9oMlW5a7E9g/D+OLjczi7/kqKA7I38rcOlPw95JqR14x6kxpn
YhrSyUdrLWL7juDnqphRRXcwTbU/u8Be23tozrlaS2oKHbzQHh8rXaT8hJkLT6Px
YJiXRPFebmB2F8nZ+OMMkhUIb9CGV51Oewze8A7sj/vUtob0DQkX+1cNObvu/uGM
A2Z7BuFgSllob/mfA3yQMHSnkwJpOZkAoHm5h+ckm3jLZUTBM7iGNExxm0iOzQHS
39jPmUxyumGIDxIw6J6ikJ1lRBtfdmGr+xJ48x5g9qZWK/mc6LrCB2zZI15JOv7W
HfJslSMycO60NKp6I3xh6a5+CaDc8TRC7jdapta3PCfNSQnDrmzxVXGJRc7uBjtF
KwZKiaWT7Jm9hRZhkBquN4Vs4zunWER1Je4Y8vyxucbz0c/lHPzJ/4lOibqFoZR7
GTn0kl9vtE8mTnv62asvTNUrqEH5G30YoG9fk0zElkffyzXd8TMnN1BV7S7csRWW
pS17eH/KSHQqqOYUL0unbbAthcQF16dxcLvtFhT8+70O168foQrD8L/CEofWQVYq
8VFYCCn3m+G/Tb6aSFBnxq9e2YKFsBl5MC+5okN2NRWWWljiyE7MSlFVPsAvjnHs
E9bY1/Q9ySqcKlHiPCSgyOKCcDJOrIc9chOVQZxAkpvoPk98IhhJgwOSglPGL5E5
Q2/2EACCMqjfTRoXQO/ygqH6KQsScoh6xTfnEqPi1VNQp2y+BSQPocs1Vbam4FmX
OMX5mipf2OEwxAlh5/qBfmDrAfhmCmoXb6SxL2027KyKk8S+fGogmO/Odwp3oKXD
HCZHXqgkRZtNzu+m6oVKvEV8tmTGR3kuWM5sNvKZnOtZ/jbAMyCkb6oex40Z2jSh
O2y9mpqQwBr7pybx47zo+L+FR4ugWamHHXqg7bXMB1ypntdXa9gWA7q8SQnwMtCT
TrUUhNtBPITe+aVXPQZIFE4HGY04fut+jojYOHE+vuCM0Nh6Nne1ZbjZPxSaklMr
puUt0a8afMHPMSl0+A10KRL1LqKBSrEeyaCDqcQqTGPgmpIO+zyPDKngWlqYl0sZ
gBUtgy33pja/7Wv5SvRadXvHDMnOdsou/RhG3EcbeFkpl5AhLf1xk2Uh2faXsDt9
7Qxo54MVRGi2e5fiaLf7E+7jBlyV+kGlsUZvxCggLNmVMw4TO3tVFNdrw5i0judl
6ayevPPmZfyLBpeyYMv9Jm6EpWnrpyOCmnaP5dnxr2DqgNtx/645SEJIsTFzDsVU
8NZbKwmAAPSm4My2qcy2UmUhFrpksgw6oTjpPwb0/4XiysBHwz9cxAtu8rLtpRC9
nK6fEVfvY8vq/p70jWrQxfK2QuC6udMKd0SBKKGImFkCHZYln5xtOSHByXRUIhhO
6x884q9S70u9fPPkw10XXGp+3fm0/5IlDZnF6xRBvgtaiqBJkgt6DHWkekMbSt7q
2oNRZnYjWvMGlNSytCCS/flcqO3DOdrsm3M7fmVPCU/9if8unXqggQJTYCBccuxx
qTFoiTCer6t0+SaGUt8KdupqJenHMvOWZQguMFL6edK+m84en3eKVzSEQMhAfvpv
d/k4o/y1h+lW+jL3JXXBHzUuvPMxqZPIe1QOBPZVI0gTQcAg4bEVwJx/2KcOYVrJ
0x/Id7Otgkltjypj36zfdZsoX84Eoeuk9VwXTKG2hMZUykCeESHfXnNLW3KDMTDc
jaJr3WcJoFp1OAws1txiSUCs5Rsh1pKZ4bpNcwQTuH4rc8F5hWAsYEp9JBVg9sFY
d4y2jENJ05BpiprQGh2Sto+HPWVXpuCOoBlvgGN6uVcA+2EP+LjG3MgLFSL+2TsC
z14dY2I9LtLluTsmoEZDx7MBjSImw7m/pJlrddBMrIrgUKzU0RYICQMhC9D4euFo
eZ51YhmSsv50lxKTm+Ux9R0WCR05bt7DAyCfDt1KhTOKLSGfrSO8kkkxoC19BQBY
EICr5xgDniLRTc5JtCuxW6B0P+EiIRjQ6V9nwITGAzl5h5MJNqVJIwfxXdL9M5Fx
suqi/RPyTwgoGZFWqyTQ9CQzaAD4uzbIetXiwlpRkW4y/S+6xaDVnzf5ipK/nuK5
IdSXy+qfAeQjvoGGvi6O3hl+IZUIIA/xg58eDDCWzacjPI1cZWqe/LRaLarVdt8U
tXPDT691gfVAl56oAkdCX5fzmpdnUw393CCY/n5TV7lYGujO5/cvXaTZiXwGaweU
w1l9VMIpjEhD0rEyB+FAneI4ah4CcBQZErMg0/LfrBkRoADbVgjL5Udt+Sczo4ZM
HH1y7pxvjdPqlgG+pjkefgiVgiTWMUSGrIzBApBwnEka7lnvKbHFOT6EVlUpDsqo
x8U3c/+GDBJY9Dog1h7FitJnM711a+vP7PT2YyXWSRneUk73RTMQgWW++c90SfHG
pTpzZa9PvezSjiRAgVp9j/+6HhlitgTAjapGnc/97XHDoiZ4I7xR9IJLVsq2wgDi
2bpbdzKHC64vWe2y6wXJ5wSYvZdAC2xDVYMdVz0T2ic/+0abU3n4m+Xqe4Erausu
J+4rBumZwOvQXhr3Rq9iWPOOx9vtfvVx4xj3ZIsrRIobJF7BmxhZ3IMTMhzLd2v+
f/pXQcB8fhKPNJqZ+mPwEU1txp92+yED8z8p1Wb/bWICxpHAT0Zb3osK19tTHARE
XjNpOEKZ+U9iSyV24RcFFZibNzUKcqnrhbeDqBokCxtO4Fc6XnKA85VQ7jlI9RP5
+roPZbUnd6j955kcMgTh6a8c+wLpZ2VtnmaU0N5pH3O9j+eUy6lIQeOL5iEcbQil
Xup4h1Dz7ltkwK5OKMiDFba3C4+nPtuH8l7fQurFtt4WgY/hbasbgL+6f06SUc6g
sS/QTtXO4g6Cv6ZNvyt4z2UacDTX1Z1nA7czJWTgujIg4KQG7hbMZy0QNYTQagGj
YmMT83vD1+nKQmJwvNDUbnVYzdpQAyM3WWfPSn6P60mUiv0/NVKXhdhT94yX606I
GzdhzVSOGyZSEFEytXU38RKDqSRViqtmhdHbFTP7WUnHf2gqSgTQATtchI+RRJRO
vjqRs7xVUqRTrp0XwYWMaG5u/veoVsb6Dez/3rI/hS/qmQ+K6i+lnh7/qxL1eigu
e2HyeZc683TJJNjyZTLQAspObjH3L9me7bS2sGGc/a89ZMHXKbRFvdQSAZnIOAhd
m9NKrfVswy7J9JPee4pvjbpp9nvPIvaujXHYVPMG2YPrb3/Ak1HdxXMBJcJ5MSON
oLpPLoD+32IFqNDVqztoA9WIGd9E15Travx4WbcokDejAgirR0qTgFcNRLNpySrf
x5fwztd8RojuroSK/jW+BYG00hn/KEN5dKwIjIsUZa2oL0ns0tuMWE6zuuf7iVE6
vjs3vgSCAQpSyosH4BycYPtQj0RlV57z/69OOQB03+4f4JK2dkcXgiBWDyfbxxfd
8Q18zVArZk/eBcBNq1US4Jstfqx1p0ayMByXkhjr/QdH0AB0bZTNQCh/rxR+Os5a
BUw+S8gP8z4S6scR0mOGfoFtUJMdGMSBNd/4GCd47Oz8bczn9476OTc22aE+0tmT
X0V5zEm9AHYx/3JkdQYBf1zC+XYLhtz9kNSc+48FPvTsVfflEYxvG0Z4poIKaYab
Wn1COtNvGSnany15oQGrYiKIlS5F35AUkA8p1A6lssYBhGWowey327Q2w0Oq74uw
++fz9A/hvG1JtXOhRH8QhZHHDXGk8nfbn5wQsV3TUTfhauokUxTtqg4rwjzGgGkq
P7jVBPELVV6uVvZQEhsuu9jUoyVmoL/cjHZOdfmuJLLkKNvyMChGjRHMvgAg2XcG
17pUx2dpWJNMRdWekw39f1Mq0HebdjdUl7TbcGQvY1Mz2WVbJA8l4VaJIkWEoJWc
ijHLQAXeWu8zBNsfb/2jy72Y2cp1eLGgPPM3IBFf3m+zamXsG6FPxM0gfk+NSuNP
ZVPIT7VlG+ibNuxzKi6is6DRDLvqRMEaND1sAOBR8NRWHno6ONdYCHQ5a88OTip/
2R2/EFj3N/O9niSHxfzL/a2ensRxfwAVRJtHMishf3l6y1XrhhEa9+XG8GWH8571
OHzfN3oSLVZgT/dI91Dr/6ZguMsxmk1ZH/Hxt7THu/z0VUVet7RDP1l8o0CZ4cdX
peuDhvAGml+88Am+eisPFM6rtEkc7ztno9MJGOBEK6isW86AP7J9hSlsWPHn8e+/
SSkT40uMvOY6DRqM/dWTFYD5g+/KpkRThXFeXPhAwyImmIClThZokvjkV6ejpIJC
hAoNL1sp1yR4vIoTinH7+u83PU2HK+uf1p5qSZN8ot1//+M3r3ZiutFlYlIm2L62
rOR2ufFMIbTOz20MWa7gVHWIniY0bxVJT8uVfrk0jeTR3ti1LbMZ0KXxRhmo+9k1
i8lmzxPNdnySED9EfDI7m+dDxVb4o3bRAu4YUgTKmBNoAC6wmM2y/Jl7eQDxIVqC
77Sq1Zj+z4+tg3+S5im27hM0Z/UbLqVSQ/PoVYvdZ2F23aeJLT7bKq5D+wwLZ0/+
QQd1Yq7veVJckjf4U9bzP/w+RasTfMfqVJNZ096KD6+o0oOWlSnjS5g62tGc1rXa
erBNDULyOEtHrPbrrD2pjC1KDw2cOxXepzHWXOCOG4B3WaxqBAAJtV8q2HrnjEeL
7jIfnCYtXPwdqyr9YQ5mBfCG9bV83IuyGLEhJ3Vua8781b3KIorVomRBmcc/5v/x
ufCMR2/tZHhVQWEzrMWM24jGXLy7bjmQv3uB97zwv5Dq+P0ebK7xCOOga3JBtprF
9oosJuwJPa/IUGmAhBSG4oiN4RodN5zCBaDaQfaCgiodcz1hiRaEl4KY3pc3I2+4
BeSQ9nmUV1IPOEnCHSfbQjvq90kQLvoA/ItyWG/75qjaF/BE3Zs4dOb4HhU2D1le
pp2pnJILxyGItguBHMcF0v34Y+zo5rLM+xI9mIZ36eIFQQT1lcKUcIP1D10hHN3g
Dn6Nu0NzGmiYlsM/QOpxLx0yXs5u+vHvclLckZf8qXhxpEyPJG8tX9aVel3sg5Ly
eoFj9Mbt7JHOEHux+iJ+mZOviQuFN/pJuN0GgYP3L3W2NS31Ipn5o3GXX3SROmdh
D/QBZyyU759Vhmh+XscZx8NGsDefVySY/rWdz0OIaJXzvFLFLE78vwh9AHaDPGY/
yaCLwReuftTzP5oFI8efyY1Hj2Of8ZV3G7Rx/I7x1m3SHMYtN8tDBcQMXcPTzXdd
3+B5zqHBxQk4LCtcM2kubRgUFhbmJlRcsgEOFH/rY0bjwwMubhgFuQedMUuo6dHb
NST0kx3pAu34T1n4oMXBOB7UnnD89VJQF1mbQF78aM3UlyX6mEYCgDIlvqrAX+5U
DamvZtN3GgKOX673SnzTU0GwJqTCuCiqxo+AY08bk0SUzyyTZITvHt1EF/Eo7V0J
wYQ5rKiik0YthpYYp9Q4wYtjKTOKy/OJ3O1LYOu77SZhZ0k9Bl/nXbUlVu+PpKd4
+mRUYBZmCdZ7FE2QaWwZwdbhnnJoJ0SBkX0GMjJs6vuONQ1VhOcgmffWXlnJCCN8
HcMoqRniKI0Vd6WZeqdsjHHLk9nOHKLZZUPGdbH6uxc9d+4b5naOBIGjjij3IT5i
spyZpil2fUHmXe6yYz2ZBOGMtb0OcNT5tGdzEyt59KWJMUtCapdnpn1X9av37afI
mpHnGpE2HFXAuEWgIL0mYsEk4ocU5qq8b2bX5SkAr8TP7xHddDLUxVtF/FhhhL1L
3QCmtCc0xD+VrYmPSXEiFyjXuezqivkRjl5JS5mdIBsU3wer8y0WGsAcLoJvGO/E
F21KYrHqkkiqL7ZhLadjFGVa9379BXVf6+QVMhW5zKz5zQ7t6MdrtsEcv/LIDGQf
H8uaR4gF9C1FLLjZ6qR3T/XZfG6b/4n8Monbnq74/olnagFXAFrOboqs15QpWgvZ
2INnyc4mgrP+8FfwL2D6So0UjUbGQK/OSRnFM8kHyGLYyMlJekiX0NmncSc6lyB7
bL0kRYy5Dau+c0gZi2UHtsBGu+NEeaD4pmO6alUhQk8eGHvc1+j52Zfv2GP43OX9
EuZTnNpV79LAKgPCHd27NjmwlvapVebL2Fgxc2j7XT7i7z6hVHGhqJ72Y6c3ph1C
yE3/1QIrxp5W9A8gBxv3dqPAFRUHJBcQVls6hK2+aXuEgaR4xsdkZOVRksXh+r67
o83sUXue2osn/vmflI0sVWwlxfW5EmF3UfRlSApb0sJKFkcGKruERB3ti8cuRB31
x74sp9iUMdDHW7vzx/DvPIfwASosUcX1Li5ig0wSZECoMP2RRoyYxCf5fEjD0BuK
5rZli8K2+pf0jZ9jzE1xevt3TexNC3Sjes4FCkAdgOoIPf6qApvKjlwnecD5Jv71
6sEErNzem3sM0EjNmQCiqvB+fcWEeCW1QMtbY/rc1xSy58XBm2w5vlDm7pAnLmU1
cdHBklvrqldAF0QDdENbOP+D+7aSNpn3NjGZY/cT0I/Bo/h7FdzIUAya9b6MZCXF
87lVm2ZIkrCruaKv06RQK7Nhe5sklWhjy5UI3bvuB2eiEQoKP+HY3hHCzZGfOyec
T+Hc+50zC/jtUDqdKT4sWRTZmVSMndq2AL/s3C8YqehsKPX+dd7jQjh3wDh4cAx/
zVOB0ueYBX8WsojcxmyTQgwBzrI6er57qENXFgdxHUcsS53LxcUdqqwicguFEeht
blcvWfZAnSlvL8nxAu+Q9AFlrES8tmNnBnBtUfKgwkMO743g4Nh0YP7BOSMTIPJy
3iOiz795hmTbBzsJ4RuN2RlBpG1jDlkvIdJUdMY+tc7lCxOQn4w6uPSJSK0wLToS
Ql32RRvOIFywoIHmQdb/s2h48TfNv4Kyd3YTq394Sn3HkSfu+VT3+RPTxPxqCLrd
3baE65ia/qg1W9BZK/H7BOTsOgV+oU6jXsYnMjTtewLyJqNpT7N/JJXv0oeP5y9n
xWm9g/qE1i0xSk5+2yq4UYtC1oHBkUWiNWcZPZu6UlHxMNegGq1H7pELu2wGDRbN
n2SSAfVfSwmkxUfVvPOqbW1Z98jjq/icQ1q6aIj+KEvp1moGNFM+VCfl0BzDPojl
aHr406r4gx36C7nppMIT+SAbK1r6ugy72cJ88mX0gEDaIp/MqQ4izB0uO2PpjtZ3
axncaOnWXPYfye15h3428GGCxnZxQZIAuqq+tuJ8IXD6dCX/0w+mLuyiv9pHAZyk
nnt0DCve7E78+ZZSlnE0Ml9Z4aMF9tebPEisICjKayMVPALSJBTpDOEkN8qaVZSh
RFdOQW9PyIIaHW925ZajHY3GQ9g9HCB9QkgpMoDClrEsuaxa0xrgU5fI7/nkCk6V
CxqomUx/9qTeYeWQBgADWx3YukaWxSF5h7phL4igQL1ntV0w0RnNSCSxlSjTv22P
f9/wnzDcJyNNm0SzdOsslzNV6L1L0fUeM0Q+SAUGsB8Uim7oBAAewnoiqxZtkn5U
zn0ADGvf5YFyxMdaKjL4AsZPX4J0sAfKdiRNVgYQcOQ7S73BHIhDO3Dh+kwkP51q
5neFesr6/LHytC9olVGo1LeKSH/SiOlQlXKsnjqUCbDWfMG8Cql3LcY5Dvg74IDt
NwHX93Y+p5lqlWj5VDoE+w4wR3JSlBGGzfH+LoVl+7FAwrYC+Oy3einmGeB3+hS8
U9dVC2gFbHTaMlt69veqI2DXwSViCqx+n0akyjr/eNd/Q0QYIUbtHTwts/ae/+hF
ac6X9c1gneHHDksJLeeSzzTGkvcnstJ3JyXH5mOcqIu+AFhrnPGhgAUpzWBMRCVg
colOPwv2azsBnN5hQDA3ZFf0bEknggPr1wqOgsFCYE+zYIUNmkarKxdduzyJbPfZ
Ng3nSULnABaw7WSwZVdBtnUrTczRrLodo/7Q3JRfNRetucypROWT2p8eXVn0kidY
cMJhEDrU74fbMDHlX032oPiH3IV+yy1i2/rLniOqKCrdAFI0nZbXDLGs4iBZC43/
17xQ+6FwPHkPdPpm5V9BpcWvbkLp50KL5bXncuxbWvwQameerWb88UuznWyVufco
Dzgh5eSrsdmuaw2HBJcy58wk1lJtYNVZe3KxDdrtZuKbP+qCsjsuJbXobUmQo2n7
lYbUTyHmc3saixRe4rubKi/eAaTIRV+NNIaGHqhD6Sc+uq64wVKQ3E67GoEeGGhf
1RRf3JfnHSPljsoMfo1vOV5E5sGLW1UPCkdlGGm0VDC7s5fOG7wTTTJTwM0a95Nz
mHBdtsXfayN4dAHIdXug/T1Ryo06YKhJZFFP0ZE3TgSPfrbBHNzsmC2yi2S60iP8
CBH38RDU6X7s29dOw8E0s0Ln+V2AlUM3J0VFd6d0D1LVZz9/uPo3Qgtc6HUVYhfP
j/4Ivn3+JeIIJ11erKcvxGlMBJ0k+/Y3eBGu4S7PQa+nhVOKLg+tR0LZTG20RVy0
XHEz/hUcVORPOt09kRBiZpHGMB99BDWCbs6mB0O0Bxmux3drFy8V4NfvL0DYaqfm
1GZG0MGE+CnAJcW6M30aqtr6AY2767G5i9VsZFBW1gNBG8CV0FHRsiHjOJisXdOq
y9cElxrwEtQIR0hsaaksctgaon/uV438q4GhXSbhAnx42iXE/nmlNxXp3EYQO5iF
Tn2jC55wE1VYJcfxDC6YX0OJ322kJG8ILmy2va0YmoHxGODV6tWnK2zaSXuWC556
i6lZDUVdzp4rZzRGjj83vlcX2Z84+oL3XftCdN/m2h6JhLaKK2JXwTphCzwclXN5
mYd5ZVhzH2oh2TG/9pep4uAriEZc9GkrzilXTpST55G5C+ssLQ4iy4BZztjLmhuE
RhfvVN3f9d1InZGkPGBkB4C20UDYilNi0tBISYz4FK4YB1Pgkz0l7+L6VFrR4Psb
1qODtkYRAmVQVGRBUe2LjtXmzVWhJKIs6C6zGtfYIKNmrb0HpaYHUQyatxwycmvi
1++X7LjyjDayC0iomMrdJhOhZ9cf/GYr3nKS8d/4VHoSf8UJa7EbFiFQ4CxCro1e
lRX2clIHboYK7cnojkuAp6TOlgxRgC7U1HCmqvDwgk34AydtOuLpU75GD7Izpla9
7n9xE5akt75x95dtTsongvVjgAh6zDpoueMNZlptboEnx9caAC5cCEtrVR8mdwKu
f+zGiKqT8IUnxfq3lp6JxI+FKsPE5isuEEJnBOUxoO9aTq+yXHdBc9+BI9QELsl3
Sn+aAkn4AzecTiZHodP0PamzfBbvEetqn5BwAnERxBafBFlxnaxtEv2dNQO7Tbx7
qVm4Geb2RMn35BVSyqEnHrGV0bJIha7TshHWBzQB8boEiisf0LSd9nAgaw6GHgKq
VXhcrbKvUJazR7tNJrrYP3d8HzrCZzFHjnIb2NDI/uVVqh5HpKwc7H+IUjsqj18E
UX4tCJRoms6L+wxcq8w/ldLCP71TUMyJuGsv54XSUluerM042NiMEmPct09jLa8+
aUK29KP46fOeh6314bYkjwItz66U6zZiO3z9tocBGjYKTLHVt+x/MjAzr3VpvEDV
kXwRtxp9jSoeQMNKLcllo72LQPVora8KnEQOC6SWjEooawhktbwcepNgXHVXldS9
aQYFsuxhijk6+DcKFjjR5XvmN/9vehXZmgf1Nr1T7R099xBI4MAmVQ4sjmuKgswi
ula+laPHFIwF0uoeat/rENjBp+rA8MEqA55z7ViXgIWRLU5K5OKpC2pzcAsh79T/
nVwnDnwS1eT9713KzXKwfiufzxMTx10sFJ/4T8LoBEqDTYx47pZYs/+nzd9IzmVe
kEgECCemTUHO8j8wf5xPA17mIa/pEwUMlZQVZIWEPgsIcKE2SNyj8GUqhrbXyUWO
9YKqr4XT0yJuR/Aw8JnkFn8S7N8pl75UyEOWp7rOA/13JbLaqxLstQ9aQNSCmgEX
+Gh9CO1BfArauTeZ7RhoZAdjSYEA/Ri8v+BA5mozQophOc7VMLC/YoKqyZRWzMsP
MyCKB9apJ/AAJe4HJi299f5aftzmiSBhVdKNlVcS7IQzxx7brTBMB/QktbmO2auk
hd5XAzju7xhvjUlqqyFq6dxnMcqtwGzO7ZbMjNyzvyZm3JsyAaQVW8SyJkUnufzZ
OG81ZmMsAUFutrAMxiRynXALBoaHh4aUESkWUSUKpD/xNKL+iIPyRC192zITJEhz
8GoLBfPrjWpBWr9sywFjN2l2rYLkFK6ir/9QZi9yKkq7jHEtSm4GxlOl15CZA/Wn
0C+hjM6ktiR66jeyOzP0c5TZZEygZwEjwHNNcr8OYrG1aXhJV3TpeDiyui6jk2kL
Czw/kPWMGQl9pFBO2sHevy0qmOsyefBx8mvtHXBZmHBe+B7nY9VWEtFQt/wE4bHA
j+JCuQc4PbmSnqXlZSDWZikJSQYelWVhNHb9Po9VZJgw0y/RSAuSGOaqwDGN0ALO
WuD2fnYnzUMKUIpDISI03Bz/akcZlFxRxusan/xEI0znOHewrRDdafpvD2JcRORw
KYxLszdreNEDD4F2k7TAgxXqIRbre0/YxygqJHlGKQrfkCEmi6oaAEJx9OH4Hj1h
wMfiFsitb0YWqnOQutv1/6nZRfTD4sdegev+8wiTPjVDIZZQhagXC525rKSFJ5RH
PS+iwmcoS7OwOVbCru219ijfA2SW9EEXEMdcOewGn158uTDcaDviPDEw37ofkmZO
Z/znJkzM+MpEqA8qM9lanyZH2XMpTC010uvB1zvoiCRMJQSQOWPE+rX3HZLyJbQe
UXWv0Stf2rOTvo3yS5gPnZ7mC+khJbu5jTBuUrOAcRRBJsLGZsQby/+m3Ywz6HLN
Xokp+M0GRIdJ3EeV1CAg1vmyk7yvFnrVpbpGAtCKD50n90eSHkLiO+nh9idzf1tD
gvLGBaLfX/TWdmNNdUAx4J59jOsjG9/o08vi2eGM+8ePLjGN3Z1D9HSFCt4crpI4
ylcuThwbPmlRwZs1PwO39YsN7k5BbnGayFYAmtNhoOVVny554M+vjCdKy7X5+6fT
j45f27ijX8JMMPpunfDOwMaLt0hiT2eUszPothKQAo+R/5S7zG3xPcLby962CRxw
vsjnhv9clkJiQdvfy1wfZ6+LJMu1wHtkpMBIaF+HgpGwabSWKipD4RFUOSR4Ad7T
FMbGv+BAYOzFySQ8Ek7vSNw3oGr0aaQKctNRL/vlISR3K7c7SW4FRY1rqYnP+Tm4
1xV8RuCF0wqzf/0X/q9fIzPzXjw9KSP7cK8mox+bUOEE5Z0TbiSYp6g15umK6Z2S
J9EAx/vuh443S7idoHqICmW377CggzY6KL0VhB+xoB/ZOunCm6WQN069AllPhqqG
n+JwNRxWqFJjokK//bN4hOt7nxCyYAL1ps8Lqt0ocbLjaVkG6SzsMzMicGhOzC1T
`pragma protect end_protected
