`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hxk8uqyoERpuufifLGtUwbcHKB7Kib5NXl0d9ZUBVOdSsyYGrd3aZCMAasbBig0n
yBnJs4JM/lyjh5KchBEjnZ4vY0nHeuPC4doWpaQtEhna/usXylsE4EEDGqVXOwoG
c0pqHR9Niasv/T6Sr4XS/Gxya4f8Hd81DrduOFDZt4o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
IqBNkhMmPBgrw6LW5tPDLzt+QrVzrob08m1Jry2BYrIdQqns15D+siNmT5kOdS+W
tKiy0eQtbr0RzH+zZeoGkYXDVdHF6A8j7Huq3Ku32sFMOjQpWNsYg6UYunoSsyq9
lixcvSbh56N7uI0DVUlrhhdqRC/do0lxWj3AdZbF2ogAfgA+dbDnV+ooEONQ5HB4
InbFP12Ge1FE7ITuVvHkW22pc8UjVrJihKgYeiLPuIMWWBS2DL7BY49twlCwkVsE
9ZcfOkutUxNSintgp4gU1RDTRR2FgtOZUDsXOPyyLPwcXeoNe9Pmbw82pJUhnT/a
qZngzCO/+tr7CKl2h5CM3fTkgqF6pEwt6YaLPJEvHBSzvl7oMXL4/65EvyquumW9
F3XlMg4kgfuhxpGSS67XdG2fEzOeuv1x4Uu3sUo+JGuK+uTGqktVGBwW/eoZnjJr
A3r9EfX5cGOtaWW1EzExCbt/ILp8keKY2ez+qwp+Dv/yjzyuhchvoaYnB2/lJ0Tx
S1LXUjsAvGwCgQLJD35bB6jfm2hiQ0fYLC02NoqD8cYFkSsYSagVT6I2mHU+9BCW
D+a8X3/U1+NNRHzLVAbUGnm/sdOk05Iwmkr24CPk4UA6pae2Vg5equgmZcy6rSjs
JmnU3nHRDauWUvc/Q41vOtIZwlNkPaQoPDNqnU24gUOuu9ez0iwR7lHyHT8D8tgJ
kZ54uAEkTSFKWztvcYlMBl3b2W8ygiLcxPkE4iVQ5vyHWVAW1mCW8AXUv7EmECUR
ThOTt5QLef94EH4DT76jdSKfbQKIf9PpapjwxgHzfp9jhEDMaBluMtC8V64Vhxdg
brEiGYWl612pw6b/94ZstHxiKS3PLmkRDzQ8GKoDkdC309DbYkIEXCVUtBDinwgg
GVfJuduWGVcPahhcQq1CJNIJxgkWzlTGvTZQx4a5z7JYSpwrYQ5c//D1tmX1pjdP
GU0pk0ZNo4mzHU7O9Bi1smA3M7uG3qkhuHZDnAj1LGIV8vByjGOhEun/+VUjxi+4
R71/DUItW4PKumZg/PM9ZHSWNJXW0GgS9MRYmeHr8F9oAd7uADs4Cap8QQnpidCn
bc5PXo68dFoP6T3M+urbqCrOnIx8vyzPKr8q3+T9hoohvfnCzeEJSzyFTTBLpGbH
1511QROa0i42O7thbtadyKD/5krUjHC/XesVy3iQo8WHni521DzsrOsYOy7GD1Vp
1a6IQtmXOVAbTTBzCvPrXQfX330NGYfL/8rcpBveYLj8ykSvGbCdt6otgrhpBhKo
f9vSTdV0xZupK/BuhiU5GrjPvMcI6km1puB+7GcrdMVqsAwBJ+85wU2SSf1rGe+8
wCWxSrcq6ugaT1i0UE44heEPTzM6z+1mMYDqi+eeHNOvhb2tOEj/NIRQzx1qFT2z
a8kKHnDV+jEs31DMWQ3hQwcRtxWn/TzPA2Repz/Gf6S9fSnUpJ0P2ESvGK9nxWrU
aCsYH67Y8ODwGrEZc6XU7DcB4Po7M2NSloU4qEs8y63HmuoF7qOa/CyYBPkPgHr6
C8Vat8XLKspGc8NiDZDfFNQyIhAAfdR0gc9ipp9sTaUsVlbDV0dxSssvAYl0zLq3
5DBUA0QXb4k55h2C7AJLMDM4iOPe287F8rOGpPLnFk9A1NqVJxA4+OW34BjJ1yeJ
zxtTmDq7skAFAREU/M9PeyYc/9cSPAA5HFptY37/H9ZIdDgYVAsNWn4HhbqCBKDD
U01ypzlSr9r4PNskPuad18yGkDpKDpXOtanXJYyicR/V2uFs0USEN7V0Rx1jRK2d
QAdShvlMKSrPY6eycfze9gM1YS7KDhPCKfnFkqLFwGzTkvK38MtwHK/DuN6VCJvY
F+0KVkf4SbpolY/7Tn6oAXAsbKpzFWCKgZJ08ynlCI3POn9bS6VC5DapzhoGWFq5
S+s46l+I578DFy+z3pvB/7PP9zpsnaL+VcrnR2aTJoSmxVBHWghFVU5Pm7KjdIF0
5dwOxfZ1Pds0RAhZr8SR+54OjJQLwzIO8vyOqR6amPDakQ+PgH4lPs5KWBLMz/Yv
ecED2Qp1VA7wDsX0Lrd/7CCf2MJnO0eB2BErITNktTs/IbxDTb7LtunKJZkq7bH5
KvPIz5/NKduWR/r2jtLcE6Yo2xqV1kazl+oCtHBsdQzO4ZE7l9cRA3IoOq9I327W
vRANaI0CkjVcQ5l+4Rdr4af5vl16TtzoQIJlEe8oOMitvBdOfhLXS6Oc8NmgZgGh
DPjFmHXqmbd2E1xh4eNu1Awc+0FA8D+q599orgMlmugofjyUcWDFicZKsz/evsJX
AjjLgyqhCZfGMlU8Jnr9H3vvWzxbTSddM/h/PI94N8QgAaAWpM1z9On7VW4jZzLs
e16FAdDsJwJqwc4ZoEPMbdNjxw0g/L2Pc0fRza6v90auQTs8WYXr004Af3bWSqUL
7zyhFHKFw1agYwBR0/LahUMhcWP+R92MdSKhLXxOzac37SKmYs68MVcOHn2L28WI
EwKZ6ACX1RCApeHK+45a2RSOlexx+XGpGBrCvl8fDJxE9jqrRuvdhYFcBDiLPctO
BG+PRWtovm1QkGFhgt/8HM+2cIMtxRo6+N0qrW+iehGdD4XgTf+4ludcHV8IeLf9
Tb+UBV3p9xTkPM2FbeSWx1tsmyrittfKdYVvDEDS8ID4h0XUYRDSXmD14GHUl2eP
XsP1aIHsLgnXPX/Cssq7oN3ZP31Y9bb+/kZzXYSjlJqI6NxTdckw9//2K0Emgk8z
If/Eg126xvnrSvQFzlBtuFskAuh7ZUxBm5FvWCFPt+1Vc7IzxtF3tOl89kb7TmOb
MZG53PsecAXHdSNG5CMj/DNNCYWWNA70sDbQXRNp3Mg+zeSVINvB6AZxusIcg9dB
9lP9YhBGtZdH2Brt7oG99L1E9e1MF+OSOn8L3Duf8uPEhxX8MnOXZlMi3WpMj/Ay
GJTs4MlQYII9sSCnjtT2eDwZzXWvx1WVCb6I5ERq2bsxetiEH1aE0KVyYt98MiG0
hCTrgqcpgUTSAcELc4UwWguDSNaKPowmJeY0aUd3mUPuF818XXcxm3pmuVN78KR5
m9YNdaw3wUXVYXAC8zQeu4JQwjayAItCFhuDoWrZ4dzhXx3IM6FU2n5qO6Z5X76T
JVzzvatDLrhyMIVp0YirFM7/TxXUWm9awnyoydASmDAuu59zal2g1wPfjexfVIDd
uNvcwGLvmCc/1SLCKPvkMoikG25uyH5H2QKoFK0DKqvASLO6ADqNzDYsjSx+YQq2
tHaKTB+FHF77gspkrbQMbU3JXwFOiC3MzuMO51udw18BqshbYGheKZLhgG9vU7tR
rab3zUQvJocZ+Af4b1hAKpRDnc0pj37qLg+3ypKra4jBwDqgx32fb4fFXvneR8tM
xiBhxruc1XQbNr6Mr14B5VAgpWOQTuAnegRdViXnUEk/c0WHr/fGxyplhqQK/RxJ
dZg3GU/68scCmDY672viC0KhaNl9bLznaFL+F2W+lAcr6eYdZF/+HvujNPN2HGIK
2d3dRhkKF3Njfk6+8k9D1lkvGz1MrjLjQJHCxxsw6g4THVbq/fGhvtiuglUEMmya
Bo7g9qUHKPNXGtIwGlkCXdDQt5FxJZzvDzOAVnUVQnvE8b/gGb6DoH5w2jU1SSRq
q4Pc9H97dWVDpt9hvq1QBPFUWLxwYPHz8re8HZbTRD+WkfTvws+rRPRejs2Ukvzz
O3mZQweLLr4ssZ99W1lz0ScjFD+72j+otgUcucGQVNvJa8aOACQuD+12pkYAmqLi
9GCTY7/SvlOV6Mt2l/ahl/S0YY1u1Wkzo87zdTIZgH4TNqbSG36iHKYWEL9FX34s
QfNDNHCIVDLEwUtVuAK9ciOSAjcoSx21hRhTdP4zlXy19l4ncnSWkLTNMwD50gnr
Rnzu/SeRe20HyEPHqMYBTbXtOHba89MIAkrgrg37+v9Fz5XDExTdC8OVJLJF4GHi
8hf4XE8JZmuhYXESNQv7yg0KaoKZmjWBcn+sdiq/raSu2NYErkwSWIeYCwipSBwF
WBEBudZLBu+wGMez3/YDB8BOFU2qNEs3bHQusxg80ElL0peE6g6Kc/1zoVAoSJD9
Z8uuLKP4Z7blHSw66O35TE1XJfBGo0U9vtiG7YASBYVGFoOattCSKO04eRmi9pK0
xPqhUNBdgJ6bCbMQqWnWc0PyljV6EbDqJhv1n/Mmr++/qZiprMoLHuVCcIAIy1ei
IMn9jrouUQ+jaqqfACF2iTOIEoHX2sKLD+A7w6karAC11lie9fPP7JChZZ6uEeMn
l6wTzCluQ9wsPplUv8BKTiwFrboR6kcGbdyY9DUboBlj94uiQuuzhPJ5aR/mmpzH
JXq+nPZmjROKe2qcDPmELv3av9yUV/xj8K73ovI0WhHJjfdqnZZ3WuaELu3637Rf
lTXU/ZLfh6tms1U3V6+zU78ihyjV1XAtm1x+yUpWmJ3JHTknZYC+ZAN3jUXhR9Yw
p8bPFEdn2nOsKDdx3QbaDWAfamUJdd8s5pzRx5Ej9uo1wi1HYpbHxkirIPwm69M8
7lTzrjEEJIA5x3cpWm9cr7SU7tT7G8tXorZWMjPrDPiHOBZvw3Wyn/g5b2iJPJ1i
cLkEKaKcuYqh7gEnXRbSVTQA6A9RWew4pCzmKNQUoyhG1NTmGLh1QCH5ZaL8zhDV
M594giPcokSSLOViG2wWgTMNxZaTvrxRcgfT+CQTtcfu9M3kH7t81E7l3caGOeud
rsaOyXg+XXuXM1ZnU+djRjC1irp+yq4FgdFuFozipsm/zAJagNUBcomdcOjHwJoz
OHeRJgKpKC354W6z0vQYupPV7jVcFV+VbsEbaYYvTrBGefdWG1Vji3jwIR4YMpm3
aMo0zQYlPokDoJanfuxqh4Wi74d7x5l/oNu4wi+LOS59PBE/XvWjkF+zz6jR7Vct
rqjJm4ar6RgG63YlsOrMRcgwVIposllIbhegZA7tQtaAOQCMn5Sm9pEpM20qhsgy
foy6FrH6T0k1y8k6/olnOpOZUYsWGVbgIicIxJ7JWfAa0uvj/WL0QwQph/bC034e
1uB3S0+rUq2PNo28C7zdM40kKfKVZ2g3Awqdae75TsJggwuzG2WlPD2PwX/LBryx
zxTBgCvtzMmqLRF9uJ17xvWQZoPMoxSSklnpZ+hreLr4MryTKnBHxwGN4QwGDI9D
p5iOd4EZtmq6YB55LxhAwPUyeOAorKoGqttvGd369my1LHzXDaBjsYqQyik5j05k
HpZyWf29DopbG75qECYxD0UnHjb/T7VUmf3+ZT+X0D1RUdWrqrjUV+roc/K7HRcV
ieUcUI/8gHUx9oBfcSalYObomTN+/w9Fd79IdCQx/vk/fWf4H28BDnKmzYzPW6gz
1dUCm+k1tdPHECFofi2dIYKtiRNfreYDup2ew5+2h9+gneWh8dPF/AfozwazFig6
0be3wFeCmkWkzYpuv+ItMqbfLS78bh/U2FLMwsJC1ga7RcXl3a0wM2g9p/bhXD4m
RiJqKSDmLWuJlYGPwJQ/HGKANBB8txbZtEMb1gE+YOuFbpLKYTIm9xA4ts0xYZlO
TBDqjC8kvzN2rS4yXMjfNPhnk3VSR5H7PIvQFZpdkxM64CLtbb1qxBrlUEHEVIvw
F5W11B3rTohUmZjn3AdWMkaNAivz5Ppk8QTzNdjT+3qp0tHynBkMSwT7t3WhwKHr
kLUo8UkqF21pQVVOwR3adAi1wPhJzqvLvRv+i5nY5m3avk+GT/pmoYAcSuVjN0nX
i2rjcO2TkBt84n5PRFJ63eeRhu9xgMr5PoEbXAcViXRTBDGEvlP4NsUAMeVdXPQv
mOpB9TFQ8W5QlrcFtmhBfHZTQ1xHcklJJMNH2n5olY8agWU6C7FOG/fCWlkFVpQg
nL2czIgFbkoWc/6qf6Tj1lpq0JQE4WdZ/Ai8KXc/JMsTZ/TyyfFCajmNnlCW58Tp
xFhvODqyAkg5efBnqAnU0OUVd3t7XMdQRa8Eu2NycWAMbnSYTsHQTV4jTZx/woHZ
2EVdRUlApr4DSmujYxAM8UHQzxDeTu029UAV6FHnz4Du7+bXl+Lt7MH2hVuHtxbM
TejQhQKaBooauUwkyxenEbBeVqC56dBAWm5dZDGyPcMJuc+uHQ2z4xPjfBhWRlua
k1MEVGi4pBFSwX0KHuAK2dXToP7I8erQemqw17Jay7lU+sa8tgsMio0GdavzMt6C
detOKvvtlybCKiBDPpzizoeIMumBi33f9J3FZIKxhp+/9JIfweUrb0bnGINEIh+t
UtrQYh8MBMiQQNWyxI5/gzdLaFjWmjywAVIfBek4uGdYMGguc0I0/7ot1uDwXgce
M815lQEViZi3VsvLh513WfMkPgW6B8YaaYnSryiJPYfk3S3QoU5wsLV1KngLge1q
lWUYC3rQa+vyRjLh81qV6OYcfQtlRMVno4nOsdG9WVZHVr86yxUCBC3waXwtUCj3
mnZf2flhRzpxhNbKCqr3bhWqrVThUCTDxsXqsT5b0r7Qy/ikdl/nryV6wzL1lSjB
KKU28sW75eowTCQ0c5maTXmLk5OvHLeay0l2gwJ/AukDCZtufAxLfPeQ41uvsJif
m70Fgdud3/pVIvd2edZqN0e5rS5qrl1MLnI3Wu78IvIlRJuTsWoWhNGKkJVM2jzO
N/kMenwqvmx7iuYkD0FcGpJADPR8Dgr/A6jjdxBE+y7uop7Y9M7WchKDyQgKd81m
d2ymUthiMCQP/S9hMi7ZOhiRvYSha3lw3HEz2lYoqH6jYrl5d2g+XXyZtYLCjArT
eEWf2UDFiiQJYThLz+nc6Z6YfKNLkcMQum5EYUQKghC/+L7Zj3qTV5M8y4JjgP85
WWwW2VAdMwfqcNFdsPAAUCIvFjNZIG27brO0OmBKsR2upfNT1gg7Qde+WOtWES6+
8qSXYzvznXpHb2785/GgCwUNJvggNCurmC3JeO72RW/UF/bRiVe1Esp0DnZj5Zdr
4NWgOyP8Ja4bOLWYoikY75/eT3Yq5o0AhZyh2ej+95ZFKzFh81TERyXiDtr7meXu
dH2Qby2yOaEalbP/eMQps6M8BmRCiwZAQbxqM0TjOIz9J13N3KqcMJoUKbl9OrwM
/ridomBDFgKOrWZd/pU9K1tong2IsMQkI/YwTcJAsAkbaxJ6js+PIj+L2uGlHAuL
ac03q12ged904jXAQnKlRJzQZN6O2WPX0Jbealwka6l7wsHwrIgu4k751KvsNnxF
pz3VUSDGzc3FiuWVFXUmWDZ61cpx9jcQEckjE5FEWlQAhOpst929r9GcNV3bi1Dq
shb4hguAqbYIphvyAVUtd/vYgfa8uKQFBpiB8fT7bkeOaxzn5yDXYPIbdojxmPxk
E2y012qAxQ0vng+0G10mlPAb2x/On2PzqMRNlSXLuTTZMdU3RIPRW3gz/pTxRh2n
Zpw1mhK2JOyINDG9oa2/OwsWRS+C09A0sDU0BZFfGm31CBu+wM0Oe1iTC5if64/M
PIKJp1MDi+fkmZrUA+/JFqKc5yAnWeQhNFJOhcWpC2oRFr6iW0ufZW3Qad8eqdHL
aDncl7CmU3rJ5+E4Jz84GJQjy/+DIR2XKSpCh9a+bwqxw3UdYjdrNtlT3EIkXXCX
jyKqsH8lPuqLKbmefwCGsnC7D9W8bGmYNHFX3sxFfgAoAm8nE0c52wYqw06PNj2S
m1ped6yC+qB1f46IyNKIzksBxYsVCFiMSwKOftsipacO6mYl0cBmj0Hb1ONtLzSZ
AML1wtQ3sJ64sqdG7e8Ko3qUbW7xB7KhHqElV7Z93EotQaj2EexC/hAVyokp2V+V
ES08ntU0TCiwBqht7fgrASj5da4w4AF3BLs1PUprEDBB+kwqeTdPvG7sBomIK0Db
7Y0fwOO4LetgGgIOKFZy+w264k0VqQAFfmJZ3qekZ07+RPJFD1bA+e+y2rxWTzdE
qF7RePXiXa/AwhYRqfy5TsvWKYd1x68t/Is0miJ0tQh8T/sTsscYI1PbftOQLV/u
2bzbObWfwcEAOKkmX/HixbHIeG/GDBWkj+PwT0MAh8hkKWUFyFPDT6lncAPBLw6z
Euc9OSp6kWUA7cfmucy8EU9RCMsWJ85DeLY8Q9EToy7Zbtnj7LTa1m8MnHDRrTdv
K8JSjTmED2eBYPbr+YgfkWInzbnfSS/26lBEU0oKSCFN8/8t1YTBzDiGoPbMPl+c
yuHteJRt4g0JR8hH9TD/q48tptK+MXY+0VjDNpWldUa8bGV2M3g87edB3KmJw7BW
g+Hw5lLsnN8w4+TZ4Xcwm9hLPVmlbmATWl+Ia+cdiub5ooEIif1TqKSd8ZE46fJB
zkZvlwLfVkHHO0M3jE5aaJiemEgZ/pGNCsPzRih/mwMsfbgc9DUNsGF10fZolVDv
22XT92X4QPsTHXlU8Prd3BcWjDvZzB+RfHP2Iy/WDSJ49TMH+7zjCuDF4mjLGlnD
Dfx6rh3//9WyV1iNqgiQlW3kWI7ZP+91INyGNVEKLuNOierzrhUKJqYSz8D0vwJT
6hLNGiLI/dlCD7bUkJNrKp5ODb5CQL7cCIXnPy7uGlcV+IKa7LANMxpVttNA7/ns
CIsa4hccoYBcE5UpWouY7U+kjWMnpZeQM4uMHvTKZBjusnNHGUDzWRKhYbS1CzY1
+lMbOHgzi339Yr50Ho3C9a5427ojo4FgPo3bLeyKFHsQm5rWzpH7Zzq+5PVkoVSm
48QahyrAuaWoB77Nvnzp8Xi4pYM2YLyK1UmzNqDiwddmX5YhWrM1cmIDuX45oqx8
9DV863EEgvQHqAEnIPb5KH5b/eaP80oTcdJIzSTCsVI+YQD8l7+pJIJMtLO0m13f
LYxZ6gXNSd4hxOVemBDGPVqFGa/ZPvevVZEtrXvmezTlU1ezfvlQLjomXQqas3Dp
MMYw465rM7MwvEf2VTRgXhatr0y6fh+dJ38jUB4b4j28fM8i1NVMEVf5eq8BY53p
2BdfzMh3TsXoWizsCXIZALZMSNYbuKASScpFidHmWkYDlHfpWxcDk6NQ55jFdFri
lHLOHRavrq1TgFoPtqvVig3wy0aEI6RY7PbW50x3il+cVUCNTIDpfh/MZF60EPCD
+vMawZDnQ7VHeYePiI6bxW6xl2lauRZhCzNDrj/Zas8+0cgmTeMXxec5kr+Xqycu
462f7f6S1mYmz8IoXc/YcwVkEScXZwW3vXD8vDOTR0Fj45/0MCbY2OKCyv3xCoMX
QMtiKv5SDVyYGLmcckQfhJ6cIlzsGdsHaOOOFuN0rvFAUI/0GeV0iWw3/9fAb38m
l6B/+zUYIILPcdNs3QXXc05RW6ikWqTUsV+XXRbIcWlW9xrAsHzyWVRr1Km5SvpN
NWhTS6gaxdQbTF2OHdgC6Tq+FKiSlZPhwXKEiFYUZm9iq0zq+jZ9sCGw7ySLRdOA
HmQEwCAC6QYOmA1dVJvqK6llI6Ylt8cNmnTzVrGd6/w=
`pragma protect end_protected
