`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aYiNkZz63al+AWRnPpelC1R/HXsbMjBNXYKF34DYdVnLOEdTlUN3fOug/qxLs/7G
kfhuW81MNJCi3k9l6FteKhx91MV2Bf+JqADPjdWrC5E/FnPqbf72kCTnxJX11POO
Cc0s59+SCB4nzovIda/mhmCB05aSy5XU6AOfMUXdj6s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21904)
YnxKWXkwJcGE0ZbMP8fzskffZ986WUk2LjGjV4UjFZFyQTipvM6bsLC2XCW3PsIS
tLVW1g0sySYLjglfWu0PecTb5S4B0y6vWPdIzj1CptSyAUS6kcUeaHU4Ukms3pOj
fYQbzLZ+f+SrGgsV1ae/gUTofqgtg51z6iSv9nfo8h+YbwDb/JIayZACjR3CNqPM
T4fbBoGOgFj78uY3KrhMhRjtKU2LSQpA5KXxUlzqSbePwwkACQjLFR600mCRbH+5
x0SINHziGXVRJrOX1qF8EM4tYGEFzM/AtIq8XMxf1NE3qYaYa4P0FLwZ2cfsicBA
rb4htCciRnTI55PNJ2k5Yj9XmmQF/XFzRS65vnkSg5ZijSlgCbHnhxi7a3lYen7h
XF8V5rb8vU6TQaKm1H2wjh/RzP1i81scrUPc+srZyDJpyBKYPHxDpue8Ie0/j52p
rYzqJDk/HxvzrDL4THe4uP+28b70dHYxLgNMICnbcjhboNJNHdBs9BrvQLb6BZWL
eMwTDcJxpnD7lzcVgM/oiy1kMviiaWmXpNSWIYmcf5MVwyavWZVQTdQIhF5aOgkr
VEtabKOBAkdS+h49xFly1rr4N4L+H0GjUzQ/Z0PuBS8F/Re0rvV5E4ifI2VbTizv
w+vSbIeQcQJlTDEScwpv8XGmiy8JIlKeSLCybQg6+263yNlX6MifSfi+eA1WS1I9
Rg0tV2eBMdMy3F2UyubQ+YL+XHo6vWNTWn6oTGSK608BeGuMQIL48nyE8AWFmwxg
9PyT9333XvdSszSHeCPbT2i9HjTfsvNSzIeS3Epa9tY1D/wE5axq3+p9jX+u9VQk
Khu84/i2unqln3TluVNGK75ZmZqJGXnZytJFrSmYS/j2h7dfXNxykfYABFpGH0NB
ZjX9D+sMWSY/UNDJkQTa28hso+C4xwEHYZQftVyoIze0pozKP2UBPCcVBlBFle02
L83sT9Mr+oFhpK4tEeEuRd0ld/sW+XOQRb3lGpmCL0nd+OZOApiLW29iug9UEHH6
y8V3PuIZbKYlb/l0ITtdaaD84qNelKZjUn9HFVSmy42tAppCi/EM1aYC4s9VjTDO
2iXc5RwidOVwEoMNaqA/EdngS8+48nVY7H7KWxJ0U+EPKJjYeX5KBMhP8BtjYDLb
0gVRVvrCHT8kZLiyu0Fzt23BxzbRYQmveby3ok8f7nvUN3SbuUSomxQGlpckCBX/
BxMNCtesbOIHb22ZL55geSQyZHJVHqsyQzyNh//ZeqIeBZwcgSw5xMa169Nsk3Wi
J0Z4f1UMK4j7U8DZpGvj2SkgIbOIdkJEO2ksXuP31oqvSOFp4EEn3OFuMqYJkmGb
gZZ/e9WEnmpikDmRFsJSoPcfnZYLZwncSYaFaZxcQtPcXgG4xxq6eK7xH/IisrdY
K+2Sh50aie5taC39a4mOO0nV9Lekl+faKA0g63x9wMymsdfgqIeNRbLU9Wf3WlgJ
JaKHsTyU8B7VgeX3SWZxnPc6LMWjn4CU49NIEVGIEKSK16/d3NVCQ5nupib9Tnak
928tpqkbGx7QIv0/DkYigWm2r07WrEF38YV0oSNqFcTZgY/YUHO4oSzbN3AzzKMt
sghDINNDG1EIQKp489sMOpD5/xub0z1iHPoSuezAzbpm1ewylYY2ybMo0WJN0dqz
WwPUEwYqgdXA33DEakU5JdlnBlg2Vrr3wOUE/BOddmmIcJTnCVtEIo0qYELkAFGz
zB8OGyMFfMQRlN/37GIyy45t021NXHX0ilCk9r8Yxjl0d3SBYjE6MYDP9HjycRwR
Z2BreM80L2HEziNUOWVsliJpJfkev1ieFH5rAeya/9EVjElqf9JCrZAH0J3Vs+M2
g1DAlq49tsqZF1wmmQptS0KB8Gl/GepILS7WboVrEeZZJ1XARZUTdwDIRyUapZZd
AiP7LsXHxlcmHjGGPqVGvT622HFbMdK0W3iuxtU+zbBtSIkARK5Ff6aYDr2FQHeh
8uyK62dHl3ZrLrV575Yu0yMw4o84Pbxl+al/lqs32YH5W6X82wOkQGsTBvBMHN43
FOGBw+UclVIshunmlZ9J0pIV++a9oufzX/QR6jxEGJpO2nkgTSsL/lqjQDVkXcud
Vs8Cjdl7nWydrRM2KInfIj9WvghjEIW0WnFa9H+O/iL28pnj3KzHHNBYRmXU2UQF
FrBXpn0xKWar66NQC6loA5WRo+ayMAOVsT6n2lNdaued/KsrfuBbywV6IrLWp/Sd
vBOBKZUadZnwQakgHmv8BBk/0P6cey1K2WOa6XQbkfWszQJ+07pV5bz6s3nxZ6iA
mTCQS0RDYStXEH7f4m0QJ5SVxj//U0s0OvDT2UzqnlaWgxxFpagUx3Z+pBWCabJI
UwTfzaj64vFKFQHvUk9h7Z2dyqndVyDRMG322THkrR9DmGXITvv7dF/DpKiAv36v
dKCaxESmu+6QHQzDJbG7tvVo71rT+mCNEkQivWbxX/AZd+VyzkfFZeUCHgoqo2z0
2LuQjf3ZPE9xbHNBbTc7lqVk7QcYCKq/3Cipg/xh4VYqyNHHug+Cv4mupxsGSRMa
9/90IXCCYbEaeLl7jQAZKqCIUJ7q/W1jU4x6Imm0n97NCwZXFH+KXI3TO0WHQo2m
m5ivkLyFLTnjdY0l7M+2yxtJlaQcC+szsZ5ckEC+sygCqXRR//ejdxkIg62L47gZ
7OpdXDT8bMug03NorOpbb8HqS7Gs8E9/NrpPr/ieM6AcZ97qS7D4Eq+iUE3xc1bp
+NoHQMs2N7/lAVbKKh8oCJHRaavbJ82/Vk80MD7l/QPi5OyUfhs50OIFtDNkiwvF
86mLotGWXlcRYrAAE9wsjXiY1fNRtjTOEHM34f1IKB2o2owgPCxvYNTmzt4bw1hM
u6Fh2L/vs2KybnrpunOW5S6pKc9UORGAPK2JKtV2c9CLBiX/rjoxL3wQRY71irOj
kOzRNbGfRhsXNO+sGRcybo+ViGJ7/20qdefRhhoaWi8iBSkCW0phONmRzqqu/bpE
lmY7lxpX9n/WOKMvtIB+vGFnlFLOlzwww5opWqjhSaZmtErfHvvMe5eafZ9fovbC
gILGsSpPCqkOhNscB8OUjg2t2/7UbfD1PWb6tPItf5iHPGWHU3Lr0aMIUOg96yuY
lPEYnqjFy5dKsPBLVKoSwbUWwlA8WSRTKIbYCPqLIDn+EmQdOwTQtT2+gak1yG7B
klYmtrwIY/BfdJBrXyp6Qa3fA2M5wERXydPYBvoXx+Fdc18wan1hiW4ot1ZPuBxO
iXs11ncBvwXkMLipsn+hLbZvs2vZq8YfJShn9XYiHduFIi95YudXWZLVpZU3Qp+a
TSRBW+onzEy8qlVmq4ct7gUugERv8Lq/KDF64V85+3ZNwd3wTlYn7/M3aFSpVbh5
5a/QkLGgfzvmYh7AR7MXEdG9dv6hc9D/HB8HUajnEjv2gmdnxw+YM7Avttz4W6Il
OabmNhYPias+bU6Gs4WGc5KSiDuZExOj2H3yPftF9uhApIeaelDDIBfXmZWwppDY
RqY+PyPAXRt0WXvxb55b9CiPFV8h5mAMkQ23v1orMqN19lqMD8Mpw3TDwtl/4ztS
H/cWfxaTk9TfMN54I0oG97pL5tNs+/Av427d7D8zBeQ8AyHkjyVqGKtPr9oabOvR
LkR7Mb0PLnoDTlR7seTRhxI0J/SXTDvX2IhzrHcyraO6hD2t9fZE0ILHmrz1hGrN
amjmS4001t3OfKdWkcGRbZNHqAxXMsMpsSAmzEU2N7gVKS2akCK5JCSAYaHmIyCs
rxE/cYZVEoWFOcBG6KIso2KPdL3OArqapjU1bZBnMsfaTIcujNuz3fGJaUJz89Q1
tLsWZjpEekkpFkSVNXD3ZNtfbqtYVmDgwrA9zXxHc8qems5eT3MdPXmacyWjGA5S
p9owb8++5mN8XmW9gXKiHY6ipPfHU9p6BFO3jHaFTfVW9cqIW8FbVMbb4dYz51JP
nS6jGJZqiqMffrsoG/lyNLhHOYPvG5+2hgtbRyr7DxJFVFqvdHhrwYeuROA0wVB0
3MhLD18U2oON/vALKyyMkEXGOPHfU2n+4OmPaXutJy2JctFTH3VHMU8+Yec7phdb
q2e8eEbI/5Oj6a3+x5yvbikpEa7h7l+D/2rj+2qJ2jd7/ZJ2KY0cinU/6vtjfzsV
TxKjvCP+/9Bxeou7YJvJmCoNJ1AKe1lqwx0N7EjPakZAv1LZvUOzuxMhOyff5GhV
bNCfAriwMZyOcMTBpAbC5Cp7l1g4gveelbUNSopiJb70juYPKseX3kq7FgzIkx6/
B880d/8QMYO+ccCuP+IYMt/N2ntvKdTLnPrX9lo0RWFSPQSm7wCKQIgeIO6mBEZJ
dR8u5HUbzW/2F9tt4ahE2NOMPp1BcDHU8hTlcJGf4yM9eia/FUNov0rpsCisvHQG
9M4hjNkbHmyqlESGTkIu/gAtiOvjafPeg2mQAFnC5tTWOsyJkWIx4LQBamSxDrME
HFGeB5vewueEMC0lLboiDipvE4HpPWsySZKgoQ/az2dj4uvcVCn6y6yLSsZgCQYp
Spjseb/P5DhKPhJkKBq6UCDIpQn2/lKaQp9iQx2xRDokOruQdBHyfnZQKdMCejy3
jKNNl06vrg5mciT5ofy+OKlrm/SxCV0DV4XJXcIMgsy4vMwzrkFWNTx6oLGAOnTu
MHJ/Q3LQBZnE0SvNZBhwdk4b204LVvSa/x5x9RrccZjh6ot23WphpBYkR0W8FHnr
5ycGUXfPnOhQx5kYw8r7ZFZ3Drq7prOBJVQRK8rXGHXb06KZ5jEuP/8bG7nq639P
qY4/h/M/TM7cReD5H/8TwqIaMryhgH/7hcf2Gv1Eo+uY8FnQU1isPB8g3/QstxNb
KQckU2O9L1+CwEkqLtIFLSpxYoK6+YLdUDkZnXDwa6EJqt8rPURW4zme3pjGEWwc
O+f/dbogbd45XQfhq2B3gt7IClLhH3EAEThJs8moDmMJHQBY2ccRAIjg+2cU46Kq
X8rj0PZ55OEeXyJJYDt6RCCKfCsG0j2mNWe30+k78FRp3WWVHmGtEX9l7xI3GWt+
NVRFj5tz2GSTLJrWK4VIR2zQzkDeMWRU3hCEaxnYPlqQohLA+FaKGDV5pBNGEpMk
GTsUMETfhAEa8PsY6VlN00msECSS+RM8TbqO9GkoEIBbIRgiktxluNFLOPdk8eXp
KVJb1XdSjIpXgQPG1SHDahc892+/qAxrt0A8HfhCrECCTYu7PWiAA1nL3tcag81N
KiC553V7URdVnZN24RsFM8y0zUD5PTMko2tu+gpaW+wv8xDvmWbYN+zzWt3O/cVO
hx2EKJerM5eiZxW1j6Xqv3XHPf0NMggbxxd8jkyJAzJYqDyAAxUukeZHWNya8pvJ
YH90n9Mr7SApwEoHDH05TG2WXJby/M1rdXt8wFuJnyxXSsaKkg570Y5ay5/Lwtyp
JHCaIDDFezE3+c13Zm2fRdJrhOHxcv02+c6uF7tvFtE3kYxRejlqOavWYvxPKFoY
JVL0jSsCKU51xw577c9cd2pvGgxaCw7rSD9iWzFB6Fzj9ozzwsST1BZXvMEx/VmD
drAk2ojYaEA4rFDcxFvE8jCgjcmsRdb6UMs00OMleNr3ooCNd8QDyEb9ItdCcX4M
GWEujoTc9hZcbOGynyRYWWsCNnzZTYcnd5rGBBqqr70NX+hv7rQjwNJEG+VELzsa
puRtd6wqI7GYAaBo+mISDcP20nbQWPMI3vIWyocjDanNEqmLl22JM6M+JDnpu6NL
5sxNVdhOTPli8ZjwtiAqxwdDLRHAA3Wv4TqzPlxPSVUDfv8BWhi6c1u39xvv+I5s
OI80k8viLfbpxbcGJVZAMm4+pLZ2QbEo5Trg7Un/6AqHsuj4LtOX8qk99T7MWSkq
sRxqi7V1KMF0ooecQ53C7+runs0ATWLsIqx5ACP2Kfr4LmCiR2hXFT6Z4uHJ8tt+
2iW3oqYGBun0HYuXR9KsBDBtMKSTfHT2+w3Osw/guCilfRhLYt3Ak/l+UkGExC+4
MFBv6MoqlljUEgfN4kOhOa6v0ByqI1kBQHYTz2E06rjctb+q6BynAd27GRyDr6yg
sfcX6rlFASOKitHXHTgaATA5gt6AJv/+F6ZBFU7TypOLoz6OgXd7YR6PPQGrAL+Y
udI+8jxsX4fpvrCnc6vKPrWW/Rc9NHOlSqhOhSUu7hKDNQ9OrPZRHvXGRZT3BLA6
VbaWEZrcCyEXmzd0ipLtT3dSI20U8b3Imi03mz1TKySywspPRkj415uQCf3jIqsQ
6GDvlOB6Nqusm9DB9zzgWLXI08LAhCAc4BY6ncEr3pEPgeFuMgRbCMK678YWOfS+
OVu15D0YWwuInqNY0ig48hj+aPBwH/DuEoVbrgUlWgqgXHK7lLLF7lfMngKJpn10
Q0j4XsJ4EptCOhQZreaRv2QAcn9Zjk1tkUPsyCP4KbLBTZrJoyXPlOVcFdPyP5cE
2bey48+Q+G3AgS5QbUNN69yqPEHakwN451bXi3/IF4u37a1uFh/XaODaBmWne3+u
irxag6UWapbTvx01nzzpaSNP3fWDdnjyvoMEq/NIyPyFUtAVMp76hwD0O0RHY3ii
ykWEhIW4k9gV+7y131QxAXbidBSf8udd1yGkTq2vTqjNi3g0gDFz4JpLdGYYJvxY
t027PDjyBcen+2LEHoFvwGnV61YXf3Vf7DZ8irABTLHBbfNp2TPS+XCPk79LDD4U
PjQLNtEcPCUkxpGKhHEHx+YpC2yVgan/ij9Pf/JxYuS4sozIgrZmP/viBoELosqr
Fgu3P/KrGeFTGMLcqsI5qGLCy+oXvxvNmyLOqXA9gCLbL2r9k0lZRspA16DFXhuT
qxpsI1K8xNTfcY1rwrGBE9VwxC3gE+CBlygR0tEvHtC1XxWYKkwBmyqm8ChH1b0w
b13zHE/i+qbYwGEBjxqhB6jItB5gU4NDk6NAHrcyIrRcnJKJ65T+U2p0GBxUsxy3
U0usJNlXubPrIHP6ikPtnXnNqgReTdMOYsRxyWM69eHH+W0Ss+nkTAjtv6fapjui
tPv6uNy11KrqXcZPeK7E4BUvxJOhHVtn5eDGcEdQDQWhQkZhWTKShSZH0LbvoAz4
pE7lqe37sHCFNDbJqSx7BQOQ6qDJsXIzhuP5R6KjBEIcDqRnHwdVOPiQixz9iO/1
4Lm0qYrMhIFmym/DI7kAfHhoAOQXsPLiyS+U490r6l8IwQiL/Z/pHhp6tREROCF3
Aj+CSmzbnGpwrZno1+wuluBL9r1yqrRKd/Z60ieVLvWH9q2DMtwPc1si4lVbxrCV
uu95NJSwg+VJrcBaT87QkdrH6WrvnJdPQi0bxxyNW7BwSH+Rx9P18rqLrJxubL45
Z61bXZQ1ny7Dlf25E58c90XG1pGWFuZFr5SVpnthRU/jKk1nYCardqmEgXPRhHIz
F++dEqCTjJHWqU/3OupOgRW9czmvPKOPKDUlSsJF2bbIPO081udp+ADfb5S+jelK
T3aI8/5UFFFvlMxDK+VwvgrD2OJDk7cDM6Uduz/7t+s6mL1dz6ob0nPvIHXW8H8i
P/TCx0JGRDPUQ3ZBIEwTuXkxlm9RstxxE2t4IgDu968IPd1fZOfGizfdnzX3B/YE
OqwCYTqtJOn+6vk88GnI5EBFKnd503vhH/4zATa1hoM5zBTGugtI2PF7iyWuptuu
9lfbm0yd38QLDDkbcr+V9wRmka3fSrpyWXyoTnOK6yEyOjBHVN+Ha4HMeYNJkIHq
SmYTrLT3dTmYTVqzwTEm5jNuW9jJuVLWA6Wj3jy/NMBkLMNfTdZhzZ6Z61dptJHq
HScea9s9jWe9vfFPYUUZEUlHLr1dhL53P6ly7q78DJPlGAwvx+pLq4+nSv/Wpp+D
x6sPvr/EUiR+k263kgJmzHCkmIiDcs3bRlyyjuEbp+G4Ad1OfAxb78wpWpQMFs9a
gMEPmt5K7QOtpBSlHOYyMdYATyFgIUJSdmqx+pIryvogLygLb+IFTMSM2fX+6bfY
/JdkXLWl0Kmg5jQ02lu+FHjQ3bcgWGoI1A1q+fXL/rUpdl6Qsj0LrJUu1Svf51n8
HOeJ+9Y1MKLtwbd0zJHum5GYjO0CmAr5lVzgOEsBVCwETO1a5DWhm1sHKZTTer5S
FQ541yhyLra8J5aMO2pqD3/+ppIAYCDX8/lM1FUxa9cxF+8jvqxy++TXIxxZRWY8
fYWjHdvX33B+nNK2ucm0y21uSypCVB7q8vOvWGN/db5Iwdj8LJ2hypNJqEMtGWQg
5s7Z2i+/RbkrEagGyGYTe6Jw/hLfHktDkiGJmu2FHf3pYdyTUe6bBaVr7yTjCY48
kfgy2y7OT2zf5YfuDwCmPQUQP42mvspZbQATY3o3p+jQmtRGOjYtrQvEafypRTnu
+KfY39ryPGYGovnF0nTRNEjbk0UY3pd8peKgl5/pyagjWPQZBspKPZ/Zvn+V7g5r
rU/90TdDaGK078iDpznbmTaZ2GiruSR7DKOVIIgzrETBrwbnTWwmucxRKH7l9LLL
7jOmqkanX5ozgCs5ki+HDbVgnkot2s9D0gTFOXGgZcVeysLo/uiaFyd4B7CEXCNX
APlWpki6zjEDhBdayfOQhgDMpiGjVh1q39AnMCNDRHRgIB67h/WibIwE1mOK3A31
LU6Y/8wI0WaPtubQCRvO9pSbgLGGCWgICGV4HOnIxyvug3Bsn1F8W8PxH2Ipr6gk
gqmYSoQV7HAUNzuwahU4ipZeJw0jgi62dTzkGfgSprMycx95Yc7npNreBznPHKPx
6ZyxfiQkY2PUKksSfQhId+UZUdanrtRPSOqx6gUsQ0fbq1L5OFhubTRNmEFvQpZt
FC2gmvYVWNVVg9ddLhpTxEgkv12sw8R7b6ucbUTgUdoIupgLgKXWpjdiBJEqvfQk
G/HyWulWfrRY33N6mvVT3aT9LT6lFZYMrUE7c3zF9MT8EnLbKWvfexPdzet8+y6H
iDzt3UeRdTjmznRTr/r68DCHI6dprUAKcoRetqGc2yPuXrjp0/P9kaDN3V5+U2t9
EKEyUZmqc7S3guFgzsjoOoeHar3V0IQdeh/QuGbekLWQcgFbL/oF4/uzmsJU5ZBO
1x8k5mhBJOTj75vIZ2y6NYWiHn8/WJtHSbS8xjfhzXhYPRxZ4htiMiWHDk90wgfY
2YtmoO6faFQXFPwSB8z99iie5zmjuFF6dpAYqYJ/kqs9yBWbdTIMTSPux8I2OxQN
c+3egM9Me9mldrSFBPeVfPLnWzkXvz6BlaGKaxdKfX12A6Ny4TgY2FYnkVFv/FtF
Braku/BJ3zc2ynwcRzdGbZR3gse/x6/kco62K9vSssgwV5/LYEv4maYdnu5Q3dQt
S6xlsvbNgTIjPwizLSgylzV6NDrf6Y4F/XuNi4aIyZq1PoP6jPhimMgWki3IdhJq
9ou9OGH182mGMRJc7YFn28A+KCV5Mhhfsaabr+u7tzBRsP5TMikMxcN9c8NAMfEP
8jBeUCS9OejLm8V016IHBVq7lDeGk5kJXjG8x1W/h/AkVibYQreUdc3sPDDsPqCK
Eo9jDw3bThteJlu3Cu6DfmuYd8Tp00w+P+QpQjyBJu9iTG/z9CtlZnuWWpsEiMXM
t9hhyFDdm3UZ0YHfU6v+YicgdzyrmrJq5vCFETDtWnW5eWsEJnaH1Luor2QquJjS
HhxdT1ZhvK0rXyt4pAdVUdFmw6ifxkx/4h+DxFpHpV8Ln15igujy6kCPVec4sXZL
XoIv/LzMY2HWyN5cAfk14IHqhEi40clC3pLPAujuQX3j3r3ffcVhvaNB0MsBM1TI
B+6CfdMLff2eeD9FTjTCGIwDIhTBxvRFeiacQHZbY65mbSkeLjHhD36kkNiRwTog
hAXtxydee574OGL3Gm326coOWZJuiv1o+m/km7n4sAI7dcFAVmBquE1zXG3y/awR
Z/pyaF09Px2IqYg67KtzN82+k/tOQcv4gMOJwhaPaKFu50O6Xwf8B+J6ZNSQQEJA
yZQTLKdBGAyn8mw087uWsnBXmfhgebuJd8u65a0G6jYIyD98ZX7/mE6vp2mGGpnL
vpYmeH/cF2cEqEDz3yOkE144/IaFXeL0uMhb7aqiXgbl6LDFAsBj/i30m0ETESMF
+v9puFJUvFagy22pDBCrmDMZCxyw3eI6Dli16k/AlAO352EIE3f+0NLH1gOycfM/
CWChwXj6EFP5VSymhth4vJb3kaeiNJRW5N6QlbH5n37maWEHxnVzgI4Xp49L6p18
OtKsQzaw0/IKWe02T019PQtJvp8XTHUUorpI/i9DFpi1nhGp3wsNzE85R7bP59bJ
SMWeUw9+Hug1RVZ2duUEhaqEUTAUdKPu485xSdQDPn+NVs9lXPqyIODJ9EzOthYb
mA3JQ1P7p1hv15wl9c1Ltem0SeS+DTsYFDQfeH2Nq2rL1etnnOQxsbJUhkdNjBDT
JWVm0+bJqNE7cMFUoE/u6ZQFShgbyWId6oh6mZU/+c7bif7U15pfwuIvU2S4qKXI
WM6v13yqYVjFKOWVBqKITdDz6hqIjcyedqDWq33syannJgNHbZI5jC+JxJ4r3jtN
gPNbQpwBa51gdoRBdV1hRQd0+dl9LbJ2NzUvIPY6uGYU97dKa/uaPv50y9VZ6fHT
NP7Dd4GfmV1hsyAPfpumlBbHZvrvopmo+OFct/vlQcIQ1kFhyigPk0jAJvRhaIi0
C+/TLJTkT75bCEDnVOL11RNIwKHLnDU+PI4tWOlolE3QJ465R27vZWI3bJkIcvWc
cWmyoCIWX2TZ9W7JYFN+Xs+GOYZeCETauX8QnN/lZRNwewU0hbiOE33IzgUXVXA0
Qi7CnV3IhCcDV/fNZU9HySoikItOqM5T6CzHlkAvaPR77GqNIYPWHVJzB8Jy/+tf
Q3nJU44xWGzueTe7/1TanALQE9+fMlkhVct4LQy7iLfJDJ6xBb7utGwFiQG1ikGu
4ghLA8iiX7UeWyTHoOg203zxe3MN84QtjcYiUQwsAic4AY3roxbRaWJTzNiM4CMY
e73ZLGkaqF8w7pRrDHrOzlFPCk/hLFC/yXQ1wEh6uBk0OiOb+W/8MHfcfwlxqAZh
Pyf5kU/VIzA2SLL+KWpIAZ4esg9/pjvPFRR620jzfDUxyJSE7I4BOlNlTkPh7UVx
D/r3bkHbom6XY/I0tQEEPtj5+bdV/HcVRBMZsoc48NGZu4GabhdpxLeK8YsQlWjZ
CNunMavih+iH4vaqkkiC80ZIRZDMehQyPaTaPXeEk9hELfrbDLKMcMniFoyDtJ9K
i/vnn7hj193xkBrAl320Z9dQ3u292Z0zova69fUsd9AJk5hOxYO4YCylewqyac4V
Davi2x5m9SUJaAYBrncmilz9NhDmKdITq1dxe5jHHFbXAiMpVDKPWmCyiIz48tKp
hNkrgAGtBft6G1zekYNakF8v88HPvwRZN37ba1yeWgK613E3ihtvQKwKi5TbTVsJ
JH0OUiIjfciwByQMVVb3osTaVWJKQX9QuxWWDDzAY+2jfvRFB4KDKXKCyLx5WUt0
21S4iawNqui2X4PYk8qB2jJy21JMoqAEQnaRPhX5iB7Vm939topolJpmQl86DkKV
rfdOMt8E/M4pCAwq3k07AlpIHj8viRDiwbKAAE36pSGpi4bvWZpHM8wbdGpfsiln
zeDoEZNqUo08XTTQusLU1GK04+KxvddhHadBPZyYm72chuRRxzIc6nO9qC13WRqN
60Jus9h1e7qxQDJiTh5JPxrwpy/Ya+MCaVe35zBda6URrWRt7I7TK5KCiEeZ3q6Z
d/KzNcvzD+5Ui141e4h5ABqX16x7wCul4pVUJ9Oe6HqZgpfCksN1c7D+BYby8Cgi
kM2OX1Pji0NI9TAL5SDeW0o2a+/dd/l9WkgmZfZLfFD1aWOYdwRpOPfLCeCH2y8E
sBfwa1JwtcApt7sdzSuwWvXQ/BOwuDJFAeMg7H3PeaH2Ha6DE0o8BlQZZPF2zRHZ
rhnOnlUxyqC/wfEvvgbEfr38gWaObGT8QQxvVwRssrIoNHbxgH5WJxX2xXZvbPFZ
PslC+CpHRJkYGEdWc8cjMzWQn/wpZGl6U785piWoZ2SGLTZYBTzr468MHdrp5bBd
g3Bj7lmZCbbawMLmaP8XD8gO+EEtnunUEhd25MVGgWySzcY/iE6BGcwIgBEdgLVn
Cxypsn1QkCPB5+qhqzybXSf6Zey12A7+IQ/TuP7dcouEbDQLZ4Toyc6on6z0vtQ4
SR3hyhHHRrXzhye91bI6TWmoy6+n1t5N01AIHMuqQ/aIlQ2MC4Dp9c3vYtX1a16t
eoqxZ8jyRgElh+ehe3HEAdLJuCqarM4Jo/8jQyTvDs6SCzZOxcr3XfzThccjlFXA
wdZobgpFqIMcHudDbQO2I+0r0lf3Y7XmM+m82juGvaA+wcaxfFBBK0ALUnrA1NI+
tvqU9/BkX3I3ZT5mHoVU6IvSPEStnu90sb0BWw5lwpVSWlO/NCDP/4sKjQf6afl2
S3CHDFWohVTPHavf1FEeZuXYVPorJzeYvJi52lIV7aGJOURQFFQcPa3+Bc4sWxDb
tpnCHdOOWaFHPEe+AHziHGq6n8kXxqNdKWWzzK8ljY1++SjpMcFr8Zp8QFG1Onv5
R9/xZoCvZCSESQfx+HW4au9XKHsFphLJr0nZTDEhFXt7RP636tN2hOCRwocA6oAX
dJACfKrkK6wdcCv2Vw8JF4Bn3MPA3yIhaQ07ZlXg/JhyglKiFCM9dZOISjl33trH
RTx4asBtb8m5nBseVcINW51gP6dEcVJZvKQFTQXlx0jsm67UU8+WgQNtVwjoXYap
QzVlNy4NPrRDfU5u2uyqgZ/4mRpVnj8+7yVQbvesGFdGaSEiV+29fmybPcMNK5fN
yiEROIgACdMADT11Ebz4bvS5JbsRak1QvbG0PhSOSPX5mkwm7XEurKbSbFYTbi2o
hORVcQ7Lizss/mRQ0EDdQ3gUoRXxFdPxXeVinOv1Vczn+mtOu9zQhlJswVAE8RdO
3zb2uSYVQV35AQdaq3VfmSSJYOGRc38tTmmX/MxV00wEAmHVBnZ+YVJqgFvTjz/a
Mh/V5bbExkGKcnaOgzo33t0U0h3JjqSI3OFL2kpFhNT3qiF+EYhC1XR8aTFmy9ot
NPrQwcTsMtxuKCK72yWVrcnAaL9oGXFwGXMmBTG4GmDoCcgLZvsDcpcg+mI6O4HD
1jr7821D9DaPGnvjUdUVEVxHAEbbkbiztz+R5I+q/tfranUVtZhkdU50/Ehw2Nx0
8MLERPPtADwitnSEA+stgeSWF4ce6MFULTQe5cRWOHD1J8Ri9+f4jr6JHPNkyMKo
pvuINMo+6ORtF/C4WJdT1d5o9k7VFDzvoE4cJeVA7F06bHhV7o9c2zrtMrvw4yGn
XplAsAS71CvSOUf+K8crrMtAd3dHQQVtfLUIdrWnjnUGj+/uhVQtiGDhD9wvP9w1
xuvIui7iLdqvC0taOyWul2LpVPoOu7LJA2+HwWgcbvZdYZ0kwuYQlmBLRFxeUVyc
se9y2pF3XCLK8JJjoJtP4435vu41DlHpggcBgtD8L6FtBDTso/RVT8EqjwULbuXm
QE72QYu22or+NNVVGnfyNPs/YkRn8Ol4hbKG5gyeUw+i32O989Ns9fRIYX32ozQ0
nK2eWhCxOtbTaMDyCEHk3GmS+OvzDfMfXAckNzZs++Ah+faUJLYtVCyiWpajU5WM
x5boxgXnhOBnEK/1HndwmodUE3M+2IW3pLvAx8PmqEpO2gx0qL+eYRDrLgaZifSw
l7rC/bEFCCXHpZFa5VPBJLJckgoi2EVLwHzC+QVntSxLKsqnILdW6ZzZgRPWaPui
Yx3O8YYzbqjgL1GTMxXStrkAQnUuwnHKQiqlW1oDeG7kALsaqehv0YR/+w0n44aa
3uAXtc6N578DhL4/ACob4BKlkNM9VF+u5D9anodQ4HzNXp0Z1mVWujNFznevaJ8f
/GESciJEZTQ6haBfebtVNishJAIQ2duOiq2sruQOg3gHfbaCh9F+ODcFljOScwcW
BBMuGcM2bSfVIXKQ5O0tVurVfjWaaM1G/IsSqo8uzdNVMNf1eHhbMbOMGbUNvoHD
Z91OGhy9TWguv5dN1hVyg2aXoBrZxucs0lW+M1RadEOni8QZJpCBGcHebvLtqKNg
mYxyosep649QkCRDa5k7W6t7zyc5TJO767qKoXAQ0G6tT4+7qXk0hQRJ/8OpXtkK
L0JNAHblQiCsrhXeOZlzOFgb2NHCv89CktC2uPJa2hvPntFLySfMyJKYsH4iJP8J
kEjLu6FVD2zQwMxYydtinpM/bIIFxP3rpYdfIKAsVbb1eIIKL0PcDt4Qns9G+JhX
ZsaKYpjAP3DMw4XXqVGGU4EboiRaSixV91kJltdlVOyDUvlPM22CtIp4mVArjxPp
A5x6b+MjB5GucmSSJ9M2RuW/gTKDuZwe6Lz9Ug7xDm+kQG8+2cE/BYmllvYpLnGT
4axj6YrIDuJKhsqe/cZxgZgE435aFxGxmFkbZqOyrTJ1EEneeBoza+vJrD2BHadI
f4Fc4fjJl9lpscM1Rag3NPhQa1qjm8HSy1ie7OANWF9a16jb7zbHCBAnuOam282K
5Mzs3jki9riikdkjGMS+oVZDUCPjfVJ1Vc1nAThiYw2mqwFLNFV6Al652MXtLCFZ
GPtUCm8NRbfv4FvfsUT4UDWQjW+lrKCoB2jiJsNujjIfmibeA5NjuF4mu6yNuhFS
K8Kr5eMXeLNznVDyy+TNwJd1e3qm12z/SqmZ6ZnDumsXMXJ0y3YkYrgepKuW1xjS
2Z7rxo3+D2AbvOsCMGjE3Mb6w+hXQVTjqK20ChTkIXS45RvlYT4IP9i5VRyae834
FLxAOO3M+OrhPTLqZ3cfvU6lasRM2nEsQw+Qj+jIUFJDiYSTBz1AVwu3uTPzJKoL
0tAGtml0LgYg6lHfFhkJnetPtCXgE5ltQQV9TNs02vnIFKfWEQJtPDfsBGNzPvR1
1EscKNDg875p48Mc/+Tx5mJov/jB4v+reiI8ciBvm0xhn8wYuDSrUY30E+cEwPDJ
/CFGCgOFj98BV0/2lS295IVc7idAuZ3GSUfQZRHWss6pw/p8DlWjb0BVERsi2Xa7
IX0/sgIfbyQ5VXo8UsvjP8Tjgvi72k9AY8G9A2SdmL3uS/am5n1H5jgo6476Ey5D
IrTbcIIQIuIgILzVnUvZEBdu2rjvlg71M9+MxkiOIHdBKoEF5rNaaR5uZczQTLlr
c4x3rFn5ttvstccspZwWYHSTzkRtN2xslROznAr/joc4j8DMOTZA+4P16K6Qus1/
1R9KGjRdlBcTU4AmbEchmq0zdhT/UntGRGMdolHXuT0HsmlFlEiiM0zXMKsfv3SB
7EqxMylCPSGHa7PCLwcQzr1Hb9uayh/ydMPUZA0EM1ol/dypQNZIKQ0Yyt8aALw9
k+n5xx6KCZnEHOBB/N+xOz8QZvAGjnrJl5s+mHL7Xibul1MdWfVN2rnHbVFnED4Q
C98ohFBdNLvopyuCgKjvMl0tcFW16id168BhAbQjEY7YNCGCXpoxod10GZFFf5LA
w8SGiQA8XJ4GwYkrFExHmGeme7umKlN/Utp2SNvbzY+RTWKla3iuM6KxaICmElfW
vGr/079f3HbUaThvziGwfKxH+nTDY0Y3i07fvpwgU6HNHAQR8d+yZcmHxZkqUds+
+3IHbN9aCKT+zOL8q1hSRCg2GLDOWwnl4GnbnZU8vQwjd3xHdOhzlQufdzCZnkFc
/bJ5Oh4sPKe+thrdryGc3oKV3/QYaLCAnU/7ZsMmqCU42BWnn6HOh0rVWc04Xrnb
qOtzkCPs6Jp253w8b2+q8/MSa7hbkuUH4VoQ+xz55AasunmW23ERxihu8iBTStye
lM0KANWJ/iRaPFvETglY6EL0vvq1kV4F7LORrz5ddjxLGc/djTk7rwO8ceKjlsV4
9wSHQ9quGJ0c7wAcD+HynQHt111/O6/XHzhG59BIyF/Dl3ruUGJZXCp/nEbxXeIb
SMcYaOc7uJvMGZI9Dmr7W2jb1uv7aqj/SqVM8hGA6Kgz5kJuMCx7bSXWbUSTFgA/
iRxRnmibCmWx/NmW0u7Q8G+fcD8vHBRtBT1Su+E+gLiy6dGlXQw90ZPX9aEBLQOk
gF16p58NrGJ+XM9q1OwXXBgeiPvVEnpz4S0AA/V03zpvRymFCHa9pnUZroQH/FBo
BmkzlpP5CQ3DuxLfGIT4OAG7Ok5yR7+FMdj7+zC6k16X+6dzfgBjmZIlNRyVXpDS
T3AY0wgweYCQhSl51plg259K6jX6Bvw35YKdA1hnrp44lRWla58RthpYL9CYQMly
uIgk3Z5Ophi9fQSqu5d3bfLlR5GEULDYdOg5aXU7cIb9pO5pe07ilT0JvlS4/qyn
HxUVUn4x3hE31eWcbhPEJrq7EWFI9CrbcWFftc0OcJnHoCPUiuiBrMH4BLyqJbD3
EHX3AwxmHwdgv3mwP6If7Ymlf9djZkZ6FpwqEFGLvkDFFxzB71dTy3nY/vV4y6EN
n15vlsRr6oqGhhHilr4QlvJIqB727arwlDlGF7ukXkJgECMfxHdY+YMe55jZuzD5
HrbKlLrCq2jbdS8svfNdiPB6rrnp3w0sVEO23fiYPgZVy/x/2y6bU8oxi/gnH+pu
SOfqoaBEoCL9/UESEJdRE6AMDxyU4WSuQqpu2YlYD1nni0bRXH+YJmd/k80v1ZT1
smxCgsC+GmavF5o5fTApILaV8NLnvZieJaIBj2bJ9KzZLO2Iw9xOqb9xyZO6KKUP
5qo4omaFk9pf8IU0BHuWtiHCslSl3BxLkfiwQoAsChQ0iZTp5QRrCxi1f/n9VU7y
N9SB/t7DLb7/7AtQPoh54pLexsOd9Gn2fhYKW37bVP4ZeyK5RYV8JJn8vybfnaf3
edO/ckJTjGuN5Gz2Js7vPbBbQgkh1ECpX87pkyfEawiBgKK+2eZpyH7Szayv7A6s
XvMxTf25mapWHJUnlL28AOt9WOgSRoBtlNsUYiS9E//BxD6oXEuxozBNTULVdz9Q
yDZ9kM7dUfrgsk8BfDquWr3f3ukZGMGCrHBSllvLWsB2aHD7Ics+FEXQQTzl7EF1
qQYFYsbUFAk4kttjQLrDqyOnvOyZUM3FjI7YX3ZUfdpz7iBniCnQROMth0Bwr6Ll
RC6hvJKW2OyNAMGotLRAhrV3uwUiN6ZQwoybizr9k5iIa8K0g7sFVsUi5HalheNN
687R7/FGYda3f9J++fhXuIsAUhAZp4Xs1XSolr8ju52SpugnqN/hE9Xv7fKq0i68
klw021rGsn607zoDb2E3gQ9g+dEJFiXP+ril+HjwFpLsC/EKRx7bDsTza5HH2vET
eDDqAv8JcXyDWE8aWoI2Rer7lWOueBSyVM8mIiVk1NHpeO/zYcMNenPsF4uUVjVf
DKB0BAALGeO0444pkek6QE5OSmb/M7oLHI1ZsGgSc89FqfCl/szDZN+qedX3Z9Gj
5prEx7ufmX2D9PV+vE0pdnVam3n3Uo+TCbjS0TyRAraqQ0vCB5tQeWfXYw7BA7dD
DVynZ50sjkCrOBmSVRqv3T77bpMKYVE6/aW1xtr1talak1dUQ+56HyXyMzIM2NgU
HldmKIGTU4vwZFOOLr0YLjPo7Kn/nTeFNj+nmtHolGVDxUrFIZJfBvUrF1IPbtM/
wiqMHHj/jKNaIvkSMWwdDiVj3fj8pkibQeVAgw+e/vXqPnbngXTy0qrSKAzUp4j2
/yYajNr6k/n1b0KjzhZb/m0AQKxbyMtl/QGN+JxKLl3LISuxgbWzKU6C/Vu6f9sL
DbbodC04ByYxh9F0ZC2bzM0CP/tuElA2FL3+8ZRvZSoQ2l9kXesvXiHtsxuxePQX
POda/qjWxqsoZYq2L4DK9B+TtnV0+HGjs8npEpOGS/SMDuijKQShOWF6qeN7znjw
h0BbzhwwOUj2P696Hq9VpUyd5aeU6OS3E40OGHXQQxMpQt4n6//nCOxJps832GML
VN6QdwVgrE/E8PMmNIn704tjB0qCIO21cDmpNXgBfmZTfYF9Qp8XacGG2GkVk6CH
+nNHOkUpampQ9QRlcN/awe4jjw8t429pKwKhVWNNO9D4d4UzrrdwKvgpiScOaf7y
iOVAIg3Zjcliu+m/Qeay4JaU/EI9RJeo/W3ZWUSZhqw70/1pvIJJAeGF+0SJKuvW
RvFmZFaxd/nUbytGWGPXrs7Xai1wJqMdHbVWOHFgAQYDAl+nOPZzDY/xA6lYr4jj
slKjFJuIVEO4tWvjDpNMlv+DcBwbNz1aVkl+8ZqwOn7EitnKignGt3FqGA+gSG/Y
c69lh+IFFPfyKJ0M0V5Lznt8TE6woCKvULyaMUhCuJ4wMlbbKiZUg2e2E+J+Rxgd
eD+Xq+pRFmLaXdczqr0u7lhBTVE/Wt4T9HjJlkJmMtjbL/Jd6anuBIOGr6TPFaFL
cPmEFMcN7re8MDHNmG63Yq4Fm8q5EslyshoClqR4FJENIy+6XLnhen8HiPbVvGIy
stzqDpUpOutPg0jfEdNxFNDh0U5HH7N/+is8jJIN8vDX3PeBvvxb7fCKehjBxla8
kboZDzK+pC9dZ5iLCmoU3Qcwtds+E3JNAJtgsbxr3UmapgzLt6EncbDjb+9kEEA/
AF6H721GZgUwuqTIOjT467bKv9QajoihW9/B6/jReoouUcF3DXB5D8lL2dubnehf
xBg0M789bzFej7lm5pN4ty/ZnoIPj1wUG01XgzuDF7BtRGmwGrpO/7ISWTrdqpSW
XjZ4Dyymfg4U3L60ZrSJ1SJLnDP//3c+lhIs9/86IEAuZWm6+hCTDZcfRmFWISxP
NXedk7J0ziI+vCBvgCyWYbLyzu+QkSriakLnBrlO36B9JbJK7vuMwP6Nwq4yBxo9
pz6HYreaDT4VOSR2Ryj7+UgTJhR9VypP0KDu8vc7+701LMmh0Oeao3TKvQPzaX2n
e6Q2vN6+fDEXcdJOthR37mdo132JAGDwB3Pu2dKCUwcU4lXhsXqm5eJJTwZQ6Y+D
jCDDGuCBH+b9ThdwFNQ+7XDdFxgvb4s/E6aODGoEoF3VrlNUVme+RzdKsoVJt6sR
AfTyWJmtGx3IuXYs1Baz8Qtl+wtW9aQBh8d58/B/J8J+ci850jXfk68nvdGS75aZ
KUNxngr5I1eXjMojxaAsvdlgM16LbAEAGodRKoU4+CU8SlqBCV8Ff0PGvduApyUH
SV7us8EoV9g4LQWcZzE+JFfbNyvlnJEBrGxBJrdCpswoHulpdUnzT5CIQGCIIYCV
6LyGOQdxUgqKC1AGq5Asw6N0iyRIqwYytYSQwAbZYX+DQagi4sH1SDU2mRU6De1r
H/eZskZVl4m+Rk2++AuZChxZhZgk1BbY0wm3DKEHCtlS9Zpzfv5YWk9VTaNxeUJG
AtcLcrrQkJVN+J6aDRT7YjEhwMsZooj6r8lPKWlgqfWEspiZ60uv4lxGMdWVQO0D
lPGdvsgS2QkM8Y668sALbpSBmGegLaM2YrTbtQUVMHZaLNZ+TvdFcFeWvHnicCOU
w8Gi6b4/AvWIcDfP0SYOQUlagLN3PfAAJT+iWtiDp7sDRFy0hdFEsZfQM8PlTa50
laxi+ujGQ5q2D4jtNBMiLXBcegrVwAhb96WvId7Vc/MHDz6gx7/abXzsYwkBdKHZ
8Gi3QMKiBBsgdj4nHeB6zmX1gHWlSl17GxHS+OQ4a+3AfNzCbejk30d0OrEKU27x
+J02uXWFoPENK/36Q0h6nDN00V8MgA2XjeBwcvcCjyubKxEt9FY+dbuww+cqmslr
edBHuOMR08L/j7bblkMqxtv6WawnM38u7vRW8OUP0/AkRSEGrw8hPLt0dCCNxRMR
1IwTbM/m13lGAYHvzhBM+6WHpsrXV75PwU15R/sg9iyF9LPzhlUCFyN+Bxe9Hdhd
4oA32Z/Jl99a6G1k7ed3eQH+gSjxSeFqHHLIGGguBKuSYwMWNcc7WmqlRk+BJUBu
JOeoZptW35CvL3JsD25Q1Sg0iLN0dSmVcayO4OVy6D29fSN41UhRpeFTXQjMnUCW
+Dya0ASpBEWmuW3T+HhAgfAahQJp+H9XLCaXUCgGd2BSZqo7U9hYrLLU7Gkm/s1k
49yceJdYfOvvQmwQa8EqG9/r3XQN8SdDz2+Dy2296aOGrsVDlFBQlNzBSWekUZGt
98VKU1Ow5TT6LcQem+pFods5exDZ4dAcYcHSUSK51XaF6xIUpYYVC8JGsISv67GV
luvtNZMV7p3BTbbiFl5KBIJ0RzBbN6D0nbPP7mirgQLYRk4/L5ICFI2gil29bfui
vTRX0XkHjgdbPYWyJVc5C5+OZ1cWNq4EOJzb3gwS1cY9lIm+LRoguG9ef3NxTaY3
hiZgrqvmUhtXpoJY/aa5drtXJX6fDgbs8c1FB9onPDDjJmlZvCiPaYuPxAvxyNvm
+WqEuLI7Bwg9MqcfsUNGTAt7Ee8TfNIW+560J6RFGm/3LGRE9DA8GCCTW3VDRBoe
iQt9yHqcAht1mB+A37+aYyaH4sF4wlCvyjki03X5qV7ehY6uH0i2vDYjlvt5EbJ0
NaP4u76Bn9hwO2w6hmF4DiPGVkKPZaLMC1le7oyQ0VONoscbYKWlC7I4bVzxHV6O
Z5op7RD60Hl8XhX9qVEE43MfE83JlWpT5bNdpbXtrrKLgTtAiXgNrrL7VGa8bUIi
nPF9NXFlHRhIoywOa6U9tf6ywm7OOwvx0l/yM44S+ax40gM2rCE22gqYadCsGnI/
Y6QnRadRMbw6Y2uLfb0IGQxla2ey8WvWfdkIqH5RaknUuOjz9AaE9rKP8Okz4yLc
JAOqXn5TfOxOxZAG0p5BJplkD0gKHH4y8FGuefsGWzby/La0jYsNJHJvfVtmrQRA
32710IMZQv3CHfqF2svh3kDyWfmZls+s+f+IbWrkej9+vsiWWAT+PR5bsBZ2c+IH
fSgUFSjZDJvscvjSFNKOt1KmWIWwPTTU0dCV99rXxfmKKidao8Go7p5CfIriwELz
tk9hD9hq133qem6A1gPjPsmXE0luTHVdIbT7d9+N1S6yVBx5tnzDyDnXRWTUIosf
enDBAEPH9XNZwkdeR9sHe3itClN2bx1TAmxL0Zv9Ab4ipWNU763kmWA1KT0nVDWC
6rP+CfWnVgPewzXb93SvYt/AjCuG5YKbcpg556e0b6g/UgEPG8X+E1wMgVEQ983d
vhKBMcHJxsfOA+Zysm42lNl59N2Q1vRMvKiFgBt1crzjb6XfaMfcQXyag7Vlqm5m
D3upqhX9EImng5TDsfE5Btg7cOYpC/cmXzF40iPgRZBjQJx6WOhjho3bgFcxZp55
5MzB1iWvpxEfIRGA+NPhH/CDaSPGztWmPYX0TKDfAHAO1dqmibTkHzzYaaohJ1aQ
Ph33Zf2t8jQ2/gMrowtV5exEBjWzKsLw1hQWjpZmSSGKoWuW2WjunC0DTlI7zYDb
8/t/nUFvm+CZMVarKcD9s4xoVx+94BSIOKXyhYFcgwdyZynF6KzkNOTB0gu2JpNX
zRApLWpsMwC1+sF1R0rgYQVHmmVurzV7GFQKteqmMsAfBk4+0yedUxmDprSpA7Jy
lF0vMA8N1kdHGmC0fIw8/XXIzoQL3wbF8Hru7j20sPKmKpUVm1nqEZiPbgyfT6BW
o0xpJHkWLrB/T8rPo0kxSH/y9aHukaSjtWztl3/gPIdV08gcxv5mj24qfY2Zymz2
nyV4IGCWDK1UKo6+A6IAqh9r8U/OojIh3WrsrOPH3s/EkxG57ztt1SQf8cRtBzYC
eHoAML6aAmezamJmYzpIJMJ+haDdDjobX67V+XUdMdSPgJAqC5SViNVoBu8L4Zw6
AWpIeMxAchD1+G9vzwVTYGzjSmaoJfZNtk60B9ChcBpTn8Te31BYAm+NEqLcn3+l
rPDeLVgOWcZkm4b/qJXf3b4Opx8E2REhqZwmBA3hO2PnMW+tOsDKP+IPdZj2gX/t
Rr9S9o/TsDrCzA0WOjPqVf7+pam1EI308gTxa5sIL1Xm35QF7yqbOWcUC6c7pzl4
3Kj1N3BXU2t4/+qNQiP8uyvy/Rvpe0AbMmGOule7PfrvxTowqLzfJ+kIl2sA4wLs
KLf/1CZ6Y1cXjFk0iXoNcTS2de5cc8SL5qDsuHSYpZ971PurJh+ifGC8Vm0HcM8F
CIgni02PX3nNpLpAOEcesUIlw6esI1WNZXBJgYerIc59/X6OZJhI54wXJE6UQwsl
XUgEHbQmsBVWPPH+caFNaJfrgm1qhqOtYCkGD7X0+NQ8Gk/j4PfKGnF14WFWSR4J
U/lXzctNcm6e9OKzUtzErdOPZGhcrCXFHuwdt5S2S4HMFSDBbRIBHEYexIEYwuPY
QnK8Cc67kADqeMUi5EpBQ0lFyqfTc/1uE/iNeXcsqnIcgBJTuSFcVIm5vJ4wcWAC
E67J7bFXyJurHqb5cSRs8vwG9sevqgyKa9uRffN1TnBbEUEA96IOwAvKfcSHxvtn
CoLTd3XAHjEcFqfT5HalDcK1Ynj2wHfFkmqBTN+5cdmKgedW1QT6xFxFSrTXZb54
FalWtr8oju5F9zcr0t10fqGi00CtHrYC4m/bsKqDuaWKCOurUVZRfUw1IhADZg7r
rcyUdcsEGOe50X+qC50rC8fbMiJfPMzMpXi3xD24Q6C/lw726hxfsSk9q5JoWZcg
jQKAOsJseZxPxL4ypeLvQnqsfCkGe7/oW+s4fD5zewoAe5ZOSKBlrRKn0WgfrP+M
mcNwIsxINDbTA5wLthZpb2nHvzZt4OdrQoK+hI5uJf26hyUsw6Efy8L7fSEy2ek9
y9gltqbTUHFm3DeAAj2OWNeBQI3LCIa1TqqnxAEFbUiSvDWfmH2Kb4O0OPNVlaS+
Vsd1o8CAu5WOTYmb0a4Hz2kULwWS/AnYaeRXxxAqXCcZMrXIs7PvA8dL/V4fMJjP
AKbOPztWHUhFVRRyb3iqC81rwnCO//ggMyOhNzTskZAYBinQ32WQfVCImpUJlMBD
DZOQErzFf4wSKStPwj1NTIdGHj2vcNvxDBOLANldPYwnUyT3AUKoUlbbd3VMdYef
5avv4kiNmvl7zuMe7tKTuEjoaXJBMYeLVIZI8ZA3oZzlytaiwlrbxbhnxJ4yN+NX
03/x6mUCspA9VA8vGPDRckN1yA+wR1lPVV1K9Vg3OrrOhy8H45y3yg/s8NrHAPiR
LoiJVyatb+zii2f6CdsY8juhelGrZ9LR6ue+g8aKJ2Q9glM8xQT6hNwFJ39ahSkP
rOPAmf5BeJ2kUph0ONN+VzmNWGunY2KnnTKrMSyujCooU3i6G4qfyUpCcPHvlFgT
ncsrfrCTLLC7tjmj8+cIw1lsXwyARlkFZyVojaqnFdhAwE2TcgsrBpDzr50XSfH0
U6CNjFzUyX51gMiwlHFmkm3Q1ctaggTpPu+OsYno8Bb2EuWW1wnRc6QPfsT9F6K8
XkGrOHiErzuuAdqXMcwznjGhqf7gnE413gwF2RFChiSwixZSPpbXkZaoU3s2jt+B
mZ+MLaIhZ3cUcoIQa5Hnj1+8T0rCh9DNWhILNR/wfBeEVE+5f39pDJWIlv17GBO4
L/xKBHyDnXkV7+6XsX0nBjuRpLXma2OxhqyUhVfbWJ1xsPdUT4gW/TMEJ6oPj41J
0U5HzvcxpnU/djDxfTg/VpNEc9qOQsifeK6WDAOcQkuZ1fWYeIRR6ubQDDMQ3V8i
FvlbK/w1rL9eRB6Kb53TmoTTOqVFi+IIE43+aeS/bNqtkP3JASN/RjySHi/T7xZo
ld2WKxbSjJEgP9zk9MYm/0DxFIqzF3GwjeVjh+tBwAA4LUsHcm3r7cDnIEjc2D1b
3S2dxhTfzfJqHIfkl02RTGOZhkl8pnchqgRtYE6GkiCze0IMowIgTB/5wQDvV8ag
V8RXq+b+cTKjgAGzlXoeCRx/kWQUUcfdOfOLu3sZbHNUMaaAfDi3gEJRQ39mQc38
LfIiTU1Y2U7aX4sWfsJYZs47mXZgy+VSD4/5X9ShD+dGb4tXSh1eWC7N3XL/e46P
tbeIrU2xvphF1C2J5RXMnC7TVX0ubY2Xfji4AD+Y+CH0yIzZcP2hhLXE68bYLTvh
rgrF6VlDtZU6AWGZKybnT8ZhrSMSaprzaA2iTAw+fzG7S4BiXAnSJ6b4/K0BKASI
nBFFJoqzZRvzozEdpiGkrWGMo/y0FAWJYHNWZ8fypwLAgb0EpTvnRYP8KuG+Jy3U
SCWzsJabfD/vr54GfNxOBacilOSyAd6U2U6JDejJc+qXz9l+fZZnAxG6h/+NoWOj
IwpeFDLbFJ7Nxb7GcL5S/FgodTNbAK2IRV9IIUnkDnqDzmnfvPVKhqPM+s0dglS/
jmNJdj7XHOOhQJVbOO1DUaau+KYSZVE7YaZjbawG4cQf7uIs6nWERhHFEZwfETCB
QscJKJqZ3suWAsU19aDwj2Z+G19HGhXXzJsRByPxpghePBMrJRFESZ8z7BZ+2o8x
aDiyiUXfhT+5OnkRyVYayQBQKcfa+b78g0Hbt0JzncSgxS0z3KP5rsT3KzbAyp9K
vZUhLtGbnlFe3ehJ+kNqiwoIUR9MIzRhl4CIwxfo3C4idq4GLUqVQTuLriTB61GY
iuGkHornW9heFOmywDqzcMvMkIvvoelmR4xJQeAdVwgzpQMf8ea7VOaHftSYoXZQ
vp/oCIBG0BP4bLeBx5zrxbt9QlvjzaPNsOiHw99LjBKvYbZPgGsWJoavmBkv/xX2
QeJ9gux2IiSxOoSBqszipOuLEqrlg3W/HFDogVotAOMon/uXm8H5VjInxw80tC+7
RfBQENhAxesw2wfkCMMVOLrsvFaV2y2cnAKHgE3peZw+yEA6kjyD8UDQGdlcaffb
y4IsEFkIG4cKEiHwuG839dwW9YeP5foQecpgdptqhIkJbN70dY1GW+8SOWwD0suX
A6yNKTp6xzT0nXDfvFWueCJ+G+Qv+0FCt1uPRNuPVJGR6C6ZtyzEnRHKtPrYpK32
FdFWam5hkqre7lTKC2+40nhcYa6PRzRbOCqJKwSMqY/Hj+kiW+WFrcZqnVCkXfJz
9+7DuisGj+ntVFaOU/AKYhCIftiivARmZ3sTq0LTm7BY7UVtQsatkSxriABp99eX
c/cfzvx1uRWnOm0uZ7jS2BB/vdj37SrRzE3akZ5HTy9dL2fSu9bafJRjgDir4NQ6
1sXbmdTKDiRZW5GNqb40OKfGEGIO27Bv3Y4FAP926mAl1AS6B0I+OjGjNvkUj/xe
CII1QdV+8B8AEV4ZhJhlWYvUwtJ6awjhIu44NgxNiYyOOWIZ22jnskT0ZHI0m34g
obLWQAIFj2BhzdFdWa7wlBARG+g3CfUg/Li+IUjuUYhDOLE+Vl8Rfcnz0+8nU9cB
Lg2NyVr1aQwhhBM6j1g1Fu1iw3cUsOc3C1Le6iXg/sewzTbYqYcMPcS4TVDr9f+U
1Is9WWcW8so0NOF/9HR0NoYtjgrX/MNtZjo/RJ176qTmXzoyVJH8NKFb/ZLXrtVm
nnJhz0wJdBF+/Ra6rcdTRH5QTR9LJeSkRPGnml6o1frFCGa5wZa4bE3ETNZPHUGd
RaX+ZMxJvd3cRLRQtAONaPZBzWJ7IHg0YwOLKVG/rxYH8j716OEHka+LICt7Ayy8
XHH3FMCAOFWJtAt7XDaB/kIiMOv0a6ikQsKN58sUqev0cxJ7kIvejU3SCk1dEly6
Iah0XS63iO7fCM0I7sT5KA8nTaZT7nLSLgbOhX3p32fvmkRuP3TjIPBJ1OUM30zW
jBDWbMoHo1cU0Gkhruoohi3NBOwTLeWXVOTX/Ip8jS8rb7XxglAq5oSDoqoGY1nF
8IH/X5o+YChQb4sMcnm1Yrts+vHWpqarlumOIOHNcBvRawGiGNWQ9IErne+KCoVb
TrVVGbTOUaKOnp6M9ziLjnSeqBHzREA+BrZs0xB4NFh6/kcgfuvwA8DN1W8AXRAb
81hviM19F1CQPX/qnEjWoo1IN2WdU0AAEEqelrttttdDEQ+///bWztsNSl2ctv6d
cMuHCIF42w7U1uQ78n/Q3zjeG+JUPonpPC29DmQBFdRKDNnJaKNq6KDMfDX4jo5J
5WiJapFPvHSGSUGtKOMvfHFGw0AcFVkonmKsRfkFs57zps/GpW0mP2IRhWYRduDw
xVjkSY59bFJKX4ezhlupM0v2E6i24sJKm9x3Xdd+H9hSpHYawmSS/OF5wTObgJ2y
FJth6I6jQDR7csiFZwAjm8BsUygPAf1Tcm7JzS4orNIDnets8YkllEjKdKIKi8JW
x+5h95De0tdBlu8XSV5YmKs9K4DBKejU/DvhNHwSguSlFnHiHfVYXkD8Gc5TxsKZ
Gr7nXya+oW0mcn4MiTw36DyOgM3t/kyIpzJjK8pIPmQNjsDvG6eUrHaCwA/AzWOt
K/ex5nRZqAdmhQE3DO6sjURtzUm5yUGf0QecFWP6ceW0swse2uDFKAOfrWxBSeXr
H6A6wPG46908cla5phbkWhCCBRW5QZfkGfGIRCpsQW+fNajB0tLm3GgKZ3PvdGsO
OtR/aFNTY5p6TRLbHfn1kogFXOgoslwa7xFSx7zOj8/ih3LOpLrH7Mz1yxSQwDBe
oAd7rDdImc4Z3ogDc3JVpOMlUhtwqusL0L7zzKH4qEC5s+ixpNiHxBlDOiHrLi3F
gudp8K0TRyrJi9WrEg/jkLxJgUSYyoi/Uww6w3mukm/NAKwDo2nfCmW0yAK+uqhg
4Ehx3zjf4AR0GQ2g7ZKz3//HzE4hdXvEqWUJ/25IUAc7xUCsJv7OxwNf0fI7ifNF
uLHukw65c1I7eGkSdCbeODFqxa6OB4ppFuqEKO/IXcI7BQsQ1oPEWst6aytbm6Yj
w3NVkhFAV8KTOFyGq6jWgzlPsT5F5QCQlYj+xM0OEmOi1Q2HzNmiaA5HP5hXsZKD
QonCOMKCKzqUcXOlxN9UVCnJMIENZUZpBZFHAqRHdn+akyqkZBaYJ9P6kuAhoXqD
xBE1saLI9B5as8XKlOJcuyGiSgp/CwZQjH4R4hCwrupOYXf8Ixq49Kzs2ckboy9b
B16NGgc25iX4oP94hojlmp/og/ZdimCU6WTTHYk7HxpUTmBUnUz9d8LQB4Lo3Wh6
yS2EKTuS0JVvEATyv+JXUug0USYeAeo6Sw+wDQFxthgW8i3KnyLjjfb2K+3ZMW0H
t05xe+IUeGpCIipCRpxTfvempLf6huBUAVGNkeeMEaQssGHdFUamVryiLlBCB7HT
8PvSiUmbd7UnmME8pHTz8kkr9MmuyquQ1KB3ixtY3iU+Lo9gfef+C163Hyc2Kezm
1PTnfQUPxpAMixQLbFdnKKw+l046WxeI9jNDh8Ww6/7X98HkFm/wlHOuAq3ThPa9
PA7GJjczOSuvYwPh5x4vQdsKm+H4tmj8duF1vBmnIJfIMD2vPZYvhUoNBYtMVM+y
FZQs/tQ+MpZydtHXYzizjow+6yajtUaHcc4mdFRm3LI9ofr+zDI5jO1gW8K4bGGj
zbdZ/UIAh25QkBe/vI9i15Zc8HCwjM/bWeP408+CwOp1MXvyfCk3BZf3CMuCD0yR
TTd+Vk/cBAUCrg2MtiUy0f9TtWdAYbNCBp7/Pw2XyyLU/w0c6EotVM1YXibcp7Xz
scfkq4kJvBkpzJ6lGy2OTSZKvy5qmYi3Ysttaf6dN4/Kht5UBwfaQgKV2By/HLGE
wQR17DkFY5FioyGLJifUbLacuYNmHxp5U5XhzZW7xum41Oxy/5J2nGCW4S3TQXvl
8cCpY8MOcwRjOS/CKeBRzMB3JIt0kW8vazs0uR9lhfZhXuRlev20ESIj9Yqd4/bG
3AeBbgjDC9p+7Xme2i/Z0TezvzX/TT9Um5fGodloPJffOCYsyHXqaHiRJXQmZ6qh
QRsdzwYctGk6n/svZh0noMCbpvHdRiD2QbX7y8WkX7DIztRTlS/l5fMfGmb5RIHA
j8o6dUA4OHdo6N+T8c+1hNmPBfK3RTFNs2IRUClSq2DL8o6SYnIj74oTHbGc3x9o
/4FFBO5WJJRsUWHkfNF0tQrXOtZtZaN+SluzvRtAt/+9WanT3IsKumbJxtLFto/5
OsP9FVzMTdkVFqM/GJyLy06mqt2QthW9zGERf5ueVrystRoKvqBVDptUpYrWL8kI
nAQ6PURgSKy0tdeqhR01AXkIjSHD9G+ZvkKhKnJt03zxNSYdGRyUEgfPznHaZ8QE
gpCJI27oH26KGHxYxYH1GjCGhT+wfbWNXQV57wdWPQ0K3G59pPGvhpR1TENVQepn
7vIxpTeUwB+CrR0qDuUQ1tlJVHjrWti4sSlr7xQr52bdyii8apoIZqOuShJn5ySg
q97TjluzAVdGZXGPIBqmq3FoQjOVZjwUNcsBHhzsGb++9+RnAXSdK+L05xggl5yw
gFp4SzhhIwrnVbvHvknO6FP0pY897X6EWaPNaAJXewYFzF1nzYpOuBLewyRA1asH
yMZ8EHZN5J7x+hDgvYxD19eGypa99SY6zBol8ZsfGrOIXC4PCHiWU5ytOdt9bNQ2
Y58M5Y3XQksbNxp7jhR2nZirztDerTFKc3mGNkxMA6kxkya2BaRLT7LNjYg217aT
nN3i9bbbyExVW7s3kD4uwjoJzSVZVm68PZPzsXWiaiKPlXN7uFk9SCo3mEdDbG3k
ILsWcb4/WD6MUGBhDJ0bdZiycuqzXN3l3E8meo2/HSvRDhvF+pdSc7lh9HhZG3gn
wKCFMxDMDEmdD5S78YnT/+DXxAfnSOhxj26FxT4Sie/WKVFTPKr3NAf9pS3/KJOK
BxR5fqU6txOoIVHXEVlz7NHBWcSXPoav8xE152mquFvdaKK3NvYQv1MOsdv3o0h9
zZV8BBBCBAU8oO25kJGLOnPk6a0I1GESGrBTbRVsv1Dwo3L+Dle2aJCAhksj7zdv
NSpxV+ZJgTCwgMb05oyYuPczT6V5f23eyZHyHOy90SkcoApwf0NSoi5tKpRWyR8N
zEwoeJN/nQPdWoZNOfOHDi969nfwyX0XyTfMpBeZkRyS8vAiqYNK53PHAioyO2a1
ZSNu5vQucLo2PAPgXugtdvaCKpOTaJtTsUiZ6iHEKZEPZ5gfOC0rR5AmLqda2uNG
LN1XHLbWn/DBliv3Mm/pevv4dCL92fHcDLTAvZHqzHqo59FgIz6G9dIC9kST2mg0
9VVAzUFW2bBWRn7hgKiUBqt1h89Md9sl5yenBFaEE1+c5MnKa+oryj9HIkgSR2fK
Iv6WWQBJ00DrV/CJ8xmUsA==
`pragma protect end_protected
