`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lDVJAMyaDgZ8hZ/kHDXOg2zDVLHiUR2lZtp5d2HXnODlkk7eHFpV2ilx/ORjrl0r
LpQvgg6xqK43eDLSvL3Fa9Wlk3GW4VkHWUp50MiLBDVc1chSWj6ioGxT7Pv/+B8c
R8LbWxqawHuP5L3J6fYk50DPR/3V410oukfDp3R9ehY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22368)
s/Fv2hYNb8wltMbNhq0Dn6TKq1CkmQfFTk8InQKybyuYXTfmVvzozVI/1sXYBVvD
0138/u2AP4vc5zvDWXLbSPc7CgG0BD+ppQ/QqPIIkmLgsexJpkom8skjxHKuo1aW
/RDHY9sB1RNnJKn6sPIuk8TCP4NV0a4Up5x4a7WHatiUMFrk5klCvOXYkvWsKhRL
1QFPIfSsl7+qHwb7161NOEgE7bN17VMLxuBZWEcI8ROte72+5J17pNki+ZjkE+iZ
4UVzolKRfUa1EmWyPItj4JGslp7KGUKNBKEf+eZG4+jYO20cPwruG/GJ7H59lqK/
XlHX1AKvwniExlWfqvN/5hj4ka/STsN8Mh+HTpEey75NYjChiEg25QKZgKdFLMxU
+L74G1FNDRWnvx2dzsLPSJbZwEGi2Xg9hWxMH09YYavtw9zVN2B4DZeeL4O+pc+N
nYZNCeAmBtI6SbR2DspfsLUYX9e76RUu2+HD0YeFOGjHBN3j0a+A8LYt0w2w4FO/
5nNSTg9vgNOx0rEWzEUyE0jUBTnu4CuM9bFD0RDjUEJAs1CI9+lK8T5XSH37JDe8
ZEegQo022uGvXj+aAp8PR+JLbHGuofsNvMR47ogm/w2rRUrdBeC3ZTF35oeDYugR
WxDZDvpidvHGZ4GX6uRdmAetbfzgMPaNAZe7+Nx38nuMGMkV5TIjlzGNRayRYh8N
MJ63K36Fz3bHZY3DL+ktAWVbDqvhTgmfLRCtoalurW+R//kn9c2oogaBZ9MA0fyP
2cGXf8BKfukr1zmw8kfX43YQ+GnoLeIGjZYCcz7Cv/uJ7zLnVihVl5bnnYIi82uH
5yapflHFFyAYWzJXxsFVrBqV1WfHWf1u1ydx34hHMC7GFpWknrQ2AzNHoq5ZmEiq
U6PlrSUDsiriAh6xsfgisKVfgE6PRfZpEUggif4E7Vxz3Y2uqOduY5OEihFMo7fq
DwW97Zuv3/EwNupLIZbP+PNOICb/SGOc2I7yZAh2diEH5qvuSdFj315WoO+s+GGQ
eKaNvRAmW8AXd9zqHVJpS9Me7spjYH+PsOXCo9o+RZ27yHC/mJNeIoYnfIRMB/zj
+7ip5LeymdFGr+cChl3P6YQDehTqZJqrTzGNKstdsAJoJIYqx2kIwIurfEiYon6S
ZvBrkusfUB1qD1z6sX2w4N0dig1HVXq/QhYhUgznC35onIOjkmueK6LtDdN2uxtJ
h/uEU3nMdkx3nQ7icOvCTW6wkqogQE6+QQkJZgQehV3y5IcqdbI9TQhL94wytuDt
rPCuCxBu9OOJrabwaw+eYiDaZctNK4H5oMH/wOaiQLTvhBjnj2tG4od298G1Haib
sOVMDNxGZfDx9LFQvmx0kCJR6tZQgXrhJBcrmSgox81YAPnpd0ANymGLfjR/+Ehe
/zo8fCuM1qkBpUNtRlv3fHEkG6c3XrGclbh2uUV4j1KVWQCho7Vhv71jZWf3G8bW
Zny++1IvImTJItqOSTc4zvTo4q7X23SXDBf9Gqw0msWpmctWbq7zLQtbF0gPXPf/
vdCOzw1NlT5JaVXvuqc6ew7NxsOR6Tob+F2KhWrDB0R/I47Lvm5E3ix+Edrm8kx1
Dr5fVrrPTCCsapul0GT+BzDHOMdOhfITMwgzzH82FvcFR861Pveh1YFWBT89lBk0
yB4WryrmMTdjPzaocmKk0hWExH0ffK4EzeeDAV7VlpQ6U+4zPPS2c/0simmCUT/+
3Lr3xRKURPSKotcaBWwHHX4c4t3YoCok5f4FfnEYx6MUaxKcLNnTRT31qAzKPe0V
g5WZbZOzKgp80/JLbc8AVbMZf59r8TgDlBXpuIyZh/sCIrLgLbTfdMrgLKCAPJWp
XryEGQdGQii4/UOgcrXDqzQxxGQF5bmhtj0Ri87dXGa9NQrTYOUxdtOjYo27apjQ
Db9Ld/qc8yKmMIQtRb3f3tAyfsGL5zPogoikLxxw+shtuGbkYcJX/QWisnt5dm4P
ifxWES1h3ZL2sEdXEj39MenC6LlQt4Bhm1hD3DNnrNWyUf0Sla8nIimsoYRnPUDK
54F7pPPaKZ40QdSBRb3QgAMOE6YujvR1/w5M8vId0f7ryav249vZPBplkvk8p7LZ
JQYLd3gZbt3LFAIy0JJVoM3yYobJQvCLsAEDxoExILZDNVP88Cjpl5sg4q9pQ+9H
pDzWCtJ5C8rclLbgfC8nVC9THEgcF7jynHPW17GjHiRJDzw43jGzQ2ctfPUdy7b3
ffczAgHtHbPiHgIgzbt8N3zfytjsW7WLd/g35KSlZbR8djaXo8V9OJT+MJ+m7FQS
RRZVWmTshjkZrB7/yhSpU6W9jLvgpnhpSz0QBQNK/jqzp56YEQGH2CxB+AM+n3sS
q2uaonHXe7/0GNXmGwrASuzyDSWY5Ih+0i6KY+2SO1Fi4nn+eXcNcJumNiWPbqG9
0nwIZCCIr+GWUgpbDyZzjXox74x3se5MbbXgbKXqii1etrT6coeu7SBEdeC+R8ku
iHEN7znbJ+TaovvhkDpSkJw2VQCQUNUrKeHNYVP7Ee8aFEoxtergAtCwVfpbD57L
VjL5LfPTQCAxTr+likD/xppKjNFosSp/hCVF4hVFoL1zt4tY53FuyOziEmp7Mu1N
xmyq97yD4+icEKioj/9ACGKCi9aNyDFl1H0NYh/CYcKrSoKjClToS9Qk33Sc8Ydf
xHU800hYD9cW0wmbOi5lMtEoIK4RunIdZMhP7I4l63Ks2rnsdJXFPc2wSPASmxQW
sLPuaD6pYjce6zMtA22Mn0V9y/uXTo+zGJiboQCYIbfzgHOCcf7VQgLZvojsIi39
Q9kKuqjI3FD5VhHTytItVkpVXKpAJMpdu2EwQjBRHVfM8tktwrM6njkJ4WMtLKgE
R1UHDHmqQKqu7E9DZGAIz+PnW2TIkzCD9FF3YTYHyneRjJrrHmuphMieYhBagc/I
cpS/h7E9WuiItVwn2rSgfARpHlyaFG+2snCe+h3SQz9HiND4myxmyLm/PkIVAGJp
vecsf+k9KwBeLycWzDfB7pVqv7aqCOj1NfgHPB3tiQi3e8zAXMjahPiTHhwXEjvJ
BiE3DCmcbPNFUglhpkampBL4jIVe9fnzM833v99q2Vffseu8lfEj+2gVVTC1arvT
BuDemK5JKYj5425sr1hd9cEnB4l8ulWSENF8a8pOZ4ijLzA0EIKkgiZ322fSaaVv
Kspl0djaY1MRstU0QQ5ncnCm18dqlFnMdrMLn9WQGDbUlA1zSvuM7QJLXD/gtEOB
XzR3qgpPUnCcww8sbrNZ/9JamIcSKwx8kRX5g20mqbkVb0qGQZBYnTnM5bdS8crT
j7LP2E7byhlyBaz7t+gX1cR6ZWuuN0pGaObptzHS/0znM8vAK85Zdz54BqHWxHaQ
6NU6fJNuq21MIy10Uh3nof+34uK10KUaKo4VKU5hbk5AXn49nT2QNtNe1JehPgUB
HvnuNzj/oncP25j7+acQsIq7gKSYBTT/tzvjy8aXpcp/sVR4ZvH214cp7I0RaAoX
egObAp7T1E+DzUb/xxFbFRvpPWXqNkGf7ITa4PKu7dsH4WcgjkmPfWJpyMvvYt5J
SAfVhTpZ91wmd9iq+T1LOsqT8rHDTEmFZm5K52K3SOIAvq2p/e/e21N4NsD7vnxA
zSqXhT+z4bJbNT1qnpNBxT/CneYRMydUUT3IofMp84/7AlNnyQlx65hlIUjisQxi
9SPlPXuOS3emQuXeVgCS6OFY1ASse7OdkOJInF5Hmf6+OHs7Rn5PI5b+uSM6vIOe
pLJVJ77V+3RLIJ8uHJ6GdChrwDYSMzqCdSpBQ3qEjAwP6/Ki2sn3f4ondjLdvBCF
6XRiLWFWye83VhVy7yyLF3uQM7mr00LraePgx7DluE7Ww1T9pRLjHfgyPFUPI8D/
U9SF6CGQlQOUljMkNW6p51mII1DbmvG47wuBizLNxizTXvHkKXCQnLzExBHIAiiv
Ql4H4zyPI9d4hcowwrgLKDgZKPtXdU2wjk9kYUl+hy6fA99gwDCei3x1TRIEuJcF
+6mh6iNqpTBLBzjbnHS9pxniPaTQAj797/w+wiHVdPo6hQqfmN3CECydWbkivYNl
9MiDhSlxwWw12uk41SwGKd7a6TmwLy9XYF51mtwG53iYO36enJ1oh8ptlAeFULYT
VNtHggYD/NOuG5kxjFaGmDbrX97KGAIl3iHXcBSf10g0byrf28+aXZNiDpQ3tpyY
M57jvzyvYonoGibc79Folug/yyqNyhS9568QsSrVmL6qjLf2loeR38wWIQ7+D1mI
RAJV5wklpt7kesoxaBWlB9F/0KXSteNuTpgYt5/pAz1fhFmj5V0o2KSDnX0QnSYC
GT3Gjut30o59TSpcfZV+usl07DRczl09ndglkblFsJhHTznO9YQuRr11rfXOsBO7
ufrL0KW8JtrYXVN8S5i3q2H90UYHCtjxvx5sAFYxizvQxFL32sBQ7cz66OnQn3aA
cfzahm6a93Gk5FznqW9pC6tVpV9JqKaabUmtbAEBI4L8S34lMDA86K53MCKzcO6C
/5DX/o784twcH4sr/+c8gREcctGUP5rpBEBOPClSkaUSFYrL8cS89VLE+0eAmfrB
sDgIl1G9MOX3c05itxvSwosrmarQiHe3VRhTAeXUTlb/Kqbq8HBF6/nXLaKL/a1F
qlBLb5/w1M7HwXnAc5RRJHQ28OPSNsB9fC3yCPg/7qZGZmnpKyylkzzEGqaWVKtJ
uq61afydYnMbHCwY5M3lhd2z7ENWRUlP6dO7AoH3rxScj4ks4mdUhCdHRFx4LAan
GBJ55oSeCEQSwoa9OOugwDT53zWDwFDtRbjwqK2oH8vJi9dk3eKHQniugZvLtnBv
BxX/h5kZliqOV7M5p2rVh8WmyLA2w7XtiT0BxljKMXgN2ZUSC0y8w3WligJtQPqM
up8vCbTgGCYYnBOf90iEkB2OnIcmEuv0q2WyJNeeuboHR436CKYU5kiolkjxDEFR
wnr/f8iv99lv+NJHe4xy/ibvEpHsMrLjhjVsOYJPl+Q70eXqmOtb7vCzTKSOo4HC
ujN1m85xldOgRz4pKNRAy/1I/2JVIlgJn9cyNBpz+NOLEDwxElerWaL2ZzfPTuAB
lXoGH1MmmxvLX3MkSRpNZZh43cJSzWyyxz1dvsHdBpIY2KUctpPknXvvE4id+/YO
gh45eUWIqWu6QyWctsBJ/Zy3LK/xufn56d5IxBf8gjZeLxr/8MOXuDH+b19iXJUT
avqI/oSk7SWgutXXQY3MecJGtOotx8KVfMaC93lJKYKAoe2M62nYxKq1VSQ1zkNY
Gwj7Kg/fhr/eNGdZ62t3rXLblojags3f5lkDtxPnclp1icr3F4wtMuyq4FyEbMz3
NZ9lINP7+035tAKM0Rvxcueag2yaGM8R/U7g9wsbIwYIpLJrWS6G6oUjKaUIST5L
fSHAGzQQ+ggLS6+dqktNpw/0jTT05Usvyy6/LSFin4QERi00o0w9uYb3sOPAlJtC
6sQgKNNyU6t8y2f4ZsTjUS83izTJBxchfD4/+t9Vl5KWJa9PILcdPJ5h5fzL1QdD
oZg+zv3G0al7wzuCjC32B4eZ/X5tQzvkWD/7vMmZjLwKNSp7cPJE46cgEfI9O0cA
1lWpWoJhExBDPbUXG6jo7wp6E7ehG+T4NN3n7QVrs4oqcm0SVLu0PhnVHmNTq+lz
5eleTZeLvAj246Ct98d7cvvUCESTuh0vxYG+kTmDkmUXauxzg4fa2iOFxjvHrlYo
zaAMAP5HJZyPT95MFLfgnWzH26lOqeycUW21M5KW7ZkCuHOY7twjfyNxf6BeIsR3
SsBh5BcGoLxifEwCFwxcyzQA4SKL2dvqxiI1m0Nj0QBb4tJM6xk7OUNKg9TLOzjm
I8u2v+1FOgikrTq9Bwmepr9YpxoGU0vEaShnA8LT8zIGQ/NND9zwow/p5XtOp3Vq
Y3d0pc8pu7Dddrtyx6oPr2vlC1ENvJe22eHlS36uSVyg3DuiSlAeQcWahyxbC/FJ
LR9tPLWwc7FRw9JEpf+a3erllU4KTR945XcCORKGfeaGDF6mBVt/AS1USbLlTqUt
jyZ2uWBhiZ1DAKbr2ZH3SFmoDJYmJ2jeE6kMhYseEzeYV1Xi82JxEqbPagz2BImk
vHkATtfQ3WRw2T7X+oKT76DwNJS2sHgimTVTyHBwnmiKOURHyaQkieS987gY11ZV
/RsAYUxT/bJ1hXXncCv0XD0E6crIWiaIIeGPc6ooMy6qJAvntEJ6axYuVtyAjZQ7
GZPBnhQk0TTOFYvPbXYe9IT2J0i+eFsNrApFEfneraZvIbAzdlYXLZK1HI6dqYC7
Y8ZXiYDEQxReoJ0ZQt9vy0FNFQkSe+ZNCfoC6niURFBDtw1lV4gGPLEmKt51hll1
CEjBL1rbYefuBZoyKzqSRO2VUN5fiLOGk1qSGEe/277VnOCmIpxlZc9WzWigVOpJ
U2O2MgvgZKzSUtFns/um+vq4FU+moL2LuaMTNQu+ZFYDABNs/rxMCztv2WICuryO
g+xgrs5BjV3bDCvSIPszR50bp9NptCwpCwYYJbnb/beBZRR4+f3pUxAt9/FcGU7u
vJHBFRu4DPSTN+TAY2k6U5eh+2Xxpr9+oziymqn2NT/AZW31GyFm02q5NKzUHc9C
uuTXArcGP9hWTjlzk5EMiBdRF7oU+LmIZZDITgWU6/ircrCs/pr6rpwEvnlLjF12
JLd/anUmxUwG4O11xq9KPUjGbRnoItIRYiTuhZGZJBJXKgVQ6bOwUqHGzTSiQlRj
S/ngsdTEVolRuSxSIa4goYUT0YB5F6LN4Oj0xXFWD1sq0Ln0en7aSk2+3w0ybDep
nhyFGf5GBN+jsZTOMLveNKqKMA/q1wZD1msIEkVLS3y5MyGEDFBAFo1jMbX/56rg
dwtOXAXW1KTb4sFrL9CKMGsa3bH5Knp7pQ6HeXYtyWgHu45kTZMRWDIPztL4C+Po
1aBwace4rM17ODzPKJ+9708xRSR7raLbO0x30jGNbBO7URa8rVwNpkydZN+xXfyf
paFrT/A39B9VAs/D375af2+W0gEvo6cOWcDlNYdObOZ7D/JbegJo59GrZgMrPs1y
Y/4WF681eXPaQioNpG1CmWaIQEAvCobWaCMQRevufCx/txKSU7YXN+3/N3wksoDc
cIUfyf0t5EC5rbWiVnLzf8sdB7kGcOob/9esJDcHqXx3AzxcI5RgGqTef/M0bg+w
1zn6W4iMf2ZviSiC15AqwOUWd6Z+6m7bvpZ3GkipbTeC4p5Ydlj42QdMAVNpXgJK
hP4hCL5Zrsu2HhdazKmdQTHBHNBZ9Q0cp+kFM54ZjNNiHItLVht4pXorVHCj+9Sr
WcgpmZlpQUc6MB+uS+DqH75/vTSKBBW+6W1IQhawmiFtsQTde1PbKN/EktuxuX3e
jJDM1citoD8CLYzQ3IRtyvj83kxZyIWcFQPxl0iUwlFSmw+UaM0HFR/kFl/IXzNj
6vUOowHuwT0YmYq6TBJMGLRcyzQIcVgWKh9ZUUTNbogTX0xoPGv5Lu7zPgxu1mGQ
gjXFeJMqfRqVL8MhjcTtvgfXs7eiv8ImRhNu3B0rhsh+xNhRwdAoH88pOb1cpgzh
LaoEcmst4uFCXnXdHGokjKfZZKlJpg4Tswqb/JoY2711LlCdo+R8EdlK/bYb3uEX
2zUWb/dSeafk2ZXvqOgI8iifH8uhhh4Xlq+3r9vTh4mSrFnDeVybcDmQXKDaHNDT
j/GUAWQSrNu+Y58Z7bju8ITJD3Rrt1kUja3C96BWO7Vl3FHWgFNPZEojoKiWEQ9q
6n/kfAIijYumo0rSpcKZIk9XcXJ1fzdeI4QwyIt+Eg/1qvoARuF9LBhx7TvnklfI
HOE3gsORsiwelGMG9Cfklk0aQ0DY0AM2KJVar1B6XhB3sLmZZC46U7LjSMEAP04h
6xjAdWjlG0O7RUOhROCHKSzJOqyo+OgIGzBPMa97B6+iMVbIMMjgJgg/Ab9ukAZk
lOW9RDhp8HeBS0IB76GAq+k8tvTD6H4Vgyx4HP/fR1+WuXtFne1Ag6pBq4Ir+ltH
v2kpXCYS8PoTaC6g14fijpG4BlyKbc9LMgo9Li/29uAOHSswm4Oai352JA/30SR/
BvtX3H2dRRtHbH1YnsKEFD9evc/1qN0t17WPNNsSLa9+FEWpoQQFz5wOKxdjXXxi
9uX5qZJbcuciqM18sfRFtM0ja3H0kG3gaNVtVovhbs/hWL+ICTv61kWwKSjQHV/t
gvn0uQgtCNFMTEjVGIxPj5si6ZhqaTvt29AduztSyRqaET4yHqAyWuhiHaEF8ZB6
Q526w+qfggMKVMOeU7j9qS1zfsOZQB6kZ0RJ2KHY8bA0x8rgzF6w3/NzNBFTj+ts
KUnpV+XT0xj5gepwfLGBs5h+GUTprGI2WGD87Gnd4pAAOUIAjRGJ0ebuTSDlMfLT
r8XUtbai+a/fQAgh0AOJke7Kual/YNGicsuR3LZGuKo+3//rjzrrWL2YphYqF7Fu
uqg1Ki3EU/LV3NcNBtS7JuCmQq4nwm8O0J8UrJrDL0meUtX+d7OCVLZaiII8tolO
/ePiKk6igNFTXzRKcV2YWpvpwNdMEagpabZkm7pRkJMFRyNvA02GV+BrLnwUwFzP
9UmZHOhGe5rN+RmnsOriz+zOvc9+V5TeeP+KGOZR6WhRXc3sa9YkH2rGhqqvtg5W
quSHakxlQVvQjy3X/kSGBf+82JOqISE95KqTAlC/VzNUqFked9WJFnO39RbnFaTB
ae4BDw8dELIWBuOUV5h+WJ/ixJfIBTGr52U52fYQeQ2Za+sA3kwLIC8LXQjD0tNx
m33z6EHy4rQlif2LWAnmD+q+PHL9NOiTnZ2ReiwqnjU2zaN37IB2KpcrrLuHfWBw
Ml3EnddBQJ1K1zsKtMgOScatQHSOxC3wuFdhGgy1iEP2njRBkBaKDUaqRcyWjENP
BZp9vrOPYlwi2VlCh50CUsqlzTBL7qFKK4jQijq2Ihtl9VYe6QVJCjvyT6tdJoqb
tH9/lNhPM+yQ4iFgQv5+3FN/JdlfMv2rDBScU2qBNucY+LdO3zs1W+hP+qLMRKE5
WqCjZBUe9oRKa7XfXXqcUEAUhRYF2NHori6QLn5kwz98QbPMpJSjQBbBZmlPWfG7
XZAUgo7fgsFuttXEJZfUbpPWd6ZPwjhGcpI9hrzeB37DyuDYQelPggBairO6PHTs
kG+cbVn/NxeSDToN042ZnfFXKgBbwZg3y0tHyyghuHpkNiY/LgghFx441GjsJU3b
IMUa9nAJbNorcX/grssxR8wGaqtGN8uRvSr7LVRWLzGuyqEk+ZG+Sc5MQqH0S/+0
u/y+f6twQ+ECJKUGyqDrPWpZmdAV79mHnlEza4lIqCvi/OPqbr+CJKOoBRTmt6kV
ZQZdH7WDU00cJuRGbjVb5eBG8lJvgWIm+HnGg9QYECjFN/CRd10Gx9EQWLjOA1HG
RKiygRPcOXW3vqtCfvJhJo3IDA73Rw3ueBNn0AyXashrG69Yr+SCJvkiKyeB7xoY
o2NELEGMLopJIWJ17+AGA+ItspT33k3dpl/IXn+/Kdyt19bLY586UKuVnS6e60jo
/z45un0fUKE0JijbpxS4cfQzU+ZObKPORGjxBd0SDN3JVhGA02T/N6oea2YlegVj
fLfC4ejzyH0sz1NwQN30vJAGvdBq8ArL0cjJC4Z5PsfQHvfpXr85BYX1VSs3HEfy
XvChzgxKLl/Qo1UwwPngLC4nK20TYlaI6nY8QBak02eLohIcDpqI+6PI/sfV9z2k
j+57RGZkbJxYlzqbWaRtkKJjFa6xEI4jf4UYK3ixiAdnxquKGaIf1yW4/wejCeYs
uaqTctPzOgmSq87b2ildZpI7NqLRbtNCyTS5KNNcDe8tKMD8YkCZc94Lyi4qpwBa
g9YTTWPTPDSSDizO8sIJyYK6oFJRCMuQ6wYIGmoBAKwwp/eLibv3UYZASLtBsaj6
w0HqDpKKZDiHZJWEeHp5KxvIYGE0s170U7beuctHGGZuI2N1tzVaC6aI9TT558yc
P2DaFNjAgVRkvfrlY6TetvoN+q2ZrZXgoFYGhVuEmUK6CWVoMWMVyc9IcT3kGESv
P/0P2xCOXPEw7pA0ZxQGhKW5cKL8KGuFqYyB06xKT6wlgiKgcCJgOJaz6RvBnlBg
oviBVC9INRwtqWx43TFh/9nZsOaT4FM0D/6T2KSTZagk47oiIi9MAW+gO1epM3c9
q48V3st9YVtmaCAo3LS4E5nU6o4yKsCVAf8I9BJ5t5zVVzl2DNs5y1HA4+EbYmom
NJoKb3ohaiuWhstRhcDPqGnZktPOPxxP+OV42YpBHrB+TgjOa1jaC2iCtDsU1O0l
doKDlz06nIHwDrm5BgqEcaUhSICIpjQSp2M0rd0xTRnVGOO7ym7X9Sg/p4L/L+ww
CM2dCrKwrfl2L/oNGy4DZWyr4d7Ar2LpDOzPMhCPnGRgLU3uc9Q70eVLfa8rmKEW
TALyHi9qE+Brqkrr4pMUqST9AawTt8yuTV/FZRjUk019Gc9RkgD5aWmMZcLdICNL
AdGFW85mtvfprwOAiHBaUfVyWPPnnPJdagXJfJpELwuE25HFDBfw9AZd5O+fytBc
3ZKQwh8bv8nMJp4As1LdavpzUC6Zr02G5N05MFBb7yOqZyCnD2hRDicpD7prP2tb
ey5VOfmQks8mI5fMsnkhEBVZcEZfn/99o/Rrt4pCssPguhSNULT3ZwUylzlGXynq
YsiGmry2pa8OQJA48hvJRk1Pl24YKho0ARzUmfYvsYFjwj/CGGpfQTYwJfJZwUXt
wuOC+Rtxi0IoBRhHxDbxWOfxdFDgFznPKUud3hAA2YNb18M0AWsC/bPgYh2o42tP
jHN5VsJApLmwZWdUzpqACBbon1bOy9H3zmwT1YQ4XQFgkyrK7XYbs8JlZCNaLMKM
Py8sMP6E0dlHU79qOOU6YYsif3mB2NCa5tJBzPhlrsYcwv1rJyhjnKZR1F0Jfjw3
h+2BkWEcZGWGM3xf0FpST2yXUZW5APaszG43rj15UfnQqpDSvnCD5jEHCO8a4Olw
StNRcJAyXY79guZwtgY/BMyBpq03QHNBbNF1XQWdvxL9Zy0lqnZz866pqJ/hf7jv
BdVn5fxhlNSAjIENzzsGvEmLu1Bd4Gg1XmJY6Pqasu8reABJNyTbi7ufoxufPWL5
W102sl6I4cJHjsCSla4uUBlfgVSj326NzNHKODrV/MIi5KL9jUJZqWPuBjLQf9GH
TtCX3jqnK6lFhlrEUUSjT84IWSB1MlK78Y6aH7UK7PTLPKAMGyR+qxQhotMuOkCz
MktpQHJNCaUUiC8n6lIRfnyn5FJ3SQ+nN3sIZT5S7dmmrzuQ1LcO9JCynRn4ts7V
6b7llVp8g/Wb+3/Qy0MXepwC8koMVtQ+740pUh9O7PIarP+Mr+5SXTwlhRQfoWOs
ZFVjKDSqsY1qnEna4iwTp/jTNQaUcbBk693bcYW7ghcEKFoix5MsbfqnboDhYsi+
5MY4O//NIvH9W+qfI6zEjjQ+Ek1MEuyIFxo+Gx5CuDLV5Pr8HIl4fOKniiFtGjgb
eN5ok/TbFyhbmrxvS461R/xvCQReITjCIqaP6hv0JKsgNTzSOCiTXd6Qslgt7n2i
0bBqeWjd/2TgLyKhglJNwOCAqVbtZr3HfT+/WLSeeMPym8GN/z5jFNoyz2bGoGXx
ABkzz6rMHyOkqTr8zpA05TsZ9jFJ5M1/VIKlgCwNbJmK7gSAs2H0iZ6Vo+7kxC2h
yJ73m5Bu+9iyle6+uKweD4DDqtDRM3Y0U4jAl0qCyfgrbYpx4147iVsWp+Z3bSEJ
LoC2/Jo8BSLF5wRQEjKqdReOvgk6R4ye2bcFiWhwIcAZudWQXmkmCRdWABJHXHLH
OOPEcuhkHEtdnEJ40gmdrBrOREJwfOTnLa9JwPL6SbIcuY3NQiGumt+yxcKTjPQW
eR/hAEB3GgAoVgsQ3jNN64VcxteYWLQ9LspqUv3vRJsTfKguORGljpJk8mpvYm6K
TtYExL2I1B+ArJuluGhv3bn2DqKPg2frfsFTMlpF67wbbgRglLYot0YpcIhtvXIa
38u2+yIfXpTEtXYB1NNRTepCiDWlg7GhYToU4g1+eAJH5jIeueFI9lBW2hDGgh3c
IhY750QXBD9Yt/uCERn2k6FO2fPjOiGOK0w8Zp1kurJN9qxu+6JOTyanMk1MUuoU
LyYR/8SFLi+OcehBjIPvopny25XcrLeVo4FSu0auQaJSZ3Z3cj4rZTQYrv6fy6V5
MHAR8qD+S4yNRi+pGstpx74/lERBKEg/tIfvBTHzxbVOPXTkoG2sMe9dCabNykam
a8GI+cu/dVbzPkHKEnyIQMgpY4m2Y5nb7s4FB5YtTQm9Fcl4wD6v1BwRJqrcyvu2
6Yk8HVDQXUsh6OiLIJ5HLsyb8BRx9L1d5y3suR7Wdcw5dNRNsKxfKvKfoE+pGif7
0goiwqcOdFdHRB9+dnRLgXWqeMlcTTR6YFyc3JjNzL+Bb9vTV27krhHq8uvzs4Pw
mNWpKUO+UR/fduIkyVurQdX8rVBU51LEVQw256K8LIP/cXKEIaaiZczyCprCWFEN
zJqiv1LauYaMp2ukSIrxSwcLG7rqkOTt25bireq1qyKMsgSvv46XLXbdV89CWXPY
sDQLSlrqJdAZVm/3pj6cMLANGNG0/TBkzF3xhjDd40NB6xyjtP36G37QwDDb1dqW
M+SCvTqHEzQ+4s5UniZtoGIEFk2F4lnEumDqyhOKZDC6gO1BtbDyAhqMRcVpNwCP
19BOrp/qfRwokZOxlQbLvutdOGinIaJhKERSLLrBhvelYIXL4jJXStVdKu2rA0tZ
GidNDRFEjgFDCz7cMrKDvzbBC/DTyHRKdBZYhjUZ0Sv4+9zRRpGWi8zu4wiNgRqr
fI19oFszYENwnqF5o79VFst+K5ZOdL9gDwG9cR4rQBWOSLpN6t0xU7MlxIk2Az8Y
nEwhUOGvUoZG0ZXLxpkBuxWHHZS6EWBW4SmnjcKM3SiXegwF9d1tFNm/ZLE87iuZ
vsZjGpSm+rMM5ibaL7RfOwjohJILTdpE5gybs1gQxHtDWgBJLUE1LJEQsb5XmLBn
XmQQIC986m7+qb8VgKNie7qAUoBE+W9PYL0Tn3m0RYnXSk/w0D37tQwxPStUfcBZ
H4yuxCaKZvG0ZGilRoDRpUyHnY0Iw7LYx30R1IjhuCwD9zTCkRxglaCtL6cKxptm
EknpIl2sQywOOoLFK0sMN8ckmgL2hEaG8aa9WejNO5uxIGGLLa9eTiGR+wxtLnjJ
T3jliOq5Ma2fUU3EYEiaUaUQwFvpgTZSUe4V8o34kTBh0IA+FQkx3o1mqtCchUQC
hlKi85c1Fcd/lGMjfglydeAAftU5tetVtGM9cGBcvfZWvYnMp76k6pOF8VM8DP7F
rI4difKWz4HCS8ZZiTtsdmI09MV+0KA3TLK0KtLB65SLr47QIMbAM3EKJEQTzXQt
qieYLiiC2kjbgoGTS9oqA9s0DnEuAnTj4Qqo7HAv9ceBh5/N8tt3BuaaSE+CWt4O
qrNO/XhY18D2A1KOFhYhXMD599TGJMlBNfcXbs5OdXMRo4zFom+Ysv3N5pNWiDx4
ymyN0262x7slfzCI8scD1RDu6UWCanbVKNhYsLX+iFh7xVWQjG2vmV6M+3iFYsMh
GFQLTuXheQ2SpdoU7LVIc8TSdoGDW4CGy2ooglrt38hYaHYcdJjlXW+W2jeSQovU
1Tu0SckGHzsFpoIurs7SvaySHofBCe0Nj/UpkrdaQxGcA+SR3sAoQeOzpLcKlonY
x4H0pXza6rI4X6GEEb5w3lD3DdLXb3O18hNIvzF6weWbq6l92h6k3ovSoq7aipKP
9uVU7b347ml4EpAHN8xWs4MPTkoToB4w3gY7uLj13hZuOhhRc1Ip5vFJCKH8oE4d
yNhrTxdksJ2PaK489v6/nC5CpOhZFVXkedCRed6gdAiQb+tKNJN+19VWfMmpjMfz
X8zPdGJPpLVAF4x674Djt+DUeE3I04RfUw0csUuzGQROO2FHo2dyfRhpX4hVVuj6
Aeutk4u2EOm0Sbs+rk/+4yglaAFKF37+/xFE2ZZOFh0P+H7XIN/VPrlbkDuvOCRB
E3bALQ6fiQyQWi1zIkL46tn2CWOAyyAbjja5pLx2rDe7VsOua9zOgGPTLr75l3uc
SH33rWLNkR00AV5yv8/rMpAZtb0X4tiHaosywQIry/aQjOl6WUV8AYkuRKxDGyVL
bVZvT6Lcl7dqRtscb+GCqaiRaoymZSz18nDiEkyDgy65FBw1SDXdVN9rxNEseIW0
hnmIvcHDXpIQESsQsnlGruuQIXX7w1eyWM5G9Ow0ig/L0aRotZ8nwz1j0tYTZ65S
mhVT42FnUiYAoA/oOI1RMs3vXZIDHF8mvwZP0KGeDm/9DLJiT6dgJ7+t3gCb95sL
Wmt2Gna2z15Eg/wPziiWIR+0a/+Rwajv3DTwfs3nk+a0eFqqdTQOJ0UOOZT/P+ww
N8fdy8T1oAJ4l4Cqlkc3yZt9PCT9YXoRCsqbaTTLHd1z4ZQe3vR3pHoMUWpa5cUJ
kLKKZAM5IBYwuKMP8YSiy3wF6XVyqmy0zJXej8SmPoSV7KC/uEH0U0bLzyjfmYA6
rClkXxYK3DA2k5wQi97ut9vw/+K/+zJQiKfGj6hj2JTuLtMncTJHDLWre7kwGxby
nienMvNQkwGaMm2r9X55Vw59dGWV2dRiN/H8OgW6Rw6AHN4I0YZDZmKR4mGbkImU
V1nuu8duC00G0jPYFeY6xzfKQl0thWyDfg/J5+v5x6vEV4vQyIPeN1voUOQCb6g1
/dp4IlJUKBe8FoUOhygn5cVoh4jQ0hTrQylLaJr/qs5m0umlOfm+g8Q6n2l3nhin
Y6d1x+YQxIalA19TUxNAIOaomXusHzP2uIl0vA8ZdVWYk0KNldZfxa/xnf8LfCEU
E/DkRGcnZpnf9mNy4OJuf2RpQELg65MDJ7uTjtwL5dDt3t61CLCbWW8Pbok00H+Z
E9d0k5nvazN6eZ+KazXxB/1NIs4vpa9moZ9eq5v0nllg0wltgBX6geiKEs7Eco6k
VBW7vJG29McC9/tLhXXLNUWvO2i9ZxL9ZFs8FbEoARQKkLcIz/nJNi87ld1SAbMm
DSNSYW/K+rLVkyaWX6VY6HgH79NmU2STMqL9VsLSG6ONsvOmPCDS+tX85T/MADSI
JZCaq/E6fCkei7kZO/zE1iv2C912n00G8wwh0PmliFRNTJ8dqu39qIzTvR2sOzVE
YgX2aULM5pL+sKrZd9AQlDMSKoBR7Hffcppvv1y6EbRaX4OuszACcTVC+vgmNjrG
HAhweUvUDlsKoFr7ypkiFnkONQ0pqZDVcgQD9U2XTxT5XFhHl/ogWvNfwu51JiEO
lvxp4q2rdyIHBKJ9o/Wi0TmiAnK2IDRHQoukkxUijWMoCLhKtpSQSM8SBdFLxYkD
DXJ0v+UBcFoqjA+4+pXzDaR5azCpQeiVmho7qbTxC60cVi7N5UV2AEgiIBv+Gkm0
WBckBoXXJALMxXDvLNPKNUyfqHuks+EMLNqh8BMc6szkUhvkFVI5vz245aLuLUNf
NS++3FhLx+ZQn2uoYK1jqTLp+So6E+S5haJ168D7uGV/zjEShuR/yGjHiWs0M18n
+ul33mfQi6LqB/x0dK10UcMpxl5BxNdfapFMA8Ys7IL0EAVco21IC1OPJaAiSI52
pka0YNR/UnJ14Y5Y4JMPcTOhdE2JR9ZEJdFubOb822VBsgL+sdIxMLWxCGuuWqk1
7w854rdNbaw5eO0SDiYftCm2lA2NWR/nO4/SopLJqlRFqxpXbbs8PXeH+nkmdE3f
8Cb3NFKbTRvcSq2TCS1YCUorHCOpMHFxG/+NDYQj4uTTdTfEuqqFa70puZtrNQ4o
eoQ6VFby9U5e1+0SGJXPxQ88joxt4usSSOADkgHFTAfrZP0xI/dO0qBji8HhSdZO
0XsaaofKo7ADYFAkG+XKMaV5rYwJ/LIiB854QvEeEMMANIlATQajjdVxGzSJBATk
NS3azmPXeZeGqYMt7JEOfT5mmg53qaD/5PWJEHn5CFVQ30E6iNd6qt0Tw4eaHAWh
BZEpcphMqAOcArTG2DvMvgLwje0FpOdmJ65jibtBQM2GYSmHrGUA7V1X/0kozT4I
GVqDe9l84I0FIoXanZnW/unldxIoGP4ZvHzhv6R58Upox4B3qkAOXYG5FiFuQ9/H
Ry5ptS4+39PxxCHTIcQWKAPeL1eRc2C/5Kyi8ZHrGeox+Iu2u5PqM4KygnI13j/I
Pcm457JfBFDlNxuoFRV4WStPfXubTTmgaZH+JwdqkewhD2scEUPJt1T369MqwpiI
mf3ZkU3UyN1cr5Hjnz9YFRlHOhcQv7hnB3Ycd+PhqHnxSf8Me4q9eA4CXKBLNrIz
KoqjjshHIwe9HV5lXXfsHjh/cpRLZCXq9Vs1OO0t6FxIaAh0sxLsufs6g47i7vFG
oeIL4hjaawxFhcULRKua+Dvsh624lbSlkWQAK//qqvbr43C8toMzZ8uwgvX7lwAC
pME79yX8X3nz8GTfM6DmkFBT/szxdMQDtRjoIpRhZkPiJe1ElndC/UoZ+ZTpaX75
i6A73Ic3fobJ/O5MhqEK7WnPsWTwambO5zehj86sXKRXjv/Ac+5pe0sioNy8UiJl
Chjoe5OR446xvaFj2r6OR+wQqYBsr00KI19GCw4cFBVoxxsSbg7mqMgD3HKYMkdH
5udI9Dnu2FiQIoupJ4T43yBApywi7GF+XGUEuCQX1Sch9VKVAnyJyBP37PtBrZD8
4WdXu5EYrrz/z+WvKUkT0LDInKJhdG4Fd99Z7deULTATUY0u0Zt9HBgaGxm4UTd6
kgNQGTctjiuPX3MyTCWLtnPm/6Q0B4Dj36TwiXo1giYmfC7HnldAuY6EdK1lgipt
Dh4UZTsx+UVb6AJJNPSfljlamWUl8wew+47joOqk6b7s8YUIdoohu6oLeRyWFOrr
YzK0Fd63Lw8uiJa0plUywNxUrJLdHv9LnMdbeQU0KZuzqq2UWcclhccp0PmrU2A+
itkiZwGhUTBdi4eFeW+QQvxUECK3N4ZlglINOqecgdKqYQOv3l3mXlpuw0T01HMx
pVSmHzZeKlwzld8FzKc2+CicVzQSxSdPoFSDgsyRjstOHeIChLA/sn2A44jnuRU/
NtRJt8wRk7C8KSEFu9wJxRfK7sjzo36KL81em44zk2FNbxWdzrEXzPN3czfv2ee+
LrL/e/jB5HQ7kdvv4QSyKiLrFmCPYaXtNEC56O06xw3jQn8opXsIAZG1w9juelj8
yJnJUYtnNvXsMZJ2PpStvIxhiBaxTx49YihHxqtY3KF+mjuuN+o84wSVkHKtctCj
HOPDXoBByIVNlHm16USJg/VbxLqVcdsT4+01mE48SqTgvNbXgJC5G8+swZdjaWhe
w6VmfS7BhiuJsXG+k0rEH5hQ9D1ivK4uLm3ybKgPIB/xxA2yPnb2zPBRMFisMHHV
/IWKZAqerMFjsAmUIn5X0ZXle5PwUIyXM7sfi2XIHYRDiDt8TCtKihovy9wMXKVe
Mid4hmLefo5iXNWZgh7lJrjm0xoIzEFRfgp6d2C7TMpwb37M9tF8Su7TwEe/SBCc
xq4r0NvL6ucP9zIfrItjWb/6ojr1pd3grGD3vpMfQ+BKqP6SdtKSJzbTiT5mITtU
9fQav3O/UvmxaPHKkdjGLXDRZzI+kNLAwxafXYrx1esYyQIaZ4tvfClA2RXO6M+W
EdPhi0lP4BD5z9vpB6jdOFer5hhBPrOyC5eCsNI8Kb1u53lTSlIoedQmJWGy+2nY
LM0TtV5lnzyeqhiD9Sw0pWOCuPqi5zpgbR7kaP3cpjNUOmp57WeAw3+i1Cm/A4kN
7py+WC+Ghcw4/U8g6Ve0WIVzeEFEG0fd1smYUPzf6URMVqm4394E0QndNoZMlYka
952FZZeFea1sIwyblS5HQBmJMsxb0OhQvIWVSV+F2Vflyjag9mobdCm6X3Se2FCP
wcUGr2IwhqvzC2NAaSbegW1P3Y5IvacoswGj0igPJAPNb+dPcgX1kjRP7IT0wG9j
W5iiUJrcG+xnxMQBnJzlKMmBE0xwnl9ALAeOHPgXpfDh7nAXbcEBsA2ZmaG2TvTo
lMZMmxZG3mSTU44xdpe0jc37hM+46nxlcTvj3ioqdTn6b05hK6n9PqnF+DNMv27h
JQtLZoGKlkNm++hz8bHwphLDUZQjcrN4ieE1Wreh3V8PWwavMKajouEtdsaCckKG
g9QzLG6At0RNm3TO0A7pOV3OxgYWgE/soSfjzMdR6CtUtxEa9g+bU8xTQtUfWCuL
VbVmYrDrMP/dP+efsHNpCOLp0FPfPiwMoNEbghlhSA4gsiDOGmL16iyeySKgsD+4
oHf7sleOSTdAuYtlZvHgtiSqS7WgWoZ4mQqCxGMN/d0RUqB0Hx7J2cyn4ezS9w5U
rTjy67orsl4/3S118u4VVbdU9nhc+ryt2CqFXs2FfugpHW40Ihn/e/0GKySeMF1t
aGnEoB4U4ih7NL9YxuTI4lO/LxGJKMGFn7+/4XCEfmpUyPMmcJaLynesOFzxVqqY
JsVubpoN8J1gjAwGGMV467qjMGSm8OfXMbCZS6UpxDvAOCAatD/F30SjTfCwK99N
8VnzDflGyVA9CCobtEl0N+NW7d3Ivqo0/51TU8WH3bpiWhrtkWiCO3Ggz/jTh6gs
d+sGGmSZ0ZPpzwLQO/E29ZxxCbkhfv3/4RF6OL0hxer6qAR8nQPSOk4VTiMl6P39
YyjrTMu0ofLVkiT+rPdMEgB1dnXsOH0xa9QnoBjCy5toZAYHFm4woaSwp2tsstM9
iQV9v+R5g80Itej/JBurLv7lq2oMdyrTZjnAUFNNsDR5v9KXTkE2QAst+fYpG497
/cQeImJwIk4RQ03dOPaO1r9K2U1r+06dGq8fZYkwNGW7xvNU3x7JnQuqDppkA+fR
tzFo5s+zAGLuXtqvoh4NZxhYXQkjNEGrb4tVQ87wEHM/O4+u2KhemGEgiD2h6J9L
y4N5JgLpRFhy8FQoFvlpsDPekQwr+HXbYXwZS7ISCXsd28M1A768asgM0/S7f0RA
wuJLzyFshBJ0ebNatGTNwsujXGsXjmQEIctLcKMOpMr0H/iNt70adJn8nvKo7UOW
KtrxPJ7vGWnRO/IQ58Jf0ZI30hnUZtgMFjLPtfwTMd5SS8Dr3pF+h8xw4q3oJYxf
/y0wNcx10cObjZQHQKr+mdwnk/cFRe7JyA2ap0YFSeEz2ccoFjwymYunaIDfD7qj
ZfQo8dOOQS0vIm/sA4mNR/BGIMvRrL1zhs7TE7NhV50OmPhUYT5pcvVjDf2d6luf
p5hAzgWDwGOcdC3uOsqtsEqaEcoW9NDPaCrDEUEcUWvzxnGqggu4BUUHDxEQtXSj
GWaMk60ACfD9HW2sjI+8PfjXG+Pkr188xQo8kSZ1pz74RRcAuICBhiptmHlItuIb
6EburKVf1t9YVERG9D6DHnCjZl0zlWaDObKQaqTc/sMDnjLk01xc9Cc3g37G0/pC
SI5q1qjRTlUmVAlaWNolXlwwO5mOYqdhhoRw6ujQQpi05pLR/+8FeqL6tzdIqY+R
yIxemU0Vt4TiT2ANxqFnLfcUe4K58HJ8hngEQhgu7ZpyVVruyr5imTUwrLNOoWbR
AMu1JLWULzSPg55Ji15v+UDimGqYFCIVYNf702RDzZ2vjLuwd2nvs6nR2AXGwt1F
qrKtkD+lHadKels7XB7V4/QaoL1nUCDx4aGnJhJcKwBo8WOKE1NvNCO2eJR6r4Ym
RhZfe0RNdoCSswcbVT/1bamFx6fh6nLEexU8wnsI/ibArdyTHX5PwS72mAGKrIzA
1dENU4BIVbLv+Wt5x2c4tdGuUc0/Fq4PFotok/XX8nMmwWwHGEqNy39VpAuNOvcv
3JCkVi+N2Emonq/Jdk8feD27TKc5FxIOBjvd2KxeqO1J0oo1XgKo5ofwQAxFIszG
4NF9dVNoIiSqs++Ram2uA1H3nzPpFDNasLcvfbOE4XWcFrK/0Y+1Yg7Sb++3jlzo
50RkIL1RsEPbqimvVmswvuWnu2nr3x9OU6EIl3K8HTpQ3BCog7KKLqC6dlDzpBp4
Z/FUmxxMXL7qsKyqpNRCKfdddzgFMex7DdrlKkqAC8EJCNvyqjy4gSvorWuscyX3
UWxi/AZRz8IPfEjMfuHgfOUvcIj0B9hGSdFc9mUnSsoL3y5zKkonSYWWhIDKw7vP
yh3/H8wc58IkDBCqvVkOOwzdI+ejpcLK8AqFWNQKku/5zK34JOII6Ot4CDGhd2Xl
yhp4YXfD47m7LeLXzP/cGkPx4rvsP2eUUdSvNuXxLK5WZCfUk3x3Dwza+htkEf5p
3965zqfoiFS3aDcf18HE+8/6d2GxuVoR/40+vgIsG4oKQBwt5A0kOMjcTSc28PXU
kyEucXMElZeCLpWbFkPz0n920eoMoM3FNnNJLFKufLJm4x6nyb4zOHC3kI/7ABer
MKoHIINoMeps7X3zjYkZ42vZ+1mAuqSUoBREC1jQBiQ1hyBV2yytPijEV7n5WLyr
vxQNXww+jsDJwfXrusM5ceP3B4UolNY47U1Ke+gnqnvcAL3Cr50T8t0VuQO4ConM
I/+U9wLQrR+cm7MxQyVfJb4cCNPn4udeJ53TdpwkOSNqaIqdoxT9YDnh5Ajm24pm
x4liGnMhDDqQZ0t1PbreDvMQD+0x065zJXyyqi6pMuD//zObZQFAk2V/8l7U7lhc
QraCq3WzhjacT//KSvU+qAxVHlQMJ4/gMxJ7d1TZ5Co8kcH7GtD8Y96b8tRrmZb0
aB1Vc5qVjM5oTqTS9eH/LE2nCCQgndcldXt04BidPaXMflkljf7oFQLSS0Mrk8HI
3NEsMJsBlnKzOESZZs5tW8kCqdB1P/TtS+jz2B7obgP7NZsP25lrMHGxsOQuMRKD
alLwpEPwDAdjxNQs84Y5I74r2dLcS5LrzNf2joh54qfPCoP/uAmWONveKKZkVKdF
GFQ3ADr8Gxd+hC/dilE7TNQ7qbTI5kvN1ppcxjz5VbZc6QX9E1CwOPrikhEo+tev
EZdtwlrhf0nxsPgD2+CcLWzyeS2azti0REM93OLjZTh2GSC84h0nAJqnOsL9PH3k
MFy9vRU9BMZv5Ng7v9G7NRnP91caJsKHAcKxXvHsdLqCyNGBrlS5UmOFWVsssYAs
mbD2zlJ97IZsu1p9JXozJl3K42Bh38jFAjws9kvtHE7xS/CqbapismiFla4comRs
cosRWR71hFpJ8JngnVTuEY0eY4EAHd8mJtTQMIsgm4IK10vFPDI5jOGBxQYqgYAB
rC77JJDvRirG5lhxANHcxmdtdzn2Q6kkDgLMhywxi+e0lExrv8B3G4UiJKevURrF
9DlvoauCSickLPz3jWNh+Ik2bpALpqMD7wFnkhxuegTc9wOMNgLTHev3JoO2jNpA
i9bIStOKPd28fIa9NHnPFYES+H/6MXOtIOJk+tctxKpsbWKYUftgYbhzn4VpHXcM
tIWKBXWQF+aUmgsAbsy+xvhoui5Zehs27SVbf+fG5Zttn4RjO7NKnk7bK/3y0gbe
4HdkJcawUZGs2Jhq8CEcrTJkNeeV8SFSDgjngfVbYCI2TT2V1WaJKBfy/C/0StTa
7n4cjQbN+Kj70EoXhliq/dlYrOlsd9+b0YhCs5g6DUToKbXvUIS4mi8YiUXvlN/z
yHETqkt0xqO5yJXm9pVP+8o0oqNhrM6fPP1UoaYb5eBXbPC4cEH8EoKYywScUSby
eUkCN/biiu/H5UKRSf+DhXjYoIXSqsOvREABn7dlowAB5IInoN0FwFjDgQgbYUks
XEdIwbD++1MtTEhd/ENBLfwK7ykFC9k77axZLefktkBdjLMN//z/kI0t86eTHr/g
9FIEvD7S1YTzyKci3w5V2t/nKPy/2PPD9xvh0rq89rj9heoZnYqF6sgNekUWkyru
cpzMxWgvHjxz8fIaIdpDTgp8EWBp06CNMEPK5WHd0Zf+kEcekKBDekDJrZO/hDhW
cj/X3/e02uFwb4eGrXeKCg8S8FOOqIOaw+RdC/t034Mv+yccokxKMUFoBoz+PzEL
EvAlRNJk+ikGzfbc5sWkVad7J/MnlSGjfcYdpVpvGEC9y4jwfdvx/tdhioVHeFFj
1kmnz/asyc2zjXrytcRVazYehRa9lskcA0Gj4suaZL8MEAaBbOY3dgjPEtUUTy68
R3EXSrSFiMhuN+ZykYHIM3aGLa5NVeAiQYeViBySEW5V43EXaqcaHW4WgHT/9f+9
vdyhtWcjGV2w9xNx1nJ2IhFPYnuWkDAZ01kD7i3R/Uhjdk5p8jZWoGyLZRhp7d3K
It5vTRRh4ENyurdpg44CxTx07rbZAF6jY+AR9trM2M49BaXAtBjtVvA8ZbhsGgJS
2fQCaaxnH1iXRO4uL9n3ITLDl7Y1ZEY3oi9eI0ky4QZtMhEmFL9K034TIYfsec1/
a2CAARBY+gmj0EHVCcARYgECBiC32F2ErNj5hRMGY8T7c/ojvt/8dmDyYkoIA2Dy
gQVUK8vc5wguGuQEF8PyVOK3ogSkZ/EkvfbI2GjTKR99x4Klaump4uRXBXV38QDB
LZHesnUE5Vb1In5f3BoMug1yjGm94tamy1l+/r6pl6eAp5irz1NuCNwus3k2eI4q
Jqf+Q6pZ4SgGDaE9tSHw9gcl2ds49TWFL6smPY4PL4AUQy9fz0qJrG2b7Kpak3mF
dWP3R/5hshcdyzmrO5oVbbs9SvJrTVcOvZ+uO3dm/V6hEohhJov5B9XSMSa14I6V
AvZoHkxRIO88YHmWi1JwGcCrW/igeDQ57h42o+9s4CvH2PFZCoAL0Ny9/nitWQPW
UYsdisR5z/rO8J3KSnh4gLFGz8w3DMGS30wgGEchnF5GQN6TB6sFefQa5T4Xcfs3
Sz5hGmR22Rl2sT4Y6ZNC0krfZlaz6h+xkzu77k256vaLZ5ZQl+hQETiZvlPuo5A3
RVjSnLPpmxyIsciXpU1meg4H+hGFlW3lcCTG3BZt45MFUfgnZh2FsNekfIiAoQvR
e02lv8SVUuGIVYXoO/zgVfxAj3eIz6xRlKLE34jj31TBj9bxLUvDZ0daKTI43Rxa
ut555HdGYxvUACwSMvLQ8KUEjoErUxqA5JTXAPKbbSfFlsonogOcfsn9ejVUoowU
yatmVH1KcFhHWou9VLVhnP2DiJPFiM3HasHHfC7MQL5d5us+e8MKB3Vvsx3YSBry
gDCG+tnIi+rwCrGvN1l/N7pfywmdSf/KMdMPFAwI+n5d9awhIcJ/DOLLaeCgixys
ssTc2oPnczsm/5uQmElNI9zLKYI0XMNreGZRzzBPO7sok4DuA6zjyXee72Gn6vD/
nCFiB0k1tcYFzMU+Y2Cb70+nrnGgkMArQXD2VXbksYZn78E5lVJPYeEY8FYISVjq
9UKeM9r4JHR2TZBozlaowoTQl5uh8vv82XAGJ3jTAwGZENcSb0MVp0FZB9U2m3zB
0gTBj/44Zw4hff5qDZgScx4Lu/ezaUFHZtt0K1OFBgjKWZdc7JH20yQRTOOPFvqo
9E0D3G8D0TudOev6W9VWw8F7WgpS+Mj85AdWqWtLdJGYDok9avAQcSnslGyQaboF
OyZwsbfaiRalcQmhMxPHZrqG70l6ELJwDy1oaBPgzJuzRRhp7mFZ5GA6d+Ye37Fk
1l7zD29IqzGgeqVW+jrVKQbrvhCcfJSr3kEyZacjpk3rNUl6pIWwQCbEyFmhz7o+
RGGvtibFuHuRGvPJPoG8WKauHuWA5Du1Pfq28GR0Uj8mcNRd46qFPg3bzE7MA8HL
xM1CMThTjEZF961Lo0cb8u4eCMDB7w5cMD2CLg9JWjkvseuw8QP5LEnoFc/H7rDY
auX/U6gHOuETtKRchiAVyUTiNtTAX/ibC9OGMdGUuRKIwZsyxBigzZS2Y9VU2a/P
iTHRTsdxp8WSjspIrYSQFwNauXK9Urb9jW49ZVSi6up2Hp38j+VJsVDK8qlJ6ZE3
t1JBwyWhQ68/zVfjxzwc4eoEG/JaHxgLvRt2FU5UFqkvttNUevZDvVgLBMH4lHWJ
HeY4EKLihMQciSQTmpm9gnUs481XkFWaBlbWFwyFTPwGGr1yPlyaiRUb8lD4yuyj
6EdQZn1UH6czxbEr5gkfqsq+mxHctd8jsY0/laessYH3F9BgEUHoW3vrSSUhM1MT
KTp79scnTipjDPxZ/7UhqwMhf6ht5SIW5LtBBnE8n0BjgV11s85OWn2bKmDhnzyR
M5BRACAnDHMoJ/ve0MWg00pm12Pk+RxzBpVyNF48T90xnANux6ja9DKYqFQd9Xh9
8OBACKJMSC7uWJAA33Maqxo+RZC/ab0T9PzrsvP3pCdmOu7JIuSv+9BEmI/ljkPP
URxkOLC/SAjVUhLJH5St7vmCcBsm0aHlH4EGMqWgsPFm1C4mM1JL9gFOkV/AHLy7
8JwE15PvYjHODIumtqvQU2jeyK+P1aFaDJQjt90ZZ+b6CS83H3WH6NeB7Rj9m8Jo
78hUNXOAsC6+gjB0XnNXeJE0IRQMx4bBI7PgR3pav49NYxOlmxAzIHiRH5Wk75IG
2tFmrJbsQNPVcbE3sl6iFjWFubulTpTCjae19rm+b19f0IrBkMe9riigk5HGHKEp
tW534vOsDTMXq7tUPDObZlSWqKQ6XD1EuTpizfHAILLNndTb0hlKFQcoTyd4dxxk
A8+isved8YYNz3Uk4vsePr0F3QLOnXDkWCPzpzoB03uYxkv9luPTWhObFyAiPYGq
j2ntiFqQCiv9NM0ydA/myCxHy6cU1ilvfGwhPX0aDJO6MYFETDsaJkoM5eAXF0G8
zgnphMAg9EZ1DERyp4+9eIwfDZT3JoBcpS5sBAMEhaH+clU+iwvprblEVEXAyRVq
uMlz382GVCRCamncrszVKBkTHucyHBBVdA/MbTAtVWTQmtp/fcFog897r5ktLPmh
brKFheDT8M4gkANDA1yekpff9jrMZPLAtnaLpmvnAm5EiDORzg/FXu4GI1IgomQZ
8s3Hys5Mau6eFgqis13tDCIbM+FXCke4v2GSTBEX/3Y3jEjG88E6h6Taw3WAB2vr
cY/VF4JcVHvqMizPjR6+lOZskUcIXjYUINEQUG1dliJHSnWdSxdjuNZxXvI9w8VC
OvheiHQEERAGs//bO4Lgr9KeSqhpj6wm7G/EZlAG5IsZ8cxIvnXNUHySZ73ezxN0
ozaBHbKOhmChtW6wOF01Q68QY3wc1eBvQXHgyho4I0EUpgq2ODFliPCwwtwitLDk
wUUb0XLjJFPyK7cfjkMqKY4w2IBwKy0WR+5LowzGFlaESmUC+EYX8pKGI+osJCY5
TAcT4M/UHUYcVoSTrI/peJT8JuBWK2VBw4LXgIqWzS4SeiQ9PutpIQTb4xXH8wRs
awDzv5R5q7WTHLZaPk9gQCU8oVe3tWO+9IHW0UbTsbSl5kLLeXqwZ46wVcLWpSjQ
c58kSqDln+6D0EesQ+8dVWwzhOX10ogcaYO91QK/Oj3IiBTNxVyyDzHA5SzUHjfw
7bZ9riMVM5VVTSddobc+b++AleEBImq10B8ze+IIX2Cf7ybd28AwNzP5oyUtX1A/
94iNIEVbJa0dR2SiVhwpWP0FJVsAFLS1JQ1I6WBPYvGOhAIXLdADkxEwQxKNUJS7
NUj7GVPGwsROmIo+panbD1z9zgOq4bCed42/5aOMP6U4Ow64F2zzo8lrxY0wirFo
3BOxKvEyDtjXddnnI1YZc1UzbIa8TtdSpRbcXZCqty6/4G+w+bA7ksXXjcf2BKn2
Xg9ufzkadrGAWc9eP/yJlT/cICCt0m6O1QYz3gvO9icF7wM5FWcQVAOoVrki8cfg
Dphxe5wjo0avbV3U4kx3F5yFvcYF9DpBJS51T12qmFIIGMgzAq8UOb/bweR1OgQO
wvIa6TJaztMr5cMnBEqs6GyXfrKJKpaudhmweapwgauCf8q2Uy2hmSgkn2eOnqF3
u2Vj436Rfdf0dThQZDqybFT4ilRklEUFn8fzVci5TgD6lxnEoc5bxWZp7cuNLKG8
+3678Mmlbom0lA4WXhDAw2OD8/syNwL/0TjGq2A2QE4PEkPkn8h3q5n2emYryM7G
cVgpc9hmUmNCe5W60IqV53wneGiqhEg4aS9QjO1f2LJ4DfpRx99qY8chKAzcBZMu
PBBhNUW9e0b+N7gvkIFEoAqSMn4s9uERycY9X+7gwyM9WXgSLn6b3iWssKK0FY+O
A2TjF6LK+i/yKOycLmUUZu60vDqJX60FgamxmLq9F1YRJ+ru6XLHQDSsioB9+K6G
2GoG8pEPMZ37pm546txWcT7DElpBb0V3/moQkTLbFsT8or8ORoCEq3Z/kcn3jCfc
U0lLKB135oIaWYfR1c35+UwAxj4WYM1ZqQVTD3yXCfJQQdz7rJQDargUiomSP3WB
pnVlCPJIDg55qEqhKm8C+5nTIXnwXCZ7dSIsMhk9VbN12pi5P5wfH8vONVrS19aX
yuwh1vIlpNkId6tFigQdQQPA2GziP1wB9OF6+5x0ZglMKAsyCItJnDTiOXnhBeq2
YS6bafWlYdIpyRdVg3/nsII/MfwLM0Bw8lFhmj8hkiOdniOUrE2UbWNoXY7kwYZB
fje9MpCWcmarpfmPF8avS3Hx8H1ru/YbQZqfrXtTBJRsqfnlbsGfaBxwKs5PzC/u
nXeqj24m4Eg7pmrKOIba0me2WNN7PPPk2ZlPF8LV1FyQddOpCGGHv6lqwsGG4n/K
nvMeB/UMseL265Qqr41cX+/FecjFaq16gTvrbisAWl7wVNBH/26BlOW11iYGXG21
mHMN2niSpcQqCcTF/Q/9NIU+bgo57O8Un3hax76aXlp38kxvVXaK0t2XlXg0Wdti
uQhhXSjBFz/+dPUEaFdqHB/HDDeR2PQ4NAUpdm3Man2Ey8l6XfjaUpNP33utSyaO
MjSDr2nQ7eF0klKGJKuDJoSZ/Fu8efSFjKvW6kMkZJsgIHOpK6xVplqo0X2XrD5P
gO9oJ/EaonmVWlZleSdiBcQcXdkxFGpm5n/YvqkkO3gKUdNVshWtO7YbFu9uyZEi
rYaMHVP18+DHHp2KHnSNE9WkU0H3uPQbzOZFwejxByhBESMASU6NU60sZwx53H0Y
wcXjKhWKIp1C1ThneP7U2PSudGC9nIbLYgRGg1MuAWJVwWErtCQfC3iNLUkA5eqs
o447mRIteSu2bniQEpkpuu6b/VibxPrCRv4hLJpCUaBFQVjIeXm/z0Dsrexte+ze
G4ajmWUO3OkkRJHAda3zUMh1cpWQ/XSuBTb/Pztmjd5eMFwkiXcTzqPfKOM49XTt
G7M+z5TvSHan5Kl9ONyy+k+iuUddGEX5TU7VNJ6GhAsy+cWFLut8xYIrTJ3cSP2r
ycAVUqnYv+2LfghgeFWbUKaXR8OwN7cs8RN/z3hzpAoMnjZdV4Q81mJIi34NMu6b
n7noai9Qo9/YXAlA/pf2UGdM55tvgfriusfDNeLfM/Q+yYIS9+YU2GEWX+ONfGdP
OxUgAW6s4StTNtCIbNTCxrf1HcgzZXUCrN6m+NhKJesp7ZEGWMHcX2pAbU5hImhC
vzsyD6d5o7tD/0cV0m/12SDzk1algp78Ep4D5AL8BFdGw6q+1p1nhUiPkKAhT+AU
QQAJB3Cm0zbMexFoLrxKdZVCSf9ksJY4bM8MxOcMBWHW8ktMH3P95mbD3FIfCw79
mSTrtH6yAGEWjXQr6AKz4XuklOagcWJ0Zcho7gvbb6BBAkRQ0CdIW3HwjaoLsDHW
JT4t985olssfNgevG+CnnUDepbIFWDS/rOMMQApebXbCwpCOStY3qgipR8tGUG4d
WassPZmH4RZ+LdrIR3w0+eApaIg3j6ZVbkxddqZCMpLiIPRZW9IvaETawOluVueS
68zNyBkb6euP2y7MSrkXgYmohAzMWJDvfK5NIfVEHh5mDTiCaaDekShJ8MdI+R+N
yelC1bzNOdLNdPiYCG6gcNEnAvuI0i6iPT77eCn/KwQQgECfvsXp2mGperx91lAF
4JlWHfYCEWfCzQ91DYfNMRGy+ocf5GRUbZqlA070Ynf1/OVMhjZpJco5HpiK4iRD
Qij1j97s/fTg0c0v3JPiMYrHy5J5ydl9Mc2VBVIzwi0QnrwPeB4xGnKy6VsaJLmD
UZbFmIgH4FUDztaj3mqar3hq6E7MJ2ClndJOL2qjctu81k8uIogzLSKxScRhVPBB
XASNuXZATZ8pXbOYqOsADhjKBLuCz5yH0QGGpagfZxeLhh72P/axSQEvtQrR+b0u
bPGr+2jcBGdM1hzNq8Ummk/v3RPfW1KnVKZequp+2AAxD5YF0pgW6ecq5p1BDXX1
FOU40loc5+kNgescQhFCm4teCjKMJ3DvvIlMh2xb6ok17izl1jevuhwUAP0zBBqf
sRc5tyz07Y7JECPZoFhjGx6FJiW46LZW9GU5xOwO4s6N/+9YOkJ31ZfLqOSZgC3l
eCY0JFBkDxPHofAF7uQAxmldBmcpbVimGVHvUJTBV6o7TIRICb6xx6EM95hcaD2v
gHTzHnKHJpUrxwJ+14gUarYOunT/BtKX3IgiHQ4AoTzvYGZTUYtVlhSCtkC2bn4L
ugG3UVfWFrbG97Kus0CSqw5eHOINRq90UsgdMFkwoxKGatCD9z1HJEMIYboIT4Ag
1eAi6rOFiBg0ecpNBwWxn/e6eB11asopTkLERYlTQllzDEoh47njC4Y1tctf3PNi
VU6FoTn+NV51Ri6douJy2U4UqMdhS13B5eHfZlBdc7HFz9SWfpS3Wa0Xs4sPqlof
WvjEZ9ohjQtNbFxLIVQtfzriJBLRWZ9qbsbWNoHbsieioNyCG9ULyilBmYugrJN+
WqGtOITEWZct3J5tvrMpKJxzhqbjM55efZu2RpEV4kYAhRbkw3IKUDPbMF3L2Yau
oRQUstBHqqQdQcwGhGeC+sR2b6TJoTEq2BoUWm1WFxV3l0lvJ0XuS1H5hk/lveOG
Nhg/Qa/gehzLKNwKC1dG6fNPefBjDPDgFBa0JBfaKlMGbCdCn4obp1HHvW5ZYUPf
GxUWjnnRZKgzQv15lL/SuGNN59RekcrvJHDRIMicb/yeMydZ9Up4tKxQlQDRHCFT
Mf03FQjcveL62USmBbMMKirE2uPZezTM79myLOnLnxlRMCRTpn046vl6NyvzLz4o
lf9VY4oAPZOtp+qjc64YVf1qtEo0Pie/O0+SSakQA75I/zhyc2Zzo2qmBrfZlrOR
eZ/t/zbDyaSdL3zuuGighUBWhapRrfEXlNz0LOOsI8n5wo9P6jJ9fdQKmAPpuBo0
3fqR2g6oJWyZqPsoKugOycDXLbkjz19WzRkCrxfEn63Db7E1WYkmlWLTP0hmgN1J
La6x+5AfsKUAIZwbzVo3XQh/dm2TEXdLRzPjtABxvR5In6xkRe1LWIleaK087agr
xYEIJc3Pm8r+U1kfcD47SLb5yQILQxAgldhSQWoEd/QZMNCdyX9e7rwSuEkmeD0c
tU/J7vXAOglr3X9f+JAmV76+D0DIfCRBMxeHpvQx/9tT+Bl49ZoZFd5ErFFCDyHm
AczcLT6zR90hOnUu9i9CwAxzsw/9aXoxFmszh0dOHNi1bRgDaWDDATFVBpghWixH
X02hRVjn7dC4ggFjlmMVNx2Jv5gs/3Zdm+KqZ4kosJk0OGCwITnZN1a1ziZJ7MJY
/1e9MYOB9EwT8gnA92/F2U916pjEI/dZWzsBEZZb5rycUoQxw9AUs84G0y66w4ku
`pragma protect end_protected
