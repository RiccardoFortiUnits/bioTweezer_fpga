`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J+sSUatVVLszFhf3AdmiGP1JgezjW+ga00e8SSBLFG4qhoFqop1qKsWYskB/iIiR
gE0dg/P+sLWyvKDy3cdO2cMLrrzPolhffgX2izrrxEMcdoOJyv07txEOyLF0ZeK5
5q3fmdc+PY6aDKULv0KaHG8Y5u7tK6+dnhP47jUaC5U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9088)
sOMaQjdx0heX3pqi3lI8H8zYoLye+Xw2gbB5qGaUz/7rgEDIRGR5SBEIpt/8K25+
EfCh6XO9Hrb7s0icPz/l/SepYlRCoP6uszE7rbczmsPVDvNphNVsJ3xvc9p2aj6u
hgnU2CJffwDTDnkv3JhL6EZBqp/qObr3a1F7Tz62lSJ/MC9+pKjcHJREI7nvQJJB
0dMNK6aJiwTGuYsmXrp5JIky9GA3KFJJcqI32VJndd4xAXOaAXzbFS8QbwuD9gDw
q2jArDKOuKxj+r/J3XsnNtYZO0KJ0NNUaSmtTOlvcKI74SH1m7LgVU2pj+JwM6Fi
7DiSp3G6v554mBmNYN/BsQIFMglFwgUP5qC9Ef0P8K7eU4odWg90jqZUnIhpnrsY
9yFeJBiHvwVy+Mj+ArXQOrotP3HXfDeDNdh0xmoHs0I/Gm9/vdJpFd+8X6hKlc1W
hKP2+wPwhjDT1EPHkY0oKdGzJYUh+xKq7d+pcIcF6aigzpBYZ8QoWDvrgjfST0lT
hN8kZ6tTQrWGMrp30JvcUkL/cqfYe42pCjdDlxZkAcPkXwhvBEroZzJ8nCSr0Xh7
ZpqcqYdCeVA/dTGNLIUV0hBPmNTzH88op8SD928HZ6S7EcSe6y76+4tNUOd1AjGz
0lHNnEAVZZbiOW6OJ1Us7uoXzavhGhwkhwEWIqvRgG/wUE8BfwVgX7IBXJpBNHdr
Ce0f+jlfCApyon5lVJmUkPegH31+sDl9/sgjY6ZcbUKXfTd9BR9PhqSnZjsE5lSU
TqipO/sRFEf3DIClTuvDTRrhsaF8Knersg3A/JlBmWk8I9hlyc6Qnxa81kmSUZ3K
P1AFhE9nDPU6BoO24OX38pvx84PkEi1FGY+YonnYi1+lQJijSG6xgy60NHDU7KJL
wezYMkZU6DYI+jO6BNJRt8mzkfuldd1WO1jc18caYxcmmtcBHlFIP/C4F8F9xesY
D6Wk3ADNW3siqQsm9+ALfD02pV95CwVx+M9TuWvNdF8V7oOQJGY860OhNekJnhLJ
CEc3KGR4KwlGQS0GUPGXoRbj94rFV5MQfjNOahx2W8XarMynypInucRPJEKfDj0D
uWqpedxeLuFfMwno50+hMQD7SAtGJKi16gTr0E/HmOcENr75x8J2BZR2pLn+c8Yi
cs4Zza+ui+TDILgijjgtvvykkRyaYYyJMlHiG6bClfdQ1X6uvl1mK03syKETVkJg
YoZ/5WffrM0zemXz6N3GX98tA8l/uSZKR6+yWuZPaGSiswSvhSeXxRwhV8UQY5kK
7zpFwi/4KcdbA5HUfqp5rGfNzECRuZWwndieeJzd43GOpGIc1FuhzJodJsNX1LLs
rqzSrAfRf7eowWN3PC839zE6Y6tDX75cRUa3joPG5cFRGbaMT0GmVWaSATjlqiE5
AqPs2ATlrhF/knJ3ydOWT7koAjEWAsfgQsNQEyC7JEtFUTx+Pcc1t6KbkrSo4iad
CMRfsHO9Y+uhuP9iSQJbwaowYeTX/6WddvbYFuzTfaV0Tx0ea/4EzG3AWQ2BWzj8
6jSYHz2E9gMhnOIv052KBB2fB7D6IDC6Mwz468QhHIq+/9R74nYp6T0+Og8OVP/2
osNQecjau0mYPEIjiJMdnBV3uJo9xEF82acarvmPw46dsB6Z29Yt8ObvNkKBLrQa
Vm7fbhoBbiggIokG3ssrBWL/F9wMXy4yAd4bs11X68LfPcf0AzONfn6qtHXSH6oE
7vdfj5zESw7zICXLplk/fICCcbKerUfajk11YnWNBkO3/Th2pjDBfuKWE9RAzxji
/KjGA98PQShTEcoh0EUfhFshs0RK+dKqraN7p9i0iG97SWHBwZpKulPmaAnPbmn6
Whhqoc2SmFdaXEGHBOMVl4wysbhRkzUSCiK/wmOpDFDzj+Oocm948BxXmZCKVoHz
fJ9H7AS40OINCOm4vB1aklVTA+yyIMdFEHmH1dnZhd2/dDDiBJiOJ5q0EhfHgfNo
BDnOLww/o2u2XECGhkthRvMzX7YpH2z+5RSa6QEYMvD1eSA3EZuryoRj90F5ei2V
nyj2EyDtnkoFyWCOVHmWc35UA3ApaEhL1GpQltqfuTsEEPxc5hLKd7T4AmzZ4JNN
YwVMrsvdyh/rKBR1b+rfvf++Xu3jDsDJtGYAIYS9GrTlK+YJfmqHr/RshxVPFpQa
N0XSadK85jY9u5+8xcPfK7tr1OxxopUk1FC+A4NcKJpXzHsPDHqiNQACIOYC4AEB
s1WYStwE/MBK8cD6A6/cIU9f/9Hi0WvRZZ7kIAEvT+4IWf0MwNESPMHQX0QN9brc
P7Hj7/eMc553PzUAWzQbaiRBFoXWduo707d0Vdpg3C1WEUmXpm1WOIBvs2/yGAav
T9pRBPPZsBYwxMZv5yzvo6CezexOp41x9E2uL5I90cNXeZtgpRz+GCgK0v20dPhx
2j3BoNrxrCMWNoZufHyB8J80Vk6T1IeatkhYFoWxjmxOGnfnopmU/0uf9JBRH7ZU
FDOB0R8ki92QcKF48qCGeuMkdSXxqZ93fm7m/8SuRwEiVF9hU/1knU0sNw/KIKwh
DuDDrCfz42U3TUKm4ayC06NlX5y8eaqY1vH9SIbUGyCcIwvfXmrxM06V1unKtvQw
DRFW6d4ArFnjq2pASPY7IdkVPat2Gqf9Vshbe3S3SudI9i+vmezN74hZZSB/lvCC
vamYUGZiGKlKLOnZIdobX6Mm7bklBGIMYw5MUGetZaUqommY3e9a7pbRVKwe+eDv
IVRZsvQV+XHrdKaRr2cGV7jIJZTZLZydhI3UNxyUrrDLGLoeKqkq6M3lkJzpM1v+
dowZMlfby2zoolRIztGQDLjeouFdq593GdQ+hELnNSuJTvQUkbDNqJA76yfjlFxy
3ViY86yKLkdC/EcQ7YHu+0eHW0UJvxO0eN6AJXiDwy0s4A7I0gQ0+m1tB1QV/wec
1tTJTwzO0R1gQfapYsiEeQcp0gECTuASeXu+lodEtDn/9xh/LmRZ+UQbXmRuDqeY
JFr7875gnBTCETUewpPCTU0Qzp+Io/UV4RWA8svLXnzLSD4UNSt5bjmeE/Zj7u7P
tbMRXFTqD/HFk9LtKL5N6Qfn7n0AWQL4CPB6CUpP/19rLDx7LGgUuVn33LM213Iq
xoa41FHyTrpuRS8lHUj0xq/XC+L0VBbu0ZGw1igin5Odfbo/ohO78wUgdNC+c+Tk
g26GH9Pz+IiOp/LmmtwwNBlyrApx7N6iX7H5yDQVFfy8lFeuUZCpCLCOhMS51Bcd
uRoHTjUFCrnG0nW8IfT4oB1kWHYLNQQ0OLkT1JCMnEhxW+Sng6w55NMFqZHCMNf7
oJ0BdxckQGfqoay74gnWmtt7E01I72W8riAV+T1g7URrBiUaU9imGhwiFcH0soR9
5z6rTJ7hcnvP2yK0tXkaWcVfmmVHxTr0h2CKrFODLGFkb/GHFctbZnuM1ckOMH/v
pdvc31wI44gQMrBEZZx0a742LS2ZqyfgRRw7ixlDRlf1lb24xZ5B/ALOEdNZEpSc
AuynVWOuvXI+N6V8p9x8TY268ktao91Cdx8wx2AVI6b8bJ64iS2lW0q2ukW0tqhu
7LKRnShGAe2yqCW7rF5AlrFLuBsufUFjITwzjOQxv9phEGOU4biXQOsCGcxucD92
7scwme+8q0vole7QPmdcijzWpac/hIxhsCKX1cjKS/FYWIuXXgdsbAMaTJByVLkn
UfHlo+qFwwPUcTggQZmLJyUrzS9pzM8KMywvxfCoUqUMXv0R1oUcmvXLNl/DH7hG
VMTfg3A7DbS/TllbEhIB9kCzNSsrq8824I4qMOMj0y1IiK9PvBkhFZxw8llG+9Xo
Jg7pwqzkXtCvsP1tYGh22dU4HsBx8zK3yl5XWjQ0/OGLJd7FiFbrG2enkmkKU6kf
HetaxRb4XfkIwTzlRlQERxg5d1+7q/76kDu2QjFcyw3swwZVcT8bVZFuDEiIGpoI
5VDkDF6wpsJhT+D4ZThN7f+1WfV3J3WYdSqNKLlp5gE2b6gfRTu5P9q3ESPEDfIT
wdDRm/cF+4HAtgV7sLg9O56o4y2zDAo7HNxwxrDHbnePjXKfGjmiQ29EmaJz+O2H
bBSdkLRPpis78Ufo6w1RsxikD3grY1OA9qVOYCjCCRF0kJGjrpX2j8qYitCoBO0q
riZAfvqoKh90dEva5wVOOjfzrm3s4tDGocodLNTSOxYnwW66kYw9kRggFNDhYNPp
QibCtg6KiCy8IRzy6bKLDdoEZRLZN2sBBdTm+u+ukCIrH7Y3f5gC+l6BcUKRV4JB
t4WplXIXRhYVbdzKct0RQZyX+Sy6FlA1funoaFtKUHyhAM8u9M3tj3Uu4PlEiuM4
kXTAf2Wh38TFD+LyK9CBIjk+EARNYOeH2t7NlpIacEJf7GwVPz4h3JOIUm1a4vtt
lvOWcmCifVzkBmAcMz29Q8H6/iqf0i58PLeq06wG7PolK2zmq8cAVY15Y2Rg91UT
Gl+UFNjELNlx+F+vvHGWbMMkvv9rY0XB4wqmrdseL2QeMY18yoZSj6lT9CqtAIef
o/V04UqyosJ36gEHPkZ8CmiOZQuWFAE5AGhR7/ncG0VQeOFJd9qKET8wmimsf7Jn
Wg+rdjCpS2u5eNu3jF5gOdB9sTngRdT0xRJTdVCI1nR7l23Ki6u1ftHxkr2jnQI1
rg6053sYKz0jw74LRbmOYcg4ysP/+VBolkqDoaX1pHBGV7iFSjdn9Cl9bN+M0MrG
+ZsZ6Jl+w8xsII7o7Y+a6Qw9rA6zWOEM7CFRAjh9Wu2fRGjHhMc6KNh8BF2UVwjP
kP+zOcGfXqI69r2wMmR/rtQkm8UuOEXAf+vn5QaxYHb2jUuiNDDQm2eJY6UjpeJ3
WeCxx0DfpeJDcSuYkUBAelAXY8vxAcO9CUAiLev1gXFPEPbg8EnIxxgmzEY0wgkx
et32g5h8ci9JuB+ZvIUHepk4e+8Uuii38hllxWK+FGASBU41fpC/NH3fy7FbyTV+
Zcv5L76PLGzrUToyDVwaOyGo7xDmZLPqk/HGVMbOKQD0xMDYGV+q7ywfAYgw8r92
vT5/Hy/PzyXi9sWMiq92gF0nyxhOVPlFwZYoUIz2Sqz0qQFN0X8PjYcAJO1WE3wl
8na+6L++umWUGDlIhsY3tQkntNrhBBr7zvxj0aUjQzAL2ha+AQeVgfF9xihaHPT/
KjQTX8+2dAL/RKbO1zDRiR7/4PmgQhgEqWP2fSuSsJT6tOTnXXeTYkBhfVEkuyPz
oNrABh3IrMMuHRB1z2ckpX0BZncYg7pv9ESxiJpGfs4lwJonFjkw5C7gh8xtJd+1
iVDWpIV+0MNZfdCMVLXYrtYECLlK5zdws/HLcz3qfujfQV++P6LqRJ+b7FLZAqC0
4EXGhXexmlM+c3JzRo86YvO36wLHEpBVwDVbo8q7hgZStDQcZ43rISf6aLC56y/I
23Dg052fe0+sT5k/adKiYlkjprJHxk4EQHhFScmnz2ReotrlmXYrcjnaYKYrBXHe
WKXIHlYWaqZv4b/zW8w5yrHWsCK1Z2AiSYF2hYyDGw/tm1tie/7GAyns9TVPxcDq
cIj9AyhOCkIgg1zYmbl4jfraq0h7YehAIrF89fIvtbResI01fmxyDEkYqzC9cIhk
tHmrC7KpvrdYRVjfIvJB0lSm/MHJCQBR7uErjfHNp2ICzuqGTG8MUHFjMOaf337X
EeSoQj5lMhpQzVNWhwgVHw2KDrI03GJprEhTCA3V4sIbHJKV7pWW4RGwJ2n3pXch
rXz32e0jtJPVhVeZJlU0bXacD5AxKb0CJU3JApQZfleThWqtwGaQm2zPLaI5hG+r
pUILa87tcNhL0FRuxjXUDW7ACFLu4CdO9NMASrBLmndaN06R13AFY1gGbI1+CjlS
E9ZaGLMdNhHsu2fEN+tshfQepleqnN1dICFSnlErhh3ST/BJrYvp0AMEORA9vWet
81Dney1jJbKhowKE1jivyZaWRXN63SBErmPxeV43o/eh+HSuKyh4LWoWT7gGm0Pf
ienp0b8FsAI2VC5s0yPZUuacm4wvqNu9KCfS6YHikMPYyTKwFq/vm1kXhyf3n5fp
DG2v0AHffeMbVTGnJ2uceiKikMX36R/naQvFITrX+n5ycEfrZ+zzFhj9xH5S6NfU
YjdQxecnlqml1gsLiAkZncBIVsYeTV+iPMKEyZiITIzd0W3PdgSNhQfw+mGfpLLC
+N+lw6Om/7lnPDcpudm9cBv6ymHj6Fs3MYiebo3PeektwOU8BX53zvC8q+Itt3kZ
NZunGYaiJJNwP50cpey7ae+jnqFIoIjivpgXDm35ACSCad32N4gU086Xbbh0Ahn5
pNlZvDX5ahWgdBIBkH/cpK0DXqUt8jzcGQxW/bKqns1VJVKk865+OoRfA+22qrIO
oMuRoRXwmxrlLgq5K00vEMe/FClDY3DZ5YCOno7coj2lLgphU+bF0xltfIyNKDwn
48JSN2IW4G1BeUaXmvgcgtmaswSKkc3M/gAGMVQme8dhcBWnRPI9wLofRewuzYB0
YlNBZlAo/jiaJrklHwW8k/DZP4viqfXguEk0WZ0n0XpqatTZg4o6HGj/4d7pdsIa
7M2Ma1qzgQBh1ogOxOWGNNK+fNOne9YPZnpZfYiYgAc4mRQW5p1lJGlt0u5zxMbs
r8xjGy/ThfiVhoYc4yNj3jN/0I9KyfHHkHZgExgIJE1CXm/nzIVYrBJ+DDNhASBi
DBdJ2S2mFo3HIKuYwnUP+5/JI1UTfU+KTMKwcBNbKVaBlqjpQcm/1rrFgxdqelpv
lgLSEhqc/ocWLpp1Ai78yumCSwEUSs1iLX34acYHPyS3s2I0Ux3reksduyCEWODQ
j+6MdT4ZH7pbBjcb6L+FSYDUl+YNQP2vZO44vmZ2Y5TqFpiyoH7p1SwefOmaWzxu
DmJJqFfp+QTpC4N72HOzaWPbK7VV/G5fh7EOLD6StNjnqG7dcpECKCtH8vJRmnwr
2aTOnMPNXS3bP08v+qX3j+YMrTE3rsJozEpdqiXkUtVNEx+w9RUZa5lNPaRCiKFj
1qyIGQdRvd6YySSr09nMyZ5kVZ/yInJkhmhBzTxQF9c+k9rSV2Ip0VzesFCjKSZx
QQ8ylgU4El0vb+ZrG2Mjp0vuIqG8XwP1hUSPCzRaD6iqGgDoEE4oYQPB1c70Rxrb
m+TwnpOGNDyJPCBXCxvdGmoF5zgRsx6h2PhfNbnkLIQOMdT71Dq/k5aekxuTVA8X
VLFe9hL08AvXzg97Uo+US/dCjF0SYF+E4Zd7SmqihCZiCI2H7bz/jyk9P9vUy3pQ
brlGjQc/BlZEK2wvRp5hQzM06WSKUeyGmopk7FYSmMfeCuN+IQT0x0n57VyOhc4e
lRxuRvWc5C/lfOpC36jlAR1mp/Jk+EnM4IUYnipw7nm9MOB81sMH43wiP/Mmceg1
PHkrGmtBF53r6HISa/EXZoGHrC4RrpZM21V2YGwBXUqLGH2FQDrXfWtgucZtKntY
+XgKcaFHGrnTVBLuw5RJbY86SopyM95bNQBKRfj8plJa8BuuIDe2Td1huuOtdtKn
Y88Wq+7NZcDwnAdfilC0SR2uH6FCNcoxLu5OGtWwsWOVUfE3+DNOrQKO8zRMuuOV
VMUd0bcaUykx22j/NGVuEHU7Th52KrBmuod32dzDOK1SrvgZM31ik3vSCt9UeeD2
8SEyh7L7b7N3N/JxbKygUQNI51HzRVa0JMs6QlHxovk75B9no7eyn+t+qVkotg+I
b5+Y2EXcJr49w8x06K31m3/BWt33afbwoAJ3ILngu2Btu55LxTAVgMUwcoDxuvhv
7E37/Y6TzMs0NzG7vxORnyYuLifBrzGLnHypgt7ltjEeIKImnonwtNxLtjDukYne
8TIT8Yni11Nz4VdWs4HydtiOS6zx2n5qn7aZ4i8XzCkioYjImfgnYK0PyY8DxFcx
iL9R7fHfCQUaSXlJlJGILdjM9cw1wjPhSX5NIJ3DZ19xFe/1msUZ/06nPYVjVXDO
DZjjF2AAHP47n8+i1lMNcfTEpWn4ayONscUn5QRkVRz/y4IJ7+HwdtNTBlv26tCX
bS1803KV3eOLtnFGL3ynskZUi3uPulWD8zlS0GI+oBKWLDBvcUJ4/VTz84yXvnA9
/uC6TQGGLvbw7UCyxnHYYxvQgPQtgi3bNrer1cmp62yGfdMjGd5VlXsICbSpL54b
mEHxNyP+sZBIXRVWICAgy0lxRhaMelmR+0cJvlSJXzMzvtKl5lzHfTYjHykK7kfN
EsMXwqy/k5O9Y4yAVbBVBq81xBYJwuFV5iX8TYJOMMeum24L6a45XRsRHYQ2uFoI
Q477HDj/rvzcuQNRYOP+cvg9jGUL3hEDbQcots4Tou9ZljGnqlIKXSdJcrRuNW0H
BBqS0ab9VtmgFeqRaEqjfhTiB6fVoa5BAQjK9hHRnK/jjpUG++j3d3BMPFUCnPo3
lGZduojekCSzNYBfcoqWrabvgLaPHVqwjFpH2vcRwUBxexFWXI9CuXi6TzciIm/K
g/joHdpdG4ZKq+6B+GPnb4/vWQroXKp1OaVicMTyGpOmWOAwnXVSwdss3b6I1EsV
+rEXDxYK79o4OmcgdbYB7aDoouyQyZN+pQVNLNoTtezgQMqhaatfR45bg/U/bg2K
YNUqvp6V5RqTznAJhnFb/+UOAI0Q0cRN93gQiiKFsHH53wVgvY3F5QWsF5gSLCBf
YC1YRSHyew2gtDVZVum5m1AlzghTjv3gk224H7Vqwok56/xklRJr3/8SB+ZZ7ET5
JlmX0wBOEoYFOlAhBqkBr6V+DhSuZH0o/fzbrCeTYSdaSF69YRNyHm48HFA1Sb5q
/unjtYvDZ9Ez+K3PbT1U4SLJrbZaWtH9tCyHZ3ZBJAA73p3wxFfyt8PBg6MXhjQb
9xIAtpWim4N4hNw3ouCWQ/VwGztUk6uI5UIwCWlbRgb9RxfQHNNOrVeTpmmxwMSX
WnhUaoB1y4GVY14rUtPWCNbWKPBVawGjFOFs0sggt7lLMu+ZeO9zuAPpdqo+KmN+
pe0Z0YfztZsM9JFhJeK6oclhZM7ghbCX4fDQzLf/uN388yrAurGz24K7bMpytmsp
6b8Rv9Is6MWQpnjvifspc1wzy13CXmmkw3DIHpiOfArHxSyu87PAJA6DEJ008hbf
iHMOEzLANgMxwSDYPn0OoN9DprWJ3pVI317kCqCDocx2PsO+EwgrQkMfcuqmTEd1
NDVMdPHtzfx9jmt9ZITjI/J+LmB4K+wifbr7RMG71AUYPj8zxD0+jG4Wqa/7unLn
0AJukMAnFjBAfyOcaC4fj+JcjXkvJ8+lnYqXrgPahQEYdCBBNoMEfE4rFRnCwi7R
4VK/D/5yKvPO5kklhyc0AizhO/edGcq4jXrITa2oOdSUko+eFN+QbuaNqNQqdzNd
fthzf7ow6EX9HVohgckj8sN/xB8kdVdXelYAZGlOontIl0vyOSUYK47NlJ2fdGRb
2y0wE29+r4b+0TPq8D4eBWtpjY3WbvVsqHl/orYhJsa6h9lunZO/wbyeCfRwENLr
Fc5e0nTJpLDDSr5q3WzWjxZpTPC3RgBTOb2M2pWbvstdiI7O1TzxKWb0N+lA3q4B
74HQ7kitzgE/ljvc3pd3ViFZbes8IyfoAt/lmtewmyqc06O31JNm2pu+MXleBdyw
0FqaN+pt4WVNosxrTXH44vatEyggLYJNBbFOLAuqIUo98EoDgeAOZ/sRqM/TkQmv
9BV1IiiH1AMZghoCe9b3SZ6RwQDjF4Xlv3GdFJZXqC6D/W4A3p8Iz3gNY4lOnBNA
g6iLKXVN0wGooYXiKasH/3HBBODBQfCLoR2QSy99NdHi08234EDODy9kAqwus8di
WIZwI/IG5KL3hPhzEeRhp0hhhvOcG+580Nf+hRBTBJVZ4YbKAh/8AcPp3qa3btoq
7whHlCNq/SvRWsvHMwFIZgkLgU/Soeaivzvi2gS6vBelb0rcFmJC72Ko0b7x6gfU
TxV60ZTeT8rCuRZMaH2TNtPsoneIDaAUPKaO5KY/GFA8/r+Q6WCXveqYHThvFEon
xIFfkS+6DiR33sfn/91U3FxC6M9fLRp5IXTrwXQ0ZeykjQyVK0wAH9e/c9OoMzHk
CV017Aym74hnubVw0ayNwULp3V8GeqkDOOhz42T0voF3lQfCYOq1rPntEkmeYdn2
EZJDRT3+WxKp67zFvyUcG0fru0zdz1cnDt03RPisOdMBqD2OgcnFtITh5hh6eCxs
G7IfIHlfG0B6xshY9a9oc0ovZUPg/ICu1VMBoLdQC2ymNcjn8j4zXxPT5ueHszNK
KNiJBdgd+beSLA8UaXj1XEEG5uyGL4ygYOTRC0ZtMFF1fCLtoGudi7xZFWM+8zeT
5HOByJTibUgtJfwQFOWwBxWoBlf/rOwsgfvqVG+AeZNXxsO/+lWItIS2FG6nXS8E
sIb+5WunmZqQIZi9PR11tljQWP/r1+bH1lFAJccU5c2O4HxuaNKVJ0mBvgaL0mtw
lIyvOYnrGUS9LNXVNoVYdQcsbZwo8f8EM+21kXhDjz0wQ0L7mWW5//hcPRtNVRCb
akYAwEhS3S3OQ6UGv0JRS6G9Y8Poc+erGIGyR2S2EPvPKqfkoScGlvZ/lJtHCEcy
giADDbrnCSMUVT3wHYAJoN6eMnMDZlaMqZ/SxbS6zjWUe5QqwCmfivUFmkKp0iB9
Y44Gs+lSy7DlxeETmbPe/GNDbu+N3Iihd2hbkKIqdDWuMtyNNXXxeHJQ4Z+K7Vag
6WSPCQ1+aRiSu0fay2Xa8bgcjw5KEw9SEzj/HAHYwztPANgUndxyv5VXNnlyClY5
6EVQ/oXOjd+Mfkr3BcsGNsZ1sYDnOdbDOekcBq6C3l+Rk/JSXFph5Vl6nMoR6K94
O5CJagOBazPPAIpANODoNOBpRCo4GuEEmNIG7TId9K70GLnboMcEd/O1NtN8kadJ
6+v5wnD1WSLeM240LkvJhP6a8f96pA9dg3hPyZBaUSg7RJx/IfrgYffQCJ1U741G
YmI6ueTLtlnUE/InYz3ohKDF+EcsiADzOL3d3lk6StudmqDHSOwafA8ZJZhQ7kBJ
nybo9SGsZzFx/RY1ZOD1CoUlLkd4K9iE/SPnWhcwH35kMicnjBj43PNzFk8xJuzL
iQVTk898ipXcxAgPblhfcRuMMUh1FsXBQhFmNlsq5Dwslxcse7Vul3zX6AhGPlj6
xV7N6sb561cHGAksFapAI9z6C4PMzzJuf23dgOSzv48sbLGEpIkYquzDp0MR0uiJ
ANPMjcGbqgNeuRoMdX1B8TNzoe2HPGw/INPH3XgKrSamjOaTluEa1ZTH6IruHkWg
7xh9tQcQDBJvN7YWRw8QKjuuW/SO13pW4e+Fq37Ag49B+TkAmsEeij/VYxUoYG+p
jciDwYSdHU5N0HsqcMmNWmIagWkB1vE5kFR/+szu50lgDLSH4qmKFG20qPQQgGG5
CWOsKtTjvHDOYRxUD6oDpDs4U14WstcSB13MTAPoH8wBYOYdTrooN7tHSKOem640
YqtCgVFFc2w0W54EgGIkjmCnx/8B89A8R/P8OZ/UnLLSnkHOYiD49uDLHoGYK6jH
lSewQ2n37MPtojMqciCzd8L2s2nyqmJuxcl/JqvoJlgG/tgMqEzwiPwfTbIEV1c5
09izAS4jSeLouiB/nfbOCqJ9sxYAmlnrwlOZm9r8f+jADSJbqFfmrXW4lpO5Igb2
R2XVFo5D7eT0KHg7YSeZIEmHR8cMhq/pxmh6bMfQ+1RtQUByp2EsRCDb53ACzmOH
5mK6oMJ7f8mzej4ZbLL/zqKDUutDaOROaQ9x95oEDKbE8n2Xw0nU9xjielMxdaly
sdhpnsYd2ZIapZqak+7asd16jXvzCYjZ1vEO+VODkjlfNp9fFgyEY1XfpQUUwK07
xx7iP7MFkIvkj3RkIdj/11E4qW/GufG3M480uvoBT9GpBkjiGvFz0hiOpBOey/AX
t8A/CmRofZCSFNrQSEWVsG4PX49VF2jg7I8GuZxS5ogAH2lSw/4gQDWLCOsNc5zP
F8W32YlGxowlk1uGE7IaDEF7voT205tlN/c/2V5Xr6XrSHSC9u57iySFn6ryCAKT
nSde/AQ1XhkGaSkraA/uAw==
`pragma protect end_protected
