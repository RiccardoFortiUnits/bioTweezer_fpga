`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hamrFBWtHURnruRgAF35EzJJ0JC6+fFFvLKEyRZtoR5PaBTl5KXdd213WIi79yW/
nbPLHY/mQSbj/bk9OtJEdY7+sejvG5UY+QiQsaBHQNgpf/wLe0mX7T1tw3hfuNi0
gFi07sGk69muKc99jqZbp+NdK7uuMfbuRENQZmoRgHg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22912)
YuEjiKHu9qr+fSp8sWf9GUCU5ZNUkzWP45mmZ1vx+SV/RqbaxSlqzZgL1EHFI0x5
hBFVzEIEcYur6cVxHuu5023uWq8DSmM5QR/ZDQ5moHzw4TLMW3B5K4F5TLpjw/zg
0IcKhtyQyRigxrshyaepuH25Ui9roUsNbliBhqklU8umbcPecdJVioG63qNyfzVh
PZrFQIwLaeJY5d06RkpO3/mHZ73Q7f7Gki/ddPxJbVCEzmehsCZyT4jXDSmel9QX
o7jqBOyN6hS54HHhEyun0nTq5iCbwd8uD1yA+r1JFxTyMILvnPg6I+LryFjbSaCh
INWKqet5lgvdbBexQjuISvjxCL8OdPOal0vXE4lFTB05HJh/ksisWSXUid9jEEzE
N9Y1rgCU3ziHPGM6Y/esqEKEFkq3bMiIYBM/BHfAMoyY3H6ebKPF+24cVf6tGMIu
TNz73ZPwdi2FVJgU2/gMUWRzi7PNz9TSryzCR06JZ5zugoVi/ufRNuXG7IQlbW1w
2vaigPWxhLKkdOXRb5mEKj7k1+QG6KSmow6d/B+oWQzsU4QnJmyIP1GdNqXSiZlO
eROkL8P1OzL3CJMo1RUKLYi1quB6vGE2ks18doOeb5cX6G2C3CKCJkOce+GBH8Ny
VSK19vP1iSXqyI5F4o9GgONPSPu84XEtO4JjSGyoo3FKG++VTLZG33+zOuFaarC4
5rx9LtKQiwA8xlMJXKzFqI9xwAVdPJaiJp+sPxBdUGwe8Rzk8PKZhNQvtlXrfzIy
+lCcIeq4A+VjCt46wgARPKlTKh2QJt0lbUqAyle0vG2OIBgaj84BNwAcxfCuHm9S
FEnqnXtTUcGhswUhvoaCjuryES40Sicbhp6cjdmRGCesFQulsyU+4no1dQp3SabW
GiFVIZ71qVXrm0cWe82VsI5YFXldQHlzes294afwp1frHV7K0F0Q6LmLrR3ZRWeG
fx25xtXQUFDH1QZoGLDYUd7y4fY1ErXcobCwFD9wFDhQiriJCco1/w3lw3KXV5FQ
k5o7lSK2be5vJPr0HsM7sMO/w9Rk8AJiKaChGdffamHk+PidMxUL9SDAYQdUNBA5
Wuu+eSSrq/2NQtVlqa7QZA6mLwy/RBDJ9GX7jjMIfMb85tIQNibwzs7/qAaGHIzT
41OcBoYso5A1F7mUItFI2+1Mj9PL3wTC1hSV8puW51Ao0PSW7pZs47xJwCW1ZweM
hYezA2gXHbH5ThgvChEgdE6ZyYiloymZCAYGPCB05wkIhLKMJaUZO5jH+rglWDra
yu/49c7NyK0uTOf1EXos8X/DYiwvxtbMplYS7BVbqILNIJSiw/wNpT8A19RniEmS
FLm/QJzLWzkOZ6EDe9+Qj2HgsXVNj/tAMsZEVaStElWtaws/DZSt0em2iHihiTvH
oBO3XSY7oXKuowZzpTaCfeckI9Qg8HSB3uqwOLp/rQg6o8m1xjSsepTr3LWZou95
+1IsyxqZf2jqtpo+dcoBhCd1/OO57ctbfFjlheYcdFKfDz9ByK3EXSCFbFzA56CZ
B4BRWdlrz/dIco0YbkWDwkNSfpkIfPc217tBvcFw4Q+2zTPGwIOSbfel4v6jFaWX
Tra0PpZNiEsQ7GUKpEK13rg98QxpYCpSvCfpYyQq04COI7Hx+vTBDhnoue4VbBoR
TIMOibjV8sF04lmVEQYiWR0URaIvK3N6D5nnvo0IFgrqEe6Zbx1LQAD5rQt7+naw
H8WCMZ109VWKuke+E6fK/E0X2GQfxD+uKdIHxfn8/xka5/7YbNDx9NsSPVEe//bD
bCsXGqgGmDLm4koIM6U/cx/X7ZyOym3axb29I9jyHcu5dIrwNLWRF+/PEG0c2qB7
X1jPPv86EMeXuwwNARjXWCKu/XzQV4wt6PuZL3Ty535kakHOVYKsN/H92Jt5I1Dn
qlcWuGtvqTXfWdEHZoTmBx7SdxkguM5fIOYJ6b39dqGSYssGoOwj47EjkfJrCq4s
LqSbPrT1JNeeMeBAz/FQ9ETikrgFRJuYodkArrZ9yr6xAki7RCwG8pduduClCuN8
LLhQ5TiLKe7uYL9icvCMo4N6O09L8vt2TOiA2cPHGPGYWWe6kBZOKf8733ZErOU+
k6NF5x7ZoxvgibM3oNp4w0m1K6a8g2aYCA8XNjw4qJ7V51SGeA12MBUrWzXs8R3I
L46W7BomMRgZbLv8i9IrdbF5hKQeH2PCgVYthRLbhmo9xK/9UuYuDOHE1f3mzv31
e+9v6H34Jzm44U+1MjTh1h0VsMLjH8IdNIYCCNlm3+L9rqjIOOQH2G0s+cNKK4Ml
6iY7IvEHtNXrssN4WD5un7fW43tOrb7XCOj68ZOdNEVZ/fQea5jpLy3+1BmbGKcU
HFXSq8jgREogNKBBQJLwE5KCH6jWLEx8zlW5sKKiErXGYjfISY59Lhg+E+GW+HMp
rPzbO9xyB021FbhoNqa/EYOUv0Vp6f23IAInuhMRTrlQsAQyV0drnTtTR8mptJ4G
FsJJ5ZAnCPEW24/DEsBID9Ru+tx/fDsD93/skMpa/Lf1kAoGx4/jIFRGxNzh/Rcm
gxZXBOn9m/cEr76Nm9hyJwmcApp5GDjwB0Dw7nZ7fH6Yv03KivVqol2DwQcYiucc
yVR6QerJq9L9WCUoXpTlstKK7vnRSTCxX1OdSynmqzfjkncE3+gbCpHETG+nSER5
vFXmtKeQ5X30GV8Ib1dfwzbs72IGBPSAqGTsqP5Hu7cBQVe9FPwnQFMvxSgohn9O
eeG9ciyF92tpAOqT1EoByFoNIo7kOQ4Z9mAy8Cra9X4MzMl0RCOiMsRrXoQAIr2y
YVaYoTlkzjDQ3ns8XQxx2lmfdR9GOAGfGDUG2S3TdiiuSVaSaKMl01RioMHOzYwI
8jXhhIrHp5nPdr0AnorLpZi3GMGCV0yQEi2YIn+OHCaSswhUx/FqzBqJFNdKAawE
dmP+vvuMgAusrt2hDQAqESaAV+gtc3DREEpLuI95YMZkYQyJoDbAtzxY4sJ79C4j
QC8NoMyqgrXMpI+CxWBxx/9IMYd1SYpkBewwlv73yAzr9XXBqNQ10p9sxNcvX8e8
aUVxAHyC9qkHZDQ/84nRWurrYcDjxQyhC3Yfa+FV15yY07wSJG+8cR0KOzBKzXlW
xXmCmkhRojOUvuFvj7vZYrllRcGLFeyasDsZkJlsc5noWbSpg+ZgdwqA4CLg0vwo
z0YpDnnie2HjJD9puthaj9V6UuIoYO1Y57B2z/UnouuXvH1XICgxL3Qt2INMP7Ys
3ZWpRWLIDjxozQ9QTl2/BUnL+rBbhaKky3yWT3G8XVp+4MwmA0idSWP5SlMUQmlB
977bLghqMJAiaE8sbq8n98YhMj/uMwTtdpHhk/U135OK95i9M4NKztkisrMr/85t
eO/RjfyihkCj4gbsFcwqaf2fhIUt3TyQoQbwmPdJpJR/1bXXaNwqTBWEYO9kKzYQ
QsaEa6oy+9kgn5l1ptBEzqOo0pliRu5y/BTuWfrg0YfYXGo6lAaRLfd9XO8Bv26r
/sp/b9SEurPS1JtrIMfcYsly8WTqlgzwraEQ0sLJd3jX9xhQwFZm7RUA3L9JfpcN
SMBXBsl38jufTJHmSFQ97ifCDQw0ob91kkeaSwUsmwcObJKg2byafCU3tAoGg6X6
vO1dfMIpVL3b6A78fwELw5g/ZUHgxxyZNQ8Yo7frN/1zqqH3OkOoyVxFoK3SOidk
1N9xqJGN9Ep/TpQ+pi5pQUzuXgUXi5NnfFkuC7dPES+/JS9SleHr/T7amxoY8siZ
VD/WEFS91YdiUpjeu1qK1J/0Uho0bfD9IJ+J39PiffrNHMO/unH7B0PjxtO+WzvT
COuS9pW0Cy6XSwK3Vf4q834cG64uDVqyaKwyU++oJeDv2dDTELc7zkqawbuiumN5
+XC0tdfUoUbXCF8pdiu0vte8XXcXO3NpX0XpS8b7E4XfTtfZcz8grK6Ad+oVw28l
mSTg1YO02uBJoRHEkxAM9Ii7xnK44G16TKNf1GEm1pQF9BbiwUrkIdx/mmnp3OMo
pstS6cendXfMEvs6AYUxApafnA+lv8rnZ94Fh5Mx1KCW3Mit8/4rAIYJM/OjB8er
AlCd0sQN3nsJaqA4UB5tOFI+wbiM9T3blocLcl+DW7eBGGt157Y1YDDL6WpJhgjx
9w6e0e5by9zE+N5Og44kqf1qUPugcKRZ50pw7bmjyYp/n/xu3VeKQAjB7np7HtkR
Z4mcrlGu07y3bsZop86ileCfw/nDgR8fySiK06rVjI8+6qMWGgCyL7ZYW9ZRPQ9+
b9FUahdnHNeVyI5VI8giItMkqrl0Oc5qNUNmHWsAhivGgF45n01GPzMzUBLmeuMp
sXKu7bf0fkYsOoHxoDPDmdnxDbHGJ/oMfODWpkVt5IETwzLIniNHIbJ+Ve0jzcF0
H4HE0L9u4mQe9yYphWf4mn9jrdn+wyGvsJ16grGTZeRtmnje+CXFfV0A7vgMNIgL
z7g6yIv+j7yLmWr3APuDLsLVf1D3HeGaiiAlq3gzYZaGACTUmaEqVirdeGH4eLIU
jU/6BQ6RdTqT8g0QkX/GgwXrgdS/B0TyK6Z7HieTiZl++Lu/xGLvY4hWzZEanF1z
X9DUjDG9nv8kHxWtFUpfHhkvLOnsti8I9iwfEiIaX2d+n7XKnEHqyLXUnJQ7h5ro
7I9gYKhWhLxK0GGM7brIuKOAEJC+YeQkK0UKG0R/IP6sogo0k8w/2C16vCH92IT7
X03/bkdgxEbmO3mYzZmfZcFhtR5nDBNtKki1XifItmLg7l5IO3VWpWshxWoCn9Wc
8VJdVNErcTlIdw45DHpmay0OZ+iCNkbgxBBZRf5Xn9i0cBADEegZ1x0/KwMRg2rE
DyQpw/mH7Hwi5lyASkR7v55Egws9/p4ph+i7RCTrpQk9mBVCz1xWj0dABXFaAVk2
YvH3C7rgXsOTBQEvY60Kho9UW2fcY0lse01VHHr5eYUgVQsv4q9+irWXGxVLaN3k
4PbMaBvOcr/rQfKi/DyLMYNNqJcgqdH4A3jeSxUHYdkCf8BFj60x/RJzAcWq+nIS
M5aKoI/aGgQUTmJ90zns12Jc0TEKIgZXWo58yuAQekdZkyyKGaDTLAVRXme1J95Q
6ANm1eW0C+9nCJgzH8GBQ9gDIND9FGusc6kLVTrqdzLoOMbnDf9N94LFlJfmdU4P
TMbEiQzHY1/ORJUgIj4lp+m08ag9LSEaU4LDXPf6hxBwi31we6M5kq3XiaFG0RVX
VHaQ12xMVxXEyoo0ra40QpZSGkX/CkczWtpG+MSgSIhNlAdRlxQ8mKDiZK59ij4L
cEzNKJerDV6iFVGpvkL27wyx6UdDTVpNKKU+FNRAexzC0kMyTClDcTookFEw6/o1
yXZBtR7YjyQrJ+tgSO0t8mwFkc+6VKb4o9Wp0PagtkFNXX0F90qwu7G6wUGiChda
3HTqrXnHsbKfosrnazTSpfsUc+cvrFi3WC9uFvupb9ulyjvA1fFBsxLSWROoOebH
SCELirxSEksM4bSaO/k7M9MHUvKR6yUUS7xV5q9+Pc5fnYfNe6xYRcDlkPRAMy52
YZiOsoeb8sv4b4vvG+meNxSSPoDQi5JL+HfsWXkr7qdle3SI2Kqx8vfkd43sSZgB
PDIFG+6hiIVsICwiaZBlpBE1O6yhMfZlbGxb9EEmnqkllAZ9A/u9D04Jo/Mv4Vxg
E8MYEKfBw058sC1mLU74Ljb3vjgrPv+x7P6fncmeSRgymBIjnwu5t7vHtivv+YyY
1GGEJtlBpy0p8GAgMUqju9mJFpUOhow5jqkj70Ng6Q0jcfux7h6OZcWt1VTh98MV
if1oY+BReK1ASYwUc668eQ46nkH+NW7J5CISc0/H5e7L5fbXEDm51cxAjRLD+GQW
0YuHAvXGrApGPIgb6E6KdiMQ43npI2/WhH6aW0Mv0pQOumpgLXQ3EUCw780IpCrl
3ZUNhGFNPlk7inDP3SJVE/rmiC/66wHK9UUzVPw28t/VopcC8b/Pxtd+7bZS0AgP
jooW/DYt57DUoZmX0jNZAQM0Apo28sXTibz8JO/M3xw1scqt2v3tfc0BM1C0biWt
HIu+eyFM/pUk/P69nv6qp9/Tqunh5LCayO+DySJZO823uDXKkVCND/WBRG1kgxhc
xlJL6jCmv6jp09vrakzRjg3KiMhJD5aYAzIvtSlM4t5lc7mXzugBz2/koubkwjvg
tWF4QD65EnlBz3vmP+GN9Q8FiIjtyL/U/RMRdqaUckKEZ1t7Bo1LEtvvfdAGrJ8U
T5jg7JrjI9M0JIxletDgLFj2DtKkyQkqJZTdLKEUBNYSa81aIReix57H4zqWk9He
QRE72zfG+Zwfm0fvFXm+HErWW4oc0mM/mcBzbAeH4+XwPH9WWpLCdhcNkliaxdoZ
w3oqxTMnNqPFBhbXKOZCfIBOrn/aO4aMzT1PpfSphDZHN5GxkVdzMysCjwg+M08+
FcFKIpC8rD0dZ0dRyTJpnhb7u3wYS0AgvcGLi1WZzcI5m4r83IghLghsqxjULyAO
0TMQ711BNGL++smCTez0i5AmNhKLqfez34IpAtpXijGVRJ2d9qHZuoAzo63aHCmJ
Vx3ly/gY0WCFrB4W2fpNoqRF6fynHggZGl3eYvmBwZNvlWeSBDcwqYZhYRsl/k+Z
MRqB5aP/kxA3b98hkbjbzGIiZ6OLeAz9H9sa60CLbLo8+G1H1G75OyTYQcgSnsFe
ruxHGOoMQajEeNeFuaQy9n+wWm242lXkwdDClWS6zu1gU93VP5X3ZbMjcmQHo8hJ
WIaA9/13Ozr5O7KDFLC1AOjcJ+XvUE6C9zOqBFFGaC9QvXqy1q00PzFgMGYObQ98
XVLGHPUQKAjJs5id0MT1oeJccdwOBTH4srYfMyFFqsICeDodDqNBw1ARPAi+pahB
arYZU3R3eEyRIubj3B+4vwN9G1zJ6p9lUJrx8xw1KeWSO5vkRipxJKip1fvCrWJo
1RjZe1WiK+DoOEfY4NGLdTFGvp8/a5/BxqKArdvR06P6Ck2IjN63Sx0xSyLnGPb5
aoWdU1UYFC1n6i0da2uhum4+/G7zqN5vrdcwDmqnUYHd1sElhIOpo3cWR+sFVXC6
GDvfn64nDGYQfJ607iOg9tO3nIx/Yq04sNLbkWn445OhNMpbaGZuEye4bvQF1dEg
2EpVO0FahlYxUzAqFLvSK4ZXFzzuOO61MPvnLgJ2PMeEE5xqDqaeh0BhsyLzicUz
Rm4zcsgaowilMjfEmBRTKg5PMQC02hCqlhPgFRP3RkdkEJ0QzGsSKBs94Q7/Tfx8
liwPFA14wWb9vhXrqOPOulL55kExfepKWWx0oJPn7ZIhkDX577gmY9UXVXtpfSl+
NQ/P+/Q1g/OZwv3kSMLdqbF54lKKaLOyAj5tTjzyDPPsSwMSFbgu20d+gl9frVPR
dhe6AeO2JW+BWlOPe7lVzldyzQHWbyRTcvL5AxgAb0GVIPgzD65Te9kSaR9Mf4iU
sKNvkCiBdAEgaCBYnp1+kQJPRhIJFElpTHV2sTVLMU2DW33QR6Ch4mYyoZAltilR
czJ/HaZDjdmiLsN2IqV7mKjv7o3rpC1qmfmiAjYNbJQweVYZzBxyLra5RZVLtWAJ
WLs3CCJtIuqLxkWLQHkjLFWinnZAn84CL0qB10bePY2sQScLmd4AZMjhRrcVIJtc
VAfFE0ssEAsw1erd36v/5uC5G4xEquWhv0cGqX/F2q+iImEuNEOJE8Ho4HQ46wKr
csmq5sq3Nc1m8dSsmwUrCml+jlgjb4BG7MFj4l+8LX3dsiqhlJYNACFxIVbqQ9jn
Ldl9NCSGx+PUMgs9NM9kqoqqauC0ad7vdswYgzIBY9v/sXdcN5NxYisoypAQ0Z0v
aETQ3LL5q6mNLpFJqSHaqlz+Xy4qm62KB2GuN039PZLDMTaA6xfHVA+qg2WXdSXv
pKABvpP9qIq8Chr7rbrQ9p28m8A1m7k6mmdL6rLq6mEBLp8UGkJg8ZLd7xC3/aBR
Bu8a8RqYehApdOTjJYPHbxdik4cq/DNzYhSZE+19iCIOT4s1wBV4Fdn1RKVhNaad
dbAk4FoJ56lAhQBOZKxu1OuTCxHRwoxImVhVSNL9OiaAIu2kjworS1Th5YK/xukI
aLF63x0eSaghPZMK/b5dvV2ENNcGEfYosElWtWS54Dq64MADJlEMXdXX+ccTDhZ7
7muvXjji9NQI8Ql0oo1hj4O3jaoqFnKNeB08LvBDkcG7yJvAwHEtDxmjgoOI7gg6
8BlZfN2mrLZy+gh/3HwImrkXCdVaJXS8vJs18Zxfm8ie3tc7KTZI0zN7tsDbRbwp
3HyZZHFstF5Vnt8ktqOHkbVhkfxLUnmrNDfvzAa02An53SiU8Al7HygpRwTgV0Jl
d+6umWUsg8sU9Lh178r2AdwumZLpJy9uYUMH7sXZKZmnPRABlTv3qZVJnhHzc6Xk
1t2zTmY9KYJIElaMVPGOUyfJMm6YRIo12VYAIsL/g1zy3scPZoEwNbdX0Tw5PElm
Syfth2NPgTDdvO1B3XlNbVhW5HsfK2QtOaOlFG6Xhe7IuzJ6lJ3VKSM5JG85JWr0
I7TbYWfjl6MquwJv1c7RL3YHAQ2AwNFRMZG/NmiBbEgDay6nQ5Va1jMF38+PcT3K
0JxZAxqOklUE52ORbt9oFDUXqmIrEEiOrXH3fpb2MKFjckKMM6cY7noM2XisPzA7
v65d9gBpvc9R2CtAQkFWqUgVe5EtlddvG+I58d4rw1txI8Wm6XET2+qVQwFF2CjS
GcR3uRqeWK7SbIHvlqF3NtynS2dpKkAOhWW4FGXBYcyoK2tojPltRWj+I1SnaN3X
YgQQMgW6j2nJOpuTuQB/nCDtW85UINdBBRlURlnWcYo/Y8NC+93jLTHvZiDhyQou
8XB2sjRXk8L7FMFtRp8KzMP6KRKM5Pa+rDaKABCWj9OiZj/OWZyfItp7DcHLjTX9
ZpUxaIplFZSCd2JiYqA+VcZUm8MwdclW3rbVRsvukbTtO5hNWUjJbnWJ0mMPmjo2
Va5Sczt4CPj2xHeas8F4iexY42pESRoLMNYBgQ0h2y0pG3MQh8kMDaz0nCzCItnT
o1gx2MuVhHqd4Z6NlLDquADQpEwBZMNh6Ulq9rv3dmsyBOim2G+u1TyMY2ZTXvds
QsJkjfGGFC6eL73yj3bu2ZxJ+4NZBRn/k5wcgH90HwSiFewfJWr3yNSpdR2C6rTp
K+f2j2DKVFqpWfWXXKR/TB0VY/pOBEZV2hjEDuheuqbvMa7Oy6H+FENMYjDAGo6r
r7Rg/2q4WpvBFU+5KjKO06nDrXH83+7BOA7gI7p45ft5+gdy2UOi1qjd/hqW0p5Z
OJeSqUNuLupomdhqBqw/k/mW7SfUdmdPBx2zi823OGNhJN+wLLUA2fJke0D/7Zdu
Q5GecNwgFrsAwdlffxZwi9iTTlOX2YobfWMUDZfYjgCfxalnM62w37M4GMwrI5hj
V00ANcm6KGNRfoPeSantPW7vFDwVrf/xZnWaxadtl0vTqXXInUWJ1q9wj0VJlasN
USZSr3QoPc/BcK9vSFZ22EYX/KF9B7DY2mSorB4MAHK/zhfVCIiA4BQXkogU7EMe
ukjTzpPuBO0vapqP//yYMKcsY6vrlgPBNwD1WDWL/gbHq8CreYc3pxT6Ts21W14i
b5r99gjUiEWvEteiXCQtT3k7i+QF9E3rNmVieVJSV1lC/HHbpf416jyKF1d68P/e
NGSXOwHE9o9gp/JA7O+D68k2TSbyiKmAKC539RfGGk0gqEOrU4W1B113Y5FPLEJV
ejFxfd1PiJSBzUwSjCHxZ3vZxuoSfo6nTAmr2kDd2P0JF2TkC1CrfkvUmLMmVbur
PTpEvc/SdONoXsTQkqVUeHGfXFForxW2oxQmFD3eJVIGLy2oDpvuhLHVyNQSF6Qy
Kx6fMEUEmHRtgTseEbQIb1ZVZyR8Ce6VIBvXIBOWhzGqTSZ8t2RxxQZ+DmuTAhag
t2qa7GV9hpVjhYFNe98nfKSu+fmZex6/FEfarsB5nyhrb1OrVfjgDOoffkDDDiPD
h8Co2TW+VvEQ1OcSj3GJj12dQ9Anpjgb5wzetSaGyOXv9lBfkTxJNxmRSSiartKs
/h968skcdyqkPmSkMhflehXwZus/RFcwAZ68qpIHJbrqLe/IUWe6EBJ2YgFwsfyg
TTnAOrK4qs1Yncs4/nZNDDZv2bcqD4B3kSSbX65hU/8VowN/DgiFSGnLuHOFgw3v
hvcfhiL7VpJXA5nijplr+VnTUmCaJtV9rjic5eyWQPRvzcViruxunVCDn3JiCOE/
kySHgRTmoqTjWarSjp4YkJxLLVFM13F0KqvFQ3d5RlVHbfd2WlBCw04mM5IwplIK
xiK/vPI+5jHBZ6VYNgYp4LlrBftnmj2GJwMc4diRGrFzTYQ/vH4x32Tg3ndcgQ2Q
aJk5jnuq0ucRmc0OF5NypQKUb47kp+Ra38t4dbf4KSiZv1omBhuDxHyBaSsB1z7e
3b0b12zQxk/0InYhuT6XVYQFgFmtEX4U01HWeuTvYo0lmZB33mm9BRg8sUdku6HF
ImyfvccK9tZ1vyvZUZSGHfLSnCEm0co02yHENEI+OLn5hWjtY1chbDNDp5GIHnB5
t7ktySkQ3sH3LnAC892vudi+BoMwnp7vFZ20Sw7Wl/M3eY8sozgmjQSZmaNG92cN
PcDElLDITXa0MTJECogty3umNtZDzK+V4EZGkyJQQtFnuBQNqHTO9Y9FNqpUMIm4
f3Z9WGwFTcyIpDQ0Qvefl0LyEaUWoKuqRyCfGM9xD+VyDMV/818HvLcHHdCbA0JQ
xwXC8CiOMynrTGB97GJD43NPqsMqUTEJw5ndDr2rHQvRWzpe1NEHvQrgXfHzoh1N
guZtPUk3GVTSzzUsnnwt/4vj2DrYvQTrEy4spnbUav2EIPPPfqwHcXPZABcGW1u7
66Z4aPWUDXkC4R5mkwvZtOmECSBtCPguwiNsil27hMf4YJjA5X1KG7rpG4pQEWJX
L6XK1fhTObW4UpnZq7r7GBtWM7pCEu2xR6dveYyx04H3oDm/fyAz3G3cIIH1YAXZ
/3GhGxGVuaenLn3v6VUXRWTwkfrKNBXL9flYKWh26EGBT94Jl0y7iH6YCoqfEQPA
viff40fWmFGdkFKlFpXjNC1AzELRFuoRHtJ9dtH21TIyd0cKc4eZrR+FDCyA3cO9
fJPoUv5HwepJ7K6/krlIU/lH5epdp1OAv9zE786hViC1VOGCvWB+zekC3hmSUx/i
rxfoDrhRTtfX6y9J3qzgGLCR8SZXOHJOUolY42flc5FrME97eLa9B7VVbpTk/LpG
di4n1R+umG/J+4Q5ngXfhvg2ej/yPqnOY2oveGkxnZyIZoaxT0G8CuAA6Ph/30LY
LaqYNpPxX0H/JdiRp2QZngPROkoAJB78i1hBhmnp1YvBQaZulo/JuswpXB629AaS
kRg0MGYeloEG8UD2s9t5LLjcJPx0UXp3+N45S84M9DomIPptC+HcjTtxDxwEc8Gn
/WiSZF3JkcdnEV15CpInoN/Jb/LzzrFL2BtTFFAoi2+W7M1t3Zwqn9vYkbeoCF29
aer+M0eEhk2ntwDT2XOHZpmVwKddIWLJaCJYhUIMLj8CmDcTjskvasaIkQP5e4ZB
ZFf01Wu/MbRSRX3e4vz2DQT2GVFwdvY69E/uS/WzeaxOI0+5aQWPxRlu0AB8tVBy
plmtFkSCAxOmhAACXkBgqFHt+2Y+Tls8N3oOCWVXRPzegtXUdqfwahOz0djCFkaM
MiT16m5NIIBnVIa1SQC+Sx1NxptiR+HaeccX2jr0ikObQhpczmcXr25/7KOHL2Kt
haGQo2TkFq/mfLXH8ugbjHaxlIaVkMYWpPmrQo78GMkkpRHVserLQgxEcoh7W64Q
oPvAn7le6O2lWTY/0zesgYy73wVKgOHzbr/Xp+5Aww2q02RmN+8lIYcT2Y4ucV5z
wjzow/9Fjd4iUu6cpZRnkH7fODfzvs7+9jKmady6yM2cL1O2PjPxuRHEr7CvTr/k
mVM73jvWsaCDUKchIkSEmUJaVzhBBQbB2poCGL898eb+pyhuylHPl+/yd5dVTesM
NNMlfybVMbigIZ7HRSrKEU2Qw68oTQV6V61Odc5+KCvPE5gN4mxrbOy5Jry9wkDS
/oBRWoRcyz2o5w+r43qgniFyzpr9cSklbZ1GB60bvyr1yyYa38ItqtqwPD2hkiWn
K7F+mCNseh7+JYcrJ6R1eg59gBUlVeta8OU3E3DCmjc4EEH2zck2jaKiFYi4jDNq
xaE7M46EJWsjuDfhbFQgrJOF4kOEBY4o7l6OX4e2tBGYOaVOKSXkESJZtC+vw2IS
yrfff6EmHKbP21XSHmcfrhWDWYoFZ6Wt1hW9UHMOkjEMwTyqn8UaNDEYCP1BNPcq
tUCYII9qM4xLCSrHY+a0G42xPSPWEolX/l5Evc282lMaGro4MCdgEx0wrEP+baAh
8H71bVseA2U32WyplAGOkh9koiX6KZlk80cQNg34xnp+TpTTjOmBIIQCsSlj4xtb
m9IIEHnhzHKGIlvwmwqNgiQR+X9CkvjDHsnicn6D6KpBwj1EkQ8D8IymFEfxCjbG
GZJIkLjau9npaK/bCXIYdf5GTOJOlKgrHeSOJU0PIzgFsOSyQKURUvij19uZ97jY
fKn2s7Vd4PPidJ7YMUZhkt5PNceajvyauvZQwywzu52dhsqJYbFAkKsGTArWjIo8
Sa8aBF9yr2e0hUv0jYXLB55TZLM6XxMUhszh949x60gfvBdX0UoPZkduiOXmF8l8
k9By4EAfrOw+IJcN2VwBsXKLPK3hSMAkOVqVGoWWEPRN9UaaRzFMMZHNEnTWhHRL
SfBR+bva1oJl9ZNbPgUTxb/gUKIU8Nd/IDKJQf8/5YRoZbdh7ldSI5lFHkezM7mn
K/Vr3Kx2aDmdZ7r/fCUzOz4KDQw9WpqyvgnQkTL4VCfr1UehLOU7lRNneR3bANAh
/kt/LS3kLbADVlzyGM5Xj3vxstv5ynXlY+blsbwuYvtA2vrzibwqmSJRFbx4MlS7
nYo5/MREJh4MtPDKiyvyj3gBgWiiimVYokl6M0HWbD4GsZ9PzQb7HdfKPVf0zD18
iXz+GAsX7ojvSn3/6xGtwXYfS7u3RO4LZsat6oQrEbT6Mwb447RJ/64iRH1ZfeKv
wDzNDQgGilDNFtClWCkMS358VBWwcoXSVzn3i6patX5BD7A8opmiWtULM/oErp4C
HLEmd+3JhgSMXZQSjtqStk4K4H+DVVP7h4yroVYI3ZkrBlAm4p7wo2vQ7W0op8aq
saz/0JLHuCwAMwvHvym0Ex3DiFF+H5w2ajm3ZjJfBzoJAkE45FUx8veH3XZGzRBY
VKlkuHx1Zppft/TmlU5co3TQmubdMLXs19g1zmnBk7sIpK4+hnt3CfezngyY2+xI
n9UJEy2d3BVtTPbJL/zNxDuzn5Tis+tCgw+TbA1khU0wncYv6fwMIpeKB16eZYf+
KAU/r+bVe95bxpzwybEcOgQUACKJ8JVLgA/by72mxuNEbM27NSTmYu1PSYar5Kyo
cL+p52vIntpPQ4ZpKg/qdYANfFVBWojb979E7BQiDaeccZ8tjVHx0+V2RjHnedTU
d51ZrS7/Z4RROHxgcKDnrJR8+UkKX9kARpYgfLbjq3A8St25SECxiWBj7+4HoqQU
eHiyk8tO/dpPAOS1E9seYjYY6+LdOs43xwVfgFuTokR91mpWMhHEx8fJ1pJgqBRA
0bAnGKLP7ger7tEPw/7BomYOCvBMbA/KwqYB29R56v0KI/NS4r4hjr+6S43Aam5d
ZoxSbLWPx6xSot3UCXa7pciObJeInuTfy0m0eOUz+L6zpA0hBkzeqDvERftI9+DR
iURaHDZtVHAkIxHdFifMXU2kxVRFl19UuVXCNw1foidOmR7krUBiChkNxg3pRJE+
v8tTPlBY7BziEnp8x55JRWuDnnImwzPOfd2iCQ4aKwXIJYeHes8EqndLAw2S0mOH
U40cfqDwixb5fUS6+wAePP/juy3dplWGwJb4N7hFlVeA1EqQXtHGDkoXctFRQSnf
2PkSkSFjn0cKajmS3XBxjsiAfdhA7zxBiCbQ0ECQB1h9jFExxIL88lVYmBq7CJnd
mVsswCSRdnUx4xD7l5pvnhV2q9ucKcf/9MIt00OE06Ebvs0xo+wciXEDEX3B2J7s
OfAZMWPluzLKqPpijejPNXOLbh69uzF/yF1Hj+01SZpDaRZzthbegQyB+2fEzpMa
sTBBt1NKesg5L/iujuecAm/VvDqhGBl55RplNynPZKi4C2MB2jIPVgMJ6O5TkChR
92W8ddwYSjfg5lX+zYdbHMpmHDtYmFEffU3AL7AxBYyRHzyGb6znuE1x6L3Lc/s7
WBlmsOsnzmOqWQW5865XTQ4hAXvvtZrFjgElAufzk2s2RpxmpU3kg1Lr0Use2jrw
E3OVf904zNcUchLpM8Kq+kQsFOvEZE7Q/XfzPg5c+Y1fEXtzQXpVfdV2P6VVp0zX
OcQMvO1R8YcVgqPNB86EYPVCnLWbfOfHSubAmvsPNbCiWML5NZS+25ha6DArXDrU
hxGTg9c2VDaNzQlOcCgiRATfNAXWs1mOhx4olqgazaaV6+nvVTer+VVaVOxfcQxc
8ARcNkFSt0aZR0fwOn+r/iRu7V47wAWQojBMh5a0Uvla8CdwTdMsQAl+NqSVc2Be
jgcmNNjprMReohBJlXh6cIZnctDvnyDFF6/pUT5IzGoVX1XoYqrdjLDEMRkZQH1R
WYjn6kJk9EgR4wW7A3heBDg4WvAkBleGtm7BujM1InPfL8t59YDVzfCcCLIfSfOo
rctS/uvX/6kkq6G8zvSvZENAvVaJq+gZQkcEk8JsmV4jKlT1ENLvLRn+kwdxJ6el
aUk0yxeA8fTLjp+9oii1Yk12Pu1lfL5bbgNqGor0SirgMVl8axawSWHbh2gBtCvu
L9hWx0mmgiWQq60G9Cq1VJ4Hpl/+nD76o7UOjWGZUoNmdNyce3rqHaWOl/1iwD1X
jTjgDkZtSv0I18Qsg4vrjDMREuRX4d2OpQaYp2uKlFu9LtRVvle3GvBy23CWKvhd
aDlrxc0VA3hVv+mpKDlsnqJxPIjKzhI+X1DRMrBsjDcPPWWpb547R4/JjKgMiG8M
kwmurwBQDq90eKAVKv2GSXscfojGCh25RlydOQDCBS5EUfTnaxvb1qYgg5UjBowW
jYNRBvdNajDs2xfPtZPwa7oj/lvjkNv3HP9+aSMi7EzEuBZieb3xbm89GEEhvVMw
C3YsgvpCgjhMH8JZef5N9Gwc7Ko4gugZTHOyXTWkMwBLJ2th69VbPpkx3685IbNy
LAR9fDIk8zDgc620DBSlY5QXn5dLxKPPy/NSZNshf1tsMB4CtkEex4zp6umXiTEA
Gc5z7q2WtEeb4hmCuXEFVTIUJLWKEGp7EnJt6ImZgraLDyI//dU/dlkUBoBkFePI
kefcsOd6nHBv3+r9SReDxrGskpMPDV/8MM24Jft+NoOhgr0mPPQhvGvjcYIkydit
keAp9JVxTw9wxaAZDy4LLeCghJBuoXgReCvYsRZm18HhFfKcFEmUQhR+dtuEvcMv
dM65b5cRYApOyGmOcO16+n30eRpxRRUQEZsLpOAEqWctIwAw2WgwjXrq1z0HjCLo
bI0BgxAgl/ruhkN+bdrcrWsdTD7zzqTmrhDrRwtEtDD73h0UDXedNPMdSgza9/0f
yBteC/C2mW4FEHzvM3jCVypLTNc9kyf1T8/KGSLLbOI4j1rHb1XxJ/QqdcU5AuXd
PRYqU9qfS1DICBlcW+xGT1cam/jf4zY2mEN+ckR8pDADAuJDl7vl5k1kTkOaegRG
tJsAebThONGq1xct7K4lCZ5vAONK1hkchAW0iDmzuOzs+pPMyOsZryyKSTRC4ryq
tRZivNPm7bGrpAZHmMN10G6vtohOVqDeHpFdd7QlP7rk6EDDDYKsSFHWGJvoNVRG
Q8UvLq69HXaRrwZPl4Z13yq2Gyx/JDdj3koOiC3lTnSkTbuGfVqUaMZO2+X4eScg
/zV7Sz+Af7UjZ++MBS3cjUzXOpho0OO6aMYYAnvK589Zq0tWq71hiUYFXHh1UXAo
7XICmC1e0eD955lnFs4q0qv7Edp3u9wRDM0aJhKSMLiG9W0HPJBFejM+luQfCjPK
8t1kPQc7zQqhcehWBCKMfvgRB82Dr6JxFpcekmhX3/y37bHGgfii68oF7ZZoQG2v
I6vcM8dL69SpdA/LASa5RIEg5Dc5doSuYktkcURg1M1tXWZKtEsvzWYAKFF31zQH
xThk7Xkp8TufhAkdzyd93Jx6uSCzM3pf11suTXnZHLchfuIYgJ0ghVphvQaXZz91
jq/5xPWWShTvkFK6kID/fpcKjoUxkhntGyix51bpJyG3uL+MTiNANGAEplsFLrr1
M0ld5qLNiUIZtl+TYBHAT664RsP7PoO0J5giLOuHvucqbvCexW5700Jr4LYr8De7
gt6cCNwrc7nagoylbieGq3rA5nXPCDXRBrSFvGgvW3NdpWUBy+3FMeU/fJwmSUoW
6ZUklotruOFV8ceLLykNL7SQW0K3X9BKp6oAhyso2l9U6dvGZ8qmEiA6MmwzVU8c
CNHaPCx//WgL4EO0HyjDspo0QQ+Qv7boWAHkcVuigyR8XAOcUQIDhVw/Ar/OIy0i
M0xWNv63VgFUmELDiDqaR0BhG3RgGal9cvah8DYlKT+AF5kbw6/yiHI7Z70HNSoa
ZKHYGI/4Ap+Ua9XOeTanU3u6Jqel3AAhxeDt1a+ybyCKHHrf0ZrcJPg6LLMvoaWW
pFbxEOBjbFNhpmXfm08zrTrPC21Ik94ZTg+Qi64KEVJ0/YuFjYaAFKJKM/4KJ+GV
6N4yY7GM5478yd+wpqEnYw/+pAaCNrT+JqJYJKtVo7qg5KC6EbbE6SQHPbmvMx/1
Ioxfr47sHN3gzSLO9U2bApOEJfDyswnWf8PcAlUcyyAS2WnXHvI/PiJH+3pTJxWM
0uZNtJb5VhRCOoi9h98NlnMhPno/gsN+xdP+g/8r7bIUO5R/08W8yNy83XkDTgN9
RNKqw4RrqcJrtzCa0dYRedxJDSfYdiGAZcGj0AKkBtL+oVhzWj449bZEwvsApPC9
hxwGVqTJNn+YewboKpQmF84wxfSiUQAFDwUgh097tMUytZZWk4SxIHrUHpETrj8R
Etr2d+LLbZ+hKwghbWybedaWW6YUsRjOY7VtWFJvhOEWh7bg/dJzf/yUONYhzAIY
diwKLw2WHS3lZb48KQVM3hiDX27H7YFUfB5s1k0EATOaD5SKmD54zHWLehRSo632
tDXZubBjgeBiBlluIPzh4RPwlT7Ilp8q53b0JFiBpOaaj9msciErnqE0PFw7AkCw
jn/LgdltajEuM4ALWDgXcWs2nRlGAyvjZmBidAmw3Dsh+iGdQC2cExIKMDC+NTOh
42Nmvp3cVSyJYzVCzfbMUvOk2ktghKt7uXxOFuiocYNNTMCrVw++lTDDUXdtelzR
CJVRRHcYq6NFZJ2rNDy/wn8esBJLHMaDpHRskn0tSneM8KNJOQebkzzmDCZqqCXs
rWORKaPuXPeWgVTx+yqNKfgbpMgKpG6BNQW8BnCncaYy4hETKDTGRktzE3ab2htv
wTo6nXdfA/iHzF1PQ8KKYBTxsm55n3/Ut/jntzMbiL3D4KM1l1VBNuzyeP4vJsS7
GxYpJG9wErghk+9g1GsuDrtV8ZkuzpLyGH0/+wWI0YQYrn66rPLHzH4PNKTp94IM
+7B/xafAbwugaGZ6GWnNJKz3pE9g2FwlvzB7N1jI0xIuGgxmTewhS9nw1blNSOf5
nCC5DonlBffHfMTF2O1VklzWODF7gSlqMeTror4mEQ+Pp6r2NQb+DtThMjEGT+11
SC/6aq1ZXhS9G033L3Q2uGnlhVd5LUcjeUCORuLX3OkJ/kcu1rRAxyPJzJKbP6o+
9nnbIbDh4ln5xD/s8nVb5cX/HLeSwfgfCz64k4dcvKbuRV3QjatSbU53l5Qv3oH8
oK5NQGo+uoHj7WNWIbXTMdljQEOWJLq9WMjiayTScIdPVF11ddYKaMR0v2qIAJuC
nvmqkHWjQIetk9Gzp1BWqovNh+mWRnGzmvZWfGHz29dB9vHfgrWZjIcfXuk2CEm3
1MTJSruxCoRPaYg5bxnijLWALuHB9E6nm06Quu3RFcx/s5EYZ0Gg+FaVn9xLpMaJ
ZCFhdhHpcMCl+2hpAo/hJd9vshrNof73nUlLAGb1/qrRjIZ357KDMsWRFoXv4MAt
Djt0aQaWlXj4ySEF4B+KIk11tbkyWwpu6P0ozGzNvRNNaIVJIoekBf040CZtIIw0
TKyiPs7LHHSJ8hSeaz7Hx0ZHc7yZksmcVccrHj8abHkMorGKZ881ZVhtw4aQROwU
BS+C7yPaOvoUEnCXs8Bw73ZU4o+af5Vxh/uSCzhd7exqwQySwJkvNGbTNugESauU
At/5Xmt5ScXpoE4/szH2D0g5YampbIMHjdq2OreJoXvhVbbT50ptDGFkmqmPZhds
n9C9Hgp3KPRjq3iH/ejY8H+fiEp2hH8XjsRFshzZHzYhU83NBJI9whCtOv6BJxE3
Wxgq8l7ap2JKkihPuUD/fA11MGk07exTdKv72r1VQik/GpvphBaqMEO6P0+1C68G
tm1c7B81X3HH80nZNfMaiC5ro9q4wsy3VuHq6nS4sHir33eAUS25i4s5KLg5WOMN
aLL6mPS0a02iDRAhwy4Aj5N1suJYCf01OxJhndcNAEr4ugt2W6wJv8fFZCfggpBH
8gYjXqMe3wSV4Iwkz8j7wJfQuPGEdBTP7YcrivALVvHwWyoFZh6KDH6SIXsnRnA/
s0rdyiCmMqR629W0hwkuL6YEez1KyJFrpZC6Errn2Wghj059xsFx/BU+8AM6Fpg1
17Fp4S/ma9oWICEhJmJh+gesEI3slLkxbqCG3KLL/KGTelAZfIsj+JdcMkaEWCmZ
5kbZaTr/xT8eJl+urhvJ+4Li0K1qbQWKN7gMciERXVkwzs9c7POkbep1m+8tw7Gz
K8C22xqo4niIuZ65k2VRb89qXqYmptaxgThazAmBATZFJYSRWxqOan7ZVkAmOBii
0GaJilDxUKAUas/DA88FdmOru9Om4RusY/0TU2lkYCp2H7trUkb5dhDYi+r3PmNL
MKfo6S1hckGM01i5NQTggSAn4wZXRsfJq1uVjHGaA/o1S0kSuaYjkNkCF6LJPJzc
qqDRddF69Sh+qyGt2sl1IerOp/nonISSkIxyCIFXjLpzqqCZZ+OnAuLr4+qrXOJn
ey+lSlmjwNvqaPIF2myjHuUPGqOfGUDUrNibhRjdtRWEpUmE9GrEjgUWPx/NGgOs
TYfEB6Fmm58d3QKjohEzCCrzYM3BfX0O6XbslK6V1PVqnWgBbUzEzwXoIA5MS8p6
H7yRAWEUN9OFSLSSL07ec0JzOgIg1jJKhyElw+lAqo/97okWF7D16kFRg/LQ0UcE
x4EpU1xbdMjlWgRUAcdxmazX2B39pW4mI8fYy7FyBKAVC/iMLY42BSgYMErv3l9u
9hnGwJ1KQapB44kjAKQNSiKLZI2+yAQq5PEvJZCNeQlw1JHpnwqt7NKBZcD3n8va
bSpaTiauBmP7qhFL7Dmw9iU5Gq4T6JaP99XP7gzKgGXhxkWj9HUHajm9Sr6JDA3q
XJD1qG9RBvsWuAPAl0ZCxq9wgniyUaohpvZMlgi016CW/E1iVeZ7r41pkGYTjUh/
X6aM57zhVSSdRHUIFVA3/f3IzSiPCfoM3I3hqCRWyvfazamo7Ie/GKqDn6pKSUjS
RI5sIMdFJOlkSRXFn3LCqxp0raaQnLf5ANx4cnyzeUouOqSnufUEXRl7qmqqNaOZ
OJkjdOk0Tv6SBolROI91UdQZpL0noCD7FX2Z0LRdA/yA+2ZceC4SSW/cL9nIReQG
2pfSd3eGZVokgkEVP24UQBXgnvMm2Ryh1Ikpi92f2R0p2mpaOTofuJcut6gJy3ha
gdz9pV12SNn0fnqeT/xyzBih04wq46elWpV+8+5db1Vnuu4ax3xwbnCHGQyrtkev
yywfGMTUuZhNlJj2WsnkRH4HAeIPXDE6J6cMp9OvvR/8bYk6UqnsW1B7PmvcTmcZ
qF0/zt82Mx2LzazAU53WzisXRmEn1+JgdLBz1OAu2MTH/Q3DSp1RAr6TtPyf+Bej
6hgvNy+k3qEts8xEcuiEaxAruU3GL0igg6c34nktfFVABue24DRgizo9qHyGzSw4
qAwXNDEg54sWB+Gk34DiPpiiuEUVO1SSxGQihRI6Z0ju0Fg1ZiwxnMPLXLBnKiRv
JY17mS+FZUaa+O6acd8RV92p5sQfQgAwI/QlDGEoejq2k1vhYTOUyExx8/SHmQYk
u/zMMg3G2n3tHr581WKDj+q2CmwWNR6MhyB1/UEU+QYr73FYZxEHRLu6LvqZFY41
7wtyU1P/DR+dkuKUpeH13qQTLNyS9GXHjNfsp+blHnP/KBvIKb2hLYBjJABZvTbM
rd5F+KpyfAmNqxiLZt9uktUm1bmJJhIsN3owjFch/lOOkYUNNfvcZf2VzvK3UvR1
AvHbSoDBiop/XIEpm5ifizsjmHwOo5L+r2rVe54ccjhCdzcHZuI9GwRhcTF47fRf
iCNf3pRQuII07n5matEupxCvcQevVZLdcBPJXgPXWE74LwytzIgB42IVjpoU9KoW
skkU1ZCNBxQc1nJfpxQ13L0xQ+3VU30AbAbbCm6Pv8uw4smadXc820QykrkPOsCb
3q2Gr57w6moaZMvDSe+mtz/CSFseI1k22ilhZTEh0EyTA/bPWEP0s2I/R0Tjn7EQ
Xh4dzsJcp3R2STs6KMHZ5vp96XZ+/JxYXKPLwAtKyGeVDplG2I4ndRgDM7KW8GBO
ee+M4uHIJkhea4Axqxu/Tlo1j/jXYoXEA9mXI0qGFUbjBg+eSKJ8BQKoswpSKxDK
45XgnunltIjXlEqRUCUGTo3eNs2L6UIYxj3b41hOqiSzC0CQZl3F78WNzbPmyhQv
+RtPZF4Wg6pGvJbx5TY2Zd6eT7rZKFWrJ9H8kfJ79RmDTLrPtWp77hbEWGVaHIxb
XjjmbT8jCZIdwgQX4zOrCpoMWQuoXLoeTryDjij/tUNweSyb3qB1wykOnW5/SV2T
0n1xWZ3g40wMwqE4hsAbxFbjk21cvL7YVWlJnC+eaKRnRtEfJszTTTxwD1APAx8q
CkEukrBvtqaPYT8QRIZKFxus4xKeR+Q3QxPUB/g6qte7/z5ooUFjH9uY5M1mNYN4
UY7TfkDeYlWDQuoS2ZD/P9JFXgonrL+3FjAF8DLBK3bEUIAxK0/st5mYU0V19oy4
XYO8AeyFCaKGxnGFyEZnNoA3CaJ9pAc3PXeEaSqrQIugnylwkiu4aJvcoIZ0S3zS
pYJPVReKfCXfEtDkykJNfqzxvExE6RB5UG1mxQjWKWIuoDIdofDC18izaqyk1KmB
o2iDdTJFKtEqCxJyqyyjx/3mlhIXLvjQ1uHiTy3ABlVhVGu9djPs7+Zwdj/9x8XX
H13YDrlWgnoDUIiIlZvKG8v7fsLjs/Pq8pccu0OGEUQLPNeH1Ru1C/Ea60UsFfcB
UfxCAZUkeib5uNULLpc07UQyqbBoLWuZXKF7EnRjb4Wx93EqOOW4AxDed0qu5d+5
+/D1XQjw4VsR3FvFWlEMhcNN57kO1v9BzVR9SqwgtNPkxnQjwT+AeHN6bsvMC8kF
dUNf0MRHNQAYHg48x1wZUGTbZCTXlL1vozaSJ0EXCr8Qh+IzLKGD6fqN02UhjS3r
MeTzqR+aG0Fje4s7FaMGGNDGk4hgwcbQnuNnEvi0UEXW6SPTmntx3TJvmI3EdAQp
vT1xuoTdMd/IFe1ZKk/OMxolViHII6LFlevzAEXDFOZujudiic5yFxfLj/+6aiS4
V1nHeIDL7T7HSec3rVfM/W2KTQ7AJC4fohUT5PI5/eLZ6fYNzYrKnlI3NB/W22L5
WdDlZm8snbDoCZ8D+oiPPbqtVC7pL3Eex085o+JhcNNEK0AIR/Fv6xJOFPu3iq8l
aS2zwXA+W5btrDJn7XZX0BEqfILe8iaDw/jv/0wdAzejudivr4Y33ymNwyhSMoMA
uMFJaMXUvQBUyyvutZOmRaD1YvwTwt1kqjoODK6FzO4Wa+QxizcRG7TCxLz/BS0L
b9D0Ii6H4zVDOzPXz1d+/f/kXFtboWB8jFhF6hSQcLdC1qd/w36u2HP5LqVypkq4
KZ2ZbyebWhzeCxpHk94LrT/Ngv1PQzhGfVKaFHtS0g0dZuC1GGAKhor7VEPkkemF
wkF6uibW5iGkZdelALOPMKvEw2Pp9lmtdQUrqR+oZTejH0Aq/nmaj8TeKa3QJkJa
aWAI9b3n9W6qPB8JiA99WdLD8AsY6bxyQCnbpvJqDkPigse02CGBn/MECpKPchsz
Zyg4rv4uWU3nLkBXZe3MoUz0rtmj3CbpAVfXjskLZ2kQFRJ45MNaoExTny2L0E+4
hYcD999z1O5/PIEe+C+mwnUjKJuMiPB9Ha2PXWymMK5DfqmG2dhYDK5ZX28p2CWv
lVpsMTg56IJgxSodafUs+3gCy2Z0Q8mfM6+yhV4JsnOiduf4iMk9x3fp+CIGDDuF
DZ8UFsRCiNVdk2wJruAjTRXkaGqhDgPfHQpZxKFZLrG7ZWcldNk6ZV4ZRv+6n5bR
1u+lnbXXfuqVAPgviMtA98hAVZ8CShrYJ3tsCEkyKfGupb/9KYjvBajd33QLUeAN
64EjunOX98bO00vgdOHlpo6XmBBr6fzWrgaf73optQihveXrsNOfmfd5isXU4eaN
v6NvY2Le9bytis6Aqhxid59UAAn3C8zmwSVNofldvhpoc76xmptwVeXElQL0KbML
/zqX/bY4Gb2tS7YumWMDgNz8GjecNJIYPs2zxMQVnABgg28XiiV1Wpt7dMnQBgUm
5nH++8K7dRR35Vj5tDY7C91vco0b50si23p8tywPLvtQaaEv4ZxNHOh7PPFESadf
0jL73dUl4oMiB3/9rPSEIPmY8IzuwGXXi+NpIzqRtPHLg7K/aw0I8X2VON/5zXYm
ZVYK+PsXoxTMGrCnFvSleiDjNzqizN2+Zpe0ziklNbcPu1pcDotrOWCnRfr4/dts
Qpvljz1Lpv2T9YOIAK9TRJHahHqqArfE3hvohdT48gbpgha4eFePEA/D7Pp9RQSf
j2a2b2tgupvWUGMn8HoDxkp/WmYr+QVkz026DWHkqx5HIuO/sv83biESl/S4of9l
6B9mQ5Arc1PcRPn8d+aRlgHfwUw5FMfiKrWoQXPwHaCPwcsaIx5zkgg6hACX7LXy
p4CH3pYFM4BQ3OSu63n+ihv/cSCSk37j6Wy4KE+k/NVoQdPfkcmTfxJGGNExuoxE
W9ja1S+K/vUmNjRQQP/HUJM12D9kPekOsKExEBXinv9GP3SOFGGjFBYIO4bNMlhH
M/iHlp9TYcg7Qmr/KoycWksBYv4oUvex5JI5UOJGqc79vQhfo+3KXLC2OfR881qY
ZcYrvX6P3b+a06bmw2rdTkag1hZfCkyJ/D/jZSyoFGuYPbCTldydzorrD7d5DLjt
bD9259GfliD7V51wNu9sApHkWkyBBeB2iKDlTogPD8Aqshu8GAInpKX96MIp0rAO
MKpXkASWco3XxnjJirAFkCPyw3vu6fVInoOyuKpOmo1aXK5fVNEhD4KBSRTCRScH
RoTTpj3/m+UFGMQ5f9Cw2ABLBq2j0io7HOIbOSkyKt2Bq6SqY9MCyLDqdQe03GwT
EjnkrFiMhVbwWMhFvpPlHmlgQxbYQ7MT7ixXptrtoTF5PWnrMMhc98XPrExJEC0m
gQMk7RJIP2kmPte6ZiWM+SDsZWglA+Lh/E6+fwYzhRd+f6bMkHD7BQ8BE0IVLsaT
tb0dfzb/6dJG7om0ICwy9qu9uuOMo9DF5u+lzrrhmnWhP3mdOiUiamsQ16Af9WTw
AX4iVYzF3T4kU4DG/PVV8krq+pRtduU2k0hEYUIhiRJO7Ymu/SDNcCQ3GcYTUlbt
XGRt7bN+gusDA+/hmGDiSLZNZA6LbadGydg4RKgi+/EpCo3iQVncaOH6OQ6SDe33
GxeVQu81QvUukLTOhexAXr1XHORt2bundLv4K3rN9DC4ZP0GzcVJdWptKXh0dVME
KrNDVdV2IJp2FA3NqNnzz+NmmRlNQN63cWBGovz8EzKgg2+CvT+IwDvTJFPbXpeA
XL3JSoKrPMoGaVKb99ROTzqSBL8A871PFwZK/+tRpXXOswgv7iJEr0XI/FoqLAuy
96rRLnE3XagJo8xzbOoRINGzW40OSQ1yT66Au9c4JqR4/Z6xoLLqcZKld5gm1Dw9
K/XJId8O7/wbQGlgYIrTJHHt8dqmQ4FqnUtmdpPzPpERtFtKSn7iUJhcQ55LkhmQ
OUqIdBQiFNbwB+hDc99gnaVkW9Nhgb3ZwNBqnlw+PdK9024VgCPVttxkP/dDsomo
3WvCV/m1SnJKl1eJtWbQkoBjWkgQUmaV12/Yhk47LMrn5mocQrIMmL/GlgaXDRWg
PHE9RAR8Ne+NOqhSS0Ch9CDC2V+Uuo6czrKu+ijip5/161z7wE/DS0I6RF7Ar/HJ
3a9ikE82ZL9fRKa+QWmr+uQodvRui6pFuYDW5RO4lwWmkY5Ndrt6Eb9zKQaA0i7P
ctgJWJAMHH1lHL/FU+oZ2qX5FoEFdL/3K6YRwz4+5KjWY3PsYWH/ICnqZG/uG3jh
Z/wPfA4v7b/xasoxXnXxcJIGH9OnzXnU7cLqLtDQovqT8tgs+HdzwnO1c8SceB0T
IB3QLz5mDybzuCVPgRiiWSY+fyJM+5iYFuWFBzDmcjNOC8i3nyUpZvygz8YWAlg9
ovmGJCuB1DSfFq9wAM17olcScqgeUsNpIrdViX8ZdQ2a6BmRBLrxEuvz5HDDUmZG
bBTrpUN3BQrKU6haZAVZZ1gHWrkT/ugB1ZTdpR1EPx2CqeL4RY/ukbAwq+KcCttO
/rizrSExtHqlG7LLVB4MiQDyHRVSZHJhrGHZzwWKQ+F9/7aBMPPX8GkO1XzCSxkr
79LI4GUa3aWTjYAzY02g0FZo8u5/+19qbsr9QvYvQe7H9YxptjtTTTLQind1cDE3
nSXXZT8tt1AAZlZBZE8jTUTfnPM3uHu+NNabaokubkazwPcOdkkOd7RIFuqv/6ow
QDZncXPARer2jZMvkK6FxbdYkxNuoZMuypKTCQljFK7BrjM147BJeoXSfelVo2V5
Sq2vX4ZbyGJT8ityGXQQD7Wed7EkBWxLXn48Ff0+ZMywIyQG1Ydohf5M3wHOUOvR
0CoOwKmfHpDirtzD/G60dqWIcwb3+kM9UkkfdCdb3qDoJYiuM1qFG7dMC6dfinnV
/hdkSSZj6A2UBohnGpb2wmH1ZCugYLXFBykWuI6pkPzEhzQqBPteXNmEm1mb7Pmu
UhtrN+8jFenSLrAtAn/0PMuPiKc4NvLViK9Z5nLLs+JvRt7iNEEurVrynBT/Cjid
IHEaTDILnPfTUmBH/3KL7NR1NEwcOLpyPdR8n7LR2rXDqFp23GYD5YegSMGgeCz6
ktupr99xCMlnW3VWk+KJhANDA52L22h7q0SM9bC3Hlo5VIsF/z0D+lzHIlCghtMT
sn5YHSxozWdoBPZp6BxyaUlhAE8/1NsfC7w+zOC940BTAorxFiOV2ErF+d7ejtOl
pEKCg2Oa4RzdQsogZfZyOZ+yzWWH9SzZc7iLmtRxQqh8GhQSZmfXXVm5Vd/f0ksi
ZRZI1iTbeHgXa6LOuqyryU6RegxPQ8oPLGF7nMA/QDqlhjXQZ9bwD6/Z80p9q+Uk
nEf4cmEYHCXYNsjzp3RzV9oysk8SIO+Q2pCaKpMb16yBBkjoTKlE4XKA/4QweCkf
hOPrZQD2M5mPK1ZYOBWyChVpthiDIUnPATen3CbC66n1R5IXwbDosoPFe/0/p8bg
AdHrLrBbgUt3Eg+gkdWgQty5Y0ITuH0om6n6jSx1hpsLMYgIYiNGljSRSHdNwaC1
yLB44zR3RojFU94j2LUP6PmVU4mXVEnjPWiS/szl6OUOlkPA157DJ5fwwXJ+n7eK
ieD3VGCZFrcSYcXSaAEZC4er7KHtrQBW4MztLPcNpdUVLDv8l+kQ63Xldjt0n5sm
hZGe4k2BQVnJF1BGF7x+ld5WdoK3z0Ki91c13No1OIZ+dv8zMt6n+berBBEQHc47
i4k3WiL5O+cpF+Jh+Iv2fUZinwzp5qyfCrxJHwFCtgN8gmpCS8wUC6+tHOSog1qj
H3u9NfQspvZJVMIKzIAOVUA4pi7SteN0FkpKm9DQ1zFU7RSnXdGTKTlPkYdz+5Sc
FGZK6f25PSe7vsxH3d64Ru6KYXSvJzQKM/0tTFGArXRJPZjmq28OXj7oOttahTy9
P8BEdZFLV1mhVSv7HzM/NX/cIR3w+c/BgFU95FeSYqq+k/Aft6ie/PdjipbeMqfu
gFygJbALjWpjHCiRhP4+Ui54i9g7al0JuSGW1qhTEd+mnSs5RYpgBv1/qppZ2cQQ
4QwHDcOA/7D/5m8zwKMsCWuhJEjR8TIIwrC8e8jhXKDM1jj/Iee/59GBBGnsnNHd
5FBEq61aZjRsBYx9OUqjNDRcmwJdIBMp/JM9RlgZrRSd7yZep5KsK5MFmogW4rMl
tCOpY5xnnSMDV4HqZ+UVPgel9qyKdLCFwSrNcXOMDi86zNQCANd5+k1azOQdPiV+
UJEicAGDrnJmViZOMqB/JnyPM1OLZIpDshDiG2xd/vUcVxdI55o9ip2RdVKUzOsi
xqu/iXXxXfdlo59sCfGrZljjgoTvDe52qF1EflBofs/YPU5QjuRpvH78wypHXe6H
LEWTHx2UfG6lvvhUXTxdcr5EoIFcwhZt1BP4xWp9k6F9znIIPRL6Q9bKXYjsyMEl
DRWCfTohdJMlsY7s07j+fKSuwXGFd+n39QNtdAgbF1lm0qXo6ctyy3Ae1WZuz4LI
gLFVpjbBlvXXZGReEZO6KQVXpv8o9JIF/THtkcHgVoTvsaKOI54NY5EmAAQEghN0
GynVD9jTStGj4exaF8T87nq/OsoyIB9XXmA7j3dYTtq7drydHIQuODscG+b4n0rh
7XJQlDRet8GhRNRsMkrF/S4gRhPeBFd5Oh+fsO6vlNh6CT8aOY2jwUtL04cHNxTi
RZGtbQFxeUoBIQpNrdYIPfk5LdSJjBJ6lNgatSQDvPMkrsMTqZDJ8nVQtD3fsG0B
pbEmyzxZWfhyM4/sRkHQPOkb8ZsJ8iHJtW5gCea7lT4YF/MxGLlD8XX8FojqIV4x
w96l2uKTWWC9v3MsntusboumMX0GXK4BA+WyzBfVpa4bgHqWfjsZ0ne5TGqj9zw6
57NAnhiMT8rvjEFXyDPdS/6FRgeHi0m4nMtyfrC3omM0d5nocsFJTSD++3t1H9Cm
m5nqutMr/KcLwZfUoxEa7O8JaRtIKgqkpUttBJ9w0dIiX+DZeUh2tidPVHqvx8WG
/T3MokYqIxE44Cq/W+qw0/ws+3ZeF4PUdRwPB+HrK8B7jftlK2bP/lJ/RUTGcJ4n
NYyu3pZTpGSprOF897ly0qthz9AbqMjQgb+SqjcSmzF8dsRFinRc07+mFRdq5Px/
6x1ugMjGM/JosiVlU5LbvMGJRZy9pTCtK4MgO6RX4i7AHEIJN6di86Akv/fBI7I2
zfQdH/7iztAXXq05SKEyhVFulGSQH/cuMI3X4OwZQYvmohJh3tJHmPgO/NRs6LW2
VVEHl+BMZ4hAhyF+jcxG1gGtOH1m87jmotxF8t+oC6SchFwTeCmhOhZUvreStAqS
OA9eAY5O01eGGxdhjsEx0JcgHWXCBIEzqBHBpv25uq872SzfM91Mpi5rwNr+SPI7
fp8OkQLRWkPEcttmDnyHVk9ZMKvO7VgJ8iiwBIPGAnVE7wYcVU6xlNSC382/RjIS
MEFDsL7FFQ/oet+glau89xfKH96H5QBsDqF2Ifv7/3grxtczVlz+43BPZD7v5qwj
lASrXO1k0Sy6wwRHWMFHG4mVbB/UIKYpsoB6qX75051AcVYNYvYzJAQDijBjy6to
AxDrPnUYJOwdxpuvqWekywG1uarKyAVh46Wg2IDjtB7D4yrVijgXnvGr8gA0AHNU
WzerVdELHShKJQdACBlw73cFCrQl1j7CTd4Nph78Bpb8Q5em2LbML0qCB4ZQQCqH
a21k/yfkq81IL89DW25ee1JryeL9OpF0RiP6VtgC73/DpPb8wrlAxM2dOnSzzkpj
cgQTN8ZB0gPKrq32z3RIZ0jrBLgVsqaW8hNRSdUY8JbEvZ59M4PrPX9js0Qgq6zG
rZDYOexg/MdFCcdOKlbnN35+zlD+wHsqHRzbsprymLro1Xx8PsmsRhwJQ/fXsaRT
DIdh46l09FykPRMbloTL3kk0gMegaE9MECHgzjgAO0cuJaKQ0COLvOx6kCAqASKl
gR3NIgZkLaMLhdg/Ia6olHIS1kU/+oNSj3WEPM4YzFzYvVN+gRunB6pcEOedaZ4E
HO08OcE/Pq+IyURtsqNNR5vg7ACJ58JU3FQ4Ba/QMULpyU0UfjlhstMLBUsiBvk+
vPPSDJsW1mBrnfawsqS9fGZipLNV/7mui4bH04PD/6u77RcWwlX22ZM/41ZP1ZXx
nKoCWh3zTo0v4BjndanYMzq1FMHtxYhwLVxjzfASV3L25+/A3NRTkMedfn6kZyzG
j0wQ8bgMD/yCL3VkHn/yX7QNm8kh596xnQQvOAY3JHwMFXP8WDoacLNpWLzytp4f
EE40wCvcj+wSpBUHWbdmH+nmAnyfFZnQ7xWtQrQVvjzs/6u/cJ87LfqjG2pCl+NC
c16L4bdrpIhQNn9Jg83FYKh+ImCP/FkBJwM+MZET2Hxv2W/Z0brjYLQ0e/Kyt6b3
YBdOWrts3gsQYKmqlPoyFXdgY+drGVUW6XBeignMhsBukUhi007kZsYvboB6xm0/
Mfonpaocy64Qc1M5/NfSX732XCi7f3a4FYwBrDtwNV5QO26L9S09RXov29e/z4m2
U1MfGX3Hvn4jaAXf3t1VxEyBlKtrhQ+iP9Mutg7ijQWWMId/rFI+ZnEnoUv0bKTv
RTBfflK99HLjcxNViEcXwYEYgfw3MDpk5Vaa0Bt9BVJimoc64i4zVQQCh1GW77uW
J5MBE4Hm5L6tiCEPVnP4UWI9hzjLUud6GTExBbXJjQGWiD6K8mDRHkIcc2boU3LU
Am5Cnevwjw/xK7+MdayAM3uiQsS8RR1MlF5Lujj1lXW1DOc/kqfgkYv2EtQtVC1P
kzOSLNnTssCinPM3SgoOAsicI+5Y/+Xf46LK82Mem5xL1RViPm7adswxnEnVdqaj
GpILKjK6i4Nzt3PxN5VjixFFZpIpeXslDOklSaPGAvy8WabZwRT6CU/JvnMv/k5j
83sWMW67X1X7438dp2DOf/YWEA1ww0EoMUsx/98FJsLB62YdkmKfCk3w0XIeUPfN
4bUVNC4ugqx0XObsd/MKgtPRbXpb7ZwMU0Rl0xQXOlqIEdclZ77YW6QU1F/ntoK6
qwsPac5IWCy4QWaoEdPqkQrV8RqgKYrDYxDW3Ht833DvnoZf/iuff88mUtcfal5t
3wwJud8I2YtJ86+lM0JB3xfhyNy+c3vnAIHXIaXjJi5UrxW7vJQwrdWx+n5rBgcJ
DODp1ZDpbHUem1QTABwcidFJMqEO+pC2IkPiKqDoby/480lg7Lq/kL7O5PY7LhHX
L1Ry0BeSbKWdV5GVUyqXIApdSJVhF4BNLDoDpRQUBUsxIOX2ZdzDExGb51VC0Xn6
PKrNZjyZyI/O9JNpll0b0KFWkxBwGwvSnt8oeygfBfQ0On3N8XNcu1sSgP7oHKMN
//KKeOGwV6wHo9AHxJDQscZz/4+zLwMl5v48i3wQC3TNNvkU/2otm1KbkEVQ6TcL
mN/Ig/78eSXjt5CKQSf7lYqbk36N25HhjCEWsXRFsvT03FM69Aap8b316ELsjUNp
TTrVD1lrijKpx44VSuFss/9zjgj0ryjZD3YSOm9VQFh4C7ZKQtBOY+TJGoB/6mej
F4a0ysKKy3V4oaVLf8xR8NqkZRV8VmCrUXqoL0778xxt/6JlxNbhz+lm4UVnNy7n
KDkJpiLZXyDb7tXBh+KiNpetqsTh3KptuAtlbqaEWFX3WRYRkvMPFeXa1scHrEdd
rtPbNsJQc+jLhz09sz2s+Fs9ZSrzeplAaZQmDwsl/3A64EoakpjVICOrIXkvsHcX
uFmzHQw8/AMN77Yci6jPde9jLT7EgSNHZhjfpPY7UqEQmHfUfzOdI1Jxf65h3NHH
uQnaUBkmswIjL8dzFuJo5j3LX0ywpQ7YjvhbpaYeLPEtaER51oSQ2IvqcwdYZRQ+
vwXD4nkNQVqQH+i8NIXitzW81OpjWGSpG/ivKxX60Ubz/AMnBHvtEeirmiiqRnM9
xYrF5021y9qC/+cUAqCqA7vUDQr0NjDtStxQNyvkmMGTeo+C/+iH6k+BD18fEk7/
wTrRgNeOJkXGQwgW0hIeJQ==
`pragma protect end_protected
