-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YIjdghvizRqj4E7ltM75fYLcd4aFLLwofVL8fv+7IEEwJibPjOwxJygjf2NrKmBW4l/Vj4auiGUY
J0wTH+/EROsV7smpf/OdqLmmOD4DZuQJkGzITib7+3oRPxy1nh9R6dUh4mO5+s7WoI7cIRFjscqv
2eL3L5ZwslwmjFUEN5b6GVsd56GeqQQHUgHyagUEJCRRbM+aPCVxPAYoK0c6sFJiAP6TQcR0Nx5i
0E9O/3RCkCQLqqV2kILzbwUo0F1HF3BejTsgeLxRoW8ppMBKaUxnPyfvIUKReV/s6hZQJCs80MQP
ssjcfVyRkyUE+4+cIn+xOLEPN11CE/Zp2c434Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5264)
`protect data_block
W4L2C3AqpFdF1Ym7sUuoCRCbccq78LoNYAY5XjuEIb270T6K2dfZdeEOtgEyDu03cH+pYfsAS+71
AwxwqKgN/ZwqlA32TKIaifAdfUXXtlAaXN2CsEiUukJtIYiGxH/BPpEsAHBOtIWYAU3oe16TJ3on
RjbGvq8mpR6m5YSw0P6KeyHYH/IR+O/lWBpPgqDPZMOUECF7gz+rMjQUaAF4RKK3xtu3kmbE1aWk
8yP0qFm8hF/TPRMcaPfWXwLdKJoru+ssov0xd9K85nz28ppozOJg16p+FrrhU1mL53OZr9Au3aOM
AXSyvhtkEZ52LPbE+bAfmP7G1aljL3Pd6ffSMd1xiUYrVLyzhHxmCKTRyvUAl9xaXP+XSarchsUF
DaO1eYHq2f+bz0XOko6brzC20juCbItmJ73pqLhAcj2jINqfCSvTc8rgcJKBnsIOZ+aKZ9UAmFxh
k0sZ+ewE/GU24HSjLIOzKa4EhcqO9RhDIWdh+0bROUZMo1PCWZDvLoA4jQZ9zeSJsqapLXstNgH5
ZUrx/OtU9WllYLsXN5INUe2PWEkCyd8t1mRzDnomaO/uPxbIOPDW61kwG//JW1rtzirvUmvB0y0S
EUn0q/UhT4ZKyqGojRw38Alr7OWXQd06A0jRKeNewNO3zY7nuZYMC0nHOIKG18BBOjrlrqwmfwIy
+FGi8etNHxs5/RgS1aVPSV/Af4dcpanjwsQad2FtLruZK3ZTwz7v+t0vC6uHR4QuWeWCJuS/3IC/
yKcC1iHalUyBzeQdo37qcsKgv9CFSoBCzkW0DruIjU9HbJLahvCH97bxBfN3VxOUYJB+7uDyFHad
bdivDjZbN0osTy1vggOpeHx0Pqihe6jOzYJxHUBq6g4R/dmmFZd1XKyu8xFC65WEpE4j9UanS0yM
yd8UC5e2USx/Al6aDlmHTDmMr7iWJLoADQUQYd1tXpXGRJn//XiwyjpBA3Nfd+8Zh0U7rkyX+I2P
pYJ+okhcdTgALS716flZO+4EEGGbIshl9n8OKoxgXkkvTCsVtX/fCfCDOBO/zu7Y0jlZv7fyb1AT
IkHpzFNCuO9x+Ryiobw750DnypFaBeQU55qJSXSj9mXvaDKYQ7HMGfhpYlulA+1yoQpAfMVqsTva
Z7Xn5Ggd2tYpdYD31u7ZkW3kmE28paJ04+FA8HPo3xlYo4xyb0GOf2J0FedJdWgaJJzcjK7Xl1U2
q6sdQnqu/z3lAHMYa4p/S1aenBC+w1lKR9tzBUgvNw6FUI7aU/7PebKj62uLnlN3bXt8EnJru6hI
DP70WHUDCFlYWGE9O3YVLRbSTiMO4XWlB5+J2ik88WxjbneBsDajDLZ1UVNW3qxgaDR8gYThmOVy
lbjUr6KqVL556/hpyGtCMIdN562I/CXV/DcRFMQv7lv1cOU2yWplLKbxrUvcPM70MYp67dePeNqO
H/f8E7rQLecVlwbyTYd0nDgI4erlaBDOvUSgV36UkD7io8u8ZOeCgjET5Rkhd8PA5oi1+qEo2CI3
R5JsEs8D3yIK05+U9wf24mpQ0P09GhgVGhpm8kclF+LlsnyyB21HeTR3J7kH4VqmYt9SM1+OHuvI
h+OeklVAu8SMJLSuexAFp50g4PxrmGJKjfRmeRDPmbrZxIjR0TgsX11/tA/r2f2jDoI/iRvfVuv1
zztN3yconLsn3iYRp2E3kJV6r4F1antjT8HUJgCde19LRB59+qgh0VeGJb4O1i2XDjzj66YUTbh2
bKiaPm8nODiHqXhXYBb+2nOWP+FwFpIGqqLvcBO0bhDgb8uLFvkW6mNIvLsgaaKDxtWpT3Te1YKT
4P2fPy+GV4S71oOqTAXIC4EmCOwQV7A9hetkXKOtlkXNKB3037vBKDWYVyFOCCpFvklaOhhHbA0X
eBibYWzucG8PWXK6ItRpi22MulPL1n4jl5/aH+KD94NmpvDQM8HMaN04H7zVa3Kxz8vX+O4Nda5B
k56O7v9Ff07Inx++3SIII211bUQGHX2HFIgj9nB6xWktKNUbSp/BM+EOSyBEGOvmzegqB9rCHbMN
7iy6aIjO4XZ3VilDQd900LURHsaSi19lvblUuDzjpipScuY9WGM9o9syVQNmZ45K9XKxF7s5ViI0
MeqBgq/OttYLxtQwmSoHOxzdtdBcrRrzrlWitK3HeCxv5kmdKKuisSmoiVjLRGcOhn5WLcafrXOV
+kmdWA70cBIrWpvTh0bdFFWw92AEsz6f87nS6dNoX2DlbelghL9cxFbtioYnbbI+p80uTQ9c181K
oTRhhnDWUAMTvDERWp1FwSE6Sfv/LjByDgx2DEnPaRXNUlO5e5xajSffiaNTdCcoT2mIrhnLZH+W
U7PcKd7B122mXtymucr7j9y5JJobqWcEjXFFAS/2BR2/unT9o+Pan4KIY9juPoMVAJ5M8HUVewtR
JWr36cfkCrF2VY+oF6Izn01i6IXtkC+8SPMRNupFWFu5nBJdHA6SJVKrMa86Cd8GVyCMir8e1KO4
ioYnwZJViQv8rWNKw0RBwh4oQ38Ww9npIfcb3K23iFEUQlTgpzPfHQ3AO58yTaCS1HqD8xYBHRHq
1mDfQMJNBNFB21DAIzWlx4KZ+SFW1hrU5uCi+/mgDsKfufKq7nNTxxN9QeAUrYY04Mios9PQ9Wkk
p8i6aFhEJCn/aroENYprqad2RBpDeDuAWC7VTQsvGbE5WuoNdBMFyNP+SdrFG0SrGXWb36drH3R6
oojuSVMOJNWxVHXFhGvnKVMY12+x65RrLgVLuqgmmaggbji22TS4AMmyutOoobadIb7XV5LPuMOi
Lc2jaM/bNp0gdHX4q63i7SGal1ID4v3tp2QP/4zj6prtSfGSbebJ9KAqJwWEmT8HcspfGIflTR8J
1SF7m1JDAksow3ZjMqZHQYsE5sMVNnfVi/QB4Aa4moFA6D9hQ3LUYVoNoaGliXHiqTlLx3M4elrY
1TrehpIECZlsef52ELPqe/MEb0rWzN9dhNt7/nWoO0xZSXySbu9d7zjDVtFD9Bi5PWxEDkjFVL5U
3ciu71jNLwEhvUnGOvxAtxSFPV1SQvN9Lw3B3yEE7/XvTN7ty8EFhWjSVwA9QnUZRokpO1c+Y2cf
OSsl1jYxpFlRs4U206Pqt6BqGYd/zZCMs3KyqO3kmed0lm5zyLi0yN4hzY29cO8d5AFDL7njUart
MlPRjs0WJG6nQYZQDS4QR0zV6m/EXo35fREF+NKtuCh8y/PbUpz9PBKnM+3sIzoZpelZ9bGJJXjB
CpSaVrpx2MwJO/j1GlK4m7PZPDR5ksfWvygTgw4Wh1v72Egtz2dzI5mp7K1NGpw3vd8513zI1SaD
scyWzV7yqlQU3bmjw5xC6YwhVXA5d2509OhMrVIHZ/6sjcK95M+4Tyc53WYN7cJxejlMyYLrWgEJ
KxXGNljgJtVYZlTDJ6HgnXD3yV/kSZYP6mxOtvhnbEPxSa4oAO960j/1PSk8rGWyNi4e4P/+RrNp
LNpOuWV98Biq8xJst2+zuRgDUNctH/DSXnRx5p/Zli2gQlhgS7WgdxPoptEykO/94RcGWaSZt2ry
osh05sniSO90zcFS4xIS0qKL1oWHPI4tlJK/WC3oCQi+wFT1Eb0PVr8xIF39v13rWuiTHYBwA69H
pDfw1/tXOia+vPRZIA4CBUG78QTqquQWNRPpOgaCX1fy1byT2ol6e1t1U+P8+AXkMT4/7JnQUBuP
xXfUMU/pFTZck7aVxdoFqXPIbhVAu5V+ZfHHC9XAZA1SzCCSNe/lMIEmEYSU8LDmsGbwGDdgKtyr
j3K+/ZQhIr1onwbEPE/Mphr/emiavfW6ewTW1hSxPDHBrN2MhhvvbZKPDNS4/DYQIntagjKSSC5y
o2xRcJZHJoOBGV5FN0uytT0zM33vjQTgs1UQQBtZv6mlM1Sb1IMWkRtsajTtkVGZ/XD5/lZ4YJUp
Y7NWkuCSa+fZMEm/lCBU4DH0qKeBPyxfu//x9Bb5PFY2I37jsKYOrbTQSLh10tr9loDUbmAQCXu+
k2jFVToHqlgLk+TPLJUddaBhcliYbuic0FKDr+R2ZGV6eyRZLxAZyHxoWL2p+82NBEAM0q7sAj6y
coXJxnNPYGROd/TzisvV1Sg7x4EqZqOPlg7W7gA2snzCSAX1OWhHyZcT42k1tVJTV+jguI88MVX/
rOQpS5rtwlgf1xkkP7GsQEesxlmKF3RqFxNpf5SlsD+moTqI5iKjGZfjjo2vJet16BTP52ORleXA
0E2oKR5vvyCu2BGsqRN569V8mx9fCcKLVXTA1JCIN81vDIjHvB/N+iw8vyTV1t9hnfIaZNmDjsk+
ZoMsmYpXGlULRcsLA9WLyIYs12kIZrBdmQJRpPXWaHRxP2OeBEz/4Kx441hwxUuBIrzoTEoVMses
kb4r4CrtrjaeyPnmLoW586yWUDISuEvX50+QS9Yqq3O7HURo3mXN0PzQl3eH092gMgI+hrfNJ7cK
Bos7oMjM2TrCwhztDT85j5dZgHPgwlN3+FEtyH1zZvrlhfzDD9kEZb1zF/6jqLam4879MGrx2+hq
rmh5cFbs4nGtdgyNa5oS+PCkaO+3K/HzgrRKQQL4qiy0/KZrNK3Z0bVl7VMR1zDuEFJU9RExs1Si
cRDW3kUZuMwVo2zJJ47ol3OkMHJIvML+M25OC/6a2G35dYY2UaFClc5x+DatQc9uY2iI07jqLsfb
WDlGJGGAFkanpCaqKJqBaDJAA2HcX2JLrMFne8ZIwjVCR8quE4S0i7UdsyBIchRIr3TOgL6860oJ
AnkhCf2UtPzN9dEOEXV7zwFxI3Mk7lsqdN23ubwnHSgWoGOtDNZRXWvjeSQPdla95TAQRsiHEZOU
EsnUtJWj8SN8StsVBuERmGH84omQsft/YNeoYMal23WuXF+TTvu7fyd7Z5xjBgfeptvePnue+IYF
/uipY9mjGoaKNdS4PkV7PUeKwTfTF3jjpghXNUCAllhM4JtWji6nJUzyyUbdK7esS3xHgpcrltPV
m94Bft/uonhBSPEIdpQ6taV3jDwoH0gWrjrOnCtucuEN/WVLZbDhG752eBPqBxRxh0bpfinw4gif
5aQVwh6kUVmj2UglMVUPW4+TOy42ri9t5J1IhT9lXQJBqsdVFcwmzYNa2vt4oeus6Nh4xwsH7LH3
tzaC73+XIoFzB51eMi6chQwgfvv/24A3pEbBotn6gFi0fk1hJw/2ANnS3qDLqx6go/Zb8etINsyK
q/jSLrHvjD/NWe9U4m3W+2eRX5o2CjCx9kn6nuE/pwjHm7YPDD9lGQXGbngLOQyZRvACTjsrz62I
feMcnckpfRvsB2kLnbzxbx2pkHH0LXoP2S3ql1vx8HLX1zs1dq8/SZ//hpbiQISp5sMd7uJI8+pC
I1dWVB2gVNi3stCe8hDBmsQ4BMWeUcuQ6K5TQBqhUCQpcUnsi4kjF5BJVs819GzPNjpfRhbWAkdL
ieWhk5xtqtfQygZ4mmUXvM2d60NbY0mfUUPp0zFpUY6e9zJmj1Clxe8gWccgHqJhU4nFEBt9qNNL
KwKkeq01Ev3ecfvnwFHsMhGcnpQzkAmYFpygjtpg/56XdrUzKhlAtbwBh+fRMa0S9U/gNMNQ5sSk
MrULXZMZFSSCxVzDnOTrfaR4GSwl5/zZ4z7lcTcY95sE312/I5kLDcmouGGK/s6prljIVnOz4Hhn
JAbkY/By9RPNBpIqbPbMbCnoA2mHQmiKBKgAaIoAFKAe0Pv2NCTSNaD1GwLDiX7AdisuBvEdIR9w
8mAzhnAffjxtINAEmhk1gksGCma4gSykeiB/PU2/EMaKKGqk1QUGKqNhdY7zXx6Yv8eqM1RR5ZY1
PNmm2QVzM58h5Ns890tkRqAy0e8suiAElIk3UYrvFRamAjb0TUlRO0Nt4vMB8XIghF4oYNju7Prs
wbj/2KIT6MbPUPFTclm93ViUuofvFABVnfAoF6yVYb830EVsf6Gq6Vi55h98k8Q79cVF/l05uvtg
b8qthrrtoTdMQN0TSWCMFcO4suOnxvDIZdgZGiPvJSkW3OThHpplGNwMT/zkcVeTlDZ1/q6k8eWR
KM8lqy5/UaulpId9B9HiYEn+wqSJhJYZAHLVXZ8JKDiJljKMP/NtLq4fnAJybCOWFzj1CTJl5ch1
sGeCDXBrzbnZwSSFNN2tDbnDBV42iUxcUE7j62+Dfz9cJqsuIq0IeaT+KjOkAIa3IR81g+93QBuC
+WmL6BsjxKqXmaRbF81rp/+SN2/dhPTz4TmGN6HKNijFVLBkEK2WGCWG7GBeySemk6NK5fWw2bN5
5qUTy0SzvEAZj/1Xl4pjj40of4ZO6OK8cMBF9Q7xY6zvZbzk0OHoed5E2ey9oY9gWTlTbBxkRBNs
dIqrOOUnHBcD4tSFgjojaDHF158p+bb6aGosF5UAMPRuq8lCirsgwc09o4zyQS9rlcNh/qqu11r4
ePWxnTUot0DYtgMe2T+20F0uwI05HJBbhCzoWYUJJ/zQCO3/hHBeYhWbcVD0zn6E/gTwWWmQUECJ
GC5kJbW3RkInPkekHCc32yb40iHr0BZ4AAElvPr9QmGY3jJWO0cQpl9FrK1jEEtRNOG90xoxyn5R
lmxLs1Wl/mSkCgm7DDYD7pt2xbntkWgzZOeDh2rh7im3E2K5YUG8iuXlcxHm7ev3Oa0btwhtT5aV
nDjODMzcnBjo4BaLQvdSO6Gi+8xVoCg8X7cvtvYDpDV0MbUO98J27L4atDrUpvw6xmhNDnq/aXTx
8RzYX3Gldqwc0DYgc3xamKLltZD+BDqS1vvIRo7FKzbD6oeW5ud5GtdL8wbO8JM1cLAQ3NPN2Qup
1RI1PjyZfrJTvVBLd1uN3sdhcZ9q9rDatp6XNUJIrbGarD9mSOWCt+eUelofXrzYv6uy0NlivSYG
n6zW3Du/rakPd9L3Y6+2dU5OiZAQ8Zjx7BsmrY7CZZAS+fXM5q7LedEF59jZXYyRU2DbWm3SuqAS
saVxsyXlZoLsRnF4fgX2v8uoqFk=
`protect end_protected
