`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ng5zTyNXe0nHhNkUKRhApevD3dIPOsh8A5lcVauFBjrl1jE+9jHz6GM+gNxO2mMF
oHj2/nPpEEwY5bo4sJQyZIk4v4NEgWXN+sfX3qKk4P1NcIIhfuc/cnxZ3tEJ76bf
2KZLsunL6R6Lt5a7KUi5DzNPRi0Gorqj300+nIn/4d0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57744)
uBVS4pDI8sUqgo7fDRidGbTM77/QKTfXmOr8i/MzfGPn+TykulW9Bb+7R6nzGbKN
sMfRKtFZWCZARCmDrhM6OPdgwqalO4j3+gZV6OvRw6a7v2O44Ij3ico4LNPsOsIF
SAf6qwuMMK9YXXlbXvdkuzdOsXCItOaf4sAT6PIHgPj+SPgmYf/GLIRsn5vRz3Qi
PkEqti/5262LpFeiHgTAE9lfRBE/n6MysdmhuE4i31OoTpDJc8gbsRPEmpwHcIAs
ittK8DiR4k08ITBzuOTKCu556NDg++//ulMbWHvJM9bQroukDLLOy2WastumkvNg
SpQc8PgznQOZVXl5UBf/mSIUEiLRQZXm/06uBAdtYURfMC89maM8t/xb0yhzEXIC
dpHVV/dhUyLHCGC6M9d3k+SKpjy+/wWxTDrDPtZYmxLHqLieHeMBsWysYbAC1S3A
7Yip3b73wR6fgyakPJgrOndTzOV5XdaJFotdgD0DPzMlOBQFpxl3Iice+T9sIp1U
Bpq4bZK3tFIx+TYc+H5i2fqvPJuHp4Sdu/4LAljSG1f7OS+covBhHiVs28AHDXkr
WKMQAr0dJLMd7KcOGRsG844S8JfxvIVcvCerWqNTsvBHYicCrvupZqGjehy3+MDG
9rcwAa0ffmkJaVN26Vr3n16ysQtZK8S++Q5f3QnS+TX0WWtyRSM6G/I6jEuazuvg
uAK5auJR09KSR+8VVmsoQ9UaEXCiaw7wZzLxUcTzfvamJUHuSbd0KPY+0bV7w0vL
dEClZTHOtobRD8aqphXGm8QIR2E4cC4RtQox7a1opMrjicbVCPnJNgeXuyBOwJFk
H4ksbnhqyDgjQnXzgF6oZxQynBN0oKBtauS82gYF7GKCzrts0iadZE2+dG/aqbH9
ygscoHoWoFG8Ol0sy6Oc191+NY5fXg/XDkZJ2u9NCzRrdYs4h2DN48VPAeP0njJt
m7A6gFnn/1zsbajaJ5uZ0cNH4+TkA3TQUi9sIRmipFAK9GbMKd5Lmn9HS9VkphDu
QKn1Tff5WAzpHH11JVhOo9sc8Oj/ID6DTIGtobhi3j0Ghxdv4JE876MSqVX0fK6R
X41FkJEkfFmn+ulkQapoS+BFuo83EV4iJ+EmCAKHUN0rue8LNfHYkAYsFJsjinYV
iKsLl/9T4AnASZtXiq+vTyDxxEZS7EUcAFNZTo1qhFrlTWrHhaLYtEAmu1pqHa+J
RoDU9Tkkzaylyoq74ggwrZ0lfo+G2iICmUQlGydt1y0Ih50WEIDSzMHxWCIQOqFc
o9zqra8ugFmZacInIRJwZN9Ll7EyBGeVZkZDs2fzidy2WAorCTopqiQnZ7kSjgQB
JM7M9/OxriqML9EsQ0vUr6fpIPDMQTxQW04/nd0fng1Wip8p2f4tr3px5QQ+oMod
Z7C/OksPK/KAFaoDALeaIW6j1F/pAP7WpxNnaDW5yxXS3Mi4hSds1oBdiaEzqkRf
EPe9KXyQcyCpx/8hYW4rBOHQhjg3bXCEAylh17sPZ/d8xI+cPMohzXhJAETC16Sl
19l1dmc4LgdacB+hVQEpwO+EsbV+qudKzz4w2J56/58LcedWdmk7+wIZSXz8TyK3
b22wUDsSFtubE2V2mooFfOyGdc2lXdH6cVw6x8p7CEDjVIrUqLEFLXfIknkN1MUF
BvajSvzf78bKhZL64hTIZ58twIffM6d1xhWNjFwE4+VP6LZyDvo1lwDbvgmkMJoH
pwD6a9nQ8ovxySSjZ3SAWqv2HY0PFZsXUHSMNoLVOvGvHYpqP5UAuTrFIe6xJb0M
jtBxp+D1+7Tg97TQAOpCqEC+mirl/FjUqGqhPuMfe0zHJ7znDVLQ/ayNHvS800H6
4flZ6OpTqMTr/3eBKuhmY3enFmvUWrrST1V1LIab7xI3Tou84ZxXuNWQmPWYTNFS
XeLF8ZrxHtOZDR8ROvRQ+6vG4CJ4yu9pQvb7R2rZev14ihg45/XQogJDpUNuZnDe
cL1nkBYp2ONfoYrZeZP7sJ3XVOiIkmw9QN2m1y/9aYqzcAz0KMW1RXMC6fxSTT+3
tDKKAFWzJqqV+8VM/MRgePrpk/b9HLkLz5HgDX2+Q/Hl71Hnk8LVX7QxIkyzcBuf
q/T1e0LQMSY+0vlHgBqTi1ytGPo9UvBDVKNRglj4Cv9mMq4kbhi/V6B6cInLPFWV
joJuWrknBlL0n6zpQL4lHdCAgKlFoWcfih5GRs5zitCHo1xHlyW8ltzd9hrbNzLZ
FxruBXFVARmg1wbkXNuncrvU2xte0Cj7kRvQwdMQu1yi+irvM6szQuu2I075FJt4
RAekyCKAeCuVNO4lxg5W7NiebVx7cuXp4LOhlgfMlbwpivFZcBqgmh4KMWPpSs05
llLzYXffRQo5wuQDmz5ThyHuhBXPSblodP14iN+Qw9B0QEY9Cd+fHaf1MBVHA9mn
ArwG79rKg+wZvQaDzQOer0QMtQBWJY4q68dxeWXU94TbgQcgM950P/cOsc84cnMg
VmWbsbDx15SSm3CfU76+fpVx6FpmXaJxiWthoHgMrGMfPZzWmMZqdeJBNE7qi416
VsFDw7NL2hhpjELgTCElO+nbeEqc630dtPCyNyTZF13NOL9n8FdCUxKUt5g095gQ
7w9C6tKXXkg9uTNDwwL/FuTfApTQXlzbklQARAb1pQRH8mZGzpsCrIIuvWD3FVBn
SYWwC5DslnyZ/QOfgAfO978/Mlo6Y10d7Okuj42Djj6eT8IQrL9eXpJ6BLnXnqfs
XwlAlQ7c1tqdnRnHhj5bHL2McjeyRbstm1go2LSj/wxqI+foSDfe8w/DgZKIZ/yk
OY1t8y4gqp7s5CvgEvVk1DfCftSra6xbzPT5yErnOC8Taa2RwjlIMLL3LPVEcB03
L9+TxJAIj2Ro33I0aqITY9kDZfmDRIvoeEiA+mtS7r0fMYzlNgSNmwgo4wfjnMVt
q2OvBxdSZa6crcndglC7tMy7BczyzLP3ob/j5eZDrgSZzriUbF4+7ytCfA3nEXs9
WXoauYJMM8YASQ2uUjpBdEbHuIWNU6IUyGS78FRZc/M+BxB0cfkuwKNr7QTyF2bz
gaHCO7ZIjXMuxk6CN/Qe7CGHxbMQzAseIUB9WpYABmeTYw2bWZ9ULcDWSWCsWP5x
H8c/FpiZVk7odLiO/BIgXjXmzbmbAtti/xUSQnKYRuOB2ldxEMJGM2XKR0bQMaa1
iCdDiWLArLkMHreyQ/dD2CdIt5+TNpjc3fwVHZ8p7pfauriReGW1SugYOMSDF60e
x4g7/EGLkoTWJ2KH3dznw8dPeAOHk/zj6Hxr2Y/uBYpb6daiqLJ59idZukskiFVQ
OKSlAoOKd5kWUV61sWtFHk+pMl5x9DiWoC4i4NqmMF2OvZ/bD5DnJlPUaKVUXj2b
5bJaSvYDJYl42gpqfiotRiSrxClaB7cQZIXBvBoZnPd2NWin3wbJTb68DquD1L7k
ZA+YiQgjuk+dYp0vEPsYsvGBI50n3MjNPH2RUNrsRovVCVPMxAoDviwUrZ33Dowb
VZYePsZUpdzRGsWuwfN8SXriRVyt3kOWCY5OXfU0BmkiYdMnmtok6f3BwG0m6WIZ
t/5gRH8GxFhvHgR6qJC4VDrFlemq+0ILzK0HyS/Xng4P51YlfFEaQlNat8RdxnjJ
/shVsOJrqA4TGSG9jAn9mCXSEcI3nMhRxD89CT3uqTuF9hpknmz5i2bb7lIbHaoJ
pBuR4WQgNEa5Vi6FrCWvtpR4apCQkItSvlZrJ5onoV0vyKw8OutCD0yzmkWq19x5
IhSVEepdk4aT5aR7Vb3v8+U1AjXNZ7r8KedFmHHxhD1ounrBAf4V0uefJMqWPj+v
nDpKOHeMjGrKzgspRCT79OYza/jmIEokISEmROzeubT3kxorkaJw3q7YHOiy5EOs
oFUz6w64LDmGiej6TKvwEI35pVy1MLgRT73LodQ/hejYAa3+8lSa7eEaYcOOmztK
C5oIh4NYt0APLAXjf1sU54Fu9LZgmzM4AQ41bHdCUcFkC4m2192C9NBkJCpLk2Fl
4BSzq2tB41L1aYLj0bTXFLC+p6dUzsyT2QnOqOd3QT9r1RtoKqvSAeMIpDmje5AS
rSgSzrUzpY/qI1unxQ3Cz+hv3TogapuxUlgJFoEmiYRrbZ3XUee7sQUjFC0layUo
1yLIW5BZN7zi7edqTeqyLp454g4VzhejkGLWZDBHrNzAY/5E5UAtQooaoUSr5wbl
bbp2GpLckeaSoAcVpVXKaBUmR3l/C7oWxuKrB07mFtyPV2wu3CaHDfVeiY8y66xt
GX1S90Ym3y727KGxP+8hLtdylat3T3qqokN4IBv98wSroLAPu7Nj5yavrTvR8Q5+
3roczGk8TofT181ykgCew/bCdep22eFO0CQcEeyXKq4zd7jTxcdy73BfA6/LUjFx
HR0oeeBXrr7c/+NrR/atUERWjYVT4CAFerr2OONFsZz48T59EfWmrO6bmOxC6Amn
wYYt1+g3sLSe1aRXMBNtZXhSeE8rgSG6KEGqBe9CtTIwPj0MRWw5IAd8dIGNZgID
2DpILV803RP/l63xntINPShc9BMO19NzvtkHlItwGHH6K7fUrwEKSV7dufTJ5Pzh
P4dk3dSs+NGSR0120Lg/mHBXQwA1GFvbhEtON6CRFofqMjW9IO5aUIyb9DMGRY3k
1bfjq5HGCrccKAneub0lDXYyshwcuLLxoK93vk7AohtgAdgPDEgRG3XZ/1pma/oS
eWsWZkLEUwT4np9K+CCQwHWevNxkssJXYm+W8xTDplVii0E58Cxdz/fSksBsXFfK
CRA9BV1he8fECKcH6hzEDPgFSH+onrG5ZuvyvTATmJPW/RvHwN9yPEN5uneOfmwP
bmjMrlYLM1QSnVs0KR+YDJFRBGxKrzY5Z6/nJKzcmvj8Awa+Heu0Y0bBxLor2zAC
TS6+74VqDXhmdYbjtgHs0YPH/ADT0zvvxFxVreCSfbO4BKR0UesMiu7gLoNzXh+A
CrwHeXY78OulrgSBSKmkosjD5c5Y7Qjl9oI57SygoEHw/waZ3D1h+JRHCdVlSjy4
/aIBKRjyk6pTSMec9hSJRo55hLId0XKZcMukL5pFpNohtfJZVECCrvg4p1H/rzXl
SnPTj2A4JTy0qDicIXr6DQuR7hKz6/HGG6WwWIUSvIF75RjFQkyj8PKNfgPvYz9I
h/EGxkrQAl+EeMpTyL4/zhSx+u400i0CVhbSC3JMmLErNeY+ynli718y1Yt0HsbM
ac0J1dBLxPVc4EORb8bfIUwJbbLYBgLTfi6i7gbFFu09v5UyFkMvtfcrFQri/vVF
RUaHgx7gsWlhJIJsaOrbE/dpBXtdG/wuqLcJhr3OndjYVWT4s+Ow3lD51KpYTrZg
S6ifZ+xm/PTl7FAS8zgeRhlgEEi5r+AhSnQjoWzedB2MJfyKneVYW6WNmYig4jhs
r22RG8grGknzLD+dT4hU/YqU2y/9jp2gXWEG6lKJkSFKSUPU1TsHNo7Lp8Zpc/Bb
KnMKaxa3yeqh2kAmFXUueAY8VUV+4P9+8HA+miXuT5b7AVKbZwha+IztoGnNPN7F
ulayniOEp+sspA8z1E98IlGDy8L+XEHEl/uiOPPYoRvDS0Vhh8rEwlsDXvxKk5BR
VcaIN+voOQst+ppFTa32wxj/iewwCeEPgXxFf3AAkKY8XMNdJ09wZD0PbGQVhg/T
ghv/k3IzbXTnMvJLAaEpmanCLV/zzyoJGH0DSmYVj0jQ1d+WxoHUEqe0AMpSiNYp
pew832hWUg/F+9KXQHhDUCAML3THb7+y+DBVGXdY8b7Tjsz+aeiwtFsxEFHPdXx8
0HyZc3t8W9cizMHkRiAHqx2mxTS5+gAit55CpvKUM3q+AufcyqEzme01GbEB1UrU
A0GgQYEjwjYGAjEDZLmdL4fOIxPgST4aZYY7+Q2ctRB4rHQ7rdH+dUNsAi1jVyIG
sUpiytEwQUIPSfyy/cbVL9ABn8lWJej1IohH6YFHEPYWt0kXFxBzi8yAfQM9luNt
4gFR+gjrvBsWNIOS9gP/cg7EAGHdQM3uakIsjY00FXkomJss9Iz9WYcwyKeuYYsV
8Vgbb+xTj9tQqZozGNXwglrOCXX44TTyIZCTM7lOO8J59PKsahcNkYHtTDRc/GFP
+TLSzVoHk3oAWcPsWrEYJqGRps7K40+CmYKBrVF/D8NBy0GLVH7cS1683ToPSuir
kijCJ5wKMIsE+TOkcRqf8gOnXPL8cbghzdg8Mwr+QfPNUvx1yrQ5RkDGvam3dQxv
SKMGs4YS4jTGHMG1BZXtKGfui07F+V2f6QyCDOLp+oRrVLsGq0HvlHzXd0b/Q/KZ
C+qQs88M3IHttBrU/xamjAnaXip/E68L3sKsF/fYX2wCrgblfBvMEAbU/1UurQd7
fIKF0TrN80fcVTvzXJwmucq5Br9LG6eX3FCje1YgrialNDzd2G228cOlfIxGjgw4
uf+muhq1KCNXAwzAjU55AFftynf1Gt9aI0JvridA4ZXY9F7cmgI1bvgYN5V77QHq
5RrcZKs6kqVQcAOBVxjae4sooVQ06MGD09EmVDl6D7caquZegsxUf9fTIl/4sXXS
bHJgtWxqkw3Uxr88hr/C/5BywTZW5FcHbL6/Dat8CIaq/6dc0n0HwzkzMPDjrFT+
yf8foN6z0lcGtfsY/AKpIOt9NlDtKIjiD6zpN7/6JyKqUsK9uH5d0eAMO9wG1aGO
8W/RzpiTIAYS7hvaxgfHFzrAWj4svC+qst26tZQPt5T86oBsRFwVXzHSecPE22IG
GBWypmNb8NXK+FFql2rSOlkUKL0d1pVbraqGv2afbtwxMXGBXbY4gihJM2B09TSY
F3U4aFa7oPr9g4xNRKvgeDw011JXEyT4NDFsM0nS5E2tMQlt1BwNdf2vd0mpYjof
UDPpUMkDlwCe6xicw/+y6mOF4b96X64qchr22Em3jUxi/PfKB1SI/veT5FRrJXJs
q1Mf2VcrkKV0G31aqZbkiuuxb/0dcnNvZ4LBqTKUmuwxNvTlBp5GOeiLl78JuOS+
JlmKkI7wTvJGROMm9r5BbtwIZAXaOf9fledzouX45kZ+5GdoVO3+cq9tXhxb1agJ
Iy+Z0XAe77SXugd6TEAcCkmcpYX9FrBME/y9y0YlcBahuhGgIzVkoz3lv9wfFz0P
RIocYR5RoKhL4GqrNZ+L4ezt9AaH4u4FYm7KqBFrbXwavZXyZUr6CazEJlMpG1iP
cLA6JtXZ4+8LL1eP7FakkdeSvbwYWrEM/9huVzvEydmKjJt2+BJ1MjY9Y3+ot/+e
nm51VkduQA3cnCzMpMciZqIX6JTW0A/Kn7id42qsQE0scczbiNEwRwoMB+vdunSM
0RwB2hCrq0mBdbizX96QDfYaFSX5nVbGGMPxLCi7YZLdrPQiXwG1NsorRahHmZv/
zD/pigxk5aSZgeg2ETCR/JKSSzSaTKKZcpB/P3UqYl6bCHpurqij9HrjA2hgvG5s
d0r/Oyla1NVQTChwYepiu0mWPd+lrbyXEIU0u8wvILwDAkXCelehuP/n9KYet8Qh
cwZSVHsyu9LLhxkQakEosxYVB/CX7pT+0D7RVZ2rz6lcM+93HIjJjSROH30nayul
1KoC9UOTTKA0ADi6GmZIdLnjBauLkKqcqkSamf2yAxaohcyWTHEZbNwZTz68MfiF
dYkiMRrm9dEvhTVp1BAqiQQxR8jTCqNByVwBba7G9/CmFM1yuPOcyp7kALcKBFg7
O8XwapMavZsQgcWnHWMq6kX7B3xniclDzz3AMk2+cr9arKdVERzUDaPHLklnRxu7
uvaoiMokgx48rLAKhAghuOVvX2jmPIwEfCX2qa4ljdDVGuG+xutNmkxXxXZ+wGc3
XqZmwaJdFjLEE/7Bd11phWNN/xYscWJTpO1vnBToO3p8N4ROXsjlzB+4bj5RzS2w
JaaUsDHXkWrAhArNwULrd7ENwK8Zcm905YHfSfZXviFv6og/ERhrOfNrF0qehHTS
cHTvbsBCF2BCG430BRpyU5RztlMijqOiYXdg+XFr1b5V6ggMj2wzPw+tpOt+QmXe
FUCNHHMNDst1uI2BFsvW31BDBUE/rAxN4WRxHLDWuhtxQXhmtlSNdH6hQNLfpoTf
qB2JGd4iNY8bg0aTA32HQNq47a8aoQwMfQ89ME9xfHSKV4vFA+L00D7d2prkodm5
7A+X7q29oOZbpaSVOALuv45+/OfO1HaugwxCtTc8cnHkJTLvG/MYOj46L603hc9E
kg6CbtPqtqH2c1p4U4CVWSMnrVRXuxTPUctCt5E7mnv1ZxZNG8ETb0xNfuhNKuGf
utIgG1zWWRtpPP4Av/ZOB3LFr9j8QXRmDcEyy/3rSpDf6FLQ530XtEfPB8sn9X1s
Uaxd6ngnBGgkurXnqQgZyvLWoPRIedZ/sg8gY1AOwEk4HFubdars3ZmWUhssArcj
k0+7bxFh9d3eMREaeSYf8stWZwCr5z+Qf3nnLMYMEVB8AJMrKRpp9JSCz0Xa1ZJb
erybaEIRb9+jfzmfuzwJAis1MZWLTFisrwVRddLbqiQRqFVOKdwuA/Mdxgg9qM1k
BfEvbl6PAZo/GhAuXsRaTJD0aBOUrY2efaApG1wtz/KZoetfFBW6sijfYFluDm2n
wM2icamLDDsUHECHT2ViiFwmH78jHlpBT/ovTRgKCz1eZbyzbQBxoQQ0BzUeooC2
OMUlEoRVY6J67P3T0fUd4DMyA1zO3i8/XK0LOv6FszIr2IAdXJ0+IFYbEReN8AaW
poafL9fgICC1Krbn5BE9lH6I4zitzpbK1eXlr8MDXun5m9EhuA1ytm1hmwm2uDl1
uq0vQ+kfWqhKaqRFK58rieWs6SujqvMxg2XJ18syPxI0N4t4hmbx11SUrUL+Zn0S
ql2HfzGD5xKS2oO05L39bZl/tBEy0S8qe+DklivwFcxK/q03cU7nDUxryYIiDPBt
TVLg3DkIE2fQRQ8LUioB5smnpEzIOYsOaS2ioFNdaCYpQYoc83CeN19x/lZRkH90
AzAuyOk81GuBYg57xfKfFYoGNdPS8LnnY78J2TpAC4x1pSU5WcKb2QQjeXwbcWpP
vSD5t2d1o864LayCrfhf5n1NWW0EXzgFEggzYRW1AARnw7/d5r58s38sIndzwpOA
YiQZgooOLEWW1C+gKz1fYIkDlw4zizf4B6x5xfP381Va4/KaLuWjFkZLEe+qEuIG
zF1xAms9/nk5KPpwGCZBr+BOrHIwuajbY2Gv/Es2d8pol+3hb+xvSFHm2bDFSorF
IKVeBU8fhjgSJvb1trppu8n2LqotG9H9hUJvfcjeLeg2iCAzvs9OC5/okRDoxU0g
8Gb5ufYoqUe/0rcIadTd132lt9pD0GotDT2BG9f0Q7rz5jFknx5MWs5LbDRYcr6/
OnTIUIo+ch5IbrDMM8WzN3VlbtLlKbuAi7FgB96UawMR6T7tjZr9ag7e6j9CPWpB
mWJ5SvVBDNszi3qAOmz7BkT55WkpxYTCvRMRHjOep4O5FkqLAsQ148AOpm+CLhUM
HvSL1aqtjw90I25nT/oQ/gNMw/8ckr+vuIlFpjJQpfZ+W89az2C1YkhyI/TBt319
Dw0GmL811hi0dsJ3Fa58PhrcHaamVyG2DY29s4PXN0Gt6+hwtJmt8M4g8jrW6lQN
lgAT2NEvPXLSOtZ2SSg0xSzwlQtrceLG1WB/348i20y/fo9Sd7WaqlWhwarnabE+
z5r53+oKk83NhD3nTDFrkaZh8sHCRaq+Zq4LMdB7vUoJssBmpfjZSyaPsWnPo/oC
jeHo1bEDGR1fLJ0NCcHJjANfDb54nxBHeNK3CSRX1LhShyb49b2/pHfBwRhMDDIN
VNsXp5Sd7dVfp0nELNIVcALc4kroxG4TdlBPqmqYiLaODHdE4hztx4xBc3QCQl62
f7z4nVaPMBs65cH0KgvWSSkhlR7XqtR6T0gbpt4AGWwi0g3VnYOCDmE+tKmeMyIM
JbSUwtBmz37Mt9RUR0u5H7WYzN8BOjLOCJfZV6gnd6CC1qJwD5vSLChgmIBdwWqD
ErOiH1uHkUpLWMyyycx3LjjCPZzaxavr1YlgaeBF2pQrWKG2S78Ov4XxEu5/d56y
LhPhibiL+KV1mOXxXpRN/zFrNaNBfJYKZ1sVQubGMxrCD5AltmSx1L0xQamBG+QV
LUbQ6H5qYBAqDtdgT/z3Qf1ICTVopHy3C2jC9yDN6L8vpZyFVI0hx1E2YihmG6gC
iAUBKqEnfZehZ2IpQ4Ef8VlBcNJqFmNHkbw4VhuDxOMfvLukS0I5GcdNyM3rToRH
sZuTtKbcEg5slcmpNH4Qvfl2UkvNYWfpsck0SF8xwPvo4xfejLgqexagPirKQgeG
EBlaMOLDq0cGRvK1R9+nSj4JUB9Q2H4NVqAnKcZUJrY8W2Cg5HSlRc8RRDgEvUrP
hmZ0hP8z5TpeUE4oAIs5MqCKyEmHOt1vtoUHU+7Hd8J58WTFqnI6JuKo4ddrI7Ay
gTCe/JeZruugbBxjbsDV3KNSYClavVmJ2+fROuIa8jdsiMiLk+l7mVTRzrtnj/q7
ey3hxOkUYbNXyBYB0uL0zDv7rz30VSUCNRNRK5VZb1xc5YqjlWWrgOa0MvAYzj9K
P+UYoaJhcq4UBtzYMczqUiJOd3X0V/DpA4o4+f5lj03+10iGRsnD+hnxYjmHkWBu
HHTyPrpsAWAjJ8Te946am2Iiz2ocmrRg1z0WkCLntad/iw9XiP5FK9pVFB/mH0E4
3UYu8mZhe/k6p1/rtGYAy6xV0puB9TJs/btSnT6/kaC9AS5V78h8binCGOjYxjGk
Uhj8GCoON+klCNAeAd4PY+yHeMoxSf/3lRMGz/4EmCDWo5LJvhjNIO98RjJz/PN/
duzt+KwmIMTnRoXXUtnU5kyGgm6YGwVcVfULSRRAjEUM/7YoDDBGyW/z9YqS+ShC
iEVsc2Ahy6N/SHeIknVjFsy11wFn4msHBOheqGWdIE7EDAS0+pMvWboPL0dtQCfo
BtmMSGroaACVUG92CSON8vjCfoiyBTSE68J0w6GXHvW9WM3cNtf94hSd+ItECsVl
bGs5YNM8uIlFumwDQ6eNjNstAnVWE5VbBw4Y6EikbDaLGz5Zetdbiq7UWOFTpqC0
IeZNB6KSHR9O6f51OUrnhfKM6wReMzOkUykUj/DTv5ESKt37HdWLNYarvH/16Prh
Ey64+VuZq59e4t+t0PK6HwZ63SDsQAGpF/1I7XorR695hObnamVX5WmPbwRQv4KB
A9TSFeodLJby4GIGcybpVdSkAxO1th0E308vYM2mRt48ETMrFXBzfFlPnLsN0wcX
tzV+fc+w43z0YrzBU3UsEYPIIrIrfhVk6Te0IWIVwMul0E3I9vI6E8QQhs00u/KK
MRMgNxM0jm2fq2Y4QHqRmeQYQgbSFdlPASKVHJHk2dKbCdOJhdbR+xkdQZY+tevc
NWV/kjFoKPtUN74nRx05oiA0ga8FaPKoE3TAZVt2i0bShAhuLT27DyefM/R3eXit
/pU3hnrlb1KFO3NKk9mqt7f9kktdPiueSPkQTPohSXIKq7Ps/ESUIzuBqE8v3GMv
P9Ecc0WJp4njehFM36v+TkWf61tv9/3uIYO6STodPVbfv8KFJyVhK9Ebz9sM9spA
/ojPtCH8NW3CJKOIaJErU1bPGikyoS5tQ4yX9kb8t8nznFeCm9l0d4wfTfkS5mNp
7kKZ7h3lKBw1TpY0lhoOInJx4q5KEvGz1pihwYZifA+eFWxxX/cw/db3hLcbJC8Q
40sapzzA+kwHSrojBZdFY0gNeNyGpxy7SnL2idBQbJEAkOIrMMqIEkPeg2tVqeSU
sWoH4mcarm1HclZtRA2EeLKrZ9o5n2sTKYGNqEK7tch1pmrHuPN9QiYaNqT9una+
vokQ4BVXx1qb8yLxCscUAX+Pfdj2Z31mFhMVOlUhfEyG48yTWFQarD/LItV6LIzX
fdYI5DL+YdO6PfcmkWXwVEDjnOPiwVWxPhXo1blLmPey2gR7ZgLpfrhFRmcAyR5N
mh7g/SpytXouj56dLom5qEMhx9jDtcVSKldzAYqmv+FuszNCmsh3785IhSIVdrzr
4p9lJDueR1sgvNc+rdu09B6IRH3tvCfTSmo3Ur9PQNYMV61UN49UxtAcegFTiPVU
3fYf21WuqcNRZdLEMnOkFTYdG6PQWYihy8oMo1xtsYC5YLcsDS8/svfkDMylvKuF
nCI+EtNVwuY8Y7w0mO72KVnA2oFWOwNwy0fBG7VEaQlaU8GiEc52oDTqQSp9AENt
OpvuImc3q7uy6NRXs935xKd4QQlhbeno2Brb5W91qGIndmdNaJHjPWi6oYa7VzGU
wxllrBQcb4ESgKN4WyEL8qliYvE+w6q5a6g4lKDEmRuN0Uf7f99OR72SyqWqce+D
aPABIn+/li9q5o54GpAD9yGozal1e9qmp96iLdwU2fXVHmRstuOEYQ0x8h0R2IiL
RnY5G/3R7Onxv4FNtcMX/IP9pnm9CZ8gkn8R7t2peJ+0x5XF1vt4UtokYCTyZfCD
jh+L2LRQwq6XF5s8MY0UUJ39AEty+saLq4UIgck+KhSTF9Anbs7E3w78GEEiFwor
NpN3cS4ICx1mfc53IrquIl8qeUfGRGVt449fvF2nV6ezt8EvkJRuKR4ECFl/QMTx
Ke/CzceD1GMAEb0aauPWPkH1rrPqHMm6jeh5Js4OrYveUTfsfOW89O+Vt+J6CHmw
cUcfW9HCfZ483GPpsyXI9tgD6Y19rJ9tlqLWL3KntA8uA6phBegY6+45dfG6lVC5
ym2TDRuISoaelGS/2MbZkOv9YZ7gUG6DNSMw2iPmSRn7zNdUUpJrWEkG0ozzbQCI
j50lxF1RYjewyDTmVgvYlkfb2pnQzBcSGCj2ESQo6FLvA/dBFIdDSMw5oftGNe72
DdB0oIy86StrPrW7Vg3he9Z6UK+TBp8XS9bo+L7IAgMEWojYgiMkhB+ohaSHsOn0
MN1k2cQY/fsUCt3zWsHJReRUBmkLsZSCHh4uGeQVaP/I1nIkicbYP4/JsdeE7GI/
8yEpOCA6+lDqTXngm9IR92Q5qZstNXQ/aZRpBx4WkTeTt0nOAx7yNtD+gGOz2yc4
dYGVI7CtMKoxyibagqjcso0a3Pj+NpufJ4jBp5wa8XObkjEqiq0TE0isDwFKQDDO
fdOE8csEoltJjA21jJUxqMRuunIEaGI2hqlOledyenPsMJ6qxRJD59hZPGHOZJ3i
xfkW2iGH295Bh1r3k9eHuVkQlkIZuux7+jO4sLz2QP8bxSVOIR3xiA314GibsLnL
GTJQZC7Q4iqVugC+ViURR3iZpSERLW63QDy0NJzWcCK71VbhdXOZKBotaumsnfzw
y19/B2ekr/UIBqnNjFqO13hiEL+x23t372wavj4jwg1Qg1KhR7btOdGJYBinEScu
n5mGo/lAe5viuabudvfZjkSxNKLx4ypc9eDIaGHsSHh6fTGE7rOKHyLtA6fDyG9B
x5KyYMT2VTF4NIkEDxcoNq/ynIJl161OcVj1qZJsBcijmdbNkWW9YM8Ae8N13KDS
MlFwvsFNMwYKx/gT1Cda44UWHn3388fJEQUD5VAQFPglZjlmKGuyoK8R2YDvrlst
OmDwpLmipSXSg8dYGxxWpxUj1r+39J8/I8LwLfORWLNHS+uplJrlmLQsT3MQ5Gr7
rxZjGMR5VwCTUpkhKc28lwOh3zF4SSStP7dx2iz5cE830HJ9z2d9J62b2AiQNLT+
Z3TdIA7/tRHtmW91D7pT0XX2b6Eri2ifX96VqcQUXiVu6tg/xWfRqm2MZ0JimU6+
5gnZVQ/znd7aDdAzSzYFqDbvLFHbRba7RYv+Ud+VHhLQOtrIV6KqxfL7CTlpS7Kj
Gk2AjIUvFIsMtO6ORnkxAVoullgPjr6fiPiP80SBHfXpwfCMUrvnFXnWUzZXZzL6
RMBE85kpMJsrkEt1Yn58ZY8sQgKpCijKL6gS8Uxbe5YxNNz4UJDLNYAZnXII0SNv
sKguaAMeMgetli+DFSi82elP+kMvRcVZmvNDTjmZITr0KZw/ctKq5MKxO7vn3HUm
JxosoQ6AXRL3xyCNTr0tmSfykVkplHtckw314amUGLHQDWl9AWx/G/37AN35eLKC
JgKwGbctdW/1Y2dNSXtR9AZfjy7fSwki4Fdp5rCiBS8EGa80XvQ16XMHnTq6O8x1
MT3u1Q0uJcHhYh5Fuw3DlKav+nin6GEbEUKD7hrGcgG7QmnnKL99Txgg2KBR7wWQ
57NAXGkQ3nirl93iPqWAuEI5Xer3CwTJ/RXL5dpZSpJp+C22rkRvadMAQockOweF
CZOenGbM4mkpXkw53Do5u4NNEquHKz6nrJHNjkCIJIA6ABr6YekGrhN6cUmkYfWK
z0xZU0gq6Ct/qMFvEhSZBkd61HZG6Bb6ajkVWJkN4f7bcvKAL2znhdXXVaMXdfDo
9dbdtbe5kqXaVxy+v3s3xOulTAREU5FgyMMlxifvM0mzZaigpBNyer28Oh9MmvBk
ELd3WYzyi0lFl+mcmeDrQqtqKYsurC0gNQOiHUYmnHE1fX1U3sHmUs1t0cRVRqHj
9uhMBmXLlDH/LY9Zc4HVoDdGBXq+QnTF6uxWlfTtqhebM2ZPkNBcdRMtHyMqB5Zk
kBbSweotNgPuB7HEmn3zPQhlWAq4q1hXNJLoBKboHj1yny+09UpPhpe9fI59rgEx
Ri9zJ40A9yYsW5YKzwTTcKlqCvtJPy/dnczF6YTHP47cgtQlHX4olA3h0WxIUV7a
Jn5Tz6oWTPoRmm/wn2GKxUTkK0moEUgnL93LYE/3xuAdEOVqRxfPlZigs1r2RXnT
aehkriL5Y9fK8JIrBBcA/ZOfW6JquUvgeZIwd6Z4QIob5h8Dqvg/39LJ1jTQ2rIK
k48IOtDU4xfyZ5SCWsodNs+R3Bn8hcldnLTw426OSHVCLS6eMJPQxrQkN5IwEw+J
rD2OnEohzG/6puZ9sHZp4K7BrkDwS/S4RA8cUBxQXEbgGP3BqD8Mxi8/ZINX3iRF
VyRtCN53lB8j7eJue0JDzC2MmdSVo+vvlloB8F4usyoTOBDE1oKuXeEtmgTCL7r4
r6qLPND5g7UrwxDAWM1gVDvppgEavDm5uXOo1cv0wuTkX+fpCDrH9Ld68YhG2dvp
B/DAk42P6rY9dFAi527xLg/luEPgLhuEHTy8PdZJNkGYis1TwW/2nRycZS712BSi
QSnCBohXcCrFVaKBVn0ICgX+3ve3oSrJGGXB25/+RPolqIUnVOjRBVkt5Ghhlfj9
P4SMxiIWWGVLKRMPn6JD5/OfgK+DCyAkiSGpQOjf69RIJWcgIqm7fHd9txyg+zMx
m0CrHSdhaITXkAkkGMGJAOCBmxqxOKsRyDoYbg3Pebyz40CI/n2hrqSSXvNXh3P7
bi+WQzkfoFm/cq31zEGerSWjicNUuQCNQ7Bdwyln3HjAJzP1RtO2aC8sqtEtvTrd
eorxhEKHKR8mVG/DpGS/k1p+416kor85YbiGmZ5RwDVl+UeDmKdk6nDsqZeWoiJp
1t+6L0gYWx3OU1azNYmoi82cdibiGzCT55maGUPJ/ZJoi9YcJ7FnctoOyH3luHLq
k5o3If0Kbqm8jqnxmeMvoTCbopcQUK0QcBnecIELfaBNGSy7MGCiNgX6ksiTYslb
sHqfK/QOY00aYRK8v+xWjoysHv9+YtuEglomsnIMpOEGvxAgFuw9m1872HFQS0w5
mJFlH0iCv9wilwYtZLm2mvCsHHaW3ZGz/3s65Tqw25/fB/A9ZVXzqso4awZ9g9Dv
9osYiqyaIc/FlsvR/WXviNa1kc39073zKvzy45OnIMTPDTrHQ5+bPmNccXLti+oL
s1RApz/GJ6T0NscffS6vMfQpz6JYgiTM/K0iT+EkG0G4v+NAeH69U9sRr95bMSpY
gOJvpkdBtKMiXH13sE0YYQAqOaldXGFr2xzLGEfJ+pDHe1w3yD9wiliBAtuMDrYE
LOG9gNM8Y9mtcRBiHYXxKaCpJJZF3lAvohlTYkhrbWYRT39LooyCU7NowxRkaEf0
6Hmr/mdUel46GjsfJkrX9rCfuDmX2B/k8hDODDTp02J7Azf698XBqHqWgiUayeCA
oaDDBl/rz0QVn0sOc9wX4NCoGww6ooS/KaFMUU9H7EPnxRAHjZfNuyTYfOSbaqKF
z4726UakohIlNxOcx7S6jaIjL2xf1/x/5/nKd4YluysHR7A3a9e865UPkQueS7/8
VGeoLT42oqc7A77uYPt4GUmc5huZu0W7q4m1eNxdXi9LCfwDczs+uN+lSiROUx9H
zunGuhzHFfYazg6Kg4QiWEWrTsuT8hYr4i2/l2YG/5WGbVMk+bFTpTgjQF/RA/Cg
p1jEx1GROcFs/ybH24rO4SwNPT8oxa+SVsikPIcQoryjClRnuJ9wD2MvXr6e/QiR
1LuRCDrV06FscCrEXuR/xyniLuWIwurLgfV4FcmRJrjIMVeO14dhHRvXS5LeADFJ
h+hG51EjRbwLpANnz/xrf5Yem7NkBAKDyJ+8o5aJSwnovtpMgMPivqdN7tWkN52I
QqtiFLFpDoYmv8KNR195FxlTd7nW/91s8NwXDEtrjKpAdpAt4MaI3/I3jImsQJ1s
j5AIAntwOo8IRI7tQGUlPgPJqMS1BzuB0Fmmf3awh/RvQlJ58oycmfkiQeIt/7q3
PwQxsXM5IxWyiNPbFW5oQgG2WHUhzVPmZnRaUKJmT0hEz5saward5/BoBcd6IS1I
tRSVXAyxpHNZQEoieSECasd2/r4hT5TnJ+l7IuHkKSPhxUUS5FcpK7H1j3Xd0tnm
Fz7aKI4ertazKZ2j2pNkjG1sZnAx+PeZiE1KnUZEDOSBTPsAa4WxikqwXWoJVIWW
jtFqFccAXTOItBrpNNn7BqotREz2miaSw249/dS7tM7kf6N0mwYNmlthqAO/rUPF
iMjnZ6g9y80926hN+S53JqyNL4YFKmUbwNPIMETT0BLA1TB42o0kYFCRJX0geCe8
QtdddpN187pRNU0RkfU6TCzdkx7GlOcO69YgQ5yyRvfwI/k+VCI0pOQM576WdOK5
pJGACEOHlImrWcMMEbiUUdHwnB8LOfsANI7BhLJqeA7kXR7L3Bt1VhhJ+hCZ0Buu
5LlA0SIQj4y/y4sMf5LyQN4aP0q/Du2gKPgQbFykALDhPqSuDBqCtfycjwzkmPst
ONGz8G3yRxA8NnkagO+0kQ7XaSWAkgTSTRR22bNyM9ZUZ60blu1jQ21WsJNq3aYV
KoVDO2NZ5eqaj1ohpZIoXvHGOLP3CmdBjZyELcJ5KQWCGg2VIQmSam9nAD65chOL
7P6CvXSU5NTcsthMSVLoeOmHvKJ/Ci82iu5+ziF4EZ/5jPP9RXLRxAYCHx5Ut3po
LgHBWiNOCV+FO8Sbsv560RaG8dJy5UvHADHgkjq1qTcKEu0fc5EyShZ0uxbAR2MR
lgEBNNdd7rB+x6KDuvmAxhT2Kk4+4I+46yxa7MVAnglI+ib9+7Z9kgqAWMo8UBA2
neeBxuJl8f0TH3PKxH2hJLX2dvjddXVu5kA5NDzJ9xoMzNuDqVJ73zNCV5j4gN0j
ubUjtX8APpyTiPzVKppN+R8qYH1lr36omJmTdfF5ERNadTW2U5pIAVP7fIB+PWrl
+4W+i9TxKaOzqNm4SIqJoRZBArqVADOFS/8BgscVX9sQu/Q0TBIsoxvW1FCOEzvy
4LaxE6ZBfUl5N77nArRI9crO0Vp8fazBNHBmyHhohwetq/wj77JyRMnHeK0gLW4/
VVqJTJeO0cHxUtiFa+g6jqbcaU6MPhCaE7jQx121uZGL70TRgRyYlrUZLy5o7btK
S+mba83Rv2VdqqqpESxnm68llsYBWHDK8lb/0oESdGEG3ILTb17gqP0bmxkScDeq
9H2GC86waX4HjzGBJDdchEBOZ9sWFB7CMbVleGBdgZFeS9NzjxN8wfIjCEPEvLP+
cXtIFqMeUsZbwhBZS5BItA3QdL0hLkge9hBOJPKuXSCbEvGoNN+dtC+GjHL9CKQj
8SHzqMNAoJQXWUfVTpp8OWzopaWnbjxBTYw78ueN6/Wa/O/peS9q14sf+LcUYDnu
T78KK73aIFFhyDxLhkZ+b/V4hdB2BMAEu6DONikkYW+gukPmrZjRkz7MXN6SNdpG
m/t9u6IYDQEWgCwyxRbVTzfQGRHV2rBgZsoeNLbLrFrF7AUp3cBeuPqKd0+6Wx8r
JPO467UxmqEhGugPDwfnwRrp89xAIAFV+r9G846R9AP6Fa8QWlR5bcz1S+KXFUR9
pX/MaR3BRpPCg+JblGU9B7oR7IHpxbIju7oiL/LpfY3+iGrafTT/qSZyr6rf+WkC
pDt09TTjMXvqol9C4xxa08vqnFoF+xHaiBnYZtd4Hpa+qybfWIee161jPkgO64mQ
jJHD0CsrtxsDNFThO27+byvRDrUnmFdVCzEpNrdoMGGp1egbOyFw0yeR2aQJ8cHB
B85YQybn8xJjLTp7x1RTb4bU3tIOgVWaG2q/el22MnNGa2jLCvsLDgHQkfC8xNSy
UUeACKfvKavnmD3ZCchpKJODsQ4G19z/QoMmDwBg2i3u1tp2ylRJmfokeHnnuFT5
1zqrxVfw9MQGhycrwytFZm7R2MpKkuUuwhUJ7uyVr0sHtHVyXyvDvzwI1LGiM0W+
UV4oCzd0NMqxWwix4BF/DU6UH5NJzpWyxuRY3NGFWO/7mMXuZcRtdXGKIHWEbz83
ySVaErG9SfXB+yCZk3Ao8WAuIoeKnUyYOM8V24fmlzTyxASssTpqj+kii13Raa0S
mGHh19qGBKrlsR0kujJn5lvwSIk+v9yitubE1wkCwMCWyoVXr/XV/oY8Xoi+cDkJ
DkYfLKZ2aRz12j6ZglRgoT9EIsVkPBUfCmAkh4fVzfmyWnV36iZR3ElPzlelzNAy
hS1LEbQPKjy0xp8FzdiObzLD8bRKUXDWvWJsAgdLriLtQPoK7QWsVI601b/irJRp
yPyDZLJLIeEQL+kq3S8sH5ZzfRcgwfVgidQaqVBBUFSNDsKTXCa1Fl+phDL37afm
ef8B5Mj54Z2k+L1mJgoZK9D/EiHwnY7pijtWcmrLXiH06ezOIX7tgJmSqXShQZ3z
A0+k/qTTLBADpkDFdHiflvCz5SNr763hsc/O1agcuzQRwqe3Swoe6HFXbhIX5udb
/RiF6YuNkQfq47ljfvQL8WUbxZvVGvOgjJYdOUq05vav9yZ2oAINTsUaC+YnQ4tO
Ik+xcyxJIVVnHB8pS/+HmFzHSHPgPfAMPGiF48YyVJDopBGh1OQnQcAtOkYCXYpH
gROUC46m/jJqoPEJs9poWh1UhirzcVMIKMfsVrdH8UNgFWhze/F5WhtozOFbqkgr
RIe1JZGxwurH1m+MU/wv5uptiKSEJHGOUyIp1yNQ335nZ7z+MGF3N8zz/iMY68p6
j/xo518Sk7VDA5YU9PftXTAZNRc9cxFtbXS42UWLxYM+trut9dxqrMF/M/v7qLZW
YtmeULqvw7DZeQeAQfmHXM+/vPlrzfX0RyqXJn5KOhqlmbq6K3ZNWSBtfgHHJMkH
tbBI51hJbVJas9d7GIyRguQvLaBstaehAYpcLmx4hoKQDA1W+AfDvptfFgWqPMhe
q1lffesD49isjMwcskUEjRdD4VGuWftWmwRoKy8pfwEV4C2+dXobnu6vjJwTosjX
h9iIJeD9SfEXbqtsgRSQrfi7GH43s3udULrYXXckXppRG060ZGJ/LTa8bk/ZBCtw
J8YwJmqkfKKhxRLzHXpBzVVSeam2evxFqF1F5nKizomZReKQQdaaKAA6nQIQS1oz
CR2IrEX9TIVsIcJb7Vi8aQzSzMX8BVC4VJGZNx7piVx+DG6+wajgxELO9+qDJvO8
ZLq4QTOoo1XxzIMpslyn+RaQJgmJ7FdzFaorhUeATBG2tN6cdikgNpftcgDR2fs7
cP29Dj8DsR400AJFZLjo/2YlzYjw8eLJQpYgV12qBkaDcJKOd8bN+PBuMr39wQXq
IAy2c7UYgdf1ebW88dGMLggO0In+jAyfg9P9HDpIqKCFjlbyPUTvxMfonVPmgNPf
FB6o94t9GeQJOJFxGxnk51ztrdMNVh35odap1o0GcmNdYseFUeFgFwQjeuRLHHRG
a+3+9R+0ZH+0tz/uABqTJrUotFkzkAmiSNBHJAkKKoD0rrFvasM1pqWCBVohsJ5V
kjr4sIoI7R56O4+ERDP/9NHn0lLoO8Dx34xzrKT4FsLdB+kaYUU3hGENSP+qbdmY
P3Jky4YgNcNNKBCGLGJtYezEEB158rIa4DpKPcknEG8Q/1l6M0AopGkU41WlbJrE
vkNEOGTjkpjotFFNe1fokJ9/KK+NmoCdbsdKk2qa1zOuVgkvGVoPqdYL4RIrw0FI
wb0RsZJjApoSJat74oV7FkOdmK7vh3x3HJSXO7CWgQ1dLJ479LOoigC9u//ea5Tg
6v8vmIDFxQTDJO513/6kYBrpRVJ+UD7FrnlEGtfSMV81u8Rpf+kwwCFbYjVI+cK1
w3gGh1cAREHXCvbOqledtiwo7i/M6Hm2Zr4GAB3426vKVNK3GNJ0a59GE1MEZexW
lqAowhcFRPGwW14x/LvdCukro+U33WdQ3sllrJGcRF5MbhNbGGiGmVkKdAZDir8K
UKbSCOsVxZ2MMYddq9fbHOGw7C5WykN9Tpvz3wvTO04V8IwgK7jtBN+KgA9tiPdh
h6b+cwoAu9akT49+lvhpUM+0i46TLk63KLjVkblDdHD1H5VxeUkMHHVu1pPPpXZt
JpwmQFB+8541pFj9mennsYqW6SPM8kSmTU1sZB+d2qBpKDhBi+DDQDRbFlVYZxNW
ufmVoGcDCrh4YsvF4Xa0ap9JwF6IZgVVVBZn53G/abA7WqZuZ7onRDd3TdOEQUXK
EL+r3VgheQnkI95536lpWV7+rYs4QVDbHPQRxGFbITkkINq46WCZJtOzl2SScrZm
aC0VD0JCuJ0fN1EVfu8WDty52Z6Z8GNcP/qoa+jL2+jxCoMJ42Gtndyi+fJtINAO
GIsyMeUEAg0EpvM+L19Pqp1Ql+0KQ6adbxNb1n10ZCvlk8WSBktYOegOREFrxNo+
r7S6uDn8h0OQALDOlxZZpu9gTBrBFOhm01FyUeXLzVi+q6qs9k3hwebOopPWK/xB
fzE0d4FJ1bX4B6Usk21i8EUnf7UM+WHbl6KzqxfXL7g/Xmhg1SG/ClLGqtyzJtBE
A1Y/dosonoCs7ZQv7xbyYseSjoWDZNYl5azRcubi/o5HokKJbQar57DoB0OZkUS+
td1P5Mk8rdCtfHd3Js8/rVdeTYqopoHN3YXpOjwj/6TPv/5iLkiNBTlrdxMPK4ve
agB2ivwqhwTcHCWll0gq+7yGvPhBC/m6i1hkgGAJ/8+pB4Wfac2H0IO90idadtI8
8JQwSiwKvXqPRhJBI08JGohIh6ZSmdSkbVYGPwopWwBSiapXCq4eT3zsuv8SlZMy
2Iw32K0zdJ9avqgpQwNc37tpQBHAU2ZlLcEmMJ1eKtZdcAzm3XwkkrXiYskRz3bv
4+J4A18BoFxbC3Umd4dH0G6PKFRingE3j1qrO9/FZTOp4rzidFvIJ+jfNJNFP9PV
AVAzEdKupCA/qhQU268BLOMObY4kZs8cDrcVWFlNR5j42JgkawgEXBOB/eKMqdvr
dUapn8vJqUhMSTV9wusk9KayYMN9Je/tU1MujXz3BHt2AuIyKmweHXJjZZL0prF4
O086HZWdx8a+2f7mz/VCDtvpvQz+vXffLqLe4x6/R/b9xqx0wMN2+DCCAMPakS/y
gyBtw/WdIITXESPXzT+Hr1JLiits8DWwTGeskONxr75ZRnAt9d5tjbtQXGdQzavC
rxo4sxpLSMM9u5UvPsgfTCbzkIR44z+7g7QTYw1YEJv4v/6fp4KR0k6+aVgoDxFP
+cB5l9i2NwGfbVKAwI/dbMoMeSvRKZyQNAATeE228h5t7xgnhOwHKd9mV3ZW3s1W
05rM1sia1mic/hrTh60ZUW8IYIx+KRrOzqsHTuR1Ih5XwNqGxN7nDzDCuFywv7Zi
52P+yqfGrAt8cplLeXVXfCLeyRUKf8qo8WzPXfw925NW/Fz0enQVhac9QYUXHOAE
tzqYsoYdsakMtf+2oHtpEhWNnLJGI8ZBDdzcAR/Zh1fzlNWPOmQAq3/jt1GmBzqd
XIVMycVUlUiee3IT6uaQBSSbhuq2eyLOTfUREP087OHDplriDPzZYhbX1M3OXIKR
9azSEKGje44mMFNaScHRG/LTQENWBajE6J8C7u4OvUzXKiCotNj8W4JbLEoqyEf2
qyBSGUpJhbSh7NzddpUcLNYVNsobD2qG8XXdC3Dgu3lC9LVjkaTORFp/1GXyshiP
Yqiy82YAxiBB51d3wpy27ZVqAsONdqYqMTcfls0EIz+TE58XxVS2w+d6dnYoRWz7
NN0qReY0/rAa7BStenR04w66yVcCmPFDp8B5eHmTDPUIQ+T5ctOZKbeHovZeWEyo
khGNZd9tWbEn2ZdYP0/yoOmeMTZAlikBE1+Kmk2vi7dtdjahywix9bi6xjiN94Ng
1wuy8np3WSfHQDC7XQF77j9xCUf0XTcMIxcwwfRrUGFdXaI0Ou/b61G7cp9MKRmE
qYAQ4wCvSv//AInCE2VZjLxbDNAVXmOqSFtR6IYCjyyIBBbrjKrVtQR9xtZEi4XB
u1ATi6GdU+LP+wd5DoCqKXdHOTHffHXZBFUJxf2I9UAffq52yaMACcOE19Y97+Uo
OPsXKzl868plfT4kmrOh0yk65r5sP+43Nus/It9lJNmmB6SrXtuFo15RDzYZwz8P
YONLL3rlhn6tUTwNh8i9x0REZ0eUbgeGsz5KktuEQqToid68CKA/W7NaXRoWV1EA
Z4VWxk9Ib7/4A6RJ7FhwaSblj55qEi9/54+jWnGDIFW7lnaTcpvbYQ0r0J6dI8G7
/UvBRqF1TISkHzXYFq4PbnIYBpADMNUeO0HfrmTtovcxc+UpW9yV8kR+yVM/b6G7
A/6vDeOuMecwKFktVi97DgbNv93oICRaIoAF3vcFM0z4ta+hCQ2ZvZC1TKEUFmSI
KkjukiggXqVKPzzpfKU/JvYzMnJx3Ek/qQxzfTD4sBnjNQhKYoHTFEUdCI5upwS+
FX300dkjAe93m620gCV3NRWKRHmS3aniXJ6Evf5bUmQ5I9ODlSHlLJjBJ1Un/dA3
z8q1SSlmsl5MZIcH5GqM4ogJCob+kgvc7ft04FuiLFxN02NUJDNYKA3Ay4XWGDDG
HdCh4zU/s/C7pmgpzjkYUvjnBr4AxVyH8TaLylhJ57Hld+vMaS6kzW1P34dlL0KP
DKDObZGrtW70IA5ZiZwG6fTJ64WpuCBvUMHGZ589Z+OfPqut8qJtwsKnJICiUJxI
tt4/i5/mM9U3+0j/SnR4cAzVeUQWkjNGgs4L9QM8OikLDeT2fTkGwbdGx274YX72
0/8inThBj4WRyrJqUGsXHHqfiibfgTb2tabISDOK5JIQ9rN+D1ZV8qpeMqgu7y5J
BCnvq+ziL571Wuw7tMOjupY5CcyvhRx8MdaMZhwiYX5SzDgloZA0uYyqtaGl167O
XImYTUvJQZ9tukJwJ126P6L8Nf0FFmmjkjCH5cT3QJ/fHgBz7GB8z2PRyL/3eg0t
DMv3CiriNsz12s/yS9QkUi8A+9qLEClLdki5EjO0ZznILwPR7ljsmqwXGMpw+QnW
Ka6/DQ9n4RrNjzZF3vpfO+aT2sbFMlMHn6VNLAwl+fBjR17vDcusDsQtFR12B3NF
LWxOhK9NiPEbNZfDCsCnmKYqqWHZTrsmnyCZTfvEwqaVOLXLgGvvmJQTBr4yNYMn
28VX8GhkQTqy07o3SyvMlBhujcsADMxB4H5qTLMNvyM1HAOfgytEWRjpFU2hIZCJ
n/eRJZohNQVFrDV5qYuP7RJDrB/HNNt79FIpyBVCAa9HPQTM/A9hSCqtEkmKrUdX
RjiqZo0dnK5S0RU9GwtzLT6hv9Ce1c4iyMmLvBgylBJdIVszNIw9ZNt7yOei4GEs
WmtZWMBFp8HJUf/wvs733KZej2KADZlfjcb6+HRTbm9qr9/NJiDQXq2mM0h3YFtd
wot9C0SOmkR1N5nko0T/bXCNJktNAil9RxncIb2rxVc+7le/EkZy2ZvCTwk+v40D
tffQrJkKYWI5h0YxZeaaeEMbzyhBS8hkrj+SCQ2I9PGyKPSso/GizF5HoToAk/To
Ea6BccihCz4a23hO97Ov0qUAxOFcNUWneepNx4LKFmAqjnbF8bXzhYcWX37NSc7l
n2kl92DuhXVWSF8RXDPYG6CCdFtWoXGfrrCK5m5E9Hzz/5ZvPeQljqdYKJUpBvSg
uxs287aqECF1HKSblWY2C5VVU7jnomnXVJpA+5f8vvon4bbpewEZt7QPharpNcL0
Gxseq/0Jx+Hmifa/BpgVG/BzDuXDNjdfDyqB9iqrBqUvI32ZAqv66ugnppqqTobO
2yLZ+VLV9Q7H+FSMiw4Zs+zY4bZpnkInz1yZQlDa7oMusm15xaxQWycQSZZYFsk5
tF1AiIy/OIAP/IPiH2mB8AtkcXekFM7r/VJElaY/4235LjgSD2FP+R+AiqOq0Ber
XLf1Ax8HzIjeGkx9NOPassZyDjwcXJ4dJqxkIrrTY4WWgiJRInJhZDnrBB9fvnli
45ko2QWAF3XcYnj5SnozZnXacDr11BtEi5HQeqCBmpHZWAgdkrOnKnBtEfXAcerE
mJp1EDUMqQuvPeKKRXt6OUtD7zy6WapSKLLRwSJ3n74fgzRIiTqncjUhtyVjAjB5
pUVrwyd8ytRrwtCDA22BBqk0PuGaJQNo4lg+wzBRvXJK6gAzKbywTCiKS7qwEan4
PSFzhmexALMU65I8zT+w0ZBx8QBHFIGv4+Ov4PfAwr4vHfmC8DeUIW9pusSElyeS
/gjbAMQ4tpOEb3wQqGVEaaVgQtGFi6nogT5naAmX5Xhu/WOKozrcFLRNbs+tHLkO
+BMaKN1cppAkXPfDKIkZ3YiLdTp1kIaf+abgLBuvWiV6x3iyjT6R5MEQ3n2Jx5bu
Y5l7vxlCE2du3y+bBX8tG8GHPRreN+WDgxc8W8/fSqNDDHLDEPZY0RIZ/oga/Ffi
IrMrKf3uLzKoNEsi+/t0DgGZj22M3ubgJkkQEyszaD+wI0wYi/Xo3417sm07t5jF
BbCP8D/z/ObiIkRgA8x3BqU73gMoe15PaWii+T0XeQsNNcA9G3skbIMVETs6bmW0
XxNr/4jiN5wkzb7VeLV//8Q99gW/mrVdz16V5SQ+uABsSyBFINFOwKn1P7684Q/8
BpY87u00fTEZTl4wT/YXfBVyMTY/q1Nbs2U1kT6wpo+92U5AG0nhEO1VCuE62qDY
QsTwWdVkRYnFK6c/G+IOzwi7wHd4me7z18zFnkFn+wGMDlq/VlBqidCbS7Sb6MsK
wt9JUv5XO2aeH+LZFNmPMNmubDW6y/3wsEgBtBFvekjcpZlYHwlk4vUB7sMcezT8
9UZhZomUbAqOxEYiJZ0c51v7aAbUzlzpBd/EKEqyMVDlz87OhP7rACte3gWuP7ql
3VqmGWXhqp2OWRhkI2cCjOhYJAMEHk/xiXx0w01PcQE/jPDVJNneEJDCkTI99ICA
qnEzAQJkqfl/MnUwwwsW+5FeK2tcCeB/POibyzWI3kty4yl4K5NS9C9hcHJZGXwj
GpCxFRpHpbfnWNY2kv3s1JHP1fxAXD7sZhxNEHtQMphdS0pzl8GpCsDtZr/llV+i
YYgDlwDJOD5v7emmO5we1fP+sVfjH8d1jNabgODZCKgBXBgY+Pr5QPqy9GDGi/qg
gl9Zn2gFOuepNjxHg7IRJUexPYrbgpVPTNpNNOlwsWQS28vsEtoDuiOzrJP9Ao1J
wmoR6VcvcWMNrt19NNJ9lDfpR7/BBYvr0Fn8KvGsGVh3WhnXPPkqXel/y87btFrO
NHA0o83wrXpzh9h9SORr49KdnN+Vnrgv6P4XDFBavzpb492yWBQQedeMdOo9Z8CI
3lnQZPJI6JrlmcKSgmzkIcRUO7Wg/H5RhLHKrSZ+xFU2tlospHE/mR1PkkRfI7lM
+XpcsuQaxDvZG1IFdVG9LzlQqlQV6MM+JtEino1rqNEm6KvBcHfDzKM4RenBXd35
lx4fXU7E/pJhKDHd0cY8fLnpiwlggrizIDfc89oDssHYl41CBqRUq145jjh61cfU
nk5nVtwV3NtGWfuOmjOhWwUZims9vMy3tkhHL0dFqmLkscuO8//fxvPSY0tnlpGm
bWsLUW+mxkTL9pOzOQSdiFzNIruCElH58J5v5W2KqXejkQPig5Kv3qqCOlt5PbRN
yfrdCJPEN8A0eazBixbvhkxpusO0xdnKN4ei67p7jfcUmpgopn+85LS5cH1rcWbZ
SoPRaDOzv/PEytwJ0qLyIGEOeAsns4FF+xXjlUPZSNOisIAXIHKqZYqGZnWOwBtS
CLLQ0gLvi24W20dHT/aY2U2hyIYZWa0knfN0H3nUX375dxrozqMt9eS6YeJ7x2QF
009HFLgAZiTKBS91e4JW5Mk94kgsn75OWEUCthUedDNMb8xeiMbkhgVmDDsZLHHh
dqBV55+kBfd27sCzGY/s+1ACQU43P8YRmQ8LL+aJX1aHrOjVACrkXZukBzQqv7T9
LvRRR2kbzKxYdyETyA3whCscXqBlaGzGYoDYiEB/kFzzQc3uDJVAgnHWAdpik8hH
v/8RrOZNVbTpzGSZQIF6R6WIg/VmSekz+US06i4zbq06BYdWXl5XgJBzY7p+CBZ8
tDt1BJ/kp3tuWe4xDre5Z8aGx21h5LK8KWRA1MfO7rJRhNwkQVD2dPZ48dtlxtMI
/iwos0OmGClLv/dbsgJfoWRRXlprfVOZWroLfa5er1ESV7xLkxdvvc7uGB146lJY
Nw0tgu1Da7mu755Yh0QSkc2Q9pl5dJRXlJpAmo3AEnxhIpQjHwQKyuSfJOuVD3/z
2fmkSfvEXPoVgk1n0YylSuK5M4veibEnAC7jWNhBvClY//tTCA2BtmMFZ1H7mnf+
REwAwtwEffcLVsrnMR4Xh1owSHEhfMzT9clxwnSFO1FDOaLt3joCArqOdvhty4BB
h7UjbG32zH7kfnKa2OHREW1yni6aJ9jrO8CqiFoYJ5nHFGzgBS+p3D0NvqQ4gaJO
7tWLO8n5ZA2XaR4Zj+0/2WSY5iydblepZe5fkAPA5rstY4u7cy8BIBPQsg4y3KKY
h/v/Z+iXuVOKX7pi8TsmRyTCe5jITN1/Wwc+IlF6+yS12bAZLq4ivsLG6+JTINjQ
F71Yb8Av4K9w+e7ZWePDECtolVEM+1h7hlaCHw7SAKY9rhov8uNrmMssmSFrCipd
aSCbkEUQTxaTdhnlBlNjjvTWGROPtkiBwnaGVgi6AKUrS18zjiI+NHsYxQ7asZxO
bYlHAQFCx/6tldKj5FIIWPSafqFwJOXWG3L9io91OoKpatShlD0lUdwxk+jIcM01
qWyikh13gPnkmJ9VuXK/krEqIWpCfqeJz3+1BZm/mm/V1xq6zSPv5ps7kC0rURgU
gEDTmwebani9mNSXn9yP+SRdnb7E/YTLaaxEfHbUsG/f3QanBB5wgiririp9Wa/h
Jkk+GzZtjlSi5/twzUTMazWUEcULtHYUNNPnr6j0xvLkNJuwNfUpcuhlaML/HKkS
qXFEMmrqjD0LG56QbjKBgBAI2Uv+RGbtwLDv95BLUJZl8cFw02MwW4zu3E+bsu52
40mBuNVI6AvXL4pJXig2xoFaFLCYEr6TAq514Jq+LLypf8o7yIM5Cu0sbbbPGBmd
rogF4UZ0oEFv2NyDPO6/P5CGkyPcjAGGhTOX6sueGOSxxojA135noU8sp8DWq3IS
kh215Kc7BblqfH2D9vpgDAn5Ntkv0aDB5+TgByiuEvzvn2T13P9TA/j196oy//vB
H9nSTAOv6wsOu60Rb1TH8csDYuuNa0iH6zms0Mwzo+a3OZpvC9Z8PTf1PFMF6gok
EDtxG29GAsK+xfaavWObGpPRJ3afLfkHVTn8m5JTZzqE9hs2E0kBC9rFv9Ea+Tld
8ro/4fJtS3eHOQt6Nw/5XW9PcaT3oLanozy8ULfdm1BINM0ZNQt3cNrHxU0/8yj2
4+Vjg9K5Iy+6/SOCIPIAcyLNIinr2RHaWm/qLjrGgVsC/7XBM4nXjy3re2+BNc38
J7uFsrz29hnd5FOoWxaot9sVKO7mrmZAvoTPPofiMq0vWf2nRcrK51LL/RzSw/WN
9Qjw9BDUaUbnsfAAUGmbIYPElennWJaeK0fTCimsT96tPXmyNREDIbJaS1oVHg9x
ukvGT4eiExYvmho4O1EfS2katxaJsDcv0Y+mHzzpYjppgUjzSqEkZMnmz+RwaArm
U+2YK2nhefaqxocirEDXEY0TQxgiLTcnNQmq7dR5hBCLB65SBLqYK8CllQ1iCX6d
YHLF4btWv+bcRMUJbBkr35jFHdVMyhM9EcpB5r2iXbKa0ZKNLQxandTe1xDLJ2FZ
PwZpegP5XkwUlhN/xejVaQAMza8IiR0dvJ4kFBFIKuApcNA0lPGIQqbm7mHWV9Bi
WWiozZ22eVO/RwsiUWCY3vJrVNl7brs3vwVS6gsoNSHoB6M4v6IqKiRfAP0PtGVi
txgOnXvrNJmRAZ1Enk2Sybhr8zSwODmrAtfMyFCM+PgbqPC5H8d0TrjZwpybuRCu
wcVibVkELrt5OS/8bKojiz8uh//DIRTNnPBbW/+2GoeC46cwtTu2+X7W9BKP+VOY
EExg14oDFjShwjMm+vtmiIZ5ZuKE4xL9GThPCsX9z8YhgTmrkASyo1VIgG+1A8IU
Ab7DI0LkbdaTedVwA9VcPVBIBuNIfLg+PmtFMGfNVX7CB2onNUDSeE0vmW7ABUw+
+/VL37oZtlVYUlESpE7adeyS1+5fj8aLEPR6mH0f7uNHqNBtkpem1O+WFhB9EHlL
JjQZD6z3NGyd9QztWFb0/4lTYBfYPnVeDE0Rooqr+1BsIahbmSKTjr5ATei3f+vM
jpJBUNamryDREBd3Tdb3veKpz3ZENl3/Q0Ggk/7VsFIXsPjOHzCVTFnHcIuiy6aw
8pne0dJ7jfcIkYoP2c6JcBUeKOZyz6WMPUmsPux0BihUcF//zJGGvxgk3axnCp3G
gIFoHIazEfcaRIeeJroJGiUMR3rE1S7tQoXFrs34aknwgE921kENqPE10Pyss1bo
S/0blq3UYhtANIOVXwJ2KdBikYw5GktR1gaAWHkljdyMMt/4Hz9RrLBPTwWIe1sm
UdVk33vc8Gypv4Yqwr/YYduyWHcpix5Qsk+MyZ7caFBnilQfegD/wZOwXETNaghw
vj0SjhRqwTdXn7Le3e937SC54h4WRMO+srUWs3Fn53iMIeJQPbYAGu9YxI/7oddm
8CuX06rSeQ1Z5mZvDIhGfId11ZGSEgpZQCyrpTc7uwoU/P1ywZ/baE3BY+lxUpK4
TyLHGh0g4EWWw4rGIhytHg+/JcD8qYXdKLS5TLXwDffgKH6XEr4TrYOQ4H0r5RQv
c3F6A1dDl/kPY4mTHAslWl6lUNpQoLVgtZqLoH0d8rFLYt6bpFOOyNoHKrm+4OC5
f1YTSV1iuZGa+DWG5WuP4tYZET/XpCXfSlsKXbAEuLzVGQQJ1bnDajXBFABr5EOw
MARmKZwqvFTCp0ug5+qex04rN6tbtLRlJF4elITyjTXSSGtBqdrg42RQGuC3uCBg
4ouL0p2zJ7CfHexhMcoxJBV3YWa/pWgxKGSDZzQkTPwI1YKeclNMi7nLvOKn55LT
Bd19mpqmowQa5+5WDoTlXVmDDS4O4vuvNmn6HFZ799PYcrNTNQ5/xwpNcRGBX5kr
WEFRdjVoxqBs6JdgVomEU9zyoa8ymRKpUsGuXfIsRA7NEg88FpnaJBX3IBZwHsSL
v0h5I3VoxBJLmlIk8ch7DRG6JkFYpGLtUA3IPtuHCzOKpVYgBVd5dLWcYHys6dl6
lYhbB4GVHoGcYzfh5/MRuATkzAkfs0SkpJ8W97XuirfHIztJGUNOG2CDjtBlHt+J
uKDhFnzOkscPFh2BQACEkWfHiNWl7v7DkOpmCcvkeGG6noo9pbSK9NHZ2BWuJxZx
pHCdcPtQMBlTgZRETYr0XUAnjaRyHZovzsf8BQctP+TfvBKhnzk+lYFq522SRczU
xdfjFPfMiFcMZ1Hoe0M+I17O+/Xq2DAR4IFzLF48r9nGfC28Ou+1QBPiEmXSEEpD
oJN27gsSmOiOPryWf5ke9LicqoLxlIjF5/ifitX2EKV5riOnL4uNCuuQI13qtvmN
5JZGs1tyj2gZrTfEXIlb2YlhV/nlBk4JIAAcBHsK8ozRgiOENrA5i6K8+HPO35HE
Z5WKZIvXzRjSLdd4R+QQ89DWgpT1JH8VsEkHc/Xa/lSj24CSU/UvMaY7TJXgTjK4
4yIveRYYKqUocY25aDenV2dT6rD9cOtZOe+NtW8V4HMeWC6fxFI4WAJFeouRG+Ck
vu7SjVZtvu40PA4UkjN4aQlc3Qmz9cFnmZHwkOkwQWwO10NUYJQ5ouN1fZOFwj09
Vj903rYP3UMp5iZaq4DhuAEKx4nCNF3d1WbzyPsCU2xPuvRInov7YWqTI28PYSqH
/wyTxIMWXzdZfsNFeBplDITuMudfkBaCs8WDyZLLzIegNgDSFVyMBCToKUqTcgoo
AoHtSfeGhU8wRdhM8VEW5CgDasLfAt+QW0vUo4C5qqDw5RLC+SD3Z8VdiJXZ3do/
AMQZYw9muMIIobDtmKsV6renEVvDh6HYtEZdcwvP2f5koBHpARXxj7JM55RZg8b6
nHsN0Kehs5X5pq5TUQrLC2olmxMYwW39dDEYxu80M3t6aQKZ7yogDC3XC5u7Zib7
vh3UCvEX92cLmoRcoMAchnKhtZ8ROO3l2V6zGnzB7X0x+QKeK8DAiFYsy5/e+S4X
BEhbmhrb4RCUCXOQGQzBmRj7DgV1uPOu9AG5J0WITL0bbr1ui9AfO54IumIa5BhY
R/YoWyP2HQosOyc3Lv+FePlpW/+vOqkcgrRug8ZX3X7AUR/1ezFi7+ZtdFE1PD+u
qibReiHtxiiGGw646QHXPoLPesl/dAjuIHkZ3UzRcRQoT1qOMeTTx0h1CDfIa/gj
d5oHZt5g3FrHGv93PPmXZNhBXQhwDoi+LaFGHgadoURHo3bTlvP1BDkRBVOgIFuS
2CUMtZjyYu31dvgjm5b6QhvvVFp1IY9CDAy0NyC5g5DHeSgPYUM+/EcGCVxJEvs2
h+K+zThA1AXvyyyGmGXKhyGw0HoauK0LhXa7mk6YomkquLcL27Z8hzJIFm2V13A5
JXFo5bEORGE9IsbAUFDw2TmEm0HM6qG5/qMx32Zgl5QStcl3Esf65+eb4sGyG7X0
OIsFkYo8Mcr92S7K98Bsr2oOKDSTvPHPLGrgOozOVeFGbPHSuTPO34qLD/NCxqGj
GLL5gzGJ48gr3ujmO5IZT9YSGUFN3o/v1jXOpL+8j6CcFMFUir18W7obf9r50ovh
HDYksuCpCt8UlSnGCg+yn734ubP8HSpwMBJxI1tL2i0NCooi7Lgk1M/Hha2Hbb1A
u7WfvpTmjjwQuapuqzRcWJBvzt1z5GYsRg6ER0d7eEQs88d6AgwQZSrkqg/HBSve
liY4Z2vdyHiJ7NzmIQ3g4adN5StUvggJTVUh9hTWzW8NOwCaXjd9GLqRRGim3gSE
ZUEB++32Wbt044llijYASLE+6hMsB15jT/c0zv+17EY4BhbHWpEO5s1XXH23Jvzx
h0NNuOQzvMCrjZj4DxyH/wfxqeoM+uZeqd3t7koGSXBugN9RbaZWKO1dieUR+3Ic
oktkW7EqNMUOaufv6CghhNAc0y8A+f5VdYatbEqpTjowNEg4vqijbvNi2AKtp8JD
PCOAz5boFHkriGq9Bqbz4riEspZrOtQfgj+asuxDGMiQzJ3gifhxGpMPLDXsFyTB
/4FdgHYurrK0SMUee7Ngz+P3ak8j0+0nPaX+zHpdU0l8o0FQRCn48Wtf1OSXBGfN
VIFz5xHDs3VPo4JZsPvG3E8yvUr2izw3JqbFYnNiNAtEYrZwXcwyeWxx+o/U3bjl
SOlVCatOHCR5u2P/w9P+BeCdj/q+5owvxMdmS4NzLBA1Cgf+H4K2tfQKo2+lFA7T
KKf86et7MRjaSrbZ4GjmiU9TLHIY2jFhino9g/C7NGlx+gY3GeeCc7c0hKljWMhs
N+qv2LTJq/qG0y22uLLSBc0RtGavmw2Q+JRpHABf7dje77HYHo5B270kmMjzD2Fu
OMgb0nEzKNC1qQAnmzyvJDlK337OSligUVpgy9H0Fmkc3fg0Ox2IysUiQ4nFnLHu
tsVcIvjMRTVfF1VrHHSTYLyCwSqOkyhjjrLnF62uoXM0NX5gH7E4eGDoKrLsNeKQ
GihyjtHyF688VjB9ikIO6EmadiXUy7HP/3ywQZc4Ntvwn698EXl3iWZK2+shyTR5
7EKe41uOxkE9dOahQ97vtQY4n4Y1F/Jh4OH5fToG9sfEiIBpiTFWEZ2CjeMNwgZd
aCNptRK0D4v7UUP35qXhSozoZJyL/Rm1BNDRWZ2kR8Qm1nZV8JJox/3DvhBHiBlu
5w3UazqbgqS66l2rENKLAV+Y5CUaax5NZoB+HdA6kI/Mhkad9c3k/H1KbJBcmSkC
AN8L/8fjSz3amZVNZAxzl+ouC0zEkouXaVuh998+xuVm7ULHh7gWYuLJYw3iahPQ
V/UAIcibFTKOO5y44tV7Z1pkBkdTG5Zveejs0LefmzPRI/2IMHO/QYPMAIdZ8BMO
T8F5M2gv6mxQ06fqEYYUKVDjuG6t/MeeywiJXhJnWTRUGKdZYz1S7HqNIEf8H0Pc
KcG1cD7V8jBrwOZZZY4KfmqUbDIMoknT7fHiyHj6ViQW+6hYu7ANWIieNsINm9I/
X4KNJB0Xw/PcRWvOCoIqWUzBeVzfQ4fgZm7ZfZjQgd6lICuwaDVVuGDgap1yFM8+
inGZZ87H1hiRDkWE0w/hQYC5iI8GWaqKdIHbV+CjO+vIVvt5y4jXxEkrr4T60tpE
6blIiWZOT/Glrmwcg2PWPy1TsIlY43zYvUXTRa3B2e8VJ5XQ+6bzG5S7bt/VPkkE
2t4dI1JV5vJWafkwiVy3hnja4v+AbPcNdBWyn2nQBY/jOhMVphBHQzbW+8Zu1YPI
njC4pINO8rfS+uYClIijuNqy8aUdHovDl/Z4P86Dnw/4XL+sAuo6hDgfZu0z02tV
Qoh0Bw0Gmosif+nnzRr7dPZZYrJCq4iqjc7c4hnxYF4iXxfFQao9Bd55QkDCh02l
Ngd59ZY89wa/DoiHAn9LcFhrmkpqQLtakZG0XuD0/NWswUHAY9YgWdu34f0vZJUl
nrYEn4UpC9wgMtI0XUIR5uVa3R7QR68wYxfE3QigCUkEOe8fNl/FiAkTez2gsOKp
N1TR7yzlNnUix8k4lK5BKjxWNFQXJ54GdEU7K1uJgDcqOmrOZIMnScEr7qIO+NHb
xrJzlTq4RXcgov23dYV1BiS1TwtgpS8ACQz9VYbTD1iXp0zssGQ8/KgIRQA+Qzoo
Z7gwT581Xyg8n/V9gTqDLDPX2FlgRbq5RUgvI7CrpKl5zE07kq3BbMj56jbHLHcr
8ap8Iizal7Jaw1VzggrbmNhVMcG2aD02kQhjIWf8v1TfWpJyZN+Os6F79axFpX5g
Ox8pq36f9A2SeySL5ry4NqaPJ14GcNT7vgC1/Qkf/IBo/2abgRah+Do0vRny1SUW
uirH5d4qXr3qBpFUFmgf7oHNkib4eUFKpUMiNJ0833lAttf9eXzCZp0oFU69S4uC
rdyROYWwPjA0W4gLYRfJQwKyoLXSIcTGzwT4H/H5UEzEPlPnfcB7d49zTK68DLbX
/YBQOemCcwbztv2/g0fVpKTqMhW2Fzoq6eSEBC+hfEb0u2dH9CthhZM+St034eUQ
ULZbd3oLKyiWOt5PwtotDvDuRtYrYR1gpOSGy0qqaQB9z0GMxTJTlEUbZ/bn5Kbb
piL12IPGdpszfqd3/mj8F6gvJI5Gx1giM7D5WdCakUEQO3rbw3HQcLL8K5oZ3WOC
C+3B2zn+REQkRpaPv8Er+887QS/IHFuGpiAbnSP7b6f4VlK7Q0/SjMZhnsZ+6ZBz
7TYoS/qYEcyTlawpTGwWWIihau2EMGPYIY3+2aEKnAczwakvflF5LPQBezw3B8k4
jOT2RhqsxXEn/+l5beBsd43EdSG2HAMze5wHFnr0V9LsOU6nlnpIjqv5vTk5guNl
5LBbBDSCcCyTzlMMvBkvoFTlP3huVKlW2uEp/5fV6xv2ZuPgqWiUoaQK4paBnpBB
8F5O8NqlEKmj1ZERimYikc3beqzANW25MDStpYFhGWmFMrEt1AWn2aCq5NgPlyGf
yS26Jc9Yud+1ak8pmAxyjwHTC7wjTfUbaMof0ltpXVEEbfdzSQqwddbYj8S6QJbX
ju7nZMIszUYII7HS68PbuCUbV9vWd10wHUGoqOHrJCDI48s0YXDT9bK1FPgiaBlT
w2szWxHnx41x74OaTDZPuyzkBN24h/rDoVugAYIR+BHGgklXIvuNRbaybLnHvyaI
Uzhc0qHhk9WQmWD3sKAcfBZ+5Bwt6gJPB9cvZqQOLWqbLtvlpSCl8/fPdVy/Wa7p
nDpLa4EYRtt4l5Rd5huzxgIMpqmwABdhEzBBLMn9dHKshVe4bq7FSKQUbNDSg5eB
Pbv6e7w47+yA6zuuh0hYeiLhZsK8YiTjmWVhruVMlQK/oKjIP2YrVDq1STBJLaQS
PLhsEhD9Sv7VWJKM+RL1sBMttHx1Lf00+AWHU+MopNbPdESpzEmlAan884A8uy4q
Tg7oYh27/tmnAsxZPQkkMte78EgVWMfzhk4Gf793X9H4yc5ufgf5jB9fIUqmJbCA
rs3bRBClyBg/8a08GK5WFYaGzH/4hC5VC+PJL9fsFKL5ht4ry6/J/I9cTaQAyLWv
BdWnuIE2yZHdfFNBgNSyDX+8oHIPnns8yRXTrUQ+ZnISJYucovJVGdJ5I5f14SqA
jj/M+L8Aa1GJxd65KiJKJ11vYT1UCekCHL0yX+uxeJGyE/BcV1GWg4I7Ykpu3ryy
5ezDAKLfAlSEl1quaCmmR5c6WcId6SqNS2GzD/QzRzlvRkHaTiVP4+a9MEkAPq8z
9vSnOYJGu30pTnD0cSmtTZWK+vPgwtv8qfgkFEatCYS3j+fsLydntOaU/rNI50/v
XaeCIkuWQciLnwhGS4EROwJQOK/sJkYm0KHMpHwITgDshxsQRv1ToRUCAbbt9JRC
whujAdh4qQm9MXeTyOc0rggNRfHskSSvUJqfUIbEh2s//m4rZcYtv3cABWPNAyiA
qPUc+6JsBEaziuHAkJSBJ7868tY+Qto1GrL6yE8SmS5S+LnGPWGoWfkFl03/re7g
KTwtGRT37i6b+F8xABX86xU5kYaC1xtMgwNz35c6qETu5Go4sPjSkj1isDTtwlt+
CTNACxp3YLVe6M3p5CKll0vlqlbING53Lj31tmzwXRoMKJ4uZQ++uo5cxHVPt+AJ
wWQkGFumKJ3i4Qh3eDQU0/YOyV9a/xmMhhWNujootkzbsSWimkZP3w+z6eSG0r48
GAQYKTdLm/uKQSrFzl7gWfY4nT2ZlsZmJu1C36q5Ek9mUwIjMBISaVlvcdbCKWaP
/a8X4OcgBsMcr7qwtngrDfsr8pvw7z32bfiaquGeiLREBk3KN6fm5SY/JD5y0Wlq
O2ysFGVtfxsUbi2pQIq1RZYEk8olpLLo8VJZfx6Tazk/loJzhjrVWpwM7tXUYNxB
VldBnt+QUzVed/Z3IFL/1uu5C2Usq9du5gDGll2JG2cQDw7WHpP2y8iLJFi8a2CC
K5VywWrbC8er+TF+arTKyn8QP5dpXabQlRT1r4cpzx+Zb2JFQGwX8nZ6jDhEfAuA
t2F4vo+sitKAyNF2yCtr9LWRKqBkuiI+nuAKT+khidg6bgRiMBHQa+Dxj9warOLg
NTMb+5nbeqzHB2BWHBv6+YAiYMTLmATQsG692Tx4yyj/U1PvNQkjYH1y695xPH+u
IbJvZAeKx8Pa5meUuNSucyTgcbgKTP1biuWQqybvgJnwObW8ki22GgrGZS37VSgB
Lcf9RT/31aoFZ67iiEbVIj0lPf/3qUwAXGwV+/Vjn9fQnrgiDFAiU0nRhkeUetx6
e+OdYOVjMNBYcMckQRr7DdrypLsLp+kPp6n6NDOl6YzIQYKxb4K23vavCgr77eR7
WaM8L7pGGMqmUBR05IZvTVUQVo7MfHrDF4Fb2cPiMbQcoYwqDPWIlTSIukXhqgDB
mgTxwkm+PHgbFWvAHZesJSXWKVsCfMHI3IZwNt79gYgZveMLm3YBU36RdhKWbzZX
kffZQTYnX/PozlIMO1tWRxJ/KOzojO2d8dsYmn5xXsSVqEVTo2NKa72iQiFMAb3T
TwZ4dmrCobD1dbiT8rp2tM8j6YPkqmvLA7VZx6ak+QscVnXeL5qkQbFcpLImYOTU
pPxQmOk2nwMw4U4KK6ACUfcKbRMpt4DXI8FX9WpYKJCxp65Gw6YsNhOQmcAjFBHU
N1DJmEai614V20qocKMWF2LShzTZ3Vk4sOjBE276vRWaH/t3jE1lCfLUPNcXnb0k
ooZ70xt8zJ9I+mnrn5G/SLdW+bp5sCR+cJxXimJSn9Z2bAOpkMLt9Q1qL1sOUXMT
8PMBNlHGA1+HtuHhTcMK2cdqKIWjF8IYjM5b3Hn4nsj3rw6NqrnBCh3pqZlwEOoM
PvXkN5UYDKCpQsau71c9ZAhlHp0/QvC9P3SR21Kkcu/7zoYmFC1lbJoxii11Tjk+
qf4UINfoFs2dENYRgzPMx85D/RwtzZ0hLP6tGN3sKzsRU1m8FPF+qGLMK0EZ+ZwB
D9NdecOW3hu5Xr4k/KUttvI74QoAv7XOZF/00XHOBlGEq7xMEsd2lyWv/WuJYcuw
T9L5108h7Yvp4COhi8hLH/ddfjfKFwppfZ3/bUO5qKgu28wQjEELFCWxiwE0Yfcv
qDYzs4Qi4p787zrNRztgeRIwlFrplF026+bZB8tSrASLnMXz/oGEggGDpwgSJD3l
WEnf38D+chr3ej86LXXKjC2emkeis8yxoOOd1B2r93kHaE1/hVmyY/CJdD4JI8XI
mbA4ZcybZvKKOjvW3TyS0Dz/f97bSZtBAWyXijNDBDylXOr87alkL/nqCUpIo3vs
ML1mJiGH+18Ehmv92Jcl4tluYRFrOQ49bgqU/P/oZ7KrnVYsGhsru9ukvOvfi35e
QSOMfHjST65mFpWFs7TXmXOyvmzfNKN7ThvG8d86OZ1zpQ+dY9I9XmPgeYSGRoRE
LZVV8KQff8WsJCtAF62fFmBBC+y0/H48uiIyiFRTxwZosYfInluz4wywo3Fioihf
r+65ZPs9WFhmR3LK5Inb1OkoFbGRHhyC5tj7GHzqyjgCe8LagpVGWQ5df6P7ZnkW
9spYVQjxuBscTD85GWvHY4/fkQ+kq57cBcsveuSNZq411V1ty+TwsUZjwm1SHKbB
u9/q7ZJ1rQZQ+AtPp5vqHCgbLWxgEzV8RdxOngPfTH319Z0hkeoi4kUNNWWTVqZL
RjGYr4MTnKuF96mCJUMzzD+jSdmT2kiPnkNPTygAmt1YTn20wwdeQeEHq0pLbGJy
Vn/4Mt8F8gnACnO3soXBa0qsuvtAq2qVybA/+yth2I7y0R41ASKHQH8KAjlwSxwd
xNQhPYRr8gQVQzWixsR8WTNPzW9LsJoB+zmgc53GuwOb3G6WnuB6307xfUHe1eE+
s4i+t2Rfj3yccsVpibp43FJky1XWJMXK/bMj0sG3dHVrGe4F0np0jtu5xD1JprIk
ffkzBMGNXUhU7sWAGVdPZ8zJJtO8kJJhpz2fC2wQjW8dwxJJ0PQlXuZpqH64RQr3
gsboY6CEHRwOVhpMUq2HsN3su6sqmp1ItMmlzfIo+qWzDaWcoix6zbZvS490VjwO
Ixz5mN7zeHJuSDKYWJNKa8uMlWptljrgLDTfR5Iw+VPJMa1XI+jPISv8heKPEF/O
qqWurtgkL+EkKhpOhIXfsltquSX2gOoruoUKruUgrO9oCRnubsqW9WPsYn8IiRRd
IhoGKPA37//PivEHT1KDqZE4U+yjekw1+CnkI87viXeFXXcMjOg950a/DDIfPX30
ebXjtWeUiQld4OYLIhzPx5lh4tj+7RfSnAzvjGnRQ+BorSK0ojXV/L8RduybcRXE
Bhg1nMhN8GtGqzjus6UVhWawL0IZiekTYdI466JFxw6OixhNOqYb6Vbv2+rX9lmO
8ydHllDmy3g2GO/XMJYJrjLm+bpEESb2TnnWgPHzyjIRQ6IBzMtVHoN2CMS22Wd3
ZHa9iYo0D45nKXoENiDs6VeX5Mrye4BsIwdhnNetmgawNi67grZl1pntGju3ED6M
GMXuiX85DLU1Pz6I4iKqcoZ3+J77Z1Vl3kRcZ3WXRTTx9sJzzEQ8uumhdy7B5P7k
OkZ6p0axIp164fiXLFigjvqHBOx8MBwYIYkT5evEbC3gPSydKqvD0A3k1rhjwaY5
V426h34lKxqwSUe2Y63bcaMyUMHoKBDrcAraTqcwsypwFFy54XOslFMdQuE5j4Jt
rJoGij0eAfpfdN4sXg2+5bfbvP6d8WY4JXKAk8RqeQhq7vnZrJWdCl3uIvNsVCC7
c37Anhcp+YfnZwTMmXATSF1BvXDd9J0GAmv0G6Bzpntj0zAwxzZSCDZRpoSvx+gK
iWpB0koiMq3L/GUcxdRSRs9YktK6GWeWsw29cQQEVURMGXNrmdxZkzagn8VYVqmU
s79+OnjoXp2kzvNuc8lQKtL9HCcevrm/wuMG92Byq0Flap//Nz41fMBPocp0HGGc
9ed5usLpP8n6xm744b0cBKnI0/dBcezHOM7SYRYOF0L1TH0UPnTJStqzynsHTAjb
XDreZLGdFWG6oTwhrT8kg07E8IS/8lNOOPAkRjjKztEUFjoDR9sjxfWyj7WinfEf
Y3hRLXNxW1wDj9mG0WsMei9ehLYEOQjeJT79vdCCMqtWzT/H2ys77tCG03UPa6x0
EKf+qbOyicamPm/1zlrGKutdCVxgFo/0F/p2yKt54RXK6q6b/ry6kbqmazlfVPh7
HsRWh9ealjl4rfHxhpAaJ5zjQbJAE78n1Of3REWsFog0OlQ+VRRvN5gLrW5rHRby
Sqxt0kwJF6kzjEWZsm6Ee+8kpgSsRphYM/j5l70YQcJu3ysEEbRLQv8H8RsXvFH0
q1jgsQNwz73Iaiobi4lobALOMwCOf6kXndPPCHJkNjB+/QCrdSCOBpU/B7gLhzlA
o7SnDA3gVS1I6TjmuFZR6H4DwNvy1Tz9HuEiR1shLF5Ti0bl2NtEDlPBAtayG2ty
++Rz8Ck6/X/dTIGgSdkJV1CKmqXr4TWVBCkOEewyJz0PmbAYDxif2XvdS30xou6a
5bMSF7RqG/SGRlQW/bY1os+PPdC0PeR4KTEykiossPHCswn+ga7w33rMESERWuoL
XGhj5M+fXM+PKlyVrjW+gV9f4FzgEwIoRa+IIpReJE/1+948dwen9ZMPv0XRngVF
wAfdW2Jy9FMqB/lJqlFV5GQ4hBk5QLFryj8a4t2VG1FfG+54V/PZUoU59FxYoFFp
oihNQgXrMptnTEgPhbY6P6j6lU9xlTVoFQJzcbmVOGGQM3cKBwf74hTpics4yR0b
OxVZxGPR0bcO1GxogRzhZlB0Wrb2lDxyjv01ipD2l+582ypYfRjdk0al1MZ0sfFn
2g6pWc4/GQ+Ea+lriyUBTzMK3x/x31ar5c7q9CmNhybmH4oNhsP+5h8VEnsIgFc/
6OcQ7q2Y1vAmrvM01Cx9mA6eK+bk9ceIVf5E3a/UQxu+UfXX+3Bpf248CYeTxECf
QqHU4rCleoieNrE+LNmYmryWpehcrvurBGF176xFTERCi7QlvOiJXjDkwkU0u1Ef
w/9ElH/mJ4TCc+9eUKHlk9l09iW64xOJV5ri9OMFOiOywU7AUmsMKA6TPOAhUPzU
p+T3Fdkjbm9p3/2/EmYcHPE8WsabU18UTQtW57zwZ15iM0BmHH+MbZaODvIaMA1K
Blk3A2sj6gIhSFjSCiHZmqRQZBYtYkpjf/cG7yiZpiKlI8+kdE/EQ0EbjIvp9IBE
/3ECII2z3dyw7c4VJShUZLzh55rR5e0m3jMbYwWgFfCJP+WWH3YTFqufW7rb00r/
TRJQM58V4hT2CWUzcKK9+Quw4iUptrgMg8Rboq5KiRaKMPR9oE77NEVAu9p3eA5c
uQW0Ez7Rj67Qv5ALeJEfdv/lx7tgQjOcJTZro1JeS+NsTEJCRI8eFCF9JCUJ9A5W
2HYIVEehQpgE0KiKa7DffLWKC5/k6nmpizTNq6OKbLI6J8sh938EezHKPv+YReqK
YW+4BBIgTo/vHIM6jge7I0dlA9YOG899gWKaT2fAtvO9lO/SfLNVm5IZ0/enIBYN
1GEuBgzyEhsgzzErK0X1m65+fDA/nNIpM2cBRC1DVe0Hk7iMpCXGGKL+GlYNks61
fLbnuxHaUZcEus3EWZCwMw5rNodu0jTUsRtY7AMJoMYrEQpbQXb2fxqwm813cAz7
wrbei9UrGjIXSmXjpyBZyRXOcL4ZBvsy2V8Tki6trzWNo0h9XVYpmrEAlHmuOWtp
sw0lrnZBL7iG/dGnPUJ4y1RbeYH560VL3z/60rInOy0bE3lrxSM7uLin23EXa8xz
W/tMzc/4ltsy/J8OXR2/ERe4L68ht2e+20QwiCAOss7Jt0JBJ2sEROr3cuY5ox7R
dvjvm1YDwr0Dlnj6DHWt5FskMtVlIhL/dxE3IwXLs4pzZbEz7h/YOrGMjTROMx/h
hNblREqRRKPSW5Vq0SNisb4Q3m83FG05I/GqVeIQ2b+g4HWNlaDP9B+6iwxXsqh9
7jgyiWyQ3p5qXrOXYImH2c3NkdYOTmgd0nIsgNZVoL9C6K7GbpjWOIa2vqkh8EYz
NsXjhi8D5iPpIa7nxm+8888cvEqvwhTd/ez9nqbVkHmuzLTA7R9aBuMAm/eRwU+n
ewr+quU3PrfQuWeLhaHLUgDkkVgpOsJ1rlejZT/r8UiEZAa37wrFdy9iaXLJDORd
/UPYTJikHR473f4wkdesXundepc0t/rKwnTt5ZVsJ3TlZpBz9R82Rtnco1tpoHWu
5WkQxu6Y1vCkPsj9lOlj0QKuvq8g/CxF37JGAnlT8BCFXnlZQ6hGTzjVn4f3aYXh
/36iv59OnevyqHn4DrlWuIKQd/P6FTNhz0Kb7npRFJKjWPwUwFt7VipTJoLMuA1e
WnIdamdibjhAcaIkP1SnMQWoP4h3/jXoSgmjD1dgBTspF6QoCh+QIy38sRPa+1B5
t5Yd37cfNtNbEBStxpGH2d9k/tKYQnDbRmpKyvIROLklHtCKUlsAYRUy/kfKz+5K
5IZvqQqYEEWW6jGRmRkLFxPaShUdi8Jk//8YcTYjqKvzjSjs9A9IOi/mVS3LgiwU
5ZMg5KPQr0G6gppzgc597CXlwXJ2jmqbfEmfjYgfImapPwdNHLZ23kjzbOqBhinO
ewvMDHvriMar+rQ/mdu3AdSeieBnrnWgseOmV5KdLEZoYkjj+BZA51DDN1+XNnzt
LE/HQejEXrUJ/xkUChB8QQCrUVxdAB/f5cf5DGqB4cAxKmbIlx+Im+1gd/sxp+U6
S4yYj1l3Yl16Daomk+y4LMdl1hhFLjHVXJYoan3Y7nE6nyCbK4OZzT0lIXRghzzR
fx1pumZ+T2sYjQWbLdkojak20DpS7zFHMWIvFoCPaAVqacMUI/6+ckpnBoFN6qLT
bQCLJ2rCxRdTh/w4HbLWL3DaL6UFImWq1+uYT9xh1liJXGijuj4jg1zt7bJiz+Dp
RSw8LeWVQw0huvBGGghr3evVzGJ9ihL7XWv1qrPJ8hGkHqbU3UbmSlKUwenv3mn0
GjU+qOQ6AlVdpx4zjBN7n8k52URy/+ef+F4u5uE9pYCUQ3LU7m14uBgPQUR224VA
orHjUc8N+yI2oEaZWXlcmdzFeSm6VDJK4WfxhEb4f2CiE5wbWSlHX9NjZXrjNh0S
ejbr3JLK1BEQovi80O85p+cztnF38pWen3L8YW3VNIEzU1Nj24eZChPNDDBmPZVh
pDjsOh3I2q6J9WXbIF/0pQI6lHkGfTqfvk75SAo0tPa1cpXJoY6bca4i9r95mxVE
cq6Npik727BoM4mFBsgIQ5uN/nb40KIj4zrEtNj4YxDr77Xvj8ndzd7xHc73EgoD
MQDK7idigb9n8VzFu6yKSaYjW9oKIcN1CWs3bz1e4mXM1ULXToRXYGHHkElnVpfX
9d/g0QebgcknqsqY9itjnpiIDlesHIz+wIx+b2iiy2UKkZL19WQ/NE7NS/A3gm//
P3MMk5Kpgcx4nf6kTdr1npbHZ7eGQfRGcsjYmEVctDMHssjgOZTGNqN+8qz/5tIf
xShQX2BeMdqmc8yFIfZSETJxORzRXGKSYwM1IqxdAqAe/kYHFFnzCOANzo8IhPe9
UO/ERCMHbqOVflo8GNREGtCO/SVgl/D9lvEldxgsDmO+b7uFHoOS4OVeTr4kc/H6
w1MSAW1ZyOM2IW6sbwpExVaqcQkmMFDJRs4zBFLnJzDFya7Z+jFkl3qQbOYImI4T
NzYOkfBSvDeHmuS5XShNkhE8DENVSBTwqgFHHz8/3hM5JM9j+w7jpzpNSYWEvmA/
9IuEHwx3KV9tVcKlzIQnut6WkFbK3EiF5Usg2lrioicOjQM3vDEkXiQI3wjWbNHH
VHmnw3l29GfmFerwpk83kXxU/EjY+czoQkm8/iD4B3yY8shI7W6rAnMIGqOa3fyZ
bVQvYGLnLwxOvicSVy+R5ey99rniWIUW5ihNM6gdck4Jqeane1JTj/tQfion9ium
PrxQWL4TJ/jmAySnyejxDbIKjN1eYVWQQ7KWMhm/DdKJt99OpfZtS2daGlRVtn5C
pW6R8RKN4DNq935PO1Ciq0CbwrD9MA7XWjpEnCfhIJe8wBHijpXzB1xAqcAtqrzW
n2qozsfiC1CIigK2i27kHkKEC0THF1xhATiKC+uHx0V3e7jiCGb73YeQmT5Jmzw4
BeUKepG4tgnbtBhviwVjeAOOUZT/vn2wLSFZOtsYFGBukwJqnzlRuSk8UbM7Ui1s
3YU1ymJbi5j/2okExh6qGgz4FCUOwecHBUnJZaUSd2waE0ll4AXVCKLQY9xTn4Rm
x8K/7gJONDiwnHqcWkXdJ/3JsCQI8/5LfcDqOpHik0tjEY8HLdV+rCXKlUIkP15v
Kr2xfrS+6AglQkklwvwp9GNsT0+KHUrGph3WxRn7+9mmhjtH1TkGae6u3NT09rLZ
TSobEW6mGXWb6R6YZICrUmbqPbLTG1HdSTST5NG3BCZQ6KUn8Wp6Z242aoOof3M4
rKdLTjDK3M9YFGLINaKZ5aHTG7ZXKO8Q0gjhzkIdXE50TrTuKqTqv45r81HpCr22
zLNVQ55RmeDHvaWu1P3qIGjtdmFMAQX7geoDLnfN0stH1Kn4n9r8zgWn/K5IiYyO
x9wtm86sOPCehLcu63mhTOWVZyxGpJ0S7AE9SvCTxCVoO231hDc2gkZ6kGqhZOMc
FDQFW0apQcGHhOT690d+G61sbDckIWyYXOX8b+N6Po58BCre5Vu1IYy5HZ4rpX24
MOsusyy3vQKMab6xua3NNB7lDaO5sim2HobcPUMptxZoRLSwlcokY91cecVaA5Wz
r+nW1GiSuHEdEwJBz1EZ10eZnBfD8+/h5gJSAI3J7Z6fxxdOLImmCpiXsOq4EtbH
ui2mGAeBIjzanxMXcYlpOROBRIeeXKFTV6ciEdZlFaHhv2uSsWGCNPEqR49s5jXt
kqY1VdzFmobVv3JbmzrdPQICioQEsqFQjez80oWhSBnLLWQV/SOf1ws5JmTSYFbM
3MWeMYfBqx9S/b0USSSeqWATI0QBewxdLj26DfezaPVv7ef9bz9PxBB4DQkPsAJu
qOleVVgisByQf9UesXFg6+8OyYFr6wM9ThY9Df2/WZENWnvkzYJwAghcM7CB8fdj
GLcqoyPFAJc3KiIFEjeHbrZI3Uky0d3Z80iRAf5gL6JHLH3c5eA/I7sEDMVoeUll
F9JpO0lpo3nMzVYEcRg6k45B6eCjGzl5/0BTRP8fTHSESe/mf1S/84Z5qRrTLoE1
lwqV2XNfsiAvScvAXA7zaZO2virSYHg2AWHNVDKKhtLJ9RtKtluuUyfKzvifS2X5
tzywf/kADUmBCwqIzYObFHb0w0lBy2jyBndAhbYF70TX1yyjIE4c8pk/8cKSPoOT
UPKvfqB2eCQw65foS+6gYpd5jKJeTi02GbRtfFsaAAmo8eh1cAAC1Mn+Wd13ODCO
sHRkp+3C0jWw3G87/4EJNKo5TuP9Xkz8Xb57IBolau36ZW5mMyOZXXUNiHgYWFx+
eqAIpeyTu9ZYEbAsq56NZloEsGwajLEP+AWEBOCEAYhY3+EARkzetuXj8eMDDUzO
hF0SDOpR1diqT7FCiSM33JWtwLS/yhJHKjkfjOiJxjkTPWa//vukDDulJYP/E3dg
KLCBWLnTnfWpvvbmOlCqGhwNWDPK3a1R+81EHdtpro45tNlt4CTDWf060nJDeY8t
vD0naa9gUteakL6Nbvb7evsJz6E5imCjROEY/+CCTi+7w6rcKfJbr/tMv4h/jR2s
SdQSSHWmDaaLT2ingp45cqFM4J6Zm1SRLUUSAfEqR+wamuKLHLupSahWmxO/tYCE
WNc0IKvmlRicuMhtL0P8LLVKJgMfOE6F3fkblmf6F5gV7Z5eP27uVhuLxJ4vss3u
tb4ajJ+a5vyz5k5DcwaGkPfpQBhMH1CSkf4k3ku+x/f3ZWnVlYuV2W6iooy3hNXb
m0BQ8Gtr8YenjcM5jFAxzFU2o0LN96F8JvMDI8kGZMXBzM/XV2PzIJ97hYr+ZIaA
pAVuoy37F2wTQgskBxTKkjbkP3xvopJAs74ipz2LMIFwfDQBuMVlDqnVYB9b8vTi
axeQXCAV+p7MKZrBzDvtRxWzotLzB+1rT4tyIk9loyldOv5FFTtrZe2Z8La6YsWO
1bH2LlRkRl1nWwwcy4Pc8ikIPZPgHc0K73CmsE4rHkOCMltmzm+s0jif1cAVgx1k
kR3dNtiXpeq9Jt6TzQTroLZloduJxIpXwwuTLSToJ+nALfYcR5mDLNctupY3JnZg
SbnrgnZt6UB3ExOgNmx+l1vYEbuEjWnKzuqfTB50v5ZRVccMuBF+KNuUqj2pbYM7
0caSUAWDrRbFsFj37Sx84H1CV9gXCT160f2aBtp+mngGiGOaOUlq2wJPug2GV76y
iBFjiRh1Si6m89v9cdpmLarnIU5Nsx1OUs1SluvuLu1RdgwfcOaQ/JbMrtRqObx3
bLNn72cFabphzMDKjEqUCc5dVIwqKMTU36xQfxp72uuFhcjAFhEZZNtxZeC4dYxY
VLHUjrXntOrTTXYMwcHtoWDyKo4+dCbraOpEY3fEC4e7oYroScOT1IpBt71K0fF3
t559ZoRDHpLu42wTguggp7N9WI/NcL2FF5Qrq67cXwHZI+coDtJ+CnDLM2D7c1OU
KjjyiVgBwC0O1Vs7ir2RYQOjb37PF5hAjIjmouC2V9y6xKFOy/Lyg5ZhXblqxj23
buicR5YEjAZ8J4XX2oe0n1Tr8hAobWRnadic/Gvr4kj1QRQ0E2qMJhw2MzI8H4wG
Hm7v1RkwtLYrLujWPjKswZlzOdqM7rMlfSyOLLZQMwfHDPkqU/ZkrK8p/gTwcSKe
1h2IAIYkdEi9/m4qP9If6W7CjUF179PZLH48ruZU9KLTneAsZ2meMELFELUlBK/q
fuvIpzjkVJwowWK2wbbKCt2RgeF1O0Kv11fOMk39E3PDxmMRbIVY/tQDu6UJUwWs
2G9kZ+nrUBIfM7dpMgWBAIY26ui1OMBDPMInw3kJNfAqrGaRXvV3l82kRg/NI9N7
+uA6T5vZQanN7KKRPv2OhvBdoIQcnBxuCqcZCJSeYjHx07WyhZ2Idu2BJa0i2yNZ
6VT6u5c146FTSK+XYFnSVdGmqcyfnKuXj2lYyyOSD8C4v/I0CyJicIThX8Ra0GZO
G1WourZmoi9TuHfj4eEn3k1RZ7aBSAIEt8X3LiTYg/D8xyXc5I21XLbiHr12GTgs
B+F4qOOotqPCOkCX1R/pHoGa7Y17pNnjmkoly1mNqNP68owljPR9mnWUBcD2WABG
KPE0EM1xiF7GiRJh1ysT7NOpmk9eO66jdJANKR1AKZBwWlxD8PZH3b84xBmio+tZ
A68UVJQ1jeG/gx1cC9FV3M92oFFa/oRRWee975uh9ac+uOjGTiBtvav7JUvQz1Tm
5plGjZ6a7/VDDLhHDtFR1wtZ2NRRmzERQA2lqQkMI9/370Fyua05w/rxnwKphDva
hG6x5BH7BRdHtE2UwDTMXPamyMAJPok9Isb0ZWMP/+wLkX5vlpPe9JA2yoRS+2Jf
BJ+XywNfLlBdbnFfLP7szK6jMEWeOrFhX8NCNXilLCyI3sXNh1kfxjShtfbS7JEV
tYodOrPvvO4wEyxyXTPF6H/qBHQyul2slBtA3jzvj/jza5brTXQ5OwxxPqmTEx4+
DAw40Ti+mIgsq7KjugQUvVOSb+SymXbBUHrMtwbJdntak6G9hfTSm81Ihxnps/y+
C239L4WkiWzHfXiTMTD/k71VWSS5ntrKqY8QerCkH5vZnl/KobU+/vkFnbMmxvOO
dk0bwx1rYy57pr3qDdlVdPRJdZ2MMCAXa6n+6YciiBraMDyJ1zS9OmFrfLneQbK2
9jo/PRyU3cum6bjLNNkZOSQw8zj3cqiyIxNFtEPGJsBtR9P3eTlzSBiup3NHGCCU
hty2rtkzFQ1PdcFQv6yjpU+E3Gj1iG4q1R0rlYvd6pA5NWiVwQj2fXqSsR8v9jGM
Tk0KiyAf2ey0RNKLTDxq3Oy32/YhgAqUIm+203hP8+NwJj7T0bD6AIms0IfDljo4
JaPh5zzu0YXbmswz9tUeKGZhf/ePgrhUxXdzFcA4bG/jJPAaFHoD1eQHGjzq4ZLI
6ymCF8+sfURsnQ1hqEedYiKjosmmn0mNRdj0aQfmYrQumZ5iROuLK3cQ9xM8/HDI
fFe0+2+1J/EdSXqCPJY+/4fkTysHuooFW4AyYLu1VWJ0IAcWA1IWiiTpWZ9leEpJ
EY9PU0azZMqs4LEmr7uYxXAXR9g5NxWqW5xOExO3HViujeHAMVyNrHtwJvrqh5cZ
HAdKlbMM3Z66IkGvvjFGLyWMZCJ3ckGq20kOp8eEz2MItlwLMvaMlQ6gIA3xVAM+
bfsP9qiBGPDQDCmQ1srC6vnpXUWha+hVyM5dfyC1sVpOWeAIMTGnSk/hgVkPW1C9
sDx1SqYl1c6e0jy7EE2K6DuMjVvbC4hbnssAEJLnvIndgndWW+KP92OpQP+ZagsT
BnRfiKlB6S+rQ4qLthT2aDWsnpdiU0BUODIgPL+TjsY5FgTG8nHHpQcLwgeH0KGj
zu5cODTTday0AFqWGj6mPM6TMI0rS2uaNpDwQlMq0kaSzL7VOP+ocWjq6p/nPX3R
5fwx5p3MQ66DzlfeYU9diNhJXrWtg3mcn+wA9m/wcCmCtEOo46YIvglJ/6OBHTXX
W6kXyRrwzGnJdFQaSTQK1PK1m2Wni+CCoYNEj8JjyX9G7cgd8ZIrQJtaZB11Ktz1
3dDf3eyMA298eiXbDdog1ez16d0gvA+p317a+1EnWjhWrJIhXU6Q02Pw9H3fKFAr
DunuLHVZpCxIssSn5f4q3bUm1q+ETtl58qVv28udNmujAH+gLZSYdxevR1RK94M/
C93NiLjlWQoYbW5uea8lS+lngi5/LPzQI6nJPpH4Eq1OkIrlfO2qMiNpJ9cme9Lt
McL2J0BptN7WEc/1LI5OOca34LuNhBNRQY9CVXJDcPz0W4/wBfFjcLpuOcsO72FP
lngoR7ayUg4DY12yr54Tg16xnL1IlDkzZt+9b2M4oKGAkqotTTFYx1pWd5UU+p80
q68xcUAMD/2U0jr4iGi3FBKLYgSUmPnZSJ8yj2+0tG8ZCB1XdBaGNPM48yaOA4O8
EXCXAS8mrusIqFMcCS0yQzSXcBUSHTpTuFJNpEehXR4vezfpwKmYOKT/C/Qbwklh
yJaLi+wPT2MWlh63KDd/JXVZchXcb9cwZmZU0BsjrWHTiSdNhET4D1T/sKg1VYA8
gVeLV2ZT9gQ++K2yuNWs5bAz65fDBgEHyJv/0IxxetfG2qkyGamsrtosIhpIPSct
1lGDFDNciH5MWCWssDgWcylTbURLzCQG9vmmFtO1IJcQZJq5dynbTnhEe7dYpCzW
gTeFMaDKD9MUSp1wDOQUpFVQJ+LZDmBbRNCld4a0kDIlmdxgXXLVi8XPBcBJCckM
UkjC0bm1KbJsmw3RRj2/9/Xzh/BPPQJ71AFOTDZW8EmNTMRSjVzixad8eA0785tS
NzwVvmv2qktUIzRh1ml1qNjJmbn7N18dL0MJiQDtTDdeIAvzyaUEQdG44HnH9s+0
W4kMm9h2djO2zhxXfIkDZmkV+1jgaiS9oZtILhYXsZMollegPtbNMfhdF8by2Kjs
pICliDgk+XmQRnCrphbgNK1nTtMqf9wVeR/g6i/EVosOuzp9n3X1E7e86D1HbAkl
pHKSig9seSSiE2jBeC1MYcZE/pGu68/DMNypGyJuaYjdRi2dAPHDt8OXMsxWJvP/
WD0ZXisloXLgUywS5ZR7IVBIGGkEE4rDlXUasbeUNGd+hnht+qWV+H9xS03AmG5h
3d/VXxPnffwDtyDCH4ttfo5p9yZ4THZWNn4DneODWCj4K2CK4zsiClFEtaHkLv9A
l8ZuV8NqCT7iaVo7HfeFf4hRKPySmQxWHYJVCEKmELNG2E+yaYyX6uwcvZRNRPV4
XjcfefYC4B2HW/YZcMbKBF2LcRouXsK3iqf1PvhjcZaBXseADSK0hE/hfgjWtzDx
UVGjX7sx+2qQyIFjw6GSgalikJs4XvbG7lt7nI2mLsGy+801DnrCKMO3R+qkpnD3
T525sFfVlx8r90zWcfXRZNparKfZFWQSnYEB3nro1NtZpbLW707IyfrtgELHYY91
qtPH9wtf2+inm8MMOIy3I5TWzxE4nGZRW/2vT06yoLIv9Gf5KWOSppYK6YdS3SG6
GkASqArwPHgyUBH7ovqhUzdBln1afAmd8mzngJnBdhr1YMuLl+T4vYeWo2D37TIa
eiOFTQ/9VtX0/ipTD4r0dtyKi8SkNHV5h3stX/G8TDqtEvkrV9WS11IghOgsLSXD
KPI7q62gXRS6DnPHuKPeDL+FiKLD8T3C/gxhaoRtF4CM0oRdqV1/SGmfvd/hHVXn
7CicYQRjyXQF0Q7Vy51GpCudl7CWSjOo/ipK8e3ZnxRqn54Dim+zNJ2VdZKtVmAR
kspr4D8dtrjS0y3Qy0uLshhfRPARFJABaRd2Jnuk4nPyqtkN+FnlL1lFbIk8It8J
eSoJg6kZT1Fdq6+AKcPk3CvWaVwtW4cCull9QUFeK40IFah1Tdw18woee//mlmLi
NNQsm7iZyHSSGITEYgRd0vfatWpF6VHdZ5i9/fytvF59StpDaHxiby/RW8KpN8Xn
Ola+Z+pwNQlQUBiwTpo6KfP6yOu8sy0D0bdGAi9BvMfYg4PRBqQlG4nBCOgIiUgP
dfvtU7q4wvujqg6AEGtOB3pp5ThNqHd8G3+xbQF+OI0LjC5voAu4SHSvhuS5+lds
vPlQappDyQleog0axAh61l82mDd+Fce2DAuTU2iUD2EOvZo0HV3wuN9bzGO02P/d
oK3T/tHGSv1t50xjmBDRZfPYD2P3JxeufTPIbX0XyaIXoU1qjfnZMhjWhQU6gdEP
gr++UFFrKSfLdtGQojidtPv0UCxy7W2sYbLb4vgV9ud0U6dORb87mE9URQvpx3Gy
TCEG9Hm2KfEuNRqV+86xuJy8BP6LNT+HTis05dHtqmdSgw9b3KIhNxys2pIEeOJ8
zizAzVCQwRdn/ejx2DukPbInh1ChH+x5PJOOB3kwfxwA0j8RgBMT99Tty0Q4SBYu
6Cgncp/6FmQ3YiJoSTnyiQ4RD4viKdSCKteCvKlriFioh2M2LBS+rQVuEVuke7ga
zpkLDKYJ9/rfWalj90o9GzasMwC89FJWLbCBUfWR3qCoKB4JLt9Ee+R+8F/24Wz1
8NUpAGmebWnEa7UcgsC9f/L/0/7X4YuH4lZY4u4/uDYCPJdra60+vvr+IhZ1kQ2N
D9DiYhU/RLZ6CQWMIWl5rgUX1Kj0eWOHJ1J4Hd2xWBphuv/tCmR3rlR8y8VLiKQ1
8EpcOvgWuA/vqjM//bq3ZGoCH6vdWwM/VUbH1Hl6MYLk/1V3vNLOaKNjhmaWwvPr
dMnROtXnjEowOAV9LfYmuXf40pFclj11iNtIXwSA/y5L24GaUGn37gbxJ7A7VLmf
pzNfsRBeIMcKGLRCSWxSRkPFvexIZDL/6oclid80IBiFU0iquixU9TKWqHAHO+HD
W3vlxx5nrWv2NndinOIHxoMaVstX2qvSIlYP2BdKv3jAqrTYOYZYU7WQ00+5U25g
iprgJlyqhlo68AH6g7yH5yGXPKEO4fPUS8x1jWg+kSqTzE/aFgnD0/o4xlqj63RM
x/a/5UT7/RLvJsQaZpPchU8V9UZ+UuHcYPE5DaqkaJZjaaG9OCuHKfFaV1ius8Rb
iS3GE0aU0SyfDvl7s8892ADcZYbSv3HHI+CKmt5mRNJ0GrWEzmNxdxBbvJjI4jRi
5HkWfOwPoDz25LC7u/j0XIhFSX7UYMEoXhh2hBCG5dztKjAPDKuScTzuJnUsdNH3
jlRBUVUuRTMuLeD56s+i7LAEpdlFhzMrhXK/mWqHNmw+A3x/1OdoRt8uJR5MbV0b
9WYuxj4Gi0mNhw6/TSMkVl1k1oT8YZp5ReTz8J6WipN34qozY+a0v2YcnYq9jfho
eOPoWrqdqGwQuQWfLyl2jsa/YuAwbjg/GWye9tsRc43ZcB60EYzyJW9JSG25fq66
IsDWiB3575MXs7YIwgkBj2aVCXEXLO/pGtYWpUzCCudMUAIxBvENDnUyB1pV2yr/
e7N+ybJJNW2qA521dqtRNpKffwoRt11cnZJnKoE8UVWXk80O2D4A3ZWUTTiHdiFm
Zpjhczj4nKKJ3Gfs3CbBK9I1oIY/04jbifPPMmrG4HBm0CqsnLpetBqIjwP5jyLG
LxgV+ZFBvrXJ1D3LhYL2UZo4tDT0xClzgJsO768Wla9NCCGmnaZ/YUPHwE8OIH6/
SOBvrtwn1oaAUgLG5Gd71G3vIM2wwx2MkS5rRp0AQgplpZMwfbuvGXct7GXzUQWe
uTjvwe/P6R5f+QLJY8CPYK9wqlBwD3MiGBm9K5RORJ+Posc4JQnHM/xtqEi8ReTP
fNKVVlcjK9HR6/SMnoz1YrOUaroT7jHdCvcxTQzyC3xBiEfb8zKWD9BMlfAetRY6
K53SsE1Bt3iQ/GmxLdXqRD6brRYz3TrVRbMq1ohMhdpHB61WIsbFK/yHl5tQMC7/
BcWAVYM72dv547RwRf2dqN0CNltwTlXRsJzLfQO65lQBQ6jzwUTTqJpsYvbzR+0f
DqGSMzNDehtgD5t0QeZMSSlhcTia1e1DHYQf8cWDxszoXXUOJHzMnhADNn72ln7A
v3cZwu/7wahPFBVuh6+wnlwfQMdhonTxTvkr7+UUfwQXZkCdV+tzNJ+vduzBVXj2
y8tsxfabV/ZuAg2RDRlRb1B7Q+gPSLklbGRv5TkdDx3TRyjftdAV/iOk8rDHkivL
MeZ0X2X3Q5HTENYu/x0u+kDHmMw3eFroTpfFuPOPXhJAPYc/nLArESB8KhdEN8+l
S7g/3H2sb9VKP905iJEp04g2Tdk51CdKP2Dt8EV/M77NS7Ckpza/y16qvtJPxcQK
ej7iHAnuDENGNlLCPNdKRdFFVSQsy4WkCvnWm9n/qVpTHYQCvVCLBy71Pbu3xQ3C
cmaAYKt9ZVeDoxw2enAMp1pcQ04vAVRDf6cRLSzcowKt2p7QxIO4rk671FXEE+be
S623G1NrYP0V3IXl+xx0bQGzOWTUJem3swBxccD9VS4CLIElOCAmzPHep9+ZyxNw
mqqVDwFd/gHKESpJRRkrK2czIvCMgphYW3JHK7nYzfFGD31ZQ5sJHI8Dtb3JFfHl
JQfknDULdMQzusxjGSPWz9aMXfFzyZ8xDQhcAXr/eDIG4pjk9hnSDBwiKC7mqBnI
WGtcbIl7J1IGM/8cJEQJegzDtNoylcDUOFC/5pAHO4kHIRDwMCVmS3XtPwTIId/n
EQZZBFPha1AC6Wb0qXqyac0qNqTNakokgbL3OvwP2Nb61od6KY4WYor4V/hX59Or
YKCtW4qBO/J+xRF5tOETzWOFUG7gvWXD8gYwQgehINjUGQSJ/Rp2eXG6kY1lzzas
5V/df+yj7wI/kDbzbXJ7NMoc5hgNniqpHRtPef+B2KVKziy6xapNhCJWTyih+gNW
d32sV9uA94egy+iU/eY0pI4WCyCuYEHcv6fPo6r7iKxObmAlDVA0y2qkOj+FgbjG
feEF0/IEymXfgXkHDRp9jDLTNweOqfSH4nD03UqgLP7Ja/EmebeNDEPCjZCUyOvu
XmTwgp8rrgZk4DBI4sbWQvcJagKPZfsGu+CtSpCsgIhzxCRvKKHnX7sR5Z+dNgXv
vFd//1t8TKk9aTcfGQOSLHMMDm1qO57xGg6IMoHfqrthOrJ8hv4zxZsPaX9AgcPO
RkZ/BtlvikCRFMvD0EibDF7QnfOXT1PSZcikP5V4OSbMoIFLrgOKYmEQx76ttDzW
fXd821L/HymuU8LcfqEnhyVg2WogeSOeqPkjptqcDBI3H+Olu/CSa1v8B7Bx+JA0
VcSfQh9YSniA0vVetwUqMwNRChm6RO2VmjhGvWUceR83Gx4rzELRXouWJ0B5thCl
2TJEVNv98k6dR41THocdf0PxZn42ZvQ/1On8tBvxTUzFtjLPBbgOjAQ5mHPldPX1
Csy6ZK3ZrQmvoNudYk4WLOdc1d7nrg44SRby45XZYVT2OB8wMRI1qlEa4wgG3yY8
bC4CgLwe/Cb051Y/R0pTdL4jZhcB5uN0p7AI7o6JYL3drqgpeMoiTLfsKtE9m0fH
/weDNbMSro8ei4yDroQ8dkXMPOILyfGm4RzWlFFece1jrMpf8+L/K3Thc78Sz91B
Cv/woXt4uQK6o+FpQT+ntzhkNMoOy7Kza0AXOqTvyMegKqo2DKZglOTOwQMhHbUe
wVWGC8XqyqpWo9h19ls/AMbW+JBVa5lLr/QFar8z/fVFWgFkQf1tPZ4l0u5wYZ1N
G3dscdVMjReDWamGBVwQKMyY8Xq/Onpg+GKI6kbZIs58HFBEzyiGO/9+WsyZH+J+
AEnA1rY4qHvK7zbFPACbELKhbHKyUlzfMLbqXm/ZVpStNXMFJDBlrtPf1bOZf2wN
eoVdZu5unAc9P7SG3aVEBJsNhGYo8RcySmRoQKZpSGHzh2oxGBa6Dm27X45jNqrm
OWDPUO0rBuwP/VcYExBafKXgSHJhrzv9BDOkP+d1Tq/LzNHxQMEz+d6w30PN5q6z
7l92yJSWGIXNcF6/T7dvJGtIgfx8ZbIq5kOAj3CsSwQlgjxQDmQpOHU5VDaYk6oq
q5hXyamc5wIi8KCpOI6HGcta+tLaHONwUFoww6SyceubhuNydvmwUpZxLllCE97Q
ILX7ElG0SVUbodTf8ek9Cz2x6Mi92znHbNNc6B8CjtQIu9BtSBCd24P1WtL3vJAp
QD1viwvHwDJ6HLTbmYlD1gkxqP8l3hmUhOKIyGBnvayMHReSqmfrXuqImUZOsKGF
pytkTT/y/HQ1jL930XsI8gW5kR16En8wx2uTFo5lyhOhBiovuGDRgxRCD69N7y1t
IxzCMF4Ucp3Q+3k5+Oc39OxtruvRoHmZm3JeWizIg7Cokur3j9XbXtVj3p/YvXrP
zOiMDFmgpNe9Q29eVRVZ1kTJn/XC/yjWfoXJGtdegvl4baClVyQEPv+IKRFGdk4v
ylhFLGbZiPoC0W74zwdtiZ/D7EqYrw4tpUEIsOs/9GB1BDanKTBD2/IeODkiSK3D
o81lebE9q8ElAXEEdid4TF/ivUzsnwca+KrV6p0TvKv5eyhY8e1AQujha3ooThLk
Ey7Ti9wvAFSkFL7jCJCO46mIUDtEOSjbmUCUlnwpeHgs6Wo1hR+1GKyxf+QpSEde
AXPwpRYEWKTod9h2REuQfJoJBXW1kA9lRL5tHSefwHqINClJGeSbXOTVgtOMoyGV
BKSinfC4adZy0b/a1+hoA2vXKb7hhSzmQXmNbCzSRmuujKvXMHz20iLbLvaMVTAS
tkHnvQghD0AnqmRRChmh/rFhFV5Ico7N/PfnFuXarLb5rCTT26p8BMrBqL7hO+k1
bXLcuWuQHBtnk70zuThkZbLAaUHx693gbaeaJ9yADDimwfyzDBzBslS6FNj7dNcZ
3MLxnHwh5MMJ5SS16A2VOEQPxwOIMaOXBpqKOIsggRZCMMg2toVDBcyiBw8ySjqJ
zGJD4sYrjuC+29x473lC0mKc4Sgcaca8STF3luPdAPPkAIaVV3H2k7P2ttAtOjth
C1C+L3YUsaX8CWgszX8Q50aTgf8oxo4NfUr8E9QCFiAgYg5xVviW4klOu8zmHr8a
XCXMtoJ64rjaMRWMhBxxpombJj/t7/HAYlASk7pvkYTp6XGnapAxqqnpZxpDk0+w
zoDFogxg3dnexfM88l1tT+936K+XFTCWEIH8qcykW7jJJo26wo96PAARItZlS3ym
RwFAcGLXKFuGiAFeg5RzR50fHv9ObMJ7vHjXHDvkmESPdhkaUFibNk4CH4JMvfAy
BTuk4XPRE5+Ze6dDsb6N5FkmBcccsaiqq6O60QF5Lu+g8XNdyEtzMMcMta9ouyUr
/Nwyvsd6az8p4rnJt5h1Vpl2RpHJBBt+TnT/UYWSORP94VeGfsAiZ3e28tXSPkZZ
hYz7ddAQfVSomrkQDyX8z3r8CJ9pn54kNyj2B7Y/o8zSis4zgHFTEp4qFYD/h0IX
vKUCV0pk4lzOmkwj140OvFQS0ma3J2zeEbcW1FPPfsz8+UnB6+Mk/u6GapqoOI83
ffN0EFAoPSEpLupIsUa4PMw5Km6h6MPh3vq1+b+NbyY2WT4ivz5sDapWH8juOokL
GEOqoTq7Jr40S36JFFbpicXkemUqIgIl6UTyyDTRD7WXYdhksnxyKygUWJhkIW03
kxCJUp+Vrj57fqyCfXRxAW/voxk6z9nGEvFVPAUmLJD+Y0/a1m+lOG6y4fSLdfnS
6fKp8rxOSJFegaFW0fX3nYmWl0S9vJBDtR1ofxSTqSZqT2tiYZNpMdQMAS3SJoyL
IZKH14zDa74wfL0U+NX8M6h4CKTEN0h6V+VVn6EWmY+GYygBAhN1PydlWBdn6BJG
vj+UosqfN2ldSPV5NgivT5Xj/OpEamdubnjFpdv5sRqCQWuOEOnCe4f49yudaK3O
X5U1SpGy/LB4nSTk/3g44MJny+KhgdRF9I2Icv3hJL+FWZ2Sc95XaFqYPsP0OdAF
zy/DJ1rHshZq/jBnqP60kqm3aNRiuCzbltDRtheRXlLhXVZmJmuoEqkC516vhxkM
p/MVaBDxXaTtxgsnmjT33s0cEYVulNVoMvlwk84/eeV5lx0HliCHoN0kZ5skDM4T
I+TZoRvaL4Ypkib9pBlxWIc0FEh8Sl3/mY5eZ42joBJ8pymPafc3JPmXkG+gGLfN
EGy4faEAiEcpaM+tSoqqqtjstyzwNCxD+/na07G5mvs0yNYLcx415a4eeyngOXKf
rikLZeAUagEK5s62jFFQMlCt3m1Mtjage97MSCNPG+nzzjT3KEUIpLTwSMBMwhpi
1GhO2fyDXIAhAO7nY9/Mrjo6SvTLlZVvnMmLS1F9zPEjH8qmvoFWGn5kwQXLd3kw
lqc9sOODJYQzD8yqi36sEe71m4gBXW442JKvFvAkQ9SVbhcSUJkxMkbcX5rVO4iN
l7Xxh3dYHiJNwLsYCR//Iilz7hUcue880qkCbgXIrdP6jNOKvq4v+QOpZfRvqOed
XpbzDUGerNGsJPCzrdSaSUPpnAhzdOBlW9sErZUPa0PCCTJPkHU3bsYhKPVGtTm8
RXycG/ehHXJnNlIz/zBIsl6WyOmLHu5XheTQZ8blI8pOkMW6c2xi30Z4JAEE0jl1
kXK/TSwJsDPVvm3YMcbad9+18aNw9Cy5mH2kNQUX0qQm96pUlT3gB1m1l6TJETUf
JLLNo05JKFy2QOyoBaMduoh1DHwFvmDlmBPDBYPRbs3Da4svjPKwiT4/DA3ADGOa
y8InPGnBYLp8a+ELavwF+hWt4d63OwVwZU+z+FWhlCZsv4zYxmvNLmt9k8P2dGdO
MzK6RWo5SmlKfgnsQ98ZtiVy+OcYhlGfpxfmWoRNehjAB8HPVKE+WdG0tuCBuUfe
QgbJ7F5T3BIUPt+Nlol5+hbK0Q6Wh1vmU2sk125deC95QDAY8zFDMw1/i6kXIsie
kMs8WW5NnPO49zOzUgeyn0QVOYPxgkHWAz7z6B5JlZAfjr1MUbPtJzO2FW8GkLd9
SZsA0MvNVTjJjFOTpjwyt1fzMopNeWky4q3MfBUE9G0AIiu0usvc6P4ER3GSAKV5
gcsj4yE92Tp4NlPW2ynkATjOBAkzo9b6Jq9b1buyMu8HvtRL1w5vhcNhj2Tw0Ygw
v7ZS6UnRZk/zZE8zM679RRwmuzy5UJabI32lBftST/9Ve9KSr/T09rLju7z11v4o
E0e5oIXzx5wp5oWec0xRl/UbofwEfjAZVsnsIN5JbIR9C82zuwi0daWuikcjtv39
8FvbdJ+R7sZejBt/MEokTB6G36yu+NfJWXnQnKbCqcM1XZBvw6KTNesulj/zCg/R
9NB/6AGgYqEYJohixWL+YMFL4DtKfbTfHm8vi1oSWxKIzt+bWPqqiRPw9rZhaWXl
2d7mOlVxQYKSxTfc4pMIPFl3k38pr1HORYAx3bV3yQ2WCTJoniWh4QcFYU36Z2Mx
IFEOOY9GrL7WpVdgWJ7gIa3M65QcV9svJY/+hptVFN531XGP2Al63m3jJzmDpRCf
GJHTsB9tw+iv2j6B0dRLDmQwRwu9vKvZ0ZGoN97fgQb3FjxieS/RdE2HIAuSQT6L
FcDepfFCKgqWXq/pVTlxOl5oi6gHDm+sPK5DmNOh647JKOroo+IDK53zuRXsPZtz
iYWvAjaQbQMXO9HT5nk+sgz90+12Wkk6NmvTG8LDYz/8EmJFTVE+0URfBkledIoV
6GCekgO9vOewB8gjy4wgGCJFINSnI9OgZQrAbcLcGniM9b2QIz1mU8aGvYeaA7Ut
6VK9FdSIW1U3jpJ/wuGoCqpAXgBjuERirapn8Hrr2NSdOyQuq5Ei+TNCcW6UwFR3
+S/fpd6poHNo2ZkhiFu/GzTtMng3n5JEuIYWWo1RJ5tTT9oEmVwomCSZpHVdMcN6
dcxjxak3Zp42h24sNnqImrla5on/q6ngvZFoFn7bFiFsutbEqr4FmNqYwTtEcVsQ
BGUHH2ht6+4GcsqHp36hC+X1NJ+JtH6h5u5TrfHubq7fXAaTOSLaF5RNOFhP3I8N
vCPkSAzSigWKm8hVZRTEG0Euwa/s7SmpM+r4Cg5qYuOWXH2wXc14r0ZfTL6BYRrI
K6KMKHuuqbThLMmMtZO8gixtKb8Sy4KO1KFwUrDn4H/5EQaGAYzVJA/ZzeQKkJiT
mXbAiuszSKuZOvGjHj8ZdhHleV5atwQPx9RCG2lQiPUGw6DrfkJ9SdgBoAQMPhaa
UaOaZUNrkodRJi+4LDNODvFFFt3sqUclocvI0NJ4EF61ZuTXeqViraS3OZMdvJgn
LFxbkdmOic+Y82m+NdfJsqKjyyl2PQsv735qSWGbasqbRQcvZF8QrCqKF585hORN
x34pRhh2qP8UrVXlF2xXY1TtU5McbCULPDmYWWycVWYDZJ49gxHZk/qvOWw2AIQr
AkuP/3hEnRQrNpPIgNMkPV3CXFKSkHXuYBTA8mai01it1gxj4AIR8FWB0EuTnT3A
pv/UIXIX6lPcs0mD5c6TxkCMlHCQ9jcOW8WmUSk/t/ZWzooPGIMV6LfIkQ5xrAam
lQpyHW6BhxmL2ptV2mVXMikdb5ytIGciajj16S58/mhfRnUoDAbH8roTPKDsqc7H
+L11eG2A8ol7eY6IoeAs54XY084iTTOTPKEuXgEmqtzZnkDeJeC9EMvcUm5awwKt
lUQG4lbb7YXtn3icq0mtjFFVx8yA46fiBS4jnRKPBGjg2ea+geEfABjel9A7Awid
+k+UuRxfhfhIgoZwGis5zvflqBRLSRFjp7A6ODEo6KFzz3+MSTDJDdunFRVLEUeO
FGjpdjPzeeo8216dXKEtbzC1W91yDtCLpK5/MvZ98Yj5AR7rFNupHZfzQJO3/1eb
2ZxiGH/YXd7mYRWngyhUykM3WQFU5HSgiiMfB90mzvrSvezfZpdqXBsteYKaSRg4
VggVJgSk7uBmzzgsgqZk91e2a10yJz5GxXpuDE/f/UuWfTOyl1Ru/qNT9Y+Jke2J
cAkh4OverLGIa2uAu1GYf8ANr1WvuZ4bITxEPbrCiIh2NpqDeSbWUWXRW5gSh+m5
ilVrxFoF7O8th7Hz4ifhjcnGSIQnDWkWBUnjUCdPYISclomgHvJDrtJmtEp6FjB7
FkCenYpG3H5mIFypXj2LLlibmHiyfOnnWOvt1wJuD/HK4KmxV8VuAihntyVSnccB
ChNNlvth/kFB9HbsxB3KzynVDvDb9nWwYt43pIq6Cv3DQ3KkbHa4Yk9Z5Fnr2IUJ
NWm6pBbAH46+/WNnV6qEgKnE4PCpbYTdrQn7YlcIQ22Em0lpBNNu7CAH+c2ZQ7DS
unVBzKXZaq/HNGKrmyo11962C9nqTYfwtpqqQokv9O8dKBnlwu7LfIL7FpvX8Pbb
vfV7wNzIbtqMIHHkq26SsVl1I3U4Xy1Mf89WiLz8D8Rm5/i5EddD5CGbeb8bYQ00
bhgFI9RHYGuzrwqKt6AD7DFf9DwBe+pzSTAneKIe4QLgyJDsHwK4bpxOL/XUAeXn
dUgTaHpE8XToPeLBnbAbZivBnq897JbLqaHtQBRId79kQRWhERIkMMIsJGDIl6zw
sAodVA4cVYJsFhUzQuKfSZnlci5n+h7i+EV9nZbrs9X4Rzjfgl/Im/6gVjo6/lTz
rB214FeL4Cq+vBW+7LB4uOYMgTovfQy3UErzYMPMhIEoIQRQcsdd+kOVy+tFEG5J
MjUTOrekMMHDX9376jBcahPh331zmJ+i+dVdq8Nmb+vkhjWRCFmVpu3pen0IY9/f
ZE7dJggz9iKV800MkBFYXoVgJA0ippAbi8L4E2j5dXW5aIS2z6vQvYOzy3uudXlU
dx/GtMlpSnIb5M4wo4v0Tt5edzLUFxEtybJRA3yJ0SO1DktjFzbh8Svyv6fAdJup
ma9J1xm7yJUCP//Tk4jKmV6b2bOTT5Iwd2WO7G1Q8YgnVQMG8r7+AjHN9Ut6cGg9
DHgtO+tA7LdEnymMcGxI4LFp4/VARLyYFYCcAnokR+ClvvmU+lAwa5ahZC2OoSHb
cxgC9g+qF20UtkUNIZnB63jzlNTRq4ZBDLW0hmOx+Uyo2TpZtSKRRwNaR69na9xM
rGiiYPHsN6LJEgsi6TMZAgQAAZSwISykdZj2KJpzdS50/aTho+maaQELwnFz+gC9
gEsbChiYUEWOya5o5hZ9RDhoV70kwYe4zRK7kPONds81utDSPAL25Nt2F8G6FMo+
NvvAH3Q30K4YsinWM2GGDo0j0XCqWgfV+A/QZaoyQg03ujH6magZdbuHtMpbTOv5
mTnC/hDTYEj5unWPS3NhblTHjmPpj2Z/LHtzxD3ToXJ8lerzb9la5UuKtYJH05Eu
jR49lWrxR6vNQ5JBtN/n8g1lgerMmLvwhsBzyTBiJQuHPckGCWTdmvsNNFfS3d0S
bJXQmQ6XTtAr4TgpHQhyQm0FEtdBvWHujyCI+odv9jFp023pwqQvDiSvjUPeBIlJ
yLd1Fub0ZrVYsUNeNMlQg4r4RV5EUrg9FOQNnThpWUyNFjZWM17vB3zk1svkjJ6s
UEC6JJFigUat7PrNGp/2X6Q/5P0+lrKsyC/gILvDW1Lj8ruxACy1H++GJOLHSSUn
V9L6xXFtCPwpIb6uETENp1oxrzc7K30JY2zpO4CfnvG4OQ6D5ubA56j2Q1t497L1
TzGH4lMi/5t0kXEMtcNVE/b0QKKj2K9FQzXA9FoiQ8P6S04NKx4fYq2whqSKEhPU
SS5IB0G6KPNDs0yh5ly3sjK+pb5oVr+E1U78G+qQh6pKz/yWDzjYFdikwGRtoFtO
rpnSYH7i9BFUb8B8fogFZvmzfZjWcecZvwtjYAuiOBVPtHH6mA/sgR6VpwduLHF8
1gb9ToKJsyy2/kITsmVhiKpXU/u6cdiDBxokkCmXvBKyWr0wWnZTGEALS+6CZwNy
140EJs55FPWja/8Emn5JssFPVbPmEoFpWUT6xOoW9u89oRka7fgfCd7bJkFvTCuG
xA3N7Ysa2YjI/GJuTm0fzWw+tTLrbJ7Scjy5sVEZui4kauyjEFpfJjbbGGevxqj5
Xe6k+vduyg5n66gYqpb1HUWl5dPHAvaJAoqYSTcdk3+QgdfRBC6LxuPmFkbzGRAg
uTHl2hcnpUJLDnRE16TYEsJPmPSWiJkDR2R2HGEqY1FkzEEm6DIzNmfg3uDZC7kH
On/2UqQ3BoP1lkzseO5wgqb4n9MEJHtNubaJ3UC0vHDaptMXRnS32Z+UMdl2E4ds
xCr++gvXvYQ2H5P2aJf6KVGxiAW2QnWEeaqWUA6ufG0ATHhYPNwMrne9e0TEl9Y7
BPlvJCgAYWAiKfQYXNEBxICKjqOSl1Q5Ms5S9EJKb586eW9aUomf9XbLKM9qNT8v
1uzWPQ0XNhTuOalhO0xU3ggQ48uUYp+WMS/usOPW66YYV+8sHSVZYvJvtxPr/S1c
TODCZtdafj8rIFdUFVkAHjkk8vEeWd9zK3mQWgB8VDIb59KNIasokpLlFqz2d0LE
L8gvTM3vCA7hdC5rzePERUxdneyeRppCpDmCbrM/1/eXlnmBVJ0DDgg94eHYSJMA
YQsC6y1153Wo//eXmitxh7a3Ta1vUcxuRCJQx1LUnnunvwNpUusbtgjnXsIDUlq2
kEOLtVn6s8EBQmkS4n7afR0F1pNhlbnvEzlAgmcVQf+7O1fkPDbWuyHPkPRZKkwA
eEMn0G3+4wZ/oRVZ1NCHIVXSCqSfk3JOvpCfN5YYb/Yq2WdZ3jRMoZlX83WPIiwo
T7FK5PPSJbAvxHdV03Qc7zSrSp3pXQ1+Hz8slTesJkrmwe/rwnHydZcZ6mT8KXXY
O3RCqRs3pUWTwi/AzJIrs1AuKB84ypu9ZQsGgY4jz1WlHEQmCQG6E9OKCgD7igN5
zXgOJdlV+jKvNzk2i3P4Fx1lojqb2nREa9VyN3/aTkdmx6CXGZPx7fgyyxXgvYwS
jWJRVBD0H56q6JKDWMNBRNfpn7A1R9+71TMbxYwj73zmw7uCjJjoDXE8SvZiL/gI
MjZoorpvOe48QBD9KJp9g+uccUwCxiD6vUbdjqf5EXrm24+cAi6LISB2sOfzhly4
7h6HZESqRrPLgYpuqeqA/utAigpQBPTPrciZ7NxkJI57jupdr3PnCnmIoxzEzH/Y
+pSHJCcDVxOjZfcpW2Z/iDY1KZDQU+j1Im/TS0b3UJn+L5cuLQaQEmhnNY5/5PDL
pGOzANkybRxQ0vJ/MwFB3mEjwMcVuyBttTUozilodG/QNUvUQYXqKjWJd9OAwO1P
xQrOhzEf7DAot6qAZ4NQDB9FNxc0tsEYMdoaMg4c0Embk1soWShLBWrFEIPbZLKy
ag9+vNyp+s6dbE0OzpQlcl5HWgxd5CXY1J3wKZztSgzpYOWKXM6etoJ/rFQCMRh8
YU/IX1d79dfUGbhu05wpa4szZDvGGXc+6KKUTRJ7TB8VNp9B3nzg3leDagHTx0lt
A0dMQynVLOTKqdDBAPNBcBijmOCdfFyWBuasFKJ32BU6Ci5RBDY8SpS6C08IgEqU
0xutnWHkwVOGr+DPZa23E0hqhWAyEn0uHyJQwnlnOLJGrZX0SzpaYrGboCHjvv5o
UHhQYfja3RSOP0gLGe1Er0m47V12bARF7TaROGs1JPv03VCTTxwGlgdT0TqpQLdc
dTFoYB3Ys7onWlX4vvF8X//GASYdQsD4M+N69d/FwJtR7OfIqcuEDAVc/hkIDS/L
lJHBxK5GItd7qOOthnERJBqW57xwkTw464QWdbKHdOUMyWTurk9tffgGksE+wqZx
Ca+z06ReQbQaZBHIwQNKJ//UrgL0jxk0agnKx0s0dVi90PzsbGTxpqCSZT9nAYe5
cGYt45k918soHE3xCHduKQJbl+L1ssi3ut2fNNHLvfgmowTEa7fVx3bAsS3i47ml
gCB+wX03O/wTdw+nNBfdkc/1VibQtVvmoa0U6NT/qtg3LXUOSF8wuT9Ev69oDAQn
i1eRtKdtpwksAgbYk9CcXbpkOX+31VNjv/jpiQPpTrAz7uwbMZCfewpqPbINM9qj
BiTiuGin75nmWwp4Wnl1Bx4F018XST36MU6OP6y16a/tfOlWUILouSP2NSRTS1Wj
x8q9MxcQZPvSpdFXFHO55uaz8KeMwjtX2/CnsXfCGI1TVZt7HiAu8ukm8BbJC/xt
53CqTeEb8W/fjbCKE098NHxJDGnLVZieotDwgjOqpefz6Kv5ROSPGWam7JjxaFwa
vMV8blYB3Tp0uHIq0mLq2j5/52oqK0C2otldCqIQkHJpegSY3NaTzPVtwx9Wi1Zu
6O8ejD2v2BZKmFFmYhwc24TZFDEVkYCr8bFIrXobI44Qd7TwpvVjm8VbC19GlD1T
qX//khaQfknjkQg262zdioqo5HxBN3pLtxoXf5i6pPr/K9+4d+Z2zpf67CpirxWX
tV9xUnMOpVTokpotJcKaBv7MLazQUMJiByqygY+bD9B57O4qnuIPW0XXVEjZs918
vm13QWaVDrEuxFhlrldCMCFf/aHz5lqB0fxYltPGT68ZfR9KyxERdTIcNK4Dumde
yrAWv4ScOrygLX5KbweVzbPmNrXELFb38AjpiQ8c7IjWHGe43+0no9yogU+nodfH
rZhB8eXlLJmhsHalezMV7a1xzhJWa7Su3GxdJeURIlRibwMkXOJ9YErVITK/uSwc
db1s83zjDCeIXGjqpGtC8fI7qhckwejU47GQh+cATbJmEE7OFEsx3M+WB87L3B7z
4/I42lMedddF0LV0iD05sltD52se7CFdBlHdtkYpj9okwqTZ0cRBDLH3TYoN9YiY
7JB4+L3Nc+VGyYza7f+eMR3AeUnHjEFqA16rIvmm70wOi2obEW7NNCiSk42BAJdO
V21eSApQrDKTbJ9I0Vqlebsqobi819p+S90qHJhudAeICQPOTm+XlRpRec/FmxIF
MOunVhtHi/gnADCvDRcaf8Q1wMQrdPR8ZGe78Iu4CCuuWmOgNQnbrPMuwwA6RRp6
9xgCrwErcmo2n0zyLy4N0rS2HUH4TIEbiTXcyFeWph2lrIfr7cH0baVdUwLO6xGD
AqgEhgdlSKH+VFQL0t49tU0e6+bEqVgep8/VSjiIULT6DDPXungE40Fngu+Onxmn
dFEM408sC9S/czp4NTGi75zwNzP0Cq7nRP3tuPa+iP3o+i5lJM4oxTAxnhmVGSku
RcBVioxBiONTo4hn6tT08cDycdJhzk5AUMWk9GiyOubShTbmQjm77/zCFeveOqwc
xJaQa2LjpOwx0+/jc7IAHPBjzhbTbGILI60uHR69+CsYZbJZBEIiqjUrF1tcUjGt
SNGSHo7n82jTLqYLGfYUGxT+WeYTgdSTWmuME1qhr7o/h99RdNNQ/kyTTXukEbAz
+6vgx7zffJ0I5G97y0VdeX90rPgQUuCwNRWFTxzEDj9N9mOOehs9Y/r8IpX6mv6k
UqTPR7srWj+ycyjdcmhSHvNX8nB6uu69s9lWFH6oCGXMj6zqD1YgtNxTUFaS0PAI
DRrsKyipFkA1SUMvhpIm2NHCUywbuHRV3SiY7kAu4dh+foyj9LCrIICODw8bRnWM
kl+74qklpzxbmYlrqTGHEYAwa74TaQdM81urqnyHXaT0rc0YpuhoirDUKCTaGLmO
dBJHaRSxpTYLZ6IkHnNpCAFSHjTS9X1CU8WB5RvP35nGQhB4SPjlYjPs3mgjdRb6
Hshe8ZLIKIX0/qclkhVYNp1R+2XjnEDJNHMNHHwoybIi3S7sOXPDyBEtGLkKZFGT
O4WHwf/TKJ1DfQTVzN/uvQoZYiExhErUwp0zqJ07d1yC5pPZO7nSP0d8P1HeXHod
g+U3Bt2j9qnni2bK5QjGMeVvJ3l/0DsVcYSixbjbto78a3J5xhonwOflOmEJKFH5
dqNtI+DRGofUu6apZP/s5d0sKlyQVEc2koIfBuoOVWsxM0ne4vpW2yhQVRKMSnAk
ZGdDdx7gSGq3rXKgNTl7sJ4cqbsmcQ54T/XQx4WeReKcctkgGLSQAi3p2YbiuXiK
Gk14LknnuviPPwC9Ux+guUcpXm7F18QfWxWXH4J2YiC3LLGaBO28u8qen4qcTcTN
g19Co5zhFWXICi4C13zydOHi8zKeoxvoSreEvcYnGcCFCxe56oDMiN3yFB2JcHAa
k78oJrpuNfVmjKEN8+GRcy3btRY2aljXgYKSLt/LZf7BHwtPZE65sx/MdAphyWNr
vWs6G5Dg4U9zo2BkXV0MKzy+vpZjTJdL5zhZYGt4oY5jz7t5XdKgR5WRPfLV7T8M
5YrMPsP9snul1TwB416eG7kCssp85AjDrhCdHHOhy7dVPm83c9todZzR8jENb4er
VKM8IZh+POswbi891lEod2cjWjO+pWZsKBKwUCGzy1azu1ii7CP9AAADOdWklwqT
YAwyu/IULYUJ8EsKiXAR973feqowzEjus9XZ/URT5AKJcarlTIhJyv8DYdefYN9S
YD6GTKKLIhT9TIS5OvwOCrjyCDjI7jcng4VrNJrva76skw84MciA4Abbi5jWjH0B
JRKvNb2JNYyv9QmXf28/DcM9UkIDb90pLx+AAFFPMcUIieMBji/hyvYoaERGpday
yrYIEQY1rP8UxmhbXeGeFf6TbFRqPhcVSvj5th7hvIWVS864ZrSBfqgSR7aR0lBh
rAZxdeDEzJ++9k8yj8LCuiGCMxYnxEZGh3awPi1Jk6ZBecwBTvB5HAm8Qvo4GzhL
ubk2SGXfnLdlgpuIb+ApROu8JWZomih1lbnrFQLV7Ynyy3N8XsYI4t0eT33ec04p
huDmSAdKaSdoefib6vUfzmrPNkLs3lM7pMaavy5/DVD3mtLV+YpU4puQaxxBWJI8
6V4NCxlClb6JAnQIyzdC5smpWPstg0ocp58PLrhWyUrNRKpdnBKGDtOiwNBuGTCA
HSPVs+n40WaQnkzxeYVgN3qaTOK1p7HYSyx1qoOI7LaYQWE4FuuRR3vYIaGNZ7dC
8/NdSn1/RuEnXBIdD6QvmHo6BStLyGATiuFf/uyi0EsTfQFWwYvjOelrznirtCTl
WKN00svOmN89OaOwc63m8qhFnHrz+osqOv15HEeQc/ud6KWAOBSbCxIOLmyeUpuC
D1qm0P64kTOAdvo24xlt4LFdHbQUMT9/CrYZEq6BaPpzkN7nf7cpKZjnWD0eei6+
yFxEHE+IRG5RMU6VjDaYqK3LJsa22IhyJUkwHIewNUPEyW5995QOc4Tl1UmGPwCW
4ITyfF6zfYnYDm2zRQwXEcpZHLsz+6wcZsbQ7G3Ht5HMabjZqS+5QuycVhia9xh9
2AiCEQqpmqe2AQ3695iw1VdIMO7hyrP8VTVr4sS6WfLsWZrMjEU1xcWverKOxy+o
qMscf62U6TcSEBOgtQjuBRLU6XxqVLrjPsh01sHKcwbq1fOp/363FfXvWNjI+U5N
0nm4M6mQCqgOYg8fTm+rDm61GYeuPFa6zbTa+spfnGrypYXSH0i2CwoK6VbDY9J0
1k+gGpSmIAtfdBK12kNb6Tr0VAE8l30Ihwxa6dRLuBY+EcazR8Tbp6Smncry/feI
yOf2RXXyB7lCtfwPW8zrwvixWvS7XYF4pbXa+W9Tr5fLL3i0k7lFeLzsAxcRHo01
Hl9B710lK7KxaeAcGTow1V4eJxpt42DM6eNZ2TFvQYbeUlQRqgZ7aInAcIW+Plt0
Rz4YeVdPVC86/7RmpmZ3H2qj74Ue9+H5C+uV+sqlHRZ9RtSci7OsI5N4JfLhBF41
GWKq86G8gdfaXfrcH4QBGsVNgezjotrYKnS9itQ7MTxqyJCrsOBE7zdfkExBsJ69
QlB+5mKRtkEqTMA+CKO4S5ZcawGeLVFNGMnE4dLD4xx3aGneIfNBoktxnMQmaxwF
wf4RCvDpbEev3TSMTshj2l5qbexEa8XiB2K3khGuAqJ6ssHnqpPt1dKolymBAvOP
ckS+9I9SFH2Tb5RY6vmClWZw/T+inHhTsqSSvUEwGrcnpbZ2EnK7INRwf0bvGKq9
oAGMzT1azMjZ9Tdz1JWy9URvb+3vnfY7eZ19KRy+1FQSSYabbdjeJ5Vi+3l1UtkJ
WoO4BQ5u7EUInyR1p2xzMKzVOaAepn1X/8GxmugjwOA6rzqFI97PXd3RIfOgVl3g
Wk2PFe3roEaVvz99FGeHlZidY8bgocoXd10XcaCezxn0SklHp1mo/9nQL/IrNJYK
I6dvr7H0a110j6wtVldIb1pd+/ScFjBNT9bewrRZEFGxsNanLT0fL1Xfzu15FsVF
7iuJUXOQjmkHTHzf/5s/6bJ1Ap85SMi5CufIF6MLLerhYpt0k/KrK5JVhCpzTwMq
Kpdak5Ee+jgp0kApgHM1NJiq1a+bflFNkcBq8XI6kRAMr3t+bacXdiQFKiScxne1
o1LTj+OuZWv5mbaxMR1Tw3gfkwJ1TQBU1ipcAtCoukXC2+5p80mpZ7XcobRiVuT8
m8i2HgQQCZJHdxvkZfsmpJ0b0xiyW7YAm1lZSXGAhfiyxif1LLiQ2RsFmB4SRxMl
3JtukOwZR2eKwj1dyNOl1LHCWN/LQpbcKkOrQf8xapDoStHW+U6r7IRnISK9lxuZ
hLCZ/mcn1mk+9Ptv89Fmr7OVIJeLwv4r99ZA0nFHKn61f6Czq5SGYVU2wQg4otXB
IWK8n48aUIgk7IDWlJQRRQbw2/45TuJGc4Xl7n9dIUrkfGehZXsgiGMEuD1iqpT1
d9AtahV/05JxG9JpfwBEbfv8yJSeBqhYARotbK9/ltG5YuGUNI243T8owezGmV4X
MClYNi+CLcUrH7yLjYgcd7hlUZYe2Eg9NlXRysaTmDo4dCdgaRhaNsJXcalG308A
DV/7bw+p0bmBV/xEsbc506NS2XKOr7KQhqLxugppyqK1Gm+0D9ukvVlWfsttREb5
oU2FUwop3xeKnM/Ag5RJtE1mpn82DgNiOUkpBJuxOifUcmfqhqKPBAfE81U4oHPX
m/94xGNqjqG6wFP84VJRa+PZkoU4WSfUlGDTeESlfCStWK8+PsM3+5BYW7KDMg44
Av9gFST0rdn3/NqJZJjg25GBOIM3gjhYJ7HjRZ9MFDE/mq1R4xZ6p3+G7hsbauiX
ASSZPXF+3ONOW3WYFmKSsANrdwVKXZUwkNlbzrFXKZao9iehVl8PzbQA4oIji08h
ls+gkg+ZLdr3QJFj7hIjouxmQPnIwPAP4WxcSX6piQlp0zQGHo6vzoVOL06PA2fb
ZH07hiChGZa9AlUVJPMFQrVj6QhZoi2RiMP2pS7wtFSLdy5zyuw6/IHe6JF3yDNC
B2BIV9Ujv4kMGfe8cX/e4UcaC5I3hTDyQ7QDrWjZe8WG4eILzEU7gqvVKWZJ3wVs
auk195Mtdt8IwLs1TvXN+bzqTedA63GR0aRDY94jwssJ5+QjGCTjKpkgLOwKHxVX
IsLdsyRKuFctU7Vd3G/jJojnOhs6iFhPANTX+UtVJ2exkN1g04P/LkTMdKFI61Rv
QzQaGrQ234lvhcvmR4EoX+68zwj49ANisS9xNLr97HZJLnxnmn0QzwpDlGA0p9Bt
sEwRWIb+d6d7MxSZOOTgrl0SuiXgd9bhVpngnzCzHx9Dr3r9rjTCKligPN4GTXNJ
aFF06TDo1AdeC4cFbRXfsYVk3p+0i92JpFTvdljCFMe/1N+ZdvOveIo7RStnlk7P
5uhL2s6JpzZHjtTLODqVWyII19wWTUWaL4FrRRF9eOX2kb6iuyrDpb5/vT9W4uGh
wntkb9CDVQUV4x7ZColbBmSRmMjPeiGgx35eD6PLn0uVsF/qp6Aw29Kwi8w1V8Yl
QXAhSjz1t+Oy282pIqDj1itDyu0tPYQ+g5gQOMp2fXn7nkRYc1BS4lmwoKGKoPAw
z8eywSvjkutHjltC/XzULedoyVA+HqtZhGEcyOzyBNTjVQlY3mIgPu5OTSTefc1s
knixSb5Hz3XrYA6B7AXpeve272eo+d0u/qpbQGC/EyraZJBKcpxcX3l1BUw+Zmct
yU7WYkw9OiLpf6Y3bsKzSNG2sKZh/XCKJ4xeAsNvIa+Gk8ee9bUth9T6F41IWvQ+
yZRC3Hx6Zv94lvimAqo61cvUSGGK5RLX8CJSOFPr0U3OicTs51zgKatMA2Oghb4Z
LNd5tnacSTpmWfwWffpCaRlbOkRd6YgSgVkn/WLl8hI7WZbKfrrrJg6OfzCpAujO
NAIycJh5pvYUfsIYSk4plChFS+7Wu9rcqQLo3f1kwtDepW5XvRS/GcGpLGrhh7Rc
Sdm+T1M6u6kAMx+LCrjSiR2Hw+qxIPqfyzFiCPGoOKi2JIGgWu5FxQsJx3ePHH2h
ZFM9fga+W1JSsacMSDy5GXpNUU6uahUIb2HQEnU2bN30US8LmCBlE/APx/HvH59f
lRlZmuDyA3HbClbMGhnV6JJ8qP/OPVb7wddUAn5RPnOwqmeOHL4gaS+zq9QKxB76
7Ochdy8i7aoOyysvp8s2ciS5uVzSvdApnDylTvIGPzqCVsbYI7yIdMxfVFbF+W5e
QHkcMigySIG1GzlulWqxwylTLISxxXIUe3BIGNmjz7RS3cgOWQD0QIlQUCiwXRBo
2bG1MyMNNQRWwn+elpnvRM3qlwnGgiYmS72uuWKbmfVu8r9c2fILuj0OppSXTOyW
AQ7p7CflblC/qxaOhcWJsViQhC9DKFSEsZcOiWCa6Xx3bEdonIy+JfzUKviVU3XM
pSsHM58AuS+9OicJQtuDoveWKQdCBC1IjmGVFvMdq7Apn6y2r2h/k4gxXPDcIuAa
PiIktli16W89Q+VSguMDylQZyY/n9cVRifDQU5trAa+CyFyMq/cR1pvQHPZa/XVG
KktC3MLtb42MpEjOAJ0/5Nx9Bstl43QJf2PQ4pkf0SHemguiWXrAcdh5KWA3PG92
HUbGO2W4RkR+DpJhqOtWeJmvJR4ML+pmO2tHpsavnmDVjdfXpXQbmsLsN0eP7jrB
+AbrmvENKI8c8LdQORYOae+9djarzWt0nou5+FHk5WfJpwHiDpjUIKeHidRwBoth
BO7qa4pspBt1fUHu6kySWREBGmjQCtokD1u8mq3sdoiHKDhjiif32MoO6j7JRw9p
uaECgaMt0ghJooyjeExn705Ct8cFDbqKxqEPhLwqkylRCGizbfSi0+aYURmbinSJ
ymsFCH91cq23oiNtTD1yGzWMri2Doe3D1uiROMw8dzdm0cwaqzvxUkRHY7b82lCJ
p3dss5dX4ToBz7dTD6ZqQU0d4HwqHfcbcrDGKmRhh8IYUYByNU0suDAV5j1qJY7z
/dL5YaC6Q0A+tc9Jt0d8wTHlODSoObzUXmfVXWYvX6ah16ALMEz1xUUp3qfCsLLT
meYaHCTHZaksnQpg3P+34bEUQv8c0qEknX3ZaCVgxEPaUDszrG6m7uw59RLn3pkO
38wju62Rh8B/4fIHuNyYym8HlTvRpw1H4pUxc7ox67RbvUkYu2Xznx5eU80FW65a
sAXT0t4A5pn5K1maQkcv/4iIShpr0x4QER+7108lvs/2VrcyTW7ZIswWdSCWkouo
XhqoJqnfIpHfE0f/YoOljnTwz+zXiZZTg1/qCmmD+vif5lYiwfa5VtNFWO1s/+z6
J5aAvw4P8aWD6TKGL/dHdVhca+jOX7v9NYoSMj4LtTTdiBeBdPWfZqxrY4TmhDZo
x+UC5WBlY0KKMg+/xxQVmtdPKNoH4Gw28E5qyPWAtMEi+GOCKs1Gfn9MdXqqoNoU
Y55wmiZDAHM7dcPLcs7oELcyICxJu9x0MGKhdMiA83r29ltYsvCEOsqdDYNpGgJK
q3+P1nJ9grr1rUr0umcy892//eYkEGg0nQNqcewNkEg+LQW4GUmZ9s3kHRT3oFvG
cZ+THPYwkWqOo41raqZDJs2QaGSqgWql5Tvc/r+DejbVpCbPQv4Bk9BhlET4D9gF
bAfnVtFrnHxV9rnF1jJphH8/kapVuErgHJpCXHG0Z7dAheH4vxX7+W3Ww/QC+U5z
ckbfKINSORWRzL/UyZuuFoqumVt2NPCl9WFrabZPTZAR3KK/M1g7mlVLEX3XMkuz
SRNyaNCXFkKCKuwZeyzNQr2qyye7vB+fdOb9bjhbh9mjsGRyw6y70eV8YPJd4tcg
auM6xwRgnDbqIECaaJ53N83TwFfYh2Nzsn0youhZy0FfzaYknY4aBn+Y0qAvPuI1
yAN/8cGhEg7zd7GBVZJXc/RchqI9gm0kJ99X21kdE2JF6IoyxFkkgqaOjNuA3iHZ
wzz2j03Y+QqFcDHlsIajCE4MCQH20sVt+jy/6yyQyLxUY6ML6LdvvO0ZUxLRJhYc
5pGb9nuh3dOuV3Gv9WPw0qkT/Ei9O8M/5PfvM+pxsbJa6I+NMxH+d0yVyCxtzZhk
lxifQ/en324TWtO8fNbVp1pNOFQRkka7HVOSxWQ8bAfofIXmfkZXFKbToZRt117F
+ywVFvGwhUF7UR6CDYm38XcPJ9DrSrhQxQeZDs6+2tiNA4xXhL+VYyAylKCR7aRc
yU1BMXJwKGxSUAu6i6TMP/NuTt1k40dJRzLokzD77W+iurzIbmAQl2vH/z7dtt9q
7TRIzFSQpnGvSORVeHYllxwSLrrSxd6xdfyD15mrW7rg5sfbAvLweAYp6jy9JbW0
VNyqM6FffNh62djL1XqP8DuGGw2ANSyl41Zm05i9xJhAhYVKFy98VVRlvBsRBPqF
+el0J0htZO/Ayi2D6uM+8mjHiEx8XL15psTuN5DzN/Kn6AU5A+sSs+MQkokKgIU9
K07GQE+Yz9UaEZ5grJZDfxhWdJSxXO7nYrmNvIYa7mOePA1q4NXRlODrl17pMAgl
HT9THmfHe0M64+1yYkJ5Nmuk8jfXZJBkn8Hobj/wwHjW9UadDgWnEYpldYcwzirB
NSr9qDNTPkRBw3IXaLCSucgC5PVsokB0JKnWF1vdLwu/eLMXVjXtsj1BnaiZhkV4
IvKgNUzJZzQQNkt2YPBgzk1hEeJQdFZbDx5u67stXKcK9w7hsTR3L85/QVi2yuMJ
t/EEAU+eV6XRYfe2T2pAcH7LMU2MMefaooiTkKEskoBSGgkypoOqKH2RIHlpNiVm
zjaUJ+CBNxLbecpVTVkbcU7EiOzWiFU4xrAx8woTO+ycwwAKLTH4exz4q5jSqIzD
YPUiWgcIVG++5sS8is4UBnRj9CkfR7L3OOyXFa6OlDdj0Va3puFYoRKKJX5SNiPx
uVTAwmyQS3NmJwgIkr9l4m2uF/Ehnf6ee+/E0ohpEIqUrf+OeC3t3DzEzoof9nrP
Go+nna0fA5ilPbiKEC03IcSoQTNyli+fPbDyRRmdQwHZ+aSpJroPVOatbxbnZuZN
aPOLo1+5KczU/GgeBubGercwG1sHQhVrmuVMsqpslKHiIM9vnvMRN2RAlc3nPvoY
vBsznAh1EvHTqACO+hpfn65G67YJV2g4BKwvSA27u+8esKqvUpPFTevXAzbTjTu7
66S2YgphldejD+qYfDlbleoZ/jiP7l/t5LQ7sVriL04SVVmh01HhkCiAJYVkUarw
5R9oT0pAChRHuHhD2nqFMMaJixmMUKygyFo3QRgA91F0yU19W61/n9/AhQ03jLgq
50OfobyIBA+X2W6k5RtmzbMTlAq0iGUxkZR8nagAOGEfzpKtezithkoJv1sdQbK3
9+HE7tfKituXjXZzdUDwexhnzBjGYqH2VTPfBb64u465Rtuvrw6e/QKJ63t594pM
frzxeSxfuzvOGTAaB6WkOgRdvY4Vf9Ppbnc+WDDfl4GMXjw+2Pxq+ocv5dZwPrIq
WE4HjtFm3Um8KYokoZQ0K2NWOAle3Zg+m8L5pMelpCOwDD4oYc8VaBqEZeOSA3bA
Sfe5Or0XJpH0h+6/LfOqpv7yj2Uy63jtBBY5Scmcre8twqYawGylZG6OIigRFSfB
MnkwMV1FbFD3I6OC2X2AgADedfIoCkDV2JPushllBNB0HYEmDbz0rdHMgiRxD3Zc
gb1rSSoo9yy62q29pzqWlwuIQ0g+Vh5eOEUAwN2DZ5vOByj89EDBjOKULnbjqH1S
e4X0LNHwV1MbNiYH5tAXLhIPXbbXw9ifT6zl9q9FdDGyoPB9MS3YopU1FNEdP74C
qrCzUM/9Dx48SGA6DgNyq5USd+uiC48EWguLAwdpYDqjZ8ZGpwnlc4y/0EfU12Bo
NsiZLsTuZ8G94LasbPxA5pDaXxUwl1h7YYYyLmz5nvVKm4U/umnq1QZwe+eqOFv9
tUIAp8QeJ1N6U+0nwUO0XZ4D9qnF3I7UCjaHvb7qbcc3wOLDrMTFPP8HUtyWnYLe
vpdSU/ZIrU/gSvZezcmIGvDwXtZphgJX03ETQxHDjDyfqREeNmgsAP7hDCtrIEhP
qn1ll/Xw8d6rROTW2V9ChZt1GoWPvg2U42V7XxOQ+c1y5kubjyZLM23MyeLku1Bp
bGWgNPndBHDSayB1MyQ2z2rDIBz4rIv/DRerC9Amoe/tsQXbEeWKjoLYTmd2oJBp
wd0x4TaZ9CYHYuF1VyWnxW4VxmghbiVshT4JkOM0ypzgLnVU1yqlK81TWiFIEHYI
bTgkuEttXNkJqEit8dmShuZCyW9PWaKAXGdp2Mayp9lpDPr/c0MPKI6yYqqbyfoe
JgSF1nYFeHcCltzTPqdqiTEi9zriqwpmm1k4TAubArCBsgd539dWvDBMMZWoZzGt
FLVH5fsnRKSqWnXtAQPGLlzOJpSaQRld8uSSQy2YWo8XWysJo8WfmYzWrlblsKJU
4NXB65zwiQ1MGf1r+I9+HEc8OMSm2E53mQViYI+36eYfsMc0BZPZh4D671aRuUVp
fnf0MTfn/hTT1xcTL9VvYCtJAbIoeVgApA/IS7hr44NyvgbEqazCtpW6pLygUqj5
ir818FLHEsAdSWfxJ7GOzXJxLATyVDgRyG/N0K+bpRit0KzW3nid7sgpk0kJtgFb
BDDjVJP4kz3ZKzVptAVN9VEhRjsFHx3aIHsgK2ejy71jrAUHSgnqjVX6mc6V4x97
rMKUx7055dJlQsP300xqIAGa+NPdYgBoHCVFMnaMH/3VMIVdCPhpLxsZtiUCdslC
5eA5S5URUdXimeUPWN8KfHnl6VeR151MydpuKRuP7UW1+nMSDcZZyrd8LWEo/CUR
XlRd2GqiKHLyXZwNmKJhABZGpQC9kyRhxQ8QoTx36EfSLvi9ty+BD+Y0Pb4/GCqt
a/aA4jxUm9PcODj6iWvZpRZLrqfTrbbwgkAoKjkeARn2OgIJ8tmPH2u1l2WOTCjt
kLhfvbYRPAixmVsrDxSZDd65LCUbCzRQQlIEYGbf7M56iRUTe3l1qOiBM6x6n3OR
69yuLxvUTZyBtP+kLvn6n3sPecD9228fLQYttvSMfD89nlKWG/SybzlE6LAOv2Mc
RzmhLvq0DNN5J09x2e9MV4L/BrMFPyarsXWJzJBfPXWQ/e72AGd3izLCceRZkamV
82+YG/wb6eTn+wKuz+/Hoz5jrzGOYt60DPdczLkwfOHdsvjUvI7GYTdQxsmQCQFm
HS4lPZHAqLMQLbLirBycJVIK9dvIqug/YxW4hcMqOi+gHzpnbOlwvIgFW/o73myt
Y25v55UeaQFcseTQr4UOy2Fp8VS5XSFxMh/KUsyhnVWyLBDa47Wo4bvxk4f6Gsde
LFFV4Tdj8ms9HD7g2ll5PieIbyGoRxZMqkeCfjWlAq9ZCUaLycXyq4Em4dusMYW0
ADqDJhYqZ/NhiNJwBzx8HTlnJP13Ws7xkslgGmtvD0Xb8ks2cMmeY8cDcbJRXBBj
mzWlVap+PC+5t499zLpswL+ypkeehi+2k1IKt0M1KUzC7YFD8tTAtMzvw27Bjv6E
6jX40cm3Tnrgn0qYktKPL6ZR0jYyLUWl7GbgEFqvfJPnAcgT+o+AquEayv/GRNhb
RfMgdEy5q0dGVF9LgTUB7zaBhm5l7oLBUAxnPjYeaVFxSKisFsfHSYVz/6rDXvTz
lUqaZ5f4f+/0K+2yrM1ueY+uvJ/H9KUCKVApK3k7oRBXLktEg4AIhIm4GqPNSDdC
+l1F3Q8xOafvNMen0SpMOp9ecAp8VQ+i3tdbD4chcvN1u92HqUiKoELVfQXcDf5V
Fks/gb5IyC9mzolOB1K7wbKrTXeKkuyI6PPdUTnK5HItNfkvQkOcz7W0+Aj4hjBx
+ttP5I9EmLmBZ40w1/Yi4B8aHjGu4ky/eQs7/gstD9bWL4nWaln5mIiHDLFhBfN2
1Vz5JsiLlTbmaIvguNelPXRBJ+su4ZRmWO6YLpoyzFchgzSE70rQ0XHdQQBttlTj
ff2ukWS59vwLnf7hNNg7Ymo1vIWNis7eJyx7sgF3NawR+C0Et6396gtuNK3NPVlf
rnthhCITyXwz1puJIhOQUxWdFBSL2yVbb3MmXsaWSXuQmbiJ5Y7JTNfuRHw7lz8Q
KmpEe1e3MGHQy9AKPUtmWU4X/VkPY05E6Bgn4xCwcvbs71EvZFK56EJwdeXAAPkt
JBk9T6LeL843mMQUc4KN8xk2BzXcX723KOoWPfsfqScnErxOiOzy9sKZ2a+uUnW8
uDdlULUADqJL20OHkNZqTZhpUhiy//6A82oS0sx7defmx5pi8AQs4zPrQNDedKIG
ffuERLix1FuHbMMLcLOy6x3Y3vH2s/1xJ3HuUxeIneD9fpQ9sdeh601cgBSnRxGp
r+ap4odOrshwjZsJimOgx2Io9NVWrCusbKlKpj3mTZJ7l4XAVFwWxOCkW1zqRYag
AC24DGynrtK/GxRVvA56GvJYOB6USrofguwoaMMYm/9LssERnbXnzZKODsCpa0CZ
3LJ4tr45ea6mnhpRF0YyWvmrhTJasEfaiav/AmwJC3kP6yoa6Mnx1TZINiuANLjR
JNtKzOd4NKE+7p89jmVgttl/h4DvG2tWtIGC7B73tBxiP/v63rl1Surp/0Tn3ypZ
dPlrhLXFmrMOlK66h4D668RsZYyQ4Q5I8kxImT3xHTKxkavF64K+3eiavF44PgiQ
pL4x7drGlbVwmVmX36Sh0watg3qv/3xFl6EdIREitZfNTkYf3jA7I53CvsI1ltiT
CixwY06xnk6CvabcG3TvX02Z90pcOxA2B0qWMG12eaFxc5ukVQVErlzkocxXSewZ
hKj9jLMW0pmjLOfEZT5Bq/NA9aGC7AQnPcYHb8awUq+mWKBJVmiiWlKAWHOoLnPV
nU6R5PkuPPHLhPJbziMnGrcTS1WknWxNKDubc9rYWEkU/LfUJrZUYtbB9It8YnMh
DgZacyitdU+lwh77FS+HEIbIil8XnbhLvAzOZuGLbhk53pTriP7Yoioqd2SqL/wo
EgFrrS71MzJcdo8TqnAPN/qlt4o3IU16tdVSN62ZMh2QXNGnGLe/WiOFrtE3aPbV
aoT+STmwIBvm7hWEbZ6e8GBxKNx0/VjflWvbklkbCPqj5dQ0kaziFmpyX1IqcE/A
/X/3NHNThTZ33D4QspmNc8ZDibaoGTDpSQ8YiMv1YM0StgRoqzWCZ5j5f2q5/lKe
Oc9M1RV38NTo9a+R8NzNHu77k+VCSTfkozB8CcnheZPjS0tnqjRsjdbjJCx58jHt
ve07tKDYk+BLCxjt+QYGj7LOlqu2IXp3guV1XBXyJ+DMsv4g4fTHFrnEF6sxXmCN
LqcOzM+WAS9V8L0zrPxfcFcRc/YrOlqM7Igh50h8ChXIMPzVSvcYCGpFC+R12uCM
w0bpfBd97T0DNkAYqNTDgcEJ9tDWghCG3on+t9W6LV1lSOOYkDgBMxjjPSjoIUx+
iVjxSkmQo7JhbhzMVFww8l1E9Y6EVqUXVjyEknI7edAEltrjt/evh1LGJqD1h+sh
a1QoxLhfiuBSMi5TDrI1BYL0u5r2Ahh+Q/qgxQI7d12d6PDJvmFVXl+sAQ4JBBzw
qMbrgtKGPxdugYD7hGzr3GIDN6yfBGBLT2SnJB+BoV8AIsuWYIgAmH1OZodJ2mA/
lVGoe0Pww4Jpqj6aN5PP0mgHm3U1iGFAk55ZxADa7Wcps0gnpfkZ/kv6QDAUx6kJ
EfGWEyXAWgu1oUdmNRyLoVFaWHryMoyTxXIrli7BEpOplRh9JN6/h0QFrYJfzklt
B4sic5wE8fqjixiaNOsJUmFnrL5m/f0tdNgezYm9meZLJ3yLNsFNO+E5GPZl87zP
OsMlN6JEkziwNuy6kpNFbytULEnhjbFTilTpNQYuoY3pqPslL/F5Qh7GNHWW+YMH
RbTUd2gWoc69/9hJw+a+BMyz4VJvGrnyJOJN1wA1ZjTQshaAA8fGhDBnm3BWq4BF
jII85YC+p2yge+HwLsiV4VzEzB5HX+yqFbZYzCCXkYDpd1hqtuW6bpFVjFP1HBb2
MskCNvlerEDLI+MWYvFQDdkkegpYhIAhvXQeXA6w8rknQc7s5fS0rc3qP+DYu/Nb
`pragma protect end_protected
