`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PYQRJsZ16eu4qxjZljJtkYMqkuT/J8bGCGJbnYwNDf+oaQKsbsTrkl2TENwzbdxS
We6FX0eqIXh0lJLHBB3+1Xg4gZ02eSmcPxOjb4gvH2YvNCmjrpI4FW6fmLcgUgBO
MgxKZVGNmUj2o+6kRDaE4IqFeqe4XdkK2amRlG2nXNQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2272)
l4reGW7fKDYewwyGdq8T+eKrGw3iYmnZPt2EkXqYO6PzHl21BzAMYBLdUx1bjQd6
7cOh5Ak3bzqyRc7f3MjFHpycmzMgBOHdpWNp2CRx8uwVe89gAFokeBAebCzDBHiX
hS9L6R1Djn365lIMtm03p1tkt2nD7g1csUKKkYDx7sfdvrNADMt1LHcySg7GBPRC
41Dg2Z/En5MaEkdxuAVftul54A9PrFl9RjHv+CUmFOptbwqNStQIeFVLAXJtBfSb
+PhQu+qxt0levMf7wNhxmMzUoZ080aAmbxIlTz3Dq71Y6qINGapTXfvWTnKOGKy9
hUfx63t5NaHS6R9E3tFc2sBLmHB8lW6kCTAtOOjvoUUPSEG3ac06gqMsfohDo7BB
N4KHs+/1/lam7iN9lS/T3kdEdsGRnGkWP13U1D5bT37gxbYBgSbodXvqZHJmVPCx
6T5wHbZgiarR1v5p29DgA6Ksyxn2OJcNDdMxJLwJGzsgKywGFbmmDi+S9uNWvWp0
rDcTsiYq7wBC43JfivkCzahL1i7C55QBk9TNa5ghOBHFjFskoKyazzpViNCmg4kX
l2l6ax7biQdSF6a5pCErn1m/x05m2VjPZ1r0EZb2G3W4zAkhPQMNgjNgM04zcPaa
Fw8Z/MbAgblqwIi11yRmL4cz/965+BoVQTcQ/W0OVKZrSozXPKWMigFFOCyu14mA
yT0dAL47QWhK2c6MOcz3a8XisIA28WlQKKdX97k0Ov5MqO7tIO8hg1mogoOpdfZ9
eGgc6tiBOieKJwevlAivK0aS2Qr+HhXOLvLv3ruqJ0unRmSyLPhVEOJ5/8F7ub+y
r6ggzEnc+24yz+X8TjT05vUbetrnChb1cVpPVIk83gLz9HAYf1STR8T21Xrdmu6U
Wby1ITjVrlrUuoauScABHY6nsuljTRrVl152MxUBKck8ttL2Qo5QIXbhLQiNmLr+
n5/pP8yAbI9XfAN878O61uSw9fTaPz7lUyqkXCp6sjuHLiWFR8FFImaYSyF4dfkv
f6iRp+KyqZw3gRPigZs+tQThk0/8+QTUwuHgj5MedHlfjEwD7ShB/O57e34Gylos
8oIjiWjBV+jYcuFeNr84SmbVkOT4ZXG24sCPdDyQ6lZ4W43spxQC/OdquaeTfv6+
YpObnSHu+mKy7eFhRfREkBpUJdDmVfHpPsjPUJ8eNVugXQ+rQLlPZ0DcDqH3en3/
xwunISqiNXRLKiOpXtvZsXlCJbX6In3l5mhXY+trYtvCcISuHAuz1AZYSFs2LfTJ
xYdPmfZ0tDyIL2oBixd85oEVvlQuD9IAPKMzMo3rEe1y5DKyf2q9t1qSh8bk/Qu7
5wITnCj7aJN5BEwIkSw962NTwM9lZp5jQCW+H2eV/03eqCKJ95QEeWfqON2brzBV
8QUem0sUACUK4ZzOKamZxB5XCiyNP8a7pE+CGQtksWgsBukFigEwPLArNpsQnzvc
2Ps0c7jAC7meFPivcJQreuNsz2RtQ310VVVDDu2Tn2CcTBpgoxYXXnzU+LM9dbxN
G/rWqTTwK4wMfrY3MqSte1XxF8GB5GKILbmWfKqvJTYQFQIhkRszUyAqXqwRhULD
iclGTVqG3C6IqLqmXajTuIvM2kk6pkRvw/Pzd6zoJpGKqTq1bxNUwy1/7az8nNg2
M7Uke+gh8VVPasorZS5fhwVCf7H/+fdvSgKIWzX76eAXWJTIc1c3yMB/vvWl7nNV
j4u2drvZkhmBKAIs66Wt3bWcXeozgqvwylckOPb1hyRhvQsBgmiHMD8z47LwN70q
fEA9WFqQK8JSnbHtaIaMDHFl+mKiIfFKcvf7xGHLKrxAQIEsqGGNbt7X1H5P0Jhh
7wfBLjcPAwEePLB2CMIGGAZCmm2fKjURlqDV7y2oJRayVoXrrBbPcKr/KhLk6/Un
svomlkCBDrVIT1p4NYsSs0i9AGQh16Stq3EJ1FIEeUTt2PnClflZFnEBRF6AypyC
zY9FIRzbU8zdC8WRCiTNU1jSPbQ0SoYTXDj70tO9xfnho8LWdVfPGCflHvZZUp83
l7ihcs9I0kOLrDzuM6oiPcE5Tc/+4fdodrYtFfmzh9E7KlLRhPG1e5uAEQ6zcJV/
rvR1z9kKUKOneKUGRFqgEAxoHfF2kSVKS9gOf16awtec9lQ6tlGEiaRaNru5L5mH
YleGzSdlxdBjKUAkTRk2WCpGMMx/OZ8uiTN1PZIXIDzSuzz9sUoZt8ZPr3Lx83n1
sIabo2jLhdhFNR7E+8jgbk6GPPohmYQLf4wu9dD/aUI7CUAo8xTKriXXHUmY0zKB
CnWa3zJhgTN+JtC0wl0+uU9Qgg8Pr6i/Jz5j12Gh/UxxqUEXxyGNMk9W1rkHQZL2
t0gAwbAqB7FOE/bTGhyUSp3BR6L2p+GjTbk5sXTThAXTDO8UgKkjKl1w1oi/a3Qy
W69GbCjxcj0+XaQiNAN5igGhYwLQAsVGFJ3JkgsGWCKEX1W02J+W1ITm38gJm0sj
6O2oZijuBMvY0cpsphw1g165O4cga9on2kok2vV+yPLaEBUxv9vGPkk8Nj+eIjpg
RtC7LYLree75i5TVkkBgMI+p16kUPP0ElguV8Hcsj1g50eM9j8xI/pXAYxiBtN9q
k2lR0uP7JZDFfvZL1WV/h/FKuwBa9SKtc4mmOobrFN8gBQJvlaaX+r2emDGm6Z2B
4DGBghIL8hnxH0f0WUxmC4FK2aPGomrG4LZtLkoj7NuwGm6a0myAhHaC2VHpZ4Rn
1X2U5DBpgJu93zXvsbaZ0jIlrbf0Gg5OUYTNnFX9hZe9JcYyscEZBUerjKZICqLa
0l5PmaRjDRfKD4fSyHGt8UwXu0fL61v/G+FGVfCht46nWJpScew0Qfe9nXfr4luA
Ft7dnNAFwDc2Bpp8ePjjUyr0oaYexZbwTwSYd6wj+24Y0kOkeQ7CIn32l0VauRtg
w+jkXWK3CKW7E20TogClVFOsPQoEUXzew1N7yL5MzPqGhb997OgSG07EyQ36ciMo
V/QI/0AlDJPmQ68csYA36A==
`pragma protect end_protected
