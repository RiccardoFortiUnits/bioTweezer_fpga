`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tpfxKd+eHCqW1p7MC9WHkamCDoR3L18Lg+M/81ILWKvddW4X2C3oL5h2Ver6QdcO
SYq8Jd69g4lKXgTqNK8StNy178PmLl9U3Ew7ExjQ9uc5UGwJMlQaPJi7Auq54YFy
fE40VTW0O+ZOpFW1oR5ESBKGyYT137J6Fkr0Eo9N+FM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11040)
0UzZkPl7mpwt12v73Tf0FhjmhJYk9ORXegHvXszx42OtADk2UI4WXpizdUCgg5U2
FHtpVzLZqm14puFaEUr9RE/jJA7blUFAkSxX/QSfaeVgKlqlmelp2lPU1csSm0aO
phtK6EqEuvnwulgyzLe/smTlPGW6FHH7La1F18fq0/bEdE13BucbRTGc7ik/WSEH
U3Ibnt1topSUNMOH1vrshzOL/g5oQBS4nLbQtUGIEpxRbZ7PmQw1Ta55h4ZF9IHY
iv4B5UUyXJd3fuwPVsRTnlo1tIXWTUreYPWpTv0hXYIpcMjshDb60ODJD2eucirs
6S/wDim5U5Mi5umLKwVoF3hJsN162zowjjGyJLHRJ0pjwJNDoLsrwQ5Y7Esbe/fF
jqyfG0pKqdA0+pDLiQX6Ze91gLHipP1Ulaat7+w85T+ng2GPfChGj3nfqyZqBikK
+j9J8JDrYn938PVRUni1plnq1rdQjmvrrXkPJ8fz6Va7NSvdhNEZTkcHzDKZVKA9
T5429Zu92ssykC7rlx1/Ws15DHniSh2dFJ/04WZBeaHmYK6FM85k4KGX7O+QQ8sR
4eBbxswWwX54VA3G9RobRFU2vzH7GeaiY/wOx9Hzuykd7L8XzMlOI94EPOJnZIcI
bdQdIsgg2JRJYmTkkn5lhyo1ZQf7o2WUP+BXE4zRg5df3GCkE/Z4348siibhw6fD
lQ4ybq1jIrzekh9XA/kejuSKwxgxovRke3GefUd9vxEYr6jBcwukCtFgPe0s5ZnU
L4t9ioJmGIo2I0mUJ9d1QzqkaIa9vSmUxIJz/ui7QXqs2jgt43iQCazG+vO3xZym
a4yWwNTusV6bph6B2pT9L6Q6OPVKuLIlM6ofEmipUsG6CShSSgjBaKcaaTJdzxEI
LrLXQ1Ujau4c9GvFRc+iPfeS4GsBO+psW1PTQOG8qp8JtYKb36sAdPRmMakTObhv
9ZbkozTRGnocyN4cJH72eozuZS/xLQiWZQJ6COhHIEdUgGea/TafFPZggWHeAjCM
slNqq8kau68sHVn8j6fPkdIkmY+bpkt6uz2QLMEGzfeZmh0l71U3vwmwVC415cTr
MG1XWYJ+Kuay1U/B+WpdgxX727H2VmH+9sYXHXcYocdyuIxcr3E5J0fdvH2e9/HD
ow+8Jz6i0yFuoOnNOSWEWHL0JVjPKcm1A3X/LmKNKFHJ0/M5g9wYF6CVqusLbPqD
Ik5js5KZJk64CbO5oA2Cyg9MaAuFyrTspC+aSsAMWdCnM8gPF/SqI9zUaK10Ff4M
A1CQ3f4YLg8LAiQ4k4snqMLGNL/nKoQ8mC2wE21bbjRp39HEdJ1z/TloB7+Ottok
XVpturzXzUx2RqneOmkYZQmurRhln+lTs37yz4QepJRT2ciAZM+RoHSexrvrbg66
iCvnTtm7jaFrnfMz/jZ2M2+qaOTAKGkWzEOZiXkez4TfPwlVa2W3P3+uAS8821ak
NkEuXdCpawD+kOUZzN7CgDoopbI3X/K3w97q7lvN4BM7/GKTRRTbKu1gypA6UvdR
IhhZN4TrMZSyY5gVb0/nt8eT7tObgdXo1chQvB1VGCVM502oC8uWFSsa9fCufyi1
mcHtMoNr6pwv7pdkEOExypuA12fYXtzhpP17iFfSmig3xXQ4eBvq9uRLtlHTEVU8
2pMAKMlzXUzzcoQJ+5FCCwiPaKz1t/TrJm00QFmNIKvAmvXsk1bwmbua6IODXNwr
z7ITCUGhPwo/3Uh9CpB8fQQnanNshg8gtfYknaNq6UbmLbgeO6Ed7d6e8sif1+EX
t6agKxkT0x06WIQB0N87pTDjarapBEdZ3TTT3cLDHDh/4hG+PnRI53ASxgk0IiYg
gimXm90gl7caT5YgDHWXUrJlRJX/W0mRzDFQNnJlMivhZn/ftytms7HArTJJuDS1
Q5mYrT8eW5H3yRPS7SZ03E24fdrP9qX9K6RfOUC5RwmtbkLsn8Lirj2SjIhTyEW8
5JO3zLYSAifalSgOjG0BK89ON9NOMBUBzecHX8ayvmSVTyhCNHZlDBPwF5DRnw9L
IMfRDYf4mRaFgPMJuRy3V9aCoko73cwLv4J29RrXRbmOE9xvUY33vm8/5DZRChpt
jUzHq7RZcMn6u8h6MdPE65+Rcuv1d9okLzGYKMqzpy1bug4uprpNJZytQe8CHWIs
aqNdKel2aGNgHPL/baQ8JaZIdV83Q3nfqVpSY2OSVy9mBzizk7DY46dxJCO2x1u/
yYNTDp1Q3mNHvxAREBix9fsf1tfaD+qso/8XIEwo5RvxTIAxbXauAC5pexS7cjrr
ChiVA41pUt+9UEO0vkPNhxLBNXW3AxyzwryQpwMUNjpZGtZ8jI4JM9xPH3H/wGY9
wOfTuysaCr28c0Lasewu3i8ukefkKNhwg2KWIcYrkZZYZS+mxB8z0S30JIpvQLMX
qQc9DZQVv8TjIFEI+gfspFA02hvRgTUexanlJkRdTotCKT+Cl2E2aM1LwxDsdzRT
GsHMg/4p2W/W0e99aZ2kDQ9outuQnhv/YVO/kvLgWrevxXyUZgvi++zgP/zBUtCe
U+X+kC9+vPQdog6ps91iaJdbbLrRHVV0yLneHgT5WxdBfM0AegGNs4CZu48tpJeW
cJe9+xQi/r8jiuC8d8a1hA74yySeGw8Gpz9WYdIhULyP/osrOaucPaB+/AocNvRS
5JZUabciUVIVMvzz1FELl3N+L4/cxd0myR9e59gb+f+twVsrlTY1f/zN8xumkDPk
U8rMTzFou3yA7szrb0/YKJtHGEHkWr8OU7K8QXHCVZlaf/4QFi7LZ35CtlS5T4g9
w5othTNvhv2foM7jtlVKdp3DRqS+1Tn/vQDlzJFub+d82vaizI82Hy47cqsVcDcb
FrfxNTw2gWj7x43yNxJdrOlW6C77JSnCLQO3GJjgPGaR3EBHQhu+Pf6E2UUStl8a
HftldZ8V1MyBNZGR9c1k8rNJcSM9xBiZ0Na4HR+VJbAT7zKq+HwYPJckYJlvrM+M
yJRRu/412BmVh0ABZYNoUgUWzb5oCqASMWFw+dCjOeROv91O88F3YWzCB5vpI3lc
OspqvLdbwkG2ENsh3Z7f3FnQByaq+/tM+gKnfKI2HdUq9h0VSewhLFLxhDsGoHVa
CkAeK8OXQOPvjgn5A6pM+2/yavDSY2k6P1FMDMdm7Ik6Ki8X6hI+D9nFsu7A4c2q
FmBe0TR3Yb3f6m3aDNbdhQyZOC8ewhSOHUacsCCVNfP4f93UjNObu6sWYvbX95eo
N0zhod1owNmUUcY49zst0lXYD8JmQIRqILrfZO6/deZVVlvMQd5f4NR0bswssU2r
fzLyx+esFKvDbxgKzT748uAm66k08wIPu/hWUUY6l1Kst6Cutd05JSYrnLbpBlzZ
bP/j/Oug3SDe9zS/Kw71UOBPXSKvFwdzK4xh8U2UrTeZc1uDn3C62a8/LEXxs+sg
kpF3JjPCUCnH8GSvfXY208ZwtC3Kv65PPLrcG1gq2zcWPhhyARvouE9yQH7XNGLG
+LzX03NTIW8kswAEtMmkR1P0xMzcFUPH23AILfyr+po3TLbZfll46KM4HoVk5D74
X8zeK4lAHy4SakZWqLR6UrHP9HzMn3V0qsKi5BPOcinct4fxxIBsgNUfyOJTdo5D
tGe5391fvDpg7lkCAURe2ejocbUIQJUnaO+372Lt2E+QKWhxl+gLgRc7zPWsBbW4
y0womxdDju5Q+E5CFL1bwb8SZ7oy0hgo6ApkkzCtc9knp5v3Dwl1mxbPkNbBFh1Q
Hi18YJ7CXtWEet8+60C3qrMul7rhY3rHmS7tFkt/yQsFmbjdlSM+FhGsrzNcLK5A
+SB2UFu0RyzyOH0ET+RkyPDZtc1WQM1EEM/Rrf92lCqo0uLS2AcpqRV8ay1w8xxj
vcLHl53ESkm2y4wnDEjHQzSSbOK9/1easx+vC3hk74d7rB5oAljXh5CZIzKca0cY
auXSSuKmvHffYd1SGXWWubDs5PX3KqNbSXKuQP6hJY0IYgIhRc2zCcg22I3wHcR7
rcO1NEit9kv2mKkVuTeklSQaWzYYEuuRFU0Ko4IOOBeWa+3Syc6m1shMT1Wj8C3U
PnJRQIIFDUI0Ao8v6mQgqlBttVggAaYW8qVRjGweBqS3FS9exsCRwfhPyHjAXzKy
1Oho0rciDfFMX1238WJgXXlCsj2hTu7riHn2N/m+JVC+CG6jHfyX1w2GEd3pRRx4
N4JJ+dRVMf43P79pdyxnXyXkxOd/CL4da5iruEkBodiT9E1ZJxN0vrULCiKyo2gX
kZWc4Kr2l9vzzkMBeOygm9KM7Ehat4h8lLNllcyA6jw2zmEn9j/XUr/MNH3bc16L
Yu9HorLWCSYW2ogNnkPfvebr5uCP0sBfS3axWWqG7r2/JEBLaa6EwJaiZ70WGeRi
73GE37uY9EGJep6zYekNbRn9LwA9/v5zlnY1w9vfasa+HZgKaP+AkP6e0Vp3WgeV
lBm50sa6JUSmdLO7IsDUJzHSUAP9TQjTVtAt2Vo8SRjFcqzQj8A6mR039gg14E5i
MgXqzPW6ZjC2u5Do77drLWQjlbZdcry7qwi9bKx9EtoHekbX5+3BYKvtOq670nNF
HQOuPRKeuFGazO6Ypjwcc+K9SGpr/I78IwuPqjl8LT8+4CMz9S5PBNqa3H9Y4WUo
9oFbONnEXDktCGCWFBWRp+SuOET9NBHRzcjvWLbQ8Go23k2DHfBbNuTzjFSfQ/3h
WAMPQi8ngJe6RrvVMMCZJrxRYusrthvv0HAkXnf8ifuhvmTSXtLLrqkT9135C2Bu
X6Eu6CavnOes3Ox4drxHCdLhIXcI8/oiQzn+6lwe9w/P7hy7AIMwRbYJ7Q6mX34e
ZNJNI73j9yzEeGYUYs7DF2WKhsl3Yq2NllFprJYVUegjdbaenh0XWjvAuoH7ZifL
SW3mPIj9MMnI5Qt3Oi216b4R/7jNip/VW00zpVHgI9C5xYtHfRtw9R17Gb7YoAyB
nnYf3WG6Cc3o4/ktZRSxuf/NmTeIFfsF/7vuqsUUDrcpcXg/r8b5oweGTyfE23Y8
Mez7ROjrGYJqvRmFPwtLM/kQtqBCrdDFsycKwXrmkM4406+zfw88z7arHqO78MzI
oVdJaayzJZYUmm5+iHsy091H7shBQQAHYoMCN8my7A3cdA5vuS3UVskYYRDJidIv
TeuoqTrE1EgaR3WLeV2N7CaoJHNiDzttNGyYj2wlmekSywiQPcRjSO2egYMHfLSn
DUDiXWfHH8ZgIGcT4GQ3UcnxraCa316X13Q3dbb9uTX/dr5AfChUmO47rV6jumAO
DolXAp/eRp0Qvwl0Bc+0ODRvChskN5C5gVJoDKBhCCN0XH6GQ7k1CrF4LSEAnrnY
Elc+6tVYZx27Fp0KnHtN1lDLOxmBhyAmdY00KsoWy78KsULYbQXdFkRvHFoXSbqc
gnyEPiR8iQ2fVbSHNVLOcvDpZX6Hs9hpemvVKiZqduZ/1hi/mXyd/qW6Ejh8nqqt
UyoQjnYrvPH/ZWpyDtDVYtDyimbZfU+7beD56bpsz7jhzSmVUaUJ4ABJLB1/0Oki
i8fpBcVu+KAK5Qxb2c244wNX36ZC0f4oYI9Yrcgcrs5PH1UWGi4CSkeloVOcIGoK
6g22N2dGclqIFw0JgvgEz2IM8WKMWIoZDEJiyzyH1TKd+1MDwe0gjxbsy0YJW+fZ
t3T4JB7OBRVHvF2YDL7zo5K2XmKreKT/A0U8lK406Z5plU9Gx13yLhlAMUx4mYpc
NN8thwuMXjnmsUKzzXq3SCne8hE1HZg25yjVVUGnRUtzm82vx9EDIPm076texWaf
qHqGGSDCYeuHKFXOrRtYALRdof7LeaPOhXMFZh+tLh0HaJiwqIuynwJ1De+QjCJk
fu9swBtUQiLL0Ko9ACTxcyydtaBpyKKBiin35YgBgSafS4UV6qp4UQ4O/qUF2AW/
xA30RMC7mnVZSDCbzxTn32PrhuYNhpZ+gsJO6Nt+Dc0MHaEE92MKjPIvfjjY1lVg
SJGnid8ctAj94zfrQoZFjiWxTY1pwfCGghYN4cX1Af3z6gtTVya9ne1wuP2WVe8q
u1Cf4wi5MJZlMogQ4BQLcT12D5qZMzBkgTc4A/9l0hnAkLibS3X8lfitmxfOH0VL
0Y6B1BVgA6Ewxeze+QqQ6HQmg6tJB8pTDaeZBYgsgIhgsyy+sxl2skqyWaLayKm6
SZFk4kOzWkuLSG0gEkS7c2Zvoy9SJhprjY1MJUSxtOR2Xo7yV6Bkohs44wBTwOxP
owAzfuMfmTUsiQ3FBrA+SAdWm1yMiApLkGtgwY+ZDnjWFG/9eI/uF6PuzRo3yIIS
Zu15S+HjkQZb4bM3sfgr7l3HgKfmFmzbecP+d20YoMspQu8Ccc0JwznJ+WJb36de
1lWVl1MLNMe9CztoV+rb0200cC2Bs6J5FBuV+8SG693OB2fC9vLGt8YsmNa4TKs3
H7UjhXg1cbyGanjqu2RX291CWe2RuclljuRkf2TWcVMYh4IeT9AxaJu36SbkPScP
NwyoUToR4KK0JDvc3etonWJHbB/qRmUrfjbb8WPIFltSgI1N8Djqs+4kU9+PmRVn
pZNIWKDR1qq5R7n9YlxXJILg2VV9LyaeVahf2Pp3QqFRMLHqNUn70D6aZfho38pR
ancEkJ8U4GnCv9qgsRTdQXqrRjP8mu+a7DmldIVTc+V3EtSZN+sfVU0lUc0jQ22k
r+0FfDlm4hYjS56MOBoKwOesZPjuBFLLnyv1NX4bMQbQuDn0vpA61n5AsW2IDlT5
0EVcs9K6O4DuuOO/pqoJB4jQJODe+fbZ37okMVzaG9yJM68Z3WkIjgx5sqfCURCr
U5U5DUkCS8WGkSYxMQzBX+ltFn7ULkQHQ+v5F1upL9ZhR09Q0kmfal+VYcipQ/tJ
QiXrdM6xK4/x7OD7SXod2/vmUg9HV279/2NDgQao0HFQWvziPiFk2SVC9AgglDp+
+9bX7syE7r3JZo+l/i7CRLFBPLWONsDzzEE3PY39rIkPwHkaLf3DCwIxrfKNeedH
57pLZDy4HTZw1oFNaCd9UQXFW6eJS8GHCQLGfRMXvlEpDURxCTeLW7RivOx0a/wT
PmYM5SwokOi5Bdz1utc/ZW+1ke1On164B8WDXD5zYypY3kQLUDAjyZud288JDmDS
jNQsiE+P+NStU1oDbovGdElRqfUDfZQiiGjIzwTrvDRB6N0WENsuFKZtgiXm0sZ5
iToUi5Ajue62Z3HkmZvFRhOOi+mxOWXt/r+0IhJh1sRP//KpJA0k+MRktth7lQV9
BKS3jwmsdLCRXDgH5YhBAYO1nlMQeFtb18sNJTAaw5MTNrHTfEF5x4Emx6fcEHST
28/quUnzs5UYQ1Kq69FpuG3GvE4FNCq3d/e5b2dDLcsrNllHgS6CoyIva+KAqX5x
c55NNLtjbkmvPZu3aTfCxNhoQvjQbyuncM3vFG/sS8E9RD0ei1mwLaRsX6xdTwiO
u1t7igNF3+0JSX3izvl8JUA3QQUBFfExGELlyv91jFWPpRPL1PvniVI3tLNxlWCG
oW+ZEsYZYUpP/ojWA8EDP3uwpwX+2QbzllVT8Ub9ETT5k8OcKla002M+N37k58H0
nv8ZvIiPk3gt+6qnpn0WiU0nAffvPwNdEnpdDNgkD32+/A1fA0QhZPzZc+fMIlul
0FTh7X6/hRAUs74br/Z43+S3jfC/N3yDKaTHMMwHxxL9B5Wsu9mcvKx+OvXPBMIn
VlGvC+ov0Nh5tPwWEBs3iaqgVUbgOCF3Hdi4J3U67IUUEk9NgAK15MChCNFak9wg
t1u53Tl2uAP93+Pc1vvTmmWKOs+r1h0NFslYgIz/r6Ru+QU4BXcF1eCluM1J+ts9
7/XvfwEa5fFIwTlQkC0USdo7zTXqQqOmv4XtJq6Mm1NZraUjcraEDk/VDHQiFVd6
Hqtbzs6/CtQXpn76AZF1U9ZGRbC7hW61wz7btMpJ/Rdg98owDo+/fOWD9SJsSd5l
KUCLBrLuSEJ+oXKee90AiCpDwEb3STC3f6GtQ/MylW2+z5/0B+WeMljChb85rDOv
bH3fc4VvLdYKxBfEst8U1BAHze8oIDqpP9GiLmXnFEmcYDk2Jg2Tivqd97ai7rYk
Jxbid3Y3eAvyKuvalMGXa2Mi1NfXlyLg4PsuBZ0ut+IM6535qNSGOfQWrtWqAkce
kSXzc6FX5FEfpBAL10gCovKOke2anwk8XhhwEqDyMbJCIBhNw0O9EfrdduZlA6Vm
VtuO/MC4W03P/gfI2tlHvU4cLejT4rH4v54s1QlgrSvpLdbeWmOFCJAMeWHrX5ll
LKIaPtA275eW4pp+cyu78vq/URgG+M4lgq+nHn6RoZQx+Oy9R/RrJ0KrUnQn76NV
sLehRaA9TMxbRmIDPtiMUuxa7/Rb5RwKxQFb1XKhX5FhEFvgvW/WUpezxn22e2+7
1e99EqqBhSSSC7GrIv3ki2ShRIPNfohYm+9cyxIzwGwjUqU3e4R23arYgwGdGpyx
yakjKJlsV40kolLno2Aex7DHnvMBjS5ua9OGNmKcCRTrg78npkcf6aHHQqi7pUsK
StVgVB6reO8ye2W+D6NCzbz0wqTry4ARN8lykX12XhJgAnRGS0JAxBokAqZsh1j7
C5TyDNVyLXbGpC8z9zKPKyuB3alZYoxyBAX2tH/mk9baylQdzLwxgKmPGl7WkamA
f1fAztJAyjmFHMiUD/BUiAe9Afugn/fnTJcyhA92JnaA+FncMvWLNB736RXBn1mf
Yna2MB3xYkoPVX1oaXI2PxgDc/QNOXalql7pBw8dzlxVl6cSZ3LYcpRU9oVi/cWP
5wFWpneCVBlniKFLv3ged5wXG/SSw4piw7vGo4OL4roskgS0GDKw521R6izEAc5V
Ntx4M0ZA/xZqqjPZ67WKwNZXKVF9JF/kdKuU2N2/YjFJfIIzGW21pC1EopXlRW08
hkTi79VytCwXD9cdper8ss74OrJCq9BirU0YWXTtO0W5vk10eeh2IXxzPLjdh+kW
JB7EsVM/4sN4BGBeRT2U9FfKAmhNa21hVCON/0ttdPtBrAgVHc0oBFWdBVsgcMtp
qWrdBRMXSvi9VUZ2S3a62Bgpe8paUSOENQT1CRgOJC5qk0dYHDLBbXFIc+Cx03yx
brMxDd0yNCSphQStE3+TLPQlZpQ4SV06CinEbTMGNAs/xIo0TlUDotdUcoIVsAiN
R71PFpF7GDoVpNmgN+G3g3p8/o5K4AA2NIUedyCsLeXV+oLACgZWDLh8lZgZoZn1
5zMxUD4GR5zEK9MS0aI+OgVZlfcT5Uhc+/YefoY5X4qtnSCr60octjPohTF4wJHt
r/68n1rQhiLezF/aZ1rZdxhrh23lO7PByqlVTB7vxwY/yD98khNIOvR3HOlPFgY7
/mdJSdCkO6+O6ke+KYLJf/aHhYw2gYrRtJRCTkwptqf1TrJo7xnAB+vqKDRrAgvz
mEGlDndHyrrmDTSb8ypihaPoRPGHM1mbn7pQbnbA76R0CRkSLSpX6//J0I+SYcci
XQ5/gV/X/Tq8PU+ItX4cElFZfiOxGkYvQqX1IhDA9btEtpdGYTN1RrKZosj8KZiD
kTX6wsVSWkQN8s+2NWnmXGD7uG7FaxDVX+u0K3w9OGw/LNEkMqTw6YsgwwutvRtV
P+4ZzAd9/xaxPh5XSoYQDMJQnEeFLbCGrDb4SK9kIHMYpUmy97bDK4Z5rdDgwl/Q
QvvJZo/upT1NVu3ymyy3ZiTYtIyFbc0CzteFj4zKxi0BYc/i2J0EpvC2Oc/mMICZ
lgBUf1A8RhonjyXKkKzJ5UiN7vshpv6iLJF3C454w1ONhtmevj4uw1In/PYxtx8v
s9r+SkIeavhDJiTclJ90GDECDeuQJfEw6r6XFIVdtgA9GyO4uIlm6hPmYNX4tuDu
AhD3UnIWEwvpXt6MB9ZKk7MAuCcj+7VeXukpTpl8crNNF81el/FOtX6+BhPWf4nh
RgM5/RGBGoboSTgSmFGfEYxU/eshaNTm9CcjUZurWvIV8qmFiDh4IRx1CLtm7Ysy
erSlhUsqMkwXf/lIYjjc9QTg7HAZkWB3GJOqPacL3r5qtlMi0om2Y+vPh8JDwzlz
CyPB+GZ574X3FEpskfhXu85zHYG4Mulj3VLzpWNvdoP0at3JfE29da2nH+vZ9tnA
OXMG0t3xzTXz9EyLZyBK+q+1pdahZ4jrfBGZqIvLXHQo84eOoJWto1KhAkU1QrMn
XwT5+s8H3IEKDyoXw4Xnqo5zayaG2vCPX/fcLgMyccXgtedAXXYfguvzxIezrxwQ
g6jJWCnOvgaIfctZM9C7F3wmkBDIpabkrQAb8j4uqjPcpxClG0HipX4YuNLd5qt0
EB9Dtg/rfHgu6u+0ZxiT2hqDNwoy3u63bbwFo31bRcA6wo3oBxvLtb+oxmZL/3Tc
iYmONoabe2iJ1nBoGi1XddDpheWBx3eAWfn29Z0PjQYbS2PPCU5t3n1VL/CJr9ZS
e02x+358cchPRZWYg2JTkZuST4P47tVZ46vuY4k5+LSZEUH6YXOYkoUuEzgBrCrF
n0h4vxbDCcdJsMP8f+ny2uDR4IKbn7t8nU4ov36bb2w1uy65eaJFxNgvz2B/WOi1
+drMF06wXP8ZRUuNieKg61eGL+/J/s6ntIGYZ0nsMqqpGtmxWjliZ6W1ETFtEPoV
NaW8NELhLaEy5Ajr/KXHUfB7IdQ5zRmjrmHYxDKBxr57JolcA2ms08KSnAByT8PP
ovZQEqqfXJwQxXr0LFAHoMC0HX2TrblswL8ERPCEcwtx6E+LYwM1X6+Hee+ryD8B
BOvd8Gm8DpH/zAPOx7jisJodB32OO0JEevMMGm60V6AJ4IWYNSyA5UHeuPdbUgHv
aKfii//vSbWNPYT7GdSUWbFU6KCVIxfPnNdw+0Wr5LWhlr7n7cl4M5KYjInqcIYj
6saLFK/Np6CJXvxjkmM9y4NpSlRnqo6zilk0rUzLqWmX7AR5rJ9M96fHneQbCwL1
66+N72BMVJRWqAHTdwbus3C3r+m2XhjLpCmAZSKAbqRZ1h9IK40rd2nyucDtLVmG
BTkYI0eZn26DQCQsWXNU8L4a1ypR1AZHAC6EYzI5to1nxyqHZqM3EL6Zvsp+QmUs
NhpWxJdtadpcfuJpINsPszmRuByHH4v20z1MqnKUZDAWcaEfVeZX4Fggb21N86uc
rR/h7u8ArCmg9pnxjafgNiW1Lbp8bk8sYLij/v9YvmR7+Ymeh8sQ1FQvCz9Fim2w
swCWRa6t6c+Ig2eBj0wxo9ixHsmcRhN0zukHdx6KnYB7neQlbbR3nYoNUVBTVPSH
UN0skato7v1ziMwAfYB/NJxCzGG90EUfzIGP4WbPas2hOuudauxOfwTjO56dkjv+
bS5qDOJDvizlUU/DUzj9CRPSwgBzimnZI/oMMcxTomPlpsonDRlRl2sz7GoUSh7O
cf110xRpLoAhg469dK58gbBPHvbDSTv0BQ/GkfE8IFpNsaz3v129rJ34wfT0afAc
0VAi6PCPQDThpP1DcPfiDeyEcYYI+ng3Lsg++78utFPch+Qgiqd47pYQzZ9zqlYZ
LS7RAWxh3KRwPkM/PV7eGGjBcbGBERX4xg+F776mqpZHMm3tHmiG8DBLj8Vv6kHB
UKot0X36+KzntyARz9j5tEr2hETrjm/LMXi8LAlBSeYGIYZINqgkdn7mHv01HCNJ
nAhaXnCDmhFuSkDmEGU8oi4vx9gZLQTx8H+H5orEoomaV+scHyDdPeU31f6gB4mf
EuRaT2hzP39+XwzYz/pPiI1FZ4QNtp41UBQK68YyAmwxGI0AHJcU8o+jpa13xByd
ENp9hRHOILC3PTq20jEMU9vbFG7aK/f2pAQMpvnYEgPzLxn8ynXpwBWwart2xV/I
VxU60wqEhGXSHVvjVKJdotXWMj0iR/LPkosbYuba1zM7xI2pUPtQagZ5jSTN4twx
0acl5n5sXpYlKAPbbZIlqJHRtWeMBQv231MLopwElFi52sUu9Df5JvtGba87YYmm
OO8uc7W/7EaHsODY0kfaNCvKkTJE5UGvwpQpncghMaLYVLPxFETFWEzDqkrOwwtM
HY8Btew+kG2R6rFeTAxov/a77pFKYhVDb7hGiT60nsXKVd80O5SpaB0bw7zrPbH9
UIWuwwD4X0CDs6kX5E8xFUkfmGgKFtvS9g8N00RFTvpTbZplG84zdg4iDL7aG+6p
k5H03uOVlQY0aXO7l5LfYfMwpZ42jPKOcyGKuNkWr7Z/W1GvwembPFvN1teHRudO
QEmRIN2ai7GBNZXvmnHd1Pue+aDsu6Pv3foqxfuYgnkX6BemAqSdi+ZUQt/uV1sO
8+tX59NShKStmiJ1O3aE23dj1Bh6IL7TdIoR1psFybZe1Hy3UoxLXsaSj/rV0TDg
4Fe2jaPB41CFHh0mgZS/TJzAE76OpQRAo/08rzJMMb7P6ocIIoMPZtLVJHN+5u2q
dod8Ne1+lp8V7dvjFZ15y94OKN+8JNoVJIAqoPCDCQ736GN9P52rttjFoHSuuqlC
A2K7YFmQovshb/feD01aYBpHW/+D8T1YbCtTvkLwfcae6E/x2x0FcIVgBcgcEmAg
LqYB5htJ6pOJkAzQT5v1n5+6dKp6Z2/ducpxDcgmMt/5Ht7uyQg3pht1WbS574tf
q/iNS7t5h3HWyXxFMGLUQ2Sy8IOzwgIywj8wvBrZS8lHJUm9iupkaH7JbSOWzEr1
PBWchYWQiR8CggsFrdoaibfObBXOXDifMlpTyy9x1kv7c8BHTFz/o0ROK4Jt8sfv
O/nyFi+sxJCwhMgj7MU3fGDTH+O3mR7EZ8FKYwe0vvTo0eBnvG1zOxiIwabDHyxW
oa9OL38aS1R3SfbY9uF255ziEPHNqwt9B/09MYtcG9rE+pnk1G5ar7FY1prpWPiO
XrKaVZ0uxOBslHTP0iZ5gNNS3YV77q7OGZuytTBU55ysuQWKgIGuGCkAFzU62qnd
3/P36Orep0qYbWSooU6Sp+Fofq57732q1eUgE2rfIpUxC1jGNfjGzcPDIBWb9/ZB
mWsWh8ksZpeIchDuWGj6FNJ4nBweItZmuf8HQj7apYsthqLihAq19ZPmWkRccw+a
Ix/yGdZjLSppU9CJyYZ0D+iojDLdQ/O+P3Bgt0Xy8d7efVriOkeKTjNnPYoxPsMP
IJjqBZiNyxQa/upem3p4mFngliz8sdzGiOp72lVcWAKHNjT51INttgNt6AZ7yIN+
6Fid33Jq8x3dOkfrUOCUYjM/V1mfIzxrFhwwERKSoCPEV0gOftGN02VSpVP+UfYD
XaHBRNaXUqGpMBNSWD6iOxQCFpSxmnjykKL4TNKTuwGoABazHPZ/MirV8309Dr5i
NMDGx2S7p0db7+cA3zg7Ksz0dbLvuitE4/TXyZcOAA/UU4Jpvc0UqdAL/G4vQ+AR
nJlNso587UD5mPG7hoE07M4ERZtSD+KMQf594NqsQUjSBfotKtvXMOXRC4NGpmRU
d7iojd575rAOQedyF9lxWwMMZDvL0cEOn3s71f0dYLdRyqtjIjxvCA5bhQPAo2eU
s1WzTKS47zsCBqLwXtWMQEGDm9UQLArTidiyzALdmsLDQX3Lj2fKsUgnW93QZK5s
TtuZt9+GsTcApArRsrnIXZbJsM3sRErS71UxJzY5P0Cfu+hx9Trz6h/efl3tkf4g
B3Wtl7OYQjjvVtIs/PQCurcIKev18GRy3M4wCU0+VFnA8tlgAInOlaBgA0T02W8Z
998B/bAFEpgjcmdBFVpj3G+uz54UGA4QSsX7iOKXOY0BDMEXgTAT6GQnHbYiIyLq
yP1k3CuQo9T+5GVEKckf7htbfNOOvJZNkl0vDMdoggBMjRzz3L5tTNVcpZNC/vNs
j6R17N8moM7EYVNK/EWGcE8XRhUhZwFwMvmJapdbV41MOzX0+3AybaSAMJ1zryLA
4zDlPS2uqBtaguEsNK+Gn01Mn11+riIXD+urNX9qqk55TUcqvqPjAJyaLOyafb/y
28LG/Tl5GpdpDt2TwqyfUvCUWUwOKR9RpRsBhPbgqZ5FtNjKGUaoNlQxZawe0o3Q
OJFnedi6+di4UE5blcUq/c8CFnFjbNfb/Q9ddrirwdsvitcPjh/Pzy6fXvCvxggF
Q5huIVYjxI4YLvC+ZZycS0wa3UY62a/5F5U8BktUPG04RTpNz+VaAaeomKYBQwG1
G/kfxRSd28B1t//gVgQ8lUnPkOTK9HvkHkF8NLudxMkT9MqycxuhVt8Fax909nJ1
zImVOHvKNRr0aZQXt71qTInz4WW6wa3LrrQpl0BFhpwqhITvWPJogvPLnDw/syT4
LEnf4xD/dVnw8r5vLefYrinExxIajW5NVVE41oAmvoY//zoNjNf2MLMiNaTNcPrs
W5ZyEn9lGYU3vEwMBEalP6oSgSX9bpCKPSLqenVniLq0wc9QAmUyn/iPmLjDi4QD
Jt6cI6bhpemifvqHXReJFL/0hwGiCccUCj6e/xP/POsTplhsgWGWR4V5B+RhoMU7
1anfB3alGJDplXzXG8Ki7RGx1OtLHghJMl9iIDoc+H4bgoF8hzEsHkegVBStBJZw
/sdCarE5YtsWvgpXjsn6ZYM4n87X6B3YVtoj8sWM2/p2IIQ9ENszLQdjm4xEwRA1
KWIsedI4CqtAmKev454ZNEWf89296KIadxyLlEQwcGY1h57tDN1T0qwzSRydhfGB
`pragma protect end_protected
