`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dCU9fmXFsqtQEwoQ7h4OZF8iP2/dX6YAJKeKCgNcw6Y5m6Z9+0xQ+GNxL3YxNKwW
6XmrljsbfhvgTYfkCkwrwTp7aQHl1d5wxgKEHHLMkpQJXHfR5527OfZgqpzktCe4
dEGPtxd++cqgg19umC8HRxej7tJ7SKJ65neS91zk4co=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176768)
kF29/nHugsxgxfKE+gIPPHXI7TlNrY7c24+YKM3fPwsvSgZ0WZL+kDnoysZP3s5h
C3SqE0QKLw45x3c1M2GeF9TBYclKjg8pAXu5UxsPcRWqV/NKDp4Am2TkyE3d5Ts6
fxUZ+997SvxCJSL1PVCmgkSrt5S8tbIAxkNcTRTSp34vyUPrmNCRH6WgY+17UnQS
ozf59m6jTe3JxEcIhWGvoTIkmHYVHPNql4hoRLhCV5w1Qh9gGjn4K7awv4SiTRzt
nmrajxUCLIHhmGHYy9BS6UEzkdv+tpf+gM7NQQhiHado7v+SoBBd9RNOE/rFasEV
MZJ6Yczxt/lFSK/9owsZ/aEfZTaEMpC/EZGLfL1BTRggBgzbB1xgtcbXboI74nMC
R9BJzEG2SHp4i98aya5GOS7lRfueQseIyBSNsjHuvKMar+KssRqxcFKmtHF+4ctd
GOjW1JKF27sgR9SXq0qH/q99w48T2xKVEKx+FtCJgfMRwNk2uo/Wvrz7QyIkJEK2
lc0lCG7Hu4jT3m4JIEHaDzNIwEaVjL2fqx7113j7Cxivkl0rRXI+fv8t3sC/eu77
p3KxA3DCkn+HOvzTBFm9jYBFiBXcNMLgeeDI+PUW1BbnswfRvn012VXon67RoKRj
cqvBaMA6aStrhi6zrXlFFwKbPHYZoaXT82QmpBsxph//Zq0stdVHbNNLYQf75lHH
upFrQqlZdEzIJf6lZ/V4HY9lPErKH9GK+QYhaw78jPRG9zN8ttsCNwzL9k+uUjk7
o+qo/cByvO4hDgCEFmsgL7o+/1mLXdrJBWqnAOtNMYqdi1u/qFjLN5KLbyq8xhIb
aerf3cvD7CVpBGigGGZbn/5Ed+8t3g6U18F8P1VnkE+UqaJTUhuT6I2ELLdt49Ji
lajGiiC7Ld8gNr0INEUZpSYmX4YxZZKFO4m0PIDyPTqFsJnVpjdO4c5YMQ4xi+yu
3aRfLKd6fpqiSoIWkPuknRu4qZCU6IUVrv9+WSlI4xnp0MY0B2Rl9k6STP2qX82d
j7cUu5eL8SkAcaIKCAGQxDFV7rnTXUhCU47lWZ6+S0QqUnXJPwkf/oWv/1IM7nKR
QWHURfuGZTV5HWjuj9HA/9Sm96diHEj2H3iQxV1SzzbTG8Oh56z7cDuorez+B3Jh
fao6irMTRbthtey6a0tVUB3CRnA4s61Te4G1M7LiudSp/Iu4HxdAj+/u6pHLgeAL
4cHIVuzRl4n1EwRPa0070pREnQ+xYbjfvCbl9uYOVOOVdX2ky1/ArS2KYh3MqyKj
LnMhKlELwGWddSb4xRoF2EtjfKL44FXKAhV/BP6cabhk0zjqAnMEKH70mqBzB4mf
GUu2v3kc7t2N9sfpGZtiHXnjOi+TKNf8DQRrWxkVDM4D0K4H9WJ/urlfh2FcMUVF
0r5wZsHv5W9OwzvwjGTBOtC6I/eg5WwPK64PJS4SjnXAFU68LyNU+j5GqdZU5EqC
XQ+U6Erma6+RaPkkzrSvkBNl2sZcRG4oH2ZAg+MjdiJaerrz6ynpdO8ewJ/jJ/61
qwOwjTfbDLE1qtj85Q8n31IkLKUsZ0J5hbBAAlKoUCD8ZMinIxiFJDIrPCoA1uq5
OD4b42DCp93gr2iJPaJv9Xob8jBmoUSKGCKrar/HIz0sQ9EluhFvLg5lmimSZDGh
AhPkmGS5kY/Du4sGXtYmvSjJE4AMjU0qejxPuBI8YaOUaJ7jlozXAfLl1Nv9ZK2u
33VuxgmBizVufYjWlUwO+Vk6cVff1dXFrZtyoyWu5X7VQuApTBXwfpj3VPFwb61v
V7U9T++oWLYwwvrsK1hcDqg9/jl4lXAdgDOotclHLaauA0oaiRW2xswjCgfh9sMU
xnq4VNSNDTdSo4dcNQbfCbRTL7H7CzkH01pm6B+AkMwjJCXJRcXpg2ZtUcY1l8kT
rXS4dtyNv6DGuym3Xc2aWpNlSHfpzbVprroc6joUq0awpVpKXzf/lO7wA3uDlxly
peBNNQ3hqm57hNVZRAhaBvIKy7neqGzm/bn+Iw1R8XMMqkF7JbTSLp3Q7lMOBr/8
hEn4I+CkT8Zd/QedYYRhGNCkmn7lMfzW2w0lo08qgWDkOEA7rB/krNqaajPeDC7i
bPYMb+FXRDyQ0hov2mChtmjOx68nJ//nC76ot7e4TqmNdShhpWj+FO1h7o4Hw446
IyoKZZrTTTgUk2ly6IejxH3ED6zcUxQxY8291SeQsw+FLZ+PHSSaEeAgvbHcM5ZO
ue0p4TQPeCDr2VyFuqRCE3I5f9IWphBX19tZ8CP1iVMRoEM/IQUt4auDaa7kGEg+
FR+7HkS8X0b1QRgF1xs0CNh/iPY6um5KnCNlCherJlhxeErrJ7a8UOd/8cQOLd8D
kI/R1dIWc/9jq/kTKBT9Vq9DHj+KRBg+UR9ZtnFtvgUT4M0szKYAbfznIsCiZFYL
XBngtBBGLhO7LZewsJWh+4DIbwwUxBgBEfLYaZ+4OwDbzxi2YcVT79BdWWibEA3c
71sn/Lq6aWLdAmwHTYGANJfAkZjxuTCZLdku0l+K24PlYZsnMeaiSbLLAhW7S7B3
OHfBCRu2j+LIG7YKXix2ASJxEjJ4OzKI2zk70npyUO0hEpaWVg0ZDH4n22Vm1Ljv
cuV1DV6sSJq3LTTv/kLpqHHodCfV64HHSh/VJR9w//BPsw1KDIWjy9r6eRa9dVYT
xp9rt7V5olc3bzzEPdfuq7/dlEGraRqPNZ7ILQfOiV3PUsdYi4ZpIUcmCucQ0rHv
lxYWLKfgBmzl9/ijXjRZXcQKKxWD9TnMeaBaz9+vsk+7jvipvitSDtd9NHw+iu2M
W6m57wXx6NXRpP1nJuZn/1OzMQGW6/wvifU8PYMmz6KyXVJgKLHEXh9h0UiFXb+q
w0/XpKZBLZ7bZ/Df9GHucO1Rxhm+GLmCeqLdmNkcxx72buR05mPqbxEAq6vfi47L
7KOGW9ETmHTqzIII8ZIR5M4z2FYIgtIOgpNz/zSxjiAZ5ItTANETDYhsQOPo7JnP
hizDcDXYib5nw4crn/HgUpz77TprmUBJlCfJCNMpj8PKNR4q5VjX4mGAQH5a0gXU
1mdCz30SWC31KgIIvYFic9zYkbqUEgHJd69hnUUrobFBytiSqx51abWC9HQlMRlu
+v0mO/a6IjCg9KZz/vBC2UicRqLsqXy/vf+EbFahBrSbGDPhBKrOXpru1jr2DpzC
UUorkzGujZfyWkBJ8Le9RJn0fBGxrRkNBVd5/gDF/0dldQfiMekRJxGCAJuO6/Qm
hhrWuDOuvM8liEfU+tg3pbcyeBR/9IpZ/23xTe5TH56VyNMr1g6B8XRnqb0kwr5y
Ltfr+uYoDNsXpMVh1XmwMW5gNGnnuPwoD5aZa7nBHSNILvM/dLL4+oqV2T4iEo2u
OkIQtJ+3+77YPHKKcgt1nhsilXYi5oJ0twh7c++o64FxpXaYkj2wFYQCSxZ+eFu+
R4rP3rENYaq/GBBU/hYCU4/KniTAUYm+L6M2VT9YJ18Wh5Bq0N68qQaTK1nXwYX5
fTfy8Ur3+Ma9q5zI/wZpW9aZj2lyFA6hYuHPn7gQL7yIR0Y1mjinXmxi3UD3UAMH
i6B2vxqbg0A9gREdKP0OmDr8u1bcJR29gPtjf+Qi/Cdu/KFR+8ZJk0/kQCu3mOKV
Ua3MBy0sW3wih9fZU2ItN2dYqGNf695RIsEfTSwQpcNM3zfWWteYRvzhrnXKfYv2
0dVKud4s119CgKfjCiLgCq0uZ1katoVl5Fa44LMMWN2CaMfgmWFipm3LN/om+oMs
zdUFDRjfb0IuSzQ4mXX5siBMJNoncvav4Drr1F/BRhCGKk69Qbm+dqFnQlqk9fXV
A/HPShXh9cQN9ZzKTeGjHZUbDt0Hr+dlHq/erUa6EsfY6A6ew5czPHqXOWKLt+lJ
KgMuxKUDmEDEIeL4riPJ+aeA0hGWvOU9qcGs+Abwb0JIQJhZbuPQCqTvm2TmlUSi
knaJaQHBKkvn7Vs/UYeXNE3UevVuv3d0M1YI0WOLphcE+ztcpmOw9UWYsMXyNlVy
YOexEqtItKRjnLoBwZeLsSswij/vp3+wWI/al5dyM39wUvbY8+Wn7m77cl25MOgg
jzlVzMMP5lPkUwKFkdNxfX4lNROYZGETzawIC0AQvVTFFkzZzyq82myhU3N2pDy8
SnUxfI8TT2dEvIKc+eViqs0ZcuGzjMJ6vO289QZAkSSPIJNTviskc5CfoQwqPeke
Po3S+ljU9XBrZ5v4iE40cwDoHFJHUa6ZWhbQ4oRgmbaTUx2xR7R1129fuDEXp5MU
gYicyMsvt3yzTY9zoHne2JiWF1/GxRpxhfv0joden4J3wSy3hYMNrrvjxqsPQqZ1
1Ub+0jxjYbe5Z0gIzNedPMlIutRW2PAjDKMGdzU70LP0ZZfZ333v4t5u2RtkY9tM
R6icmVxauGqsJUD+mws0dtQ3QBYsf1r2MRXOVrlRNBCRd1+DDT1JT78ZAu5q8s5e
eYybzOFL/Mi0uxvycN9jBfWd0q5nN6XaL692fJi2IPvyPipBa45p8VYL+ITTWS8s
jjN/8iJRATJA+VdzQadxZfLgnLYAzzTyPPO9txWthhA3bBi7bcappRoRfrsvk2SJ
ypZjj4op2LzVjL0a7G7BFmbRlJPflQAdS+1kVP5EUx0nOnrQ7WP9/72tMvRKQl0u
lLe2ER3I9inCRqlEEVjJ2h6aJ1tZvjlqeHUVnPdCjfznMa/8I8C1eU6uFzepx1KW
mSVC9CjnSDFi/ieEJXAxsp9y2eJd8PTslTQdgY6gCKdYvK/djG3w/fzY3Jp+cS5t
3rN+0HygN2k4rcO4E3qFG+vy5NQTFI67bC/Iy2aLq49L7NvagrGfeALAcFQ/XKBC
7dVrzpjomU7k3wsOczImtOEKQfaxJVr0zHm3huD3Gnw6D7U75P7Ns2laSQFVzuvt
kgUNJwJj+wPvmuA6nIFWXZJt9flE9PUaXeuNhsZYk/cU2Y75N2uEx0XiHRVq5IM+
LRaarGXB/hj5X37LcR78d5Vj3WiPylft+gZsgw5N0E8m6TRjcrLh8QmTo2dBwcKY
gghGEr4q1yi/4NSllTHvfpQJaeWHa84H+i5HZae0TrSb1+SvM6vjbbw9dNsBv5+0
HQ7ueatpgT0FeaxizXa0Dr1k8GguKlkkx3s2XvRuTi85jzzh9fgeSRyOtsQ4P0ZM
ru8Y3NJGcGF9rNzo0+46JIVPrzRggnLX7yVV5Rd8mUZjvSe0a3+eoDdRJrFR0MY9
0GvRBld4M+qwWG4u8CrDZnuUrLDVCH4PFdL9TPM5c8Maal64UZyvC5U5rARHBMYE
6gebwQisBf/pMt3G5Nt+EpSEkdzTyeNShnvH3xO3OJp3dx9oy1pfH0gEZR26kme5
4r53MJSoMy/lnt89h7SjDCO7/7aFMDLpQgOjlkzgRXoxjVLew3R/Y33QgdzvHfMz
vwAUkqbFOicglHyYGVnxeaBDWvKN3ScRz+w4NPOpgDZ6uLjHBO9HzVNdhO39ej69
e62XfYjPTZk62RaN04JNzhlpU4y2Y4tl7+Fg1ClzcDZ7CWnHKsiIHj497xIb+jsA
X1TspITj+p4/CcMn7luJDR5eMS9cR1G/wFuez6WPeq20fxN1ipvbO2neJwobAm0t
MxJU1/PfEKlYuX52R4GCti1eU9wLCamto2L3twno/XHEpzIMqa3s9ALvqEF9Vbyg
aYPnVeyuT9shArdHCVXjZuQGnln8JQyT7TI1UPq43Q8OooqW5x0BWwOUXIf/u797
O2Ql+Q+8ckt+olifOs7cmZ+bs14Qm7ReNNiICXGPsOP8Dr8e+kjihkqs0UHbmeKG
KdAYmkTZTdj8Rn6kKdSe54cN2VLAjFNF+1BPTINJVqbLXqEtt476r0D8Su2rSFda
TNhJ8wwIgGGUfwJSLtbBk5kJGL8s0HdX+Ean9nAg4FVqaxuDi0U9ip2JDe+lIrxH
HowoGzsJmvZNvDxxqRYBYq6yMTeXgqjudk5OxI85mTZHxY/OgpK5DRfZss1vNbb3
S/AindMRD8Brp7pWEglC4maadMiugYqZtbD97WkWF6wENyNchOwKit7tyqHY6pBU
UTuHYy4dT8+Z9vqg05DBTdneEH35ers6GfS3ddkTZGpoqQ4GCBW/afQx+D1hZsl+
Dx+/3Sb/uiqe8s6W8CA78Rxc9sijsJRLYB+h3Egjr8PFcfkV+dFujNE5pisACX5E
HtzbP72btxhxyruarSeAZgmCoOLU50gHx6jJxwvjKb3amHf8u/zXxsCtT54+YL5h
FyTj47O/Bc0MonwK+t62zxkOjmEzgCkiWG+zsLDIT2sO2+QVPXxGzkMnVT5BQJL9
EMkaLn1VzzmLOgVCshvhLD0I0HsB4HEIF0moLAVjf2YvuRv39ojkGAwubP5w7/vg
BVAeb5FyW/9atAMIDi+RYyZXm/IVBgyeiOprCHRSBF1MXrkEm5EDw/9KLgsSDQ5a
+UTRIdXVgVp2vP056bcz/kpBfrfiKNhfnavXeoFCHV1ZwMvy7RKgQcFGx2hck0m4
NoKChAsuEyvwHhY0fTyqX/m+Jm6z3cJwpAHqdC3feVT3+9FuKQ9BSgyflwzUxG/U
ix4B/oddFQKlX1uSelx1oXWQ7xSkw4deCrOUwvOKBqeWOFb/n2Vc8LONS8FN1Z3H
xzuoyKdlm39FmD/xIBhdP4Ol/ZXjM21VNdbDZPqMvgignZn1NF2ncWTjEp6ApQ5Z
PBcikv/0b7rfMet2V02C+INYIq2ehPY1rjvW47c0Jp+T/vOmleoWN84OPNhsRy3Z
4/vAPbqoznS3Ax1kCWwXWUz/ErmCUCERzI7EH28AJBrjeXc1YN6fiZAH/mBw8/2C
O0BJuwpQio6Xoz04Xc3ID6aqcrDfTBVo0MgdiK6FTMrfF87igs1pn4Sy9hqbtKUB
tBcbH0mT7MndblFohZYKvOXN1bE+Fki2mypj93uBqAdA6z/uz7hAOXoALYRk4ORv
OgcNfb1nr37y7cCT8gF69I/fYFlvqHeFXQtQOnNtj9/p5ddVh+RBxK6UB04o0bhh
EtLiVeebK9Ns4ALfD2B6wKRmHOpnJ79oS23lNH+s/gsPcBxHeC/aeNSMvjGg9y+a
NcqRvdXkzYi6MzSNkgTdJoXIxZQrHWFEGgoi9XIbw/E6qpb+D0COMsmkLgo6Snsv
ieY2GGA5Cz5CFwqS7dKfvl12daL0PUJ6H0t9gegbSxPbXM9c1+qCCKQucV70/6OG
cFvlSo7i05c2MdfJJNQne0ePFZmtyQK3gGE4plgz+lZKUR0SZfFtYCGxwUr/E0NF
BV7/F4U+8GYhebKtTTqiTAnnUg0/RjRo0bNsOdHXCpzi/bQE2Jz9YqVIf3y9QO6i
gJhRhjWqNq6k70k7rV5lT5VLVFjTM/0pdt/JRTOdkBzSJMsWIyjngquV0IhIzxh9
wGqjZk0+G62p070ZcDudqKnf4d1eJjRMSnvBsT47rVIAdXG+2fplRyHodAcOi/HP
q73vFwh0N5tWyaCSeFEiRLleoEeq8XeNPMfx0jydhyitjlEv+itdf9Pv4tTVs1sY
HnNjIJqkeST8TLAgobX1VR75T+QB54P9zmFbCPr04i0xr9KXu5sBxA5QHpqnPBQy
nkhg2QIAsrncoK83BHnpWcDt8YxzFEQj1d8uieK+fTtONvzUxs4wQfo9V6nZrFK0
3Fmi793xqL3db5C27caw/5MAUGrU6oWUe+8ab6GLAVlZVlEoNPXAvniXeu16KBcj
DZJns1ztzTHp5ZpjnA2MU/MWV/FOTGKCoPvB+g+f7yYR1Pm3MlAtG73yKwDemIuw
rrDh8AbfNOmglp5t52OCtJLa/WbJoUjPsWTgWhcIxfibF8fBQpFGDyzwUUTSb3oK
V/HEgbEtLx/n9jflcMmW9qM94X3KGsuDxC92cU7fADekySQqsAjCutWh7UY7fQGb
rX/90oy2mScbFJuqS2UW4mMDonQmT8rqKEpm9K89oRd4shabOg6ezrM/vPAYrdpz
7RryDF6fO+4swsbcJxsiKGBH2h94ShwaPsTqPWw8yIkEcFVBsfk0STrAiGOyhKky
4Pgubqrt0nE9ss3bG4KUmwT5/J0pksRRb/SnXv5aFsXS1wt1BtDh5TUN+u2VhjNI
IgftOf0+qdj8qXT/lSQWVM5tBO67ly5PCB6nmDVPHFx637iO4z9SF7DWX3XJ2s3I
/dmF/KAqFjNd6xqtuceDHlpMB+10sX9EkyTYCrhVmg4RIu13XD/uYvUBzklcfOkS
WWUEeZVF/q8Z39nCnCx0+aGeqM5qWPirFMLVuDV8jdDyX6TyO8NYQfsFwvZ7GXSb
FT19/SDKSBAO8r9/NXkWY+6137jJhUs0BX13wO1K7MnlqW7xsFS4Epn8XBHwLiId
TmRGThzuO84LqJleiflRLulFB2NQFnPJjc9A8YxBoMoWuWxtaxpaxG3VSIrpdKSS
Gv0x3odtS6wmCmlnFg80gAnhUxehVe5GiwTOyjqu2/cdsD2MRJYNHQUfTz8MK0MY
42312nYT8o/5Ly27zxdHumnVZBN8rOOM2hhdKrXjeB2Ygqktze2v+pfBQXwovlv4
sEu/OPoca3yjHnfWA20NQJ/LotnItydmBCsxQCz+uhMv28GpQyuVY04yK4Vl+4Cf
oKvI/2PJ0dplv51k3MkZeY2NLqVlsmMr9mH79zttGXIW3mTbcCbWZ6BpNA7k9XzX
D/SI0PJ/ui5rNNZTaJmpnmNlvDT8Nl0FWx9eRoRTreEXajmEj2MLl4WlEoezQCjX
XIfp2nsXbPL4qrC31kRI7zJHCz0UdfxEN6MAMg3PG+1UsIY2hEsD/anqT/96xTB9
CfW/Ji/g3YwvnrsyfF/0yomU0nFXT89sB5zwflCi/bDu1DjEurqin5JBbEAR3ksR
gxWg2obzk70wf0uTXtBcK+lUtfdiT/So0659RaiTlcTpu7VMsZa+F+jYfzs4o+YQ
DUKxM9c3/qEANpnObeQ/RzVJN6GvQ9D4iphSbfo25+riLYZk8AnRWlyTlr3KZdsq
3kp0grKl9e70DEQWwc1ue+TdU4GtzIniajHHY1H+sXCw/VjyM4ZOK58UL3RuV5Z/
jfdXeZs9feSfoEU0gwTXwflGh8odoRcRf7DA/TW4sJtjIzJPynVoU9xiUIGN3qU2
QGKW21AqR0YDF/eJwn94/jN8MIbQlh80AnVtG9smdaBP4ZKqFfUf9NcWhQa6luBr
tktoZFJzZjafdLk4L9MmQkpsqIJQQ2qLxmE0oTXVXZIMjjCfN2AKg+XovLdK0lfa
a8P0wWZzcZT2qEpsoyWOxdb6KhMXbkrJGX/N2EIN2eCmOXR7sqw76ahdOrkCysfq
aN5NE8PkpjLIXUtQmL/zKWRDtnICn740I8HiUTl8GFbvrXXm6yfRfZviirgX9Ft5
jDfVknKA1R8RZDugK36TgfnPP5tPtKkezqoaB5F4n5/od+lv8VqOo2fl8RD+kMNy
874kI6h5zaez+mFBIMktMPcfUNJm6feyozR6vnbbINbFK9kaLs2fDRwVlscCOdbl
gj6iakU9xv+rhLW7IAjUFzZjeeKu2or0gQ7p/2veJFf/NkkHNVUgxRRvDY+E1kgj
MAXJ+SzK0BjqW0LSIs75pwHw8lBCLL3lwhVOtJdLCAMXnbTsobFLygWAz7uKdrce
lOOj1EWJuVqsIq01w2yLU6vJXpiGtWVexTtr9eS7YdvwasMw/rEQy7KjR2ZcGF4N
DgXEifJ9SsmSkxztzIcZoXupphKcJ6uQcCKmSNJj02tMbruPoyTtyf9d3eFY5x0r
DpZP0DSePgt4dABZMfJC4W/3b7tXk8YFwm3Ug3/RLXFyLS3MvOusY/tJ7BmlO5XQ
U9/7rFA7k0qByVtLSWMw4Mr/XTEVVZrs1Bl5vekI6IOL4rF0xE0G5sqKpHg6zBcO
t1U+Gkqb8/LhODB5Gy7K3edfrdONNr34k09IKRE8iynA4EbanG9nCM8i1w+Nvol1
UnZuG8PtMngoAdBS22vTOl1nP/eWvDmOENxeI4alGHmHFnff5MEPx2u3o4hzM/de
vI1tXCaj+sZj5FDNoh9scfBp1iOhI5JJ5Sd6cd0a4fpteXvaVbZnvndZ2UCBDyJE
K7a5dlTa169U/ncUsDjxFGrImk211EhmrrCO5p3UruUzyoD8TdplIUVG/WCWc63t
t5FKU4kN07rt0+SxfAEx24fwyQC+hX4Bk0hJUo2sk9izfXmh2vh6qMj2VZW4oTOI
zscGM8nzvxskUIpXYeLX5wpjS+tWJ6ZhCeFsj2zQ2VnRMzRWdUQlhF08jHctvMQB
KVAIOIKowa996af1t7Ggzew+XDCCgKOlwk03PDKqOZ/v6BVHVywY6JVFcW4TIdVy
4wcn78F8iz6UoXIlYeZKcFvb+3UogkdqjVMb1usikb/pAc3fUQhguXQ8IUgF1ZaO
K7d7s9KBhX7cKGfEhbsztJuq+NAusbIvX0XaJBkQGnfOxoBYTFWhuBe8TLKPto5G
lUIZ5QZb4Vc62Ksa9gPKe8vcnqZyHkhylZfmEm7aJleyB1smAummU1Xtdag0OVFB
pN00wEZ8LhZOYInE595jGLGkPAuEfBcQm8hTFjHULaPsTDF138gb/1NoGE6JQ+9v
opio9mYThzDJmfRXzDH5Z+3j7acNqATG6cRBkLvAw/j4Nje4BlZmqWFKiADWp2+j
CMRKu2BVuTczWAz+wWSqkmL0NOfBEmFe9HMtty8M7gdj2YaYV4bmBTJANKbqQTIv
zoU8XxHqqy+/d26BtkdMbngRt+UPPERn55rPF/atXJMIQ6OWQuI7V2lCp8p6khxn
ble4NAiMGozZAxqaEBV6bQSv+Cfs9MVIp/Z/7uA4z3Me7HPwrZ8NAZ+UUzbiYYKF
FgCZ3JYHep6mhvP8esewBNAI/ekoJfBQmfFN7EylzCxVyDRiTC1LqNem1pdi76nV
aO5GrIZ8Ye/ruyb7odwvDKaUQ85L67R1g95GiLZPrB5pGE81dKCj6V7LXDT+gGn6
ZZYECPLLPLuZfFt2YEVIeGHBvJrq0q1DJzukZKed5v41qnD/eFb5NCiGpIAMdcwM
KJRmcv5Q2Qbwa9wq8pl2LEKknwnunV7zCvctvdFiX28Q547Hb1jIBR7s3IiPTcPE
8ogQ0z/w3iqTcewVyQzQ6Fo28Lyt0xQyuE/FHomaPw5SmV9Ye2lV+5brsD2WdvhA
vg2o1gadvDpeDyAbZwABtW5EWMl76wL/JhAWVmwaTmLcHLBtMqO8n4v+Lzr2bW3W
nD7RH5Tx6KmSel13kvZkia6Jii5kbin91GIt5JKZAknRFzwMPc7jS/BSYaztTgee
ihsLy7o39XmUh3A8IhOUuaf8gCNpQoIfsnTOjR+1Ou3CGn48yosCgSD1hJcdckx4
pejEIKHUksNylcxzaGqCzUvER8P2NhAJ/5FSHHtTFsxCEpkV3x16uDtq6sFT46fW
O2nSHAhL9ueyCQjWycS5nykwKm3jftBP2PmHjjtJbrl4XxczKBF6JkvguT8TFq3U
rYZKutwlrJ1LOPv/nrcBVfA02zrKlHP6KfpMJAguZaXX+HavxToPTWHtdLs9CLM2
yv1DtgYPZmMoeH3fYcsKaJ2AXh4suTtHVzZfMezZj91cP5Mh8ChQZiiXKubeBFeT
K1OL7DWvyHJxX/Hkia7HPqVgq9X4nSnB+PO82VEHr1fs7XIuik2p/L7r4UuEm+zA
kwKDDLfY3s3W3aTKNGi4yMaGZOBlRRVyl4ClYCXcA6MnHklMa+qSp9m/4z26TcU0
1uX0i7sg42ajWG0nvPIl0D9GNBoxC11gN4w/MDLbjviohAkFEE4U5nH2o/w9C4SJ
hk32FGkooGGVgM+EujgzMg0ADIx5D4Mo4qzj84MmQT48eQ95ywMyTy/+SJcsGC6g
do5uSUk1JEaL/ShdwuDfBjRmcYv/V0FX/nfDHI+qUawc1N4nlXGysctC3b3QEoPS
0c0RAqYWe1OkttaLReFXrjGW/G5gL+BQRe/HuSdcS6NjN4Yvv6h/yHIVaWKlkBcO
WKraNhYxkF32zPlSnz09ULxHhagmphnU7xKxgLJ3H7fxlU7XtcgDEFvNa05VD5Z+
mtzFG/6Aq9VgWQSCYtMhj0Lp0Q9d/EWb/rxoHppGeIODkGYfKDPHien/mTIS85ff
PzCHsLbsT16RZqNTLVS3EQcJpTajgaFN15x0qXUqbmIjkMw+VWrBqnA2XPtNQcmV
rHBS2dWbUe7f+X6ZsqpydKpmaq+mlR8iW8IK0klSdgLFI4lCE1sfHT66pWFE/ij9
ykbfvlMLOsyyae+PtbhbohElHYFyz3bI5ZWO/qQtEKja7LF/KXp7WFrPPn0cgloT
pRmlN+kratRqiGDIrUIXBhWK+7wAOdRuCiSuS/3Z0LqiKxQwQobbtG2c790TwOLJ
CeAvmAEYl0E6+F0DNkIB8yWDVsLhCoPsQr+Sv38wReT4ai9Tzc0X6TFqnjCsJmGH
6uBlcMmOXf+KuowP+Dkyh2xtn+rnLZzmwX8LLRN1YycL300B+Nw9yZrnwJDGIPDP
nhWqL9iBRJTlQpZfGssvWofd8R5B73Xhp5QG/hlwUPtQ0ohUcJL34svZNYfwGoLP
YoVhDNFijjXt/ImYX7RUVbuBI6yHigMRTHFYLygTamI5ui/Z68aZpv3DQbIwoXoJ
kht/ai+tFUnKCajKjF0GYou4w0e7x5sQkYwh0FQisAl2RsqCYo1h/WfMRnEgzGHf
5qz99dKSG45gO5kyXZ8Pd7RAIcdMRUhdUlYHeJsHwqi/C4c4PlyKCaMiCaDPudyz
yGVND1PKa1LcHhbPs8lub5SRzoQI0xNskfl72zkbtuNNJeGs6toO7auqplpMmWmK
0Mk6rj0oE2ejiF6ziHSrK37UBof6M6enWA4IpAwN2Kn05fYxM/YK1JLrylq62GVk
Soilw4c2Kvocfw8S2R/iftJEwjIoToLVfdvoWHJCLlrbc7iTr5F+VI2cd6npUcl9
CJkcfd8mOIXqCSzHh3sLXioX8jjRZCqVQL38jBDRNpvmvR2msaPSvQB2V9wRHyHc
GBee8aKyZM6Z0Gj/COdQDl8oL5I/3+r6t9CtAZTfiS2qd5TH35HVd3APYhwhNNUo
i2yej/62F726CQlvJ7I8UF3b8NFcmxODpnXX/MPlmy8dykoe1ahjCyeAEv45JRi7
nxEEAauqCLxvt20zSiHjb9i/ovPkIPeqJWTz8hJeybvt4o4Yib8RxngTUH7Mhbz3
bJpUMYv/LYuYmvl0+uS9oYYRzqaczr9hsx4wkdDr0ZnJH1o+0qmtD3nPHSo6gpe3
opH81KPOvhYLS/nOCVyJBmfaBKgDrZUVtIuTotl4IFrwDbE+iNQyXS+meYlvlq0/
AkUuMd3tHaqrmhTJe44hCjWAtfOUX+mjCAEDiOUxVsTF5G9RPzCjRd+j+OPdirH4
e4TNz83NU5tOJaiWTcm9e6FNKs/0fWVujOMOjq4vhXgfhr3zuroiQG6Ia2OKi1Ey
TNMijJBqR+9Tty9UCbc6qPHFOkfs9szjk8nk4PM0bNgywS+Kjxr+M6GN5u5Ih6Il
J85syiJ+KMMYxdImxALzy7FPE5DX3pOMDjs5mHMz9oLPpR9x8ElWOMZ4W+6ERqD7
Y9VA5qfCrHtT72rwGoDfjbJ/Mv+e9KVAkaLiS+hQeKLaY4MP1Ay7Ct2cZ6sBezif
wsDs9f3M2wKq2b76C5BwQ0XBHMPkDgVeQ8S3RY+MDdau/0pyRUT1UqGPCx1lk+vB
fi+TecB8hVwpTYusqXfAJRGXsdwCXrGEBBsEEEfcwyO39mQCmNidYrx/HSQXetZC
l2/kJR3ogtTErRbNp+UU6SYweFuqeB7wYCWflmS2NwdNyRySDgvM+A9GUEppAPnQ
p0CYXmz5qDoxvWnknF/rjg2GqLaXl2wtEt00pzCodNERBCtXSoBtxllFiUZyIsem
uhDYiUCEkcpLeN+zS8WoTrMlYSr7WGROIQ6VlhoYdEeDY924/UT51OBpEAK2fwq5
0Orp6cyf2mUK0CUhU3uY5FXdlZ6rqz526oHjJm60COslCw/jmWGZ/i1xgCBqn8bD
Y4Ko31DOeNsXHv2lkbQSNAKPNe6PXtmN8ms/slIU2DpxvLBZn1kdSJ51CrDpAIHb
wcfxWZlvhHokJKjYa49FUTXUq5iZkIBpQZqfryrQ8wsuiy5gXYJkT5o4ywdupOcq
31wpYnaujjg6q5grSQI/jgC+p3eNyAsWdpx+ofJn263KLMWwTaz1sg9u1TIVA8qn
mdrPn3m/lzJ/FM2H9uhQmoBu8TFkwqoTMnH7KA93z3n1XNwmgF7ljnkHPaqOcMP9
1G4KOVTbM/+8KZ9Us0K3LhqRotUZKoBYMHZyYiRntE0a55qT4y1kjcmyTBEt20xQ
9PIAzWp3Ee3ZPZD4p4xfl903yz3jXJxx2R2K8V8rRqQ4UmXsS6+7R3VDo0KGEVoD
IbE7s7YN+Oys+1RWZ0CkKIpxpJ7tbfDCqUeXeXXczHx1MXDnT2yYZlIDCf+EH/gO
5Cx4V9hztsMShv1TDi4PSMjWGa/CHZStjwqBa9EdTBwRhMKMsXLRuU1QmALzYc9W
bpn/Ok/kBDid7cQJnWjQA+7uq3r0D0b1UGAC0ZdgACGXON0YcG3VvIuMPKm34P4b
AMDgoie2b8xn1NOXRPRQxpAHQn2syhpxMYO+cRP7KHC4sh1nI+MgeE/1qoqPGx9H
PwW4b/9m2tneOmTw5pymIzlivPiXhWml2ASmWXKcowMWLZrSwi94+OA+tPDwwOIM
MKwfP0qTLyNEQPW7JODZ2GYnjPcOYxN3sjlpGAL3PInn7RfUeNGzxZW6crQ2BpiA
yedj7YJMhLc+oCHfa9f/1tOJwFewedoewCfiH2xPPREOcPbmQjoHqqDVE/lPVpoa
2eQNJlrXplBWpGSY83xJsgJr1bb7tg/E71/UCk+3jQKfMiE1wucPxtR3dOlZSHWs
DSXn66YfUyCOwLZlTtzCJzRyhOiGyaCw1pGyYMsRZz+jzyPZ6ME30ERcx6/YIm8y
BOvM7kxI2KbXxuT8Zh2/ud28fUV91MrX7V7AvglDp0G43L9JQ5oScDOpI9yhQEA7
fFtYXvrLRKkU4F6PkIEhk6zpZY4RY7NEJbclRuPH9rpjsj83nLkxjlHd5JrVWmaq
iALsnhWpdJuXz4SYxUSQ8Ghskv5GjRtULKiESVu6SgbPmxwWzOsxZnV4NBJ4r8+R
N3A14l7phMlR9997Xjf7SZFvSSpecXukPwNz/P8sEOmGzsO4Klm35zOVWC57v6bo
mlMXZbt/5gRmtAEFR/WMQP4i9YaE/UGUG8MSrSBsq4TPPbKSuIgdN5DClvA2xM3m
z1sGaHk9/i2gREnXKXDnoVWlcDqYB6OUumvlDLwJHMc/tTiPICaf+hzbdtlNJNo1
rulQivXPBgR7aZ3IM3fqk2CJCkP+iCuIKevj2SYBbi76Whj6kV0LnsOncl8e4C0G
G4OenQ8AjTlGVzNr0mGhjQTPIy6kKPZe1fXHsGkuyi7N9hClUFN6W01qlQH8vfH6
U2dewfYBe69RKXshcN/mVeh2QFaA7B4I64DZpNVtB6axD853HfNMljE84Uapht0V
b79nbCQkPtLDoHHkzlIPeG+1r0w1xlJE/Ej35yD0dnRk5vnP/K4UQ3TkM742wMdQ
7hMYtcR9iciDPMcr1gAhonaHdhGphF8VTCiRdU2HwCb/fchGdJXEw1y8bLNXBqhg
F8VmQ6WZ8Op+ePXsFFebCnFNspdn/YDFaMSGT+d6ZyDAjLMoI+oennQfpPj1gw23
GSOPZH8wGjWmxa7ap+BHPM3mbF4OYWIUHDXk+Rpkf03HY9nppsCSZQQr3RyEsvbp
cy4BcUygWii0eCfwV16TRwiSZwbsitjnCLXXQhh417+qJzZD2V2dhbO1yk+NOxKL
M7QeLQWw91pT7BOtJgfshXnjGvbfweN9OMpwex9kOSdbqfDJLGytXVaNEb2BDLjg
SKm36Gw9hbcX/uHR3dnxMyltVIRBtq4cnKNPx1SgQlHQxi1jVApNcjrQ34xfL053
rRV/2VzxD5aq4PLGanTzD1ysUZu/aCGfrY6X1MavBTYrDcG2m8GtYbI/smg7Anrh
pJSOzCupe3xXvV34VcMJzcLdsdNeglkx/Wou4QkGlRQygJHnmGkaTHeFq5VvT/jt
C5C9yJTyo1vSxNDjZea3DqWVXr1avW095twdOYal0v6afy5dA9MvRa0dVF7Cnc2p
zzGbT85AxFjeojqPsO+jDkcbwD3YUClkk6/uBD38ZvLgOv4RQlTXYvcJo6H4C86j
WShOcWZigqHaN/cpcIqQFv90L4C/R+1kzu2yKTLs0j1PGUEaEciqgGHQxnc6gRsR
2yw3NtgFMvDzF32nYvIk14q1MTTlnbRZRluJnGebZiJg8ikJuSDv3Cjiyq0J2Jjq
IPRr0AW2YfWp8RPetw2QzF3VW+oYx92TzxQ0kpORrn8w8JX+AR+O5EODrO2igKrv
BNwSS1B5aVwfoI83kPDUnBTQFHRXabYAbM9QXZ5uNqOULVZrQZDi3uj5FpBltkxm
YifgYg7jlObzgrRDP/nqFTJCt/6AZdZrPFaXTNjhoGlXtBazyZSDNAEX6jL1NFG2
EI4QkDlZnjt6gSsenOhnrWR+M1NFBYQly6fo43B40fBIYvrHazuvRUjKGcnrZTqG
/orq9//oIfJAB5+QEQi990kZrmsovDQ5KTzHSOikvWvy8h2sVMR1zx0/aD1uquv5
NVdc9M1HcbIhqGCtGffWAa/Rnfb68dDvPVVC+lYiF8OqKkR3gcTQeNggwXAtsTb/
s3l45wFiTp0rhmp9QeHVeA4IFsrqIq7XnP2RaI7aRJcVcxCT9ixW/wYCs3S/jrf2
JpFOcz6StEnRBL+yFHalgKDhVHOwPi1Qf3Sjx+9Wq1OMyfN0PYAv4zjITqBtu9ER
cTWOshnlSgY+2C+CS34BqTNfmx7SLZiOJuuIGSOGUrVGdlRGog7JMGz5WviUHyjw
xaEq7alGTykHEPLMIQH30EjKPEvJiudD3z4fsTDjGMrhSuX+L7CwApFHQHqzMhlf
pxtYY/fek2kZk/6VZiG55pg68QrS8HZn8OUBzD6htSDYY/PZSP6rt4F55UXjSvMs
9yHhwRp8eutq3uV22+xjyNGtv1xpHqzf2KoGD1Pfv0h21md9fwF8HFNdVOF2u+xc
78/Kjs9s+S19Zk5jLbe4I5qcQJRWK8lvqRVDp4qFjXuq77ZaUM1e6J1JtF4BtvAy
3xvQLoYm/gTE1Ccs51YGKNVikIjB/Hjwn20D24VVUq33FWCqjdPwZJfewcUdd1bo
WzELf4gX0SZp7ULyP7c6WbK+ajEnUDVFWof122/Bh+Ch+GRujrv+mAOxRGrPTlmI
UZ9fxuPHpq7/tIPt678mrqIqUb1SE6NC65rjEPq5zoTRhcjR5cqHvT6oSi1yfux0
lqxVjmSq/liIA0u7L/tIeB3rGv4ilTvL1Z0hwjNBb+lCSBNxxFu+IqCLBL4XjaGY
hKu+YBCYYqmXeNR71WBuJ8tDOWr8LlCz+HmeLRdimJUIIboE4DcEDXk894KudgnZ
UUl6FDYfBBYaaFWKADW/oqi6HE85dM2pF55KV637HenOY852i1gjZzSTToK91M0T
6vES1b5cpP6VlCxn6GLZmb3CHvbUCqkBk7ASwZ+je+LIYHgrlKgC98nL+lzg2Fx5
TGnLQbD+Pk8BYuSVcPzXPqlKU1gD5JzgHG8iTySpZ3EZ9aq7zHsbA/ZF2qvwq/sP
XbLEyfNmttlI4qe87zvY+AoPyPIM1RlveX1CIyjtxWgTvzFrf5aNHb3lW2qLl/bO
R4Dems4fa2vQbhf9pfJNz89Ur63YssP72a+9u/nqTAt3A0PQDttaNkFupQkxTkkF
fxm2vI79DOU6Facr1rjDgK5UFVcm5k1mon6L1Gqkm/ijmxSOHU5XBubZsb2L1y+P
u+HmGqEI63NwqjuhDfG5MG40KTL8D+J9fzHe4/hxZthTPPsmZGrtzlEZ+bVlI4mX
RdW7cVAJ1fD5YigMEda1z/jv6f5BpBdRh81mMP3W3J5xXgbX6euNpWi4zUxl/VXX
dsXzSdgo7sUDB7f4sBV1aBM91IN9HBE7O9Dm/l1U2Hy0MY8K/gOOtxYJY2KlZefI
rspZMkDb0dTREESW2+EFfT6l8QQctl9Cj0biUUOkSKCXXXCbI6nce25LCsId90x+
MlZ+J8XiZolnlBVxrMaRGbRTNGXJH0DB3BMeOcbto7vlQc6TYcvNjNr49EYzavl1
mMps9PMlYhLDYuUU9yDLIzq/QbJAM8YUZ0Fz1zXJwALLixINlkZ1/fdX/Qs+TrD1
XZTGZO5oXxqCWPNhx3fipEJJX23og0KVZlOXikcjBSjVfIV/KWAU4l9OoEcr/UwO
LiA3Q9LylmtRDyuHU57gd+fUBrgAi9a1pAWfuG2hnp0/eIrR8ZZ8Yz5EbObkfhqc
MPzqdZwPEv9NzGL3Z4UpxRQDo4y8We2ADq2qcK7shtLBi/65lvhLesWciitnJg1I
W82AscSUXAQhWRrziy2mhRr0RYQORCAPpD5x84UnrZPqE5emTWLAgP6RaSdqxxkG
A3mG03fNRpSlw8CQTAY867g2SQP7Rk4PIlEN1uRs2aFa7uBGfJtWnzUsj4jDiZor
gF15pfdEGlTtiU43b9ploMEb1EIQ/mmbZtPkLYUD0vLZH/+M8cYzvRc8b795L/dB
k+3oyk89RUMQIiszFmlDEQWSFWs8GAHyZWgUUOaOg0bJyPsSua2aYQov1Lwh3N1e
YdbNC6hU0xyKmoJC06hKzfr97TDgYfsyYyWmXkcVhXKkXSDwcZP1ywVaLgq4Bx0+
tdXJpdLfyUa7IasjBfcW9Qv+oL2PsbslMfDWMqqVz8l1htw4nzjLZDdWcUUAHRY5
MJ6Bd5JlTHD4rXG5SwJaZ7QWaylkJxhIhMBob49AwO7WBWHLc1KFkl95lC/2GE6m
LvQUp0OvY5qd7CKfyfCwzuDkWCY1ZcRgeTxluDQaesaZzoykGWi5p2e8cu2yACym
nqzS2fdD+PD5tXA4apao6cKfRaoVB3zlZQYW9EzEwBjCLde5qDqmKRWUE7/do8mO
TvIGaqonadpo/hqb6rYzQoBlVQDvp39rrgme6oYZogcXuiqgmtFAb4/cmoe4W2Bw
mrdwJi8fXLMypxA+zAAmMrb8UbIyuvUdirqjngYQN61bGVtKzlPKzk476yUImy1r
kDz7XfpeeaYaHojtPOaDnW0qDzZVxcVAP1SFZx9oJQPI3BCbzsTDsOTOFPMuyv1V
rNnX4eewBb9rjeQ0V9fmcZlM+A8wzjQ1T+U3DGhqJ+di6t+ZiNL4491bjWSTK7jr
4Bxy3oWfNDRG5KtyYbyu+qH9OqGdnDvRcjgZovyDtSjQwtC0x1jS/tmDTwXswkZl
JUVtsozsJAHGAXg1Ct7sCIlGGeDq1QuKmHXNnSLuNto9OYJVCMzJb19BH+cLmMCC
TLoUjnmdaPSDUA55BzA7Df/FBO1u1wjAsQf7C4ZSNsvKaMkLrhBcAjEk7+bntHyB
AP/MOZk31Tw9i7ImoQi5iqHp6fvkvPKN9nvmOotlz7TMgnUxsv49yOIXOHm5byyw
48lcAWXezAO+Ppq8sKqIcnEnGVmA6Ii3xulONeGXEQtNsd8cXfUtUHjnb4j3Dldw
C39A9LYEu4dFRnCi+qXumbqQeGijeJaohBY7X3HRbDOxNlaUiXKgaYvAH4PwxnYh
K/V4emsf4QppkXJ5coOpHMmqSOxFTAs8eZ+XZXBkqhaiYAF7SDfVutKQEp89P7rw
Wo9IDefigRU/T6SkOTWZh2Ey7lLPv2cVjIRy6CXosHsIRxh9FXF+lYPURa5wecx6
NzTyEk3k2KmKW1eu4FF/GXWSaGYi1PLpuxmy216ivqjptOCNmKzw1eqRPxlT+LpA
KI+qhydMlF4Pp7T+rNRk58LM4iDj+II4Nk2zATb1LC7EIz5cKOgEBbCtSFBUf/lp
dx5OkdBDbQLL0aWm3cF2VWQweXpJSSVn4SdNGzgTxz2k/bTBDEOThcoMMJ13fWEO
J+E6+YwLCEoemQqQWM769wKes/ueCRKy/GjzWnVaG2BkM34SoQQt1WqACSmKC+uO
rMgsNhYLPyydtuPDm+APy5Wq79dRg3R4hmQqM8JUJTcPlszviyMWt1bsD1nI3oDB
ww47AZAQ6PJbblXbbrGqWwTC4cD0E7CWcSncMdBAH2Y7tKQpaavRY6MiF3/JmzL6
7GyyzK3l4OiL36vkQmHd8b3tKbk//fjNUEysysDpImGaYgYwtnxanUm+idKMpIL4
zxzy1/0viieSjPg2OREKhJz7XhwaFpjzWGOmuEqDBh3DAUv4v0IJh//ZrKV1uSTR
la1wpw7WAMoGPhrMiKEmPkWQ2L853PPhKguLIj/niZxdLQsbgZm+dutPoukIEHQy
c4s8+q1JD1z0rQWKJ356VpyW42Q+pKEi8FnZB1v9YJLdlAT62fGg3n0tH0pfEdnm
ROfWn0y4aSsRE9IIMK7BOVtE3lddNeggPiKErNXQxiSQH85wbD7smSy6VYd8sUxA
/T2SEEwXNdootIS2JCr7t3ZXWei26/CGNmCotHzWeJ/TK/NFnkayt3XkEC+yBy1U
Zo+SQFRUCOJ9Zt33DkWsFa1Wxq+nYtTg3JDpgr+Ygq7VaZuU7HEw2n1zQLq5/OxF
wpY7XO3CVrqoJ4wV5W/mCP7bmDm4JCp4TPp9rgzoV3HSFjhgHmPdo8RACCEE0sVn
16/C/DTrfZGFoD7S1hYguHY96qwWRADB0pEoYAuYYFn6/j8eMoAbNu6Pz2L4PXxr
SS3bPtZ8oBefiGNXQTPt4kKRFUah4ogWEBrVNtvQ/BwgpJ8re4kVRhzbV9y1XHD0
XIyiCFnW5HjubimDJwb+qY8pItgJbfQ4sH/CZHLwGC2cG/k60oBQh9mxa1mdqGWy
AJVTWfnWgiIqCJCIjND9X+WsI8DCBAZxdUWzMSSkZe1eznAT2309kiZGI3C//K4x
vnfukCH8pMhT7z/qG3J43ZtKlEf3VSFMxCr7idIeM8Ah4G8Uj8w+0QJjpikTcFnf
sqOlO6MJs4tE+WCynLIvoY8EEoBIZDZXmeUBqPop0LJweNofm1/BDcRwToLe4FKN
JNkUcTqkrjZ0qZz2Yez5SPVWJR4kqQwwAyU6mdO0S6ULVmSF+tHNz/AUe3O8CFLt
wrikYlsxtCqAY+y95VwJGcmv178AxtKtWOl/tcdvDoI4wxPqcA5KLzISR2rqe78r
p+7jJWg8bInVqfPdWFVvO50fFIVm/D5otOzgaWb3u1Hc+wSEXJVOSri60H8J9Rwn
JaNbuGlE1D2x61T7w3pbi4bgn9Fyz/ZYY4pxNEobnO2+CLhWf7av/L3DHDb++j6g
0VgDR+wf3QnbM/qG/HEqt7Sp9zxYI/E4nXc4uxwusX40fMfcmWdbySvlD3VDATz8
oVGLiJ0KlhC0HIUfTYCuBd3Xk4StIleOVK4cpv47P27ZiNPWLPhTHDH24OOFS2eJ
ZQJLk40CY+Jw+vxVdf13w1gR1OfS6I4rIbn/acGBdveDJS4H5egOQGP9QdnPWz1C
lVuxMbY7/Fxdf+a60WXD1YHmydXZkCCCKhYPwpak6jWFUtFnnnfwSDpHaMrzaFVR
n2SDKK+gEvc0BFi18osxRxLIAnYC0jYbC5uVvNYU6mH76066V0RFs6mwzmm4eJHm
DUTjDuqxsVc01HoaDOXLrEqrSM/ItUNrDb5ev8o7asEBD/hSOnTF/iVowLWvRm/z
ruozrNVugnk1xlPjrPQrAq5wETWanB1v/+eNrEVZztyImvlPmiJgC9Z9oRw0jZ3Q
LLiIWrttPtEZV4IdMb6+pDyD6MVuP0OcMw2bdkVUwbHkTVzG72CiM/7AQlkhJVhE
+WKQnzSHamx1xhQ/KZQrd6cTUCKpchdl3Sz499E5w3zm97uUKuaKai2CenWTy/Oz
kvoyYV1p2mnSXwhtkA0PKvSn/uaDuo2gPAUWErrm0cRqJfKnC8kcinhcR87gW654
JhcFqpmolj/DyqxroV5QzjGW+oVlBIZ2K1DB/meLyv7zqboqfse/jbQEuFCxKu3Q
2xIcV9jJLwurakZexGHzyKWfAPfv2suCbQIJpsI8VK+ie7AAi8SohNCYxoLWOh61
JstVPBohfQHQ+qATDi6en5kPV4QwyqzgDdnF24nzhvS9dhBNfTaDhlw480zQBSzu
+9krB5AeJo4WPuqnig0vLHKvhkJbEjzzt6jheJSVKorvWp46PzPeNjijbrEuE9bP
t2ndhFPB4ovcQs08mCVjYZFESOqXujU1et363YFD39KKkmiWlhXddPe0E0RjTdSw
Sln6tq8/C7mHqzJlENu+bS2kIiClmlaFa6bHjURgHjd+kE3BApyf4Wk84rLde4bJ
mwZSRNXe46yFnI1z7EWE+YyGJdmTTG5RoU3RyqZ5iwOv24CW8BfPVbY8B1TFd3X+
nNZgYWQMUwNTdmi+vzo0VibjzZGGuto0Km6lnRvLshrxRH2T433C9HQUuGL39BL8
tv5f+uMuSFXhXVtvhNhM/T3gCMb1VaTYPba8EgSc6PFCG+ODv7M/o4OGZVvinFXq
hNdIgyHYCdAAvIDC5gnt2uZpCmeylWoKSRJcvlD76cuJQNTWXtnWpQM8eKJcTg2a
nVlzJcafwHL/LGCKoDiJwhrtbbTt/Y8vB1lLMwrsvpRbnm/7K9YL6JK1azrRuVK5
oYSVPPrqO+msITSVWRvSlYjuCgVV46v3Lt7oZwyj/ZRd2E/gbpjl5rrwytGXvOFz
6LIcnowiCWx6eSLeYXmCEIr7Et2HD2OBbbUEWz+K6NfC9j0Hh68UksgLoBpDTNvZ
toFYFgrwNZqy+Q8XUmvNDCrnxGqm046ejW8o9S9/k0JwUoIwJCcqYrVJL6s+7dtJ
rwkfkC0+X/4gr9C7fbTD/SKLYtbvipbFt8p5aEr/Qn3WjjjqKh9SzNqbG9GziVpx
1dD5weOb5uOal1lxf7E2ok5BiePXR9ufDzzTLRIpkquVmOh9YaqExB6YrCLT9L3v
eLb6uOaa/rcR1cFS35HSCMr8xh1WEZM8V6sgrAVn0nOZdcGWMpJCkyxuCav40xw1
pcVfeUr5jyBVZ0GQc0xLQmuwHAkNxDln5LFKSswov9PO9psR+/X3JyfaiXsyUwWs
EQmVswmfiOnAVllldkxiC0VRyO06/V79/FdRyXCmuLBsyTr0TwzoegnW6MTy8/CC
UCeYdQZ6zgFEVALeGvEnYmfyVOu12Mb5VFc6Q9NESQzCeVa8DPaluSj8mfhNksIn
bJ4dQYBRStWdAy/2Ne/9llhfrccrf/CdskediCacgbwLx6NxrqzD952TynTnu55X
qIcAPXptFP5uiLO3BpFcvcSNkJxTpiwlQwJ0ybAu0ggFt4oDhPY20CGuXXPVkJdR
4G3H2DzhonsWl3GK15taZk/zpnb5Z5qVxdOazd4iq78i3tEwJkpMIW+/iUNfd3WT
6kKA9hFgPovQCfBdeRnclCRCe4CkDlK+p3/JVrC0pze69Q4fnJaNEEJ79tdEpnS+
+rQ9Idf013yS9xf6bLteCiZlIpULlclcTk/R3W7wqNoyJhfWDYys4EbSiuHP/V0w
X1gHK28570URvp+jjvIkBaBZWa3UnAQxJfBkHCTXpLws7BISf+4f4kNOhd5U7LHP
4gy346tsRywLQkvf8u07FDC8ZtT8qeW8i2lMLrv8bGhfv9D2ysniT/E+lx5t87jy
lZ4diP3te2fLDbFt04dh6m7+dw6VTDZz4/Ss/01KrKKCm4ENnBK7SUk6/vXRyHxz
vYhH+HPYFqGyAYWUMnDin23EIWitUg7KeeLC53uNR1I0TEX+Mt1F3ZYKK9UwMbQB
kdGEBurUA/7gpXdB3aIgpy6+gv4xp19ANkYmEUyNT3WxFICaNYYcnOved/PCBKeY
G4LP0+GJaMs8vTqayV82m7KXoy602AQsnFrj3/5HlrqAW6sBc209UtkdudjsCpbt
YmYok8GqQEY1jGtsLHAPaQtEB9u7J5R1KX5EpIX/nehD0dQql/wsqqSc1KBTX98n
PcBjP4jHkd9QqdLGoOsGekM0MLnHpld7wQEN4K5pTnaDvFlSfpDle52zUq/CNAvC
Kh3j7xhCH+WqYWxn3bT4miCaL/zf0W2D+blfjR9aFBQji5XQOvXFExUPlAriNkPl
WDhWWLYijoe/KT/5rFdl6iqUfTMOzP946p72CvLICltB4FzNvd7A9n2PcYTchFji
r32aMc8TwlIX35GNAmOT58OkUN25tw9l3vHxS8QtFYBn6mlFkWEsJMvuuuOxGpiw
NqTU2sxdtN+qKBZO45BWS3ydI2wVWPr7G8rstCtYwVrvj2tHebUJFti0V4+4Pb00
BKTtm8iwV2oAeaSzW+6X+w0XA+SO3xnEw0vP1Z964UC/StPCEgZzpeHpn61IkBH3
ocVw8FK1gHdpAWGIEwWAR/WYiY/apzXJs5hv4g36eWs6erJJyZAv3JBke1E7Hp6R
i/3bhpHR/N3vRjeJDLvQ2EGAGMYZrK/WC8jqzRZhyjL1B9OlDJaiJlkVKY7+KfiT
Z4IrZAIfrcBb2DtMWPqT3A14BDOEkJpLzNMiZ05g1NMrCKdqh/sZA+O1bIlqkK5I
WAEkoqffpKA1um5HTts0vHCV/ZsCa5llBCpDL/RZcZe25Ea2W56zQ5ldo5yqWCZN
52Pz8sRnrYrEBZzjyrA8YBhXnUZt1tXCY8RQhLavDSUspp7A3vvlAcD+D9qKQ/kD
d9bnbRUFmHvyvZCX7Ik6uzu0opGSTOx4kQYe0Nas3YufvfTQ/gWzik7tivgycjPX
gTvISm1sWT1SOF+kd+VT5XAV6H07iSYAhpVfpXAmjcdx+ctEpfhHtqcjK7AieZsU
nIBzM8HTspqNlbNONlV522PFt0ojOiTRNrx2Xy6kFiP7nERvhH5c5zzzHVBatyMv
vb0aQt2G5Nujhxpms/1+TmP66FUAqcTIn6pramUfYjRWC68apv/lT1pf9qlwr5fX
A2mJdNp0LLAYVdJp8m84Og1pPhf9UTluM9TJrDYeqLy2dEdVq4/+/xTgkjeWTigd
spPNigFj+RBrULMO7qevl2nl7rMQOtWcxodv8NNTV9nmN7vsmOnvldBaGjbj9lTh
WkEmZei8mVylfsqq4eVMnpMGGTNnXB3Y2ZXhcRXYGDM7uPPbz5D5NfYVexN1NKKK
vj9sfGxWe4vbSCkKUN1J4RS7JFOTvLOC6vfY6WBcf0f26R3v7WslpLH7w194xnev
bCY9akS50rIHDU3+okKeyTVTGy4DSB7OX9P3xom3gICx0uYFN1nvXGrqBCblsYLb
/fS4bBtz+6fYrmDVvgsgNiUEUMqwThPOdYFJFAsPTQMStwKsTfHZz9a0V4zKxXRG
Ncs7PIojR8iJmgN1PjCKLg1uXISz0ljvKzoXF++fFzXf8S9QW7h82o4H5TTCAi12
twQuQ+e+cSKGFn+kQIfnAx5PwBFI2KGBZ9qB8Erjp9FJxTYsb33SmT1RtYT4QaT9
x3IWuFqIJ8vRfYfn6RoGHEoTOAOOJkdu20grLXNP6cjfaUZ21ma+r5ZwsrqxVCB6
sDLzBpJVLcOsPWuIoDa957rnd9nSrr4sjEtmZMnheMzBj5lWgC02mEGJRNA4c0I/
QEnVhv4x92uzOSnttXX9RVhtjfFuLLTgvr/R1cJYtcv9DHcAUXmRlo4+E+0wngTf
naogZ2Ts5PeTNwD7aFyrSlGtiShHF/Mo47fSDvC0WXEdfO5sf6Lkzi53l5zImC7O
nv+YDR3Qnzf010pIeb3LadiWcO4a2y5DDV7LCkxbOzxiA66MveZvXB2o5V6MnDYt
zhF8KIUQ5c5VDDe3u+kxHFiP6N+6dtrHPS+81NJbVSnZiYs/EkbKV5ShdF+MPE8N
n4QqN9vAe+cYlVIh3IvZbQgA94LOdgZKmC/2aKu7ZDZ8ztmQ27pWSAsaY8MGl0CV
2/lP58/D4qHUwM00qDhI9XYJjSrgO2LDh/aN57U7Md1mf+Re5vOFHantxxXMKC7e
NBNYBhgzSJFgTpPTlyGInyp11oe3hEso7lZNI4aeUE+bPNTNayjNivXtX+E/tRn/
Wkwz1nUeoOLBPtx51MoNEzC1fDKn0tE5tG0xpHVcZz8GUAISw5uEpd/QIN91JuDt
UalA0FNont4pRSzcnmw3xO02Sm1uoZganUR3nrNGM1VnfEXleOngYH8ps+Vt241f
+EmDdN/tJj3BFu23LsfYGpWPQH/Q5TZ2z/JOyNa/t60NBK7StUlRXlfkUBo+3ixa
95SuvfuZTiDvt6QZzXpgGoQsz29EzfJnPeOVPmRPJuRwpkiMUglo/CaDyhdmpL+z
1IEqLh8L9KsmkEgiJ5oiOPXDMsxGEn9JPJgeL93/qIIT3VOFJxNcpU2EeLxaI1YE
OjXuhgD1CdTGCQs+nS2OZsx+GMDqxBTQblYhjx8cM3/dHfXnzlvpFcT0rZ9NfYad
qllcrkpgPVEicJVPTeuU24kXKLZqRAQuXHzSJpWe/4g1VJvM2mJ8mcp/zEC9RgYG
jAKBLveIkskA2nji6484GJybX8exBPTf2rF9SeSkcKHBfWhXZ8TUV0W0ZwrGQcyD
FokbeQK2Xak25mvilODLnL5ApRg6jhUnTvC2xBdPfjYW0eENOJtZtiyv7k8MMp3c
cIZoQ6th3AjrEuz/mvijyM1oiJv4EjiIoPNQBbk70rx7zEoRn9nzz8ElaGlqervT
a3H9ncWfFNju9iBQQ3aHRLRuLBrA7Gx5lpushHbPeCdZ641perDtqgfb/vlSK3YX
lFNozWwgfbmHfJHYNFusOsO3y7WU0YqUPcbZ/pp6WR1G5I0Xind6O4Qj4D4O1qcc
+sraz4G8dG7PE5Hi5ES5TYF7bg/5PiA8yW3YeJqYo1Q8QbSvZOJe1cJgb258uKJ9
J5B/bKEaC2ObyLpQWXgUtjQnbstPVRgs/cVV5ImsVvfqOVF1bYOe9rYyjOALXZRr
dbFLoobX+4qHUKqAxFugFTeZWJ+TP9XmyUZ007onI5lHU/iOmJI3hsHlC3K5+KGd
UQJcGz8b92CmsbCdCmUnIefk+X0Q0FrQ32xepcFphvwnC0224zlm7dItPL99nPQ+
xNWZxZfC/ssp/F9QRndGoomS6/Kl1OmoV8NvaWYKapI8EC3zsz+1LOEnjoZTbqiL
gyTesOP3/PqbPe8+U+u4atnL5Ew3PIwBIIvY+SxaeOohw0modnMwRym1hc1ZbNbU
s7z0u2CF0cXzJJm9LWcNs9srXhRm3Ts+olEF6eC9mLGy7wZqtJ6o4kyGtPWBdXdX
iwGzaOabyRpcDUxRkbLB+nw4BPFRZ4fRZ1LQzF0v5PN4QmjVbgVPNllq+rKvhqW8
jX1BY+gzWb2OcdVOw2wOuDMKp4E+XasHnzqzQr//BXiZyJrJBNr070x2gOp6iK7A
fLLKCI1vl27x8ut0NPWYAqcarKX15fgTwhpF1laVes4fa9+vKGLrg2z28zx0k77Y
QBl+k657qjUywBHf+zPCG5NWHmMOP9hOxz6WHp69m/K10c+CviRvXg4kvDbQ5f7m
Ix8b0nnBxZmZeiCySxeZ3fBKaSliS+6tdK98flp/d/ypyExDE8jLavAI2u0y/vwW
G0FAmXKNWmaB3jttwYb96e1HGNDmvgSYKI1e+375goRGzYQ8kYJKXCMCJ2qY1jzg
ImYuEXY6AHuQZKu9bKIY0FsvgmEld9gqg54jy5yplKacnC2U2/7tKYe8dliEEEav
Z/3J/R56TzKcOvMA0+4dlETyn5/UrnZV0xKkH1WJ+P0AmcrkUR4nuy0pL7sXPhFL
nohK1pyPLbTJQ/de4TFTMnfm3LIv0tRoooopCjK+P42B1sW2Hrc8ro7aHQh7TUCh
4p9jQlZv4PwI2VkCp0aK+WBoEhkTD938gHAf9fSf5SGIGeSWEDbK0fFJ4ouXDy8k
JWnyXIHmZ1HXb/hpfjGtShqbeOGtFzj6Z0SN2BIN/mVo26BM9zWa7L4Ctux/NlDe
aY6pfadrOXd0+R0tsuGku1SP4WNGrqT3aLACleW4mvae5J04pnmJY4Id6i8DiMYF
Mc6K1UqOTa/vDKCDQJD1iHEHG8WjnooWAwPpmH+6hTtt3z1G22eI25GWn2FEq9DT
lbwgjD+F3x5V+V7Ryqmq9VaeZ59nx+MN+LxevjR8ypubK4FlOXkwgAvWQzs2lGtM
4YIYaRQdt8oLQEv9uURIpAULVP5d4EYtFLFhioRlK+i6/SvtgYem3JUY+wLp7kz1
Rjv+4tQfTh5CmP8yP076g9cFRcWKoZvkaVj76gYio8S6ZYnOuGEattTlQtnxc1F5
cpbcRUCQHXii1nRqdhz2Q0BG53BLJxY1ZuJW+Qz1vF/IvkaaLgkpmdOpZ6Bek8Wu
4mpXW8Nq2k+TTGo8n008nEA9R8RfGsRtElUfJaMmmmcB1tmnj9F+Ij11N0pNtUjQ
BBfoE0C540RXxK3CqmbINSKx5uJjfT5YLYQIZQsGLKK4jgcEY3HiKFX806l8AKTa
8xqxxM/WXaF62mhJ30ADGiPt5SUaWeBz+PPXKKRs3uXZqdrb+WIrJb52rS0xNZBl
dfTdIK8O1mwhnSyfzfmht8jkI90xZLspn8WUzs99r/xWwcjjX2nFXwKGMHgVlIlZ
8OgZYe9tX6YpR7MANfaiPgDGLIKIgLTLN0uJksUulddcqq5gZn/tKAw8ZHB79TXE
kpFhd7w9ZjWcCXzaEDS+2d4lgM5GU6u31plHq8hJWsvl9qqX5uF2JgeH8+Uzg7tM
Pj2GXTN69iQdWLPwLhDu92hJQ3UfgeDf7kE6Awtsotrt7i+JnAlanzbOHipdKGVj
OKpKshU33Bs6fX2eVaTkOz9phRmhM6xAUZ5yu8noc1tp9PwczbKCZ/ud6Uvrj5fo
NzTMUJM1Q0SD3zYqEN5LQZmhW4NRHR4NSWONBr48yoU737x0h8AlML8w+C9A41FS
gujJ4z4/aBJpxf4jWvk6WGSHXdRI7Ug4893AAFURechryyY3spCTtlI6FaAuRZu2
OnClcKLVF9wk6BDN2l/8oqEU+0i8MO5G30dhfIDd/3QXgjS8gsMF7SxgGFpqSoKi
wJzipRAXDgFExQrCNE15TUNhQd+Bm1/GRy+fZWJEJCP5wGLLEQKAePmlZV594mxw
llZ/9SeNmxJ9fHewtC6gyVozvkFvAI58e2Knr2X9Q10K4lxCJizDlCI3UPPxaQwN
+sNq1B7JDwW9DlvU+p5777FSs45MNGDcpqnAnZDKRLLFhDPFnKiTpaEpGnabkk76
XxLUaIPsDvn2CFnOpp8cGDZ3v9b9j//JH7wdneTzwY1kTwY1+zfRw06XpBIFxDv2
Y8STBtlIXCX3heu8ZXMfovDNROH8qxPKLNfZTf3AAEObWnBYVpmVYgGu6KG7teny
6gwJgC3UpBc+D19wPWJ0qS46SXwuNK8bTllDGQyHaGoiJfeQxgvP2CHvRHV2bffu
B69op+uSCtX6ahKIYhI2qLellBnDS9+fPQhB6xxWZmoJY5cwijqZE81imLX175O3
AZuMQ1hTBqwdxbwa4ZKPnhgVYk3xousQYPEFwoC5Le6lIt+U+qYuiVYIyjloOrgA
N0eQzyiFEkOUc9oWT0QTjxLF/YEQ+4hGW5lalQzMJnRtl+3v65MmGG9PqiqatJMD
2jcVHqDpTHVFhvyujzGDdihrkzWgnkZJRVTr9XDyMii6hT3qqtxLfdMpyjFAGTn/
cUeEE/Wtwlp2ui0P6vtNzHpNPA+/qcIQOc2v+tIvoRCWEXCSm+3fPMIol01LlakA
aAB5fiHalddouxXoqdNWFve8U+W7FJnlb7aFQbkEF3CRkzK8o49QjveFJLIdjBdE
k9EIpPchkfFhBq3XJRzbUDcx1QGK5CF/Ds8D/lNCOxW0UKJc57WHj/Cpq8hZ2cYS
wesUkxh4WUqne4lHHJNo+h1Smfr7JVvpEOpWiyrbibA2z167Jbqc0GWOMULytZ56
xj424hGJCk7UQsPX5r26znBuOn80uyMWJcLYXlLP15eZIKe252P7X/1y+0ykCNfN
ujjif/XenyEiu6ZBZrPRyhqFlY5OMo3/x0FOoFQ4cgMnMJAfytKKxg2jw2Kp1Q9r
p+PCbW2hVn5UVry5WRc6FhHRCIq74dM4nla7y47HnPng1yiUWX/CxibXHSCngRA+
PjdHGxCy/aICewh+QGaRJHOQmGP6xB7xDKTL0NGW9sMZsQO3G28QDRgugBpSm5Yd
ZGmLveJiTJrakGY7+gll80CTcDfF+Nahwp/+jSAz0sHJIBhKcOnnU5cZkRn53vHn
Nnb3OfRNlxuDf0g7dLAzsI60YDrlAZaS4uf5VVXxQEWRlyhAnJWqD9k5yxMEMBlB
Of97GFOkWIYdjy3+bC9atF2jogW8EY71GQVE+fgfRctRsXjflxgIXoXDHop0Hv/o
nd9bcg2UVkdExFlQVdE+Tf5xQKhXGbtyD/Ppr7ULUkvEiW9F5bEbrvQZfeCdtACS
eRhpU5kqoMaMKBUvWWAKqotdkJrg79Rzd3lE3EiiHwtZ45ge9CVVilNG8HnvRoda
qASEmkeGh8bJttSMwiZgY8OIKjlSUS1FyMet3TSavGg0DLOnzVT7R0psQj7XwKQN
KPLD334taDa8M6n0lpmHocelnRl7vdNAmP+Y+qFZ14HQud1rnOQkz0WcsMDTL5gh
UBf9v0JNVk9nkmjfhr3mGP4ZggP3EJP1p9YJeJ1s67WT43VS/4z37nPrjnr2EtFN
zVMM5bibw9RBQYA5Bpsgmc+ip8/I/XE0xrxdWDGIUkkG7Rx7NwhXofS/mPFpgJIq
1j0YwcLXK6djB9zeV3LGuzwjuPQsPahMZz94QZOXQ56vwu189eBWkLUVRHtsVgVI
p3CBIjJjIw8thznIV8DWCfkqBYiHz0ZI1/pxTqvUjwoIWRMISyqXqCgohebWr0VP
LN4h0t4+VQG6WK5lZx7+/INur91DasJV5uynG6Gq22c+SftGRSo6cIRUA8Z4KtcG
CygSomP+huNYVnMlhmGEwKNFrq0nt1tGuoVT29oDIyGz4b3vmXPDQbvl6Y9FCSZK
/0oMM17nY5PeKePqysD4TDeA9BaHk49BaM8dbpqt7SUXKIRU8uERoP4brI6g8Nw2
8O0TgyjEnw/S/MRujlGyZgs9KRmmtC7ytO0X5BqSsnrR5gN+DR/K5KFUUbaa4KcD
srnvXu2jGqlqLSTR8wMErfv0GlQ5KOhX7uFC+Rb6Ytesb/JDp+A97mV048XPgoB2
nDir4saFe81cmMA1NVWRU+N3gVgrP3LEuFksUocJy9ItHybDvLtIKXOmn5EK+y3v
9ikAasUBs/OP5dCAl7YZ+PSeVe3hLy9WsDDIEhVq75E4oLzNsVGrP//H2KFNetAW
uRkU8nDz3+ZWWIF9ZwlAVRgtQjr3oszwPVyLhbwqFd/3RqxaiJcakT9G6vSJ1zM/
uhZ7NWd2KeIfBrFL3zrrwIBqDSq2nDQfEUKqHt/AHFo590cqLnNlkdtPXmLxnU/B
YrXMm73deV8eFt+oT1jgfwM7kNqwejN1i2Mh2V/CCIEsg28wGRilrQ+UYO82fevX
OndI6Hy8l1LsIX/u470j0F1F3Ss1k7tZpzUY/zduZX+/ZKuxj9f6YWUF2yuV8MXM
rMgWv1YLrvrKQH9lN30KQZzjl7oVGWXC+VWXfNDZKnBkXUbB4+VFWOj+/04odwdD
aX1rPWk79jBRMnIq3X+MfjNj/pmquVHvBAEL+YIWDr8YYxhdlHcMJE0ZuojqeCI1
xyt/CMKz91ps3BprTjVJxQKv0KFS7ZeX/uu1eMBNxc9GEN5YcJeYxyAAHcYCGTr1
s4vjQ5ZbuKON/YUtmXmpxaxdDhv2y4GatTqvjIdFbzKWM3zY1E0lVO+tEYVve2rn
3TuhcCQ4OJhwshTJQ4XyXl6E/8m8nyvKq4iKKbz7vGHaEJP8aMg+ud1FJ4fqP9vu
K9vz3vp9kB+FJ4GDrCkQcTp9QmzPy1mGA8mNVANJSrC/3T3H2WowhtQrUmBHRL42
6aqgBIfKIZtXQ5iR3lVxwSHDSXZhz7qbanBwyiZJRApIt67WTuB5NcvSCEbrKfSP
G0LDFL5EM8z1BybipC94tcZ4zHUwkr+jklJyrjPQ3d6X8r2WumXAC+nXcy6TM9n+
52qiHaMuuFHaKzd5kNuumiOkIRTJbgwi1h47DyEk6TEvy4O9ZHrSJ3+pyMaMNGeb
wtl1Viei8IWHse2KbZx7FHKNBFm0exbv7bC6Ym6ENmF7wTWVftKQxFkCCKJ24S99
c1++oiGq8YM9ZEmErsXDlIMbNUlMoyUdmAFR3JmS7Dhelq9Rhv9Jc7OUZkAIFeNU
EglqruEtORIw94r3fcqRTLJOOR/L9r32rKTY1WR8dU6f2iKMno+IypuS8tMlIfA5
WfpNvAKKgbKdhKikcHG4JKkKYhCq1w17nr5Tqza1U67+KfYjbeNQIFXoJ/NR8ZzD
pgtdUiAHlAgeCpitui1SMSPK4ziKXDr4YSdKP9Q9GA5nwRSlTCwmHieh6ianQhGj
EvMyK5jSropidyY1qt2vGuUY6WpPRpYboOdPm4F+2xMs4sueCu/IBSaMmzMeWufu
4HkQ7DzXGHcb3mAUiDQq1pZWN3Vcdckt/108anIO1JQZBrUaSaPTr6poO2ze9HsQ
AHi/VA7nXnq+ihYxAnbNFL2D804L+FXjmYoC3KITYCy023ySuIHHKPgVTwB9hIrt
1J+WjXxYSHL+5b9jxSp2H1hOrzRp/21KncTKMdMg2SZgYNS+h4wSALcp3nbs6apL
kEYHIzmp0RlwzVm098WgE1P81dr/qVuykZnnf+GOZQiw2vgtdTQh04k6oXua1hZZ
2JUdPwDpw39n/ioqBtaWkiD5O2TViYIR3JUIMwKguLeda/OIgFf9GCk3COGsjXHX
rX7kIDLiQOPFL7Wnw7n+R3WrUPZk1bQwEAen1olgs3a3OcRx9m/EGadJfAp0nMwS
WeFmX9rYlDhfpVkZdciwLTfpEnYKiastirDeipUQ8TiW7VTRNpwgoDBQu+0du39U
4c6EBftEg8GaPLT3XxsCmeLGsSN2H8fZURn5bIYn7Ixq2fHttRKYvl1Mingxeyu6
z+/ecmKD9uhs80hDOLtG7qoyasg/C1CbpG5B/+9t0sZZMeLR7Hb9tWqly7IFIlZi
d5HOofWM4/98e4TfI9m88HzbliD3dbYD8bzCnjN7uJFFquIma8hADw6R1awtUnMi
F3R6RtN/41Cl1X2RJR8RCWiCLL3MLYJynLrnAU1K+QyK898yqADKMd3VfNjd7D4p
/Nepypn7DewDFVk4bJbED0o+VzU8wK4vu6qPbY8itEhB5BpByOWvx6bEjxRli79z
H6/lOPFJpGp/G9/zmcRUlFhQPSg8thFHDpUN6G4/U+c/Lm+MdmGL25qHOHHSPRaX
wA7i/U+WPBrCPVHKr/6/+6dhY0BFYRx3RvJYPwdNEsbX2M1MyHvMBsWueCHQE1WS
QHYfpaZ/8Y73NuyC10gLf3es/RlDa4NZdvgqjIXqQtCYJd3W0mObJR2FOnyzuWx3
Vx5O9/Sf4cmLARqiKPcSdYKUtSMyda5QZSGxAc5mn15YHahLrT7amyf6XIfWDp6s
to4uTsaCBA5SfctqXjkU3CfwJj7F7X+MtDZTJxIobmQXhgnR5RtQLsZUTZ6IMdnh
O9UCN/fpIsFtxOV1Yv4sFoJV+UcsBIAXdlAHb8U71KF5AZlwLPcQpN9wOEYRbass
LeGnLaT2D1QIFmAM840KHBDM3UORAcp0jDb13ZLemosY7a9yPCRU81UsprK/Gsfq
xhAw2mgU7yMxyGFLAb+BQVlBAU/UumKzlCmLyPAqUqCFBtNnLloodu89wGnUqO3/
ovl2p6RG0TIU/zN/PlQm3Gb2I/M7RV9hemEfU0m+hLCiAVRF/SWu+d8Ba+D3X5MZ
/dS5tNLnJkQhCtoLqMfJyG4pCnNAChzktt8HQG+HLnlDtyMmO4ozi7eZB93gBTE/
aYixJ2c/jpFoBbmzomhIWXDjFv4M8QDgjISMbNazEPkPaRkumaf7SbSNzOKfxF9s
LCM0wFCfay7DjppL3x7UrzUo+JtzdmQRuWNopZ/ey0nUn/hjipqAU9tBazUqwj2h
EUimehIIacyX2OdwkWcamOfcB7NKnycLA53NMS7cms8m5lbfF4eRSwRtnjxgfV/Q
nxZxdoW1ztYC1GNEWaA7oLrVFnL03DyZtCvTP8ND+JJP6MspeLdq/Savbv9uN5c4
xnWIZE3FWvkzGZvf8ePXizkG8d+8q2lRk+O57WoYj1uz9vh6RYU9FNKRuSrlNuQ5
EMimJytwmdIwVD8uSY6CzIWCqyaKPJ6HdidIg+47l4ip9PhGn41eoi4aaTW9HF/9
meZCs+tp6QA5St8SHuH6n32G9cwIS22H3/2YfaBAxQERHWISy7g7llCPe6LwsiTV
P6bZV5A0Fkat3PyLjlHVmoOp9gEAEpblGB1VExyQ18pzurRaVblDG6D/trVw54Ch
+lhPNKSjE/iQSTguOs8kB/0D+23mH0pAH26l0Ydp28V2wNtGOfYuxsPY4rW86Wj3
z/JJlgGrC0d87oghuqcg3MlIVkAguEzVaB3i10zPaHHYUEH2u+QXTNOKkwQLJvkZ
xFop7tiwBWzstc2fNqXhCeOUcooOWBMqMcCU/Azi8b0N+LUrmEolqN7jg/DWuMrL
DJK01gUqcwKBH6pSNz09ZGQhrVyb4lrHUTSJbL6fIKnD2utcmyBDYLfjTZdY2w0B
rDkgHeqr55ptengJOf1bthPKnNGscIRytt3Im9/JfRtRsFUVIALCDf+T2Z2U20CX
vJV4vLX7TKHs9SMMNfpcI3rvFRh/QwISYBwwvgTCoMSaT1tW/5tdVhjYhHYRCOPZ
TXKH1CW9wMjQ6xQs8tIJ9ayZ20SRyjh8gdNYLtvxOR8jgUgBkvoKELaQxehtGFVe
l6BetTTESGhwsajvc9DenzX3OkJIaa9SmnO5Pf9UcGPKGdZh0g14yPYpk4JXlXb4
uNqJ80GD/w6hgNfHfDxkaBBmB4UwNN14ifbBpqZ5Lo9uLtYYQMUCYt5rqM7HVdJx
RiwXDWcr8zi7jFYN7bZwMvx6kZjO01EQQFcjr+i4LreZT8iVRvs+3F2DnnHvje4G
XJgz3R39ihVSEeLeZh6ppHFXavh7pB1TM6L/y0z0KVNae7Oegq0jzK/LPZgbRYBu
A49t1KrLbLNNIaOHMyj4BbCws2f7Wk/zqZOKiJQz2GpqNmoyfOov9aKCbc1dNLoA
oUrG2T+P2sHJL1h1hCgWdsBQaiZSBhUp3+cd4DxN4CJQII4XTfv+FjtySlY/Uk6W
BNNUpM+R0TmN65fGqTw4JoetN52oMBq0/imUwLOvCsBAgU/K9M85ZPz+KXNowuIC
uxPNVGWLsRYVrJxBZY/mPw/Wzm6gwF33gkW+SrmycZTSwsQJGMKFI+TWxp15YfmR
ADoZcONlcC8IFiuUlO/3xwQWPVUudn6smPDkYlenIK//kNH2Q1t2xB4RdUkoXVDj
FwsLENb3GhSqc1/yFPOwW7R8rKa14UFey6ClYyYFoD4he/n9Ug5QntgnhshWGeQD
RXvDK5mV8Sc0UwVtyfuallv1C2K55k5kjxBxG5aM23pY3Sb9Sumjfgrd3Uuk9nmG
RyzjFUS63UNducZ8H5+efZ6oqGb8yZMXjWWi9T5FEEutJ9lJFcU/8cfDYARD07J4
AQaaORYFhaLyFiNJm2MXXDy4q5gG1iYC8OiGgko5BynTSWE7BKmhfIBKIKZ/otgg
Bp6luIOhYBcra5NPKLwk18VW/kqcJpWbm33p033Sd5oQDqnf1b5bisA+KsE8kkem
j2+Y/QRCC3zrnuhWOV3h7uJqvlZUKWY0/AvQHq6M8dJDFrYEZs6miF5+/1YMbLcD
P7e0oya6hOOzqdKOvuFMZGpjFHigXweAEd+BKBPr1NMJkV7AgAg6M35C9mQsaCDK
NIpCK+KGirR7gK9fjWbwwbIC+XdYkBF1dC2wL7B4DmVBQ3jEwUX5dc9M2zrSq5yj
mMANoVNTwyhXhFRPQLmXDyKKy3by+mBdP5LR2OCtz1554E2j/4I9kB6h62NJrvw2
tfSqsv8q9bjvoqnzy6j6X6brVp8+TfSiOhJkDrb4YOdfVxSca0RfvJqhK9COkbiG
b1ybtX51uSOWdTjczAaHxCGmCh4VM+3mn/zzvNwiTdUzlbUubXTFdyzYKUunYKpD
R1uzo+ZxcfVsJnBcr0XUIw+3Cam2TjppKhkMPW2EfIDNros1hQn5zqbF/8M32563
snPcoCrOHw9u5EuCac5jmbIJWJ8q7boUydLkU/Jt9QkAwfJUTZc9lpT7TNovbPBF
f/Y590FtMv4jpPlDSDYTuGrKTFEqf5PKJ/YirpJ+LBaXhmUS9nz3cgIByImjA7/t
Ylsauc5cvlvKnRwpfBR8gAUYKk7/XBWSyz7q11gJNGHX5XG8689HrPCBISSBbXJO
X0Ep8/j7s3C5+I8lFFmRZRjewVMbHQxgZEG2yL6B94lbqYPCH/0dn462juX+JpyN
PR//kRxCCS3gMe002gtmUwuApkh6ouTqDmAUuQ7/nMCwhA1+gB1oYHyaTyd2FZcl
6sjntIBN9UHdmpHo0SqTrYFwADwIFcwd0JLR2ks8kjHFbrRfmLv3/Dy4GgsZZ05c
lCJI/o0pNxwaQRmT2OUsuyRPIDJ65ITSinFU+d0opMrezKwj2WF1Hyn960oxSRoo
5iqfko24HEaQeDncmmIpze7NOx8/RuxqrljJEc3V4I7bkOfzJ/f/3NisEhESmGWJ
HDfi0AbAViStHub4m6TnskPHRFjrBfwdFXJUNSPmcLLtKpoUSeja9RB+fpfxFQb9
PAZ7szV/HFFNvcmxKrqMWhYqmM8pFJcL8j7OTMm/0dSpOOvIQ8va/BuRrEfQBpk7
M4WPa66uXEoYL/++iO/Ua2jCScEfqpcxtuNCHGWwuGNvWrY/AvUrXQ6OLErXbk4P
rC7VW110Sp9n0+yHfFUzEv3HZWGjNqa98pwzIh/V/e9SbJnFN/bns9ALakn3dPfe
1malsLTSZNTh5hPTtLvFdS0lJEFXPKNNV+HZ+2MbiBAs1UlhIe2hTzYHmsxed7AF
ExIq2oa8dOYfbeWWvZK71Qiq7ZCxyLEjspOlPK2y9ooKLM7SQ/WfClzule7MKegu
DhXIokI/jDJnA8u4YDG089XZtw9Ecrjv+y/30Q9bcYbUWj0lISR47bpsNl3F07up
ubL0T/jrHxGSw8jnnCn+NAUtk71yYjbMB8onXYlN1gxgEc3gSlZDMpk3DD64m6zt
+XBFFRv1A+1vEVclICtzM+sdVa3m9E5QXFU2rW68jWau7CAc4UFvfdcnxqRelSyN
h0M1v0PmMuFhRYIWkK+6ci779rBtruMMphdSx/xRQvstZoKxtKjN/rjzGhZhWF5e
ZrNomtiJesFWh4u18JQdtdWu8tOOdMNGk6wSH9hvpO3U5he1kphkd0KF1f4mW8/v
rBFGwsB81I2d13puh2T4FCkZr/hgZI6WLg/TI2gFksDqiXnQp8wMDJjaSelqFVIV
33RHYvoRNghFhpxyeeexXFp9ZiRI8fyaZkCB6vuMetdczq4LgEAJVt+WWlFhe1Sj
D70D193n//O0jdQ5LhKqncpnteo29Qb3sHVA7F2QyvhA6n0G0XxduAHUzJlYUyPn
MCgBUtqQ/64cUfqtojZGUmFSfVwQp31UXZX+wm+YitOxor0d8CMyt5wJBNqylvm2
vZUxcI4lbK3XKqFj9hyOLxNo/P/KJEHF6CjkxabZrSlpbp4UKpAcwmesqXSMv1VF
ynS9lzJwMP82y1B4mEIAlUEJWiFflFfSPiPuJynOeZ5KW0eikUEN3khaKu91r7Qg
rIVx25XonxfubPMQpgKYiImK8z9ESxIy1Ky3UZjnyFVdjUz9n2my5WtUmbfrPSC6
kpdy0j8C3XK7HLoVRNT8TEYmQs6YR9mqC920OWczLFPBf/KADOPobfutQxHtmOzC
eNXJXqgfTLEjcSylhCmU65ZHgltRDVRD0f/U4K8zxGEcQzwJjwNlRGyfEZLrWRut
Mx7mT4MtIv9DIQYuhIIpsh8+T7OPZUuFEWAzEXoqakcC/gLAymp1l+2HNmmXvfMG
Dq2GsTF5hhVYZ43fbaVFnySZP9vCysO8gvdnL4B0MvuCHT50vihDWJL7Gzz8xYQy
Z8h1L4aXQFdVbM9AcGLTdFuvddsV5PSWukKZiKov3K19XWoyieZvg6QyayQGfwao
sacmmHwLAVllJV4AUfOZAfBmEC0E+rNEkBjefd/YTJSGocSdvP2Ma7IeilyLbdB5
Uln5swNlpc5E3zHX4Ui5XsIXPLEqgTgKePikjnkaGhL+p4DdqCTGcyTl2Ev5v0GS
cIM5c9iUxlYSjdhZJLrTGmv1FkUpATg32adF+aO2yBWwgX1FNttO3k9yF6Z4FGvB
v+/lR+YPZi/j3djebzYVlf4Dyc1pAk7b9CJlg5qB/2x7Q9IxL9h9FEvbhnQFjGe9
MZSb7giqeFIwT+Q4wvU3wUX9UYeWWfRHJ4JyP8TCMOng9STwO57Bq91blrbr5VBh
JtcA7h38DC/B7GOEE4+vtjP7zer0Rzg0db+1ikri9LHJxLbP8PHPIN7b7jHlEgOP
c8y+uyvJMNZlbL91t3tcTRKGoVdyN6hKFf7tJQUzo9yyYutgVJMOT8o6SxbscC9c
vOqZS9SoXithXjMvnoFZ4e088ClQXRF453cOdwAR1W6+nPXUIjF6HXIO4XT/XLCH
nMWKAiFPL5qJ9igev/ZWcFCZebk4ca/RHiclJisDkcudKA5yGEUxFODaAAua4zgw
T6wo6THzs4+tXRirgBYM5nfAuZZT2YjiIc2JoFk1pxn0htw9EeVEnX35vrisFWrT
x4/9ye9udyQhEAnTQieEUtNXc6sCex/oyn2IpEpsf1YH14OyxZn85l2AD/NCm07Q
G05PULDXXman2LFY98/1yUB5yvRYTc7np0ugDIAOXkBottZXpDLQu2lQychCIgP8
y4qCqRxnNsdWGvdD9jmSruQ5BBd9a2WZauZXJKK+e2hhiHrm5eE7KNn6hQrDxRhv
ZAkign5syARW6yijTMsiF9HYFrda/IGrRHjX5O0eItQr/S+X40kT6bdhPEA8mwji
KRVliFLCzf2CxthV+TWMhaGjcwJGve9o8/CNU+8+d8ymSh25pehL0OUUgg+b/12a
jVcrmur3m19CvaxgRQ5hRA2ncQgOzfQu+81njfNZp8vQQNup63+AJfRdVHbMuEgU
2u03/zp0aVBJWiueWG6tCgeDO3YQKq2ZzVvGiT8c4NFGhEKHsGt0XXxTQD75887g
ZGvFMu7M+AybpVVzVJg+bBqVor/cic9pLOO+3V5b+4MtdWjrqZZ7VOr2ZYTCN6OL
0thrdyM0Q6dpTxj71ViWuQv1fEC/hcmL4Ja3FwsWSExSrJiyMlrzzHmefeTk+gFv
eLSGTtWwMrsT730lzZdAVGl6/fmXE1Bg+5BHE014xCVrGyR/VVVjpmtIOAJCh0T8
CG6cI5TDKwA0jgbogjSCMIvEsNCkJyNlgBYTJJrhUhcjsC+BEqwa9fStjg/tcVN5
iYbQgTKjwt/OVG979gRi9QPjmVphGy2NtKNXWoK4hXdfea3aP0DDFYh0jcCfui0l
1fCre2xlNH2rEhz0ZuFnRunBpjiBvTwBCabDAqAWUxYfr1cRd7YRFM7P9ct2QOf1
dyvBtuiBvpGy3qAFdzvgKUpt6Am+G9K4BzRcOmaTg5HzYrtQlDQXzA2nJVniMR62
sG+Nur1YdqdmfHoOab67t2tztpzmnQ5EbWAPlejLyHkFBzVdFh1Y5GmMxhlvXdO7
pCJ3p7ITWugAHPc+/ULk5+ukgwoRcZkajLmLcKz89mdKZhatJbu4X2EaeeeT4x9+
dsKpLm+dhuhtaizhcF6vzuhxXpKc5NULJSpHtjayioTk0MmlB7HldSKGpLPzv3jl
p9IVX65a/mtjxdO2PRhty9FlOY63pHG1oDhDUn850lgS2K+kV1NERjpFp7bzl1TK
sDKz28o4Y+Yk4+/ABKv8MJGvcsfYusFHsaQXacQF8zzowBvmxk85WMOt3j70fdjV
x+bgbefx6DQaCU8CW76qLg60rA0oR3H3xmH7LljxNWSk3TijryVKuhePMLiD2v/o
3SI1GsbpVaLCVk9db/euZBimLq1aPXeGspXQfCJXBW7WAvuLUVaoaNDUwNzMRekJ
njjhoZ6z6wa//QAHemPN6xGkNJGcTy0HQHfXlbtI4YL0iu7vW+OZCKJnuIXEley2
Kj8xw+a+Z86s78OE36+x+cQOE0jqEe6CDOggx3ps9IstjGceSuNiVGvsqfcGkUYI
nDcmXqQog3gfGwawTGkVqEd+Bp4VHjw7HiZnk15C7bnMCMhbBn89cN1k7Ctk4II2
RAfuko/FmHqKsueH4LiDb9d66htMnQIh3EJx5RaCfIzIfmGgdcBpIZmHy58QRUBY
xM8kOvf7pFvgK0vDp5YUaLMq/zjNWWgBqyG5messFFQreII171fmJIxoCLaYxxwO
KYhaQc5Y8Z0BicpZ0RtkkUdJ6LbA8FaUFoKFkMZ7gNj/h+qIFThbYviOonCYIidF
IYVO1DVOjZzAM1pRY0BdovqJFrgXO9jwRDReTxO0qP5v6qJh6AXP/VNIrZp8dVem
JgyKkVYLD3ZqKQXBClXjz/voKICi50mw30GAjzcqXciI80NoQHxzhH1yUXQy4X/9
N7mu1iFcL7uAEYt1Xdjq14a2THkACxVPMnD9P/Z/5v8kyt02tynpPKCdm//7lJ1b
yBBtmb8FNhjHDjEmazHeQW7SdghTdpPSmUqrYUHIYl7AFlahzPyxySiU4nQz/xvB
uW9xIcs73sOBV8QR4zAZFyaT6Xk5Vo0GRntBOexpuNz42GR766hKZZKe8YvPQdJm
0EG3TcjP33PJutPtV28QJIV4xIbpkPSqzLCWXP9oSGOLOTqkuY+9BsZrStkemg2k
UhTlZK13Jwfl48Yx0mULTU6pp7vz57R7ILK02UXZtLCFqmoo6SJdZy7iyUuF4mER
vy6aslDC0QJ2sg5QFTdYpo7QgoM1ve1SR3bJesiPqeUmG0Qox+rOqHSadzqm7q+V
Xb8tptRRoS1POKp08eaFckkG2awKrOQYpc19bWFyAAsxG4PmlB6ld6YCL9R2C8J8
BD15oMkYNWaEKme3nFxecAiyzvYr71QJgQ5GzrX7j2AK7/HcSWz9k/g7rT9qa7rU
51b2KAyZLMtBa82j57zP/rV+A3XET/17jjNQ6opKn3RAN3iwaWgQqn/QyYVbjN7n
peYe/kQ9NA3JTylb3GkkLXH3660gLp3BdOqbTq7ay2wkT1oRAdqxrSn8n3ZtTx2o
PsFNbdr3Oe0tRqwbS0fo/uw0kHTimWtJ9Etpw9LxjCeQOvZTcITiGOhuS0IabZG8
wRxfZGpOZmYVnFc5JQ4vbboTDHXbFQklGkkYMsk5Q/T87rm/zvYrG/cvT7mzRGA5
MS+i+HKyXZnpZDNI611mJdkMdW7S0sNE1vOL4n9e9GDVP+IvuqMnPdRLs8tYqZRD
iFdODXZJ8j8PM9Y91GhXKWHZCSo4/wXK36WoZEpP87cK3k2+nJsK0vMLxtj8At3q
QvVViqi4pPvUGEtlTz2XjY9UydFiUwoSRAUMlCMVYiwWnns5MmnSqhiEm67P+MCX
RGRsXx9v2tFYiRzF4Ex7CcdNU+kRz6G2mGWNCTdZoeIo2z93VovkrjgEnCeEx3Rs
1kU5ZWB93VA8wYRMJ9JSLXUny3/8zuHZFPPuUG4Y9JdOa2Z9mAu36oBqebSH1czi
BxKAMyWvZUbIyr2JcYdYVg3qABrS1J1GsjmRcQwX2cuXYPVkWKs6oThCnE02TF51
Sy3tzhcLDiza/40GWSwltXnpOmDGvg1WmyM83CwmoRr8nflF9dwEY2GUXT06UFwz
2sQIKHvF2lfpK4+CQEVj3gpAljfJ9v7T7yKr91TZA8433Ztkdzpbxpoz8a+hbji+
PMf0dOsSM3PUYIbJR7USK9uiu8aP8EcyianRc0SlBMMlDxEks42xFgP9nXdoaqSI
tedPT0OcbfFVqiQIrouIPfK9++jQpJe2sAsp2XXVN8BXnh83Tz2WB9JsDszqz722
8n3i0wDqL833ByAjxjPJTjCuukM+qU4zWJYrDvZA31gvK0THjfKq+rAE+LdSllRq
IKXIj+RKn17xa21BkdG0jDHsRapZj8MonrYOlQ/tVsvd6GkshXEWoVx2xTe/c/WY
vxGDARliWM8MGW4DeiPj/bSsp3TI1+9XaMi4rBtgV2LqpW1BJA4YH0/yf9vqPn6i
zzduZxNwnRCAGgtnEMakJyaWO6EPi/pC+VNnp0959WsiANEO2CkYNJUeMPeofW/B
LTsvcV3mVyY/uoj33JsZe2d8Tjd/812b6773bnX88e6ONmw7MQeuqb1JURn0gw21
GXuuzCTDbYDz2yefAY5FGcFGwJk3+USTr9kK8pdoxXoCJoenHgC/GWTsg5BCH9Kt
gwe1cvQF1cTXOK2N6fPfQzKfllgnNzsS6UsR44FgAIzuSpkBE37+H/BeGxmMXsjO
XCj4ea5x6tPU4rKrpKxPkjIPrlnRK1ZoSfQUS9u5dT9rZukbU90dNjUPw2YYTu+d
dTMCoykqVDGga8rcm5eh24WPOnOCusxiDH4DF8Jy1wqzz4Fi8ClZXvlU6w0F3ZKP
jtkPY6bwZK0xCP0GldM0v2WjTWkVtOWpmUJhOFBqjQgyOo97QWY3vPgxPray8bB+
pNCcaAtNeN26X1MMPsZiYBJb90WGpz+h6g2RUOQ02K+1sTZ7s4sm1st9dChcp2IT
EbegmnKdhyIO3Pl3lxAYSfri6W2cjFqoP8CZSkgJjYf5KNMXtKlF+X3RBTJ50xWF
kW1PlX9A9oJxy9wWkZzT981EutlPViLrPy3xndtqozzkIZ3YxhoMcI+ei86th4DN
OxrPL+cmrL3/tQh98WKqDYB9/LXbTihSw4E6L8Bp33TBcDEjdgzGYMhI12MCTE+3
IxIlL+ZIZ+AuOvdyDzHG4NU+TZTXX86lr+BTKDvSWgcs98JcxCZ7aF75ZJiWytv9
kEI9NgytfPfvmL3cyLQx7hqOy70tyOOYpqrkovkuFGIkAM/0rQVdRGBEFrTfLQ3q
5wv/WzumPR10lJRei1cXUZIaFx525as/2n4SCS0sO5y7ETDz+23iVJKMEdJh3LAr
cLUwND+Ht00G5N30WTyCLgQpdFxen4y3vijqE0USOM8/NW8/bkVmnU66AGUj4zUy
cMvO8EGWrpOREbSikfd6DpAp4KVAKnUR/hb/5cipHhwrtHooPiRvwkeKB0ZTtizP
61cmgP1xsFclW+L8vWwOsNJyPQRCObp28taME0bi27u7HRPsiYo/3vBxEmJ1ggY/
l2CTsHGchOCtKI7NGPxMDDwPw3qMEV1yFnq7kof+Ppuo5ipnjwhh9kqTc/LFBmnh
cLdKjS4uRchpzi56bfJ4bA1JCa/sw+fyqBVfjpLOXpsLAgVujgKlOZOYr1isLJ+h
/1VDMZlbV3hTC/CRmQxhPR7oIqTcPMVh/5rohy5SqDlhwp15aRnU67TVltLrG2uN
gIPkrrbRMi28FYkj4kdnHuRDaRAQLqvhQp+3YMQm96CdkWawJTx3RzynISu0spDW
QsQElGYua1YnHGxSlYzsbjgsTHlZsQcqCZesWRwqSZ+19FmB0TXekiEy1wrQo47v
rfrYasB+aQuZqma6vsagz3BQNnCPtlfXyvFOnFZD1pfTifdl26ZiY1rCwr9FKeC0
+/uOmHTt/jZ5RaSHB955LQutLW97xtIDHjub+ngRecoLt8/S9ZM+u7PrayWfkgi5
9sFFVhkvq5NkWEGf5taapR2SAuUqraAaoHjhSFAPKK3S53Rub2lgV2lM6A0cegPE
n2y4cgvy3rEk+BJpdWuFSbgrgCi0Hefo8COORk576oHxVWXAVOzlRpZOmQiSVvqu
gQfCtnTcX+7g+nAHhXY2wZpu7WdzhayYPvdbveXJC2uCcLXkgC21oWscZr0HGtBa
/4wiOLBgWogWTNtlWfUXD/rgMflNRegADlQs6y3XRGn/POBQlNjzDspt+M+Bdf8A
lKjGuqjEpCo9Rup61dcK+jsDkM4SAG9nn86R8ZPwVPw5AMIMeo375+bfgX+AZRA2
dtGi6+L5DchArq26/PquUgdP/UOf/1h/j9zvdJ7LCenNj1TP5u5deZoRP+bYUFDk
kf8R8BwF23IWzVbxS/EQK1gXZXqTmNNkGvsP6XQLztaQSUA6VR18CrkURMRwL/C2
nCR0CNI5jMX+3tXCpKT4lHPNhulBdXKW1HM+ju3agDStF6e2KPMeULrAZy7C3aRz
Q8rMdy1vHPtuHuUdjBcJoWz4bLLKMknjULQW7JdIu1+E46tUYDc+z3wiIUGXdmEz
60nm+NJ9mAQEVlo3CZWkWvTYvmYPgkgc41eT9SzqlUsTlZFHeuVNgQpEVrgr/9n7
mrIqkbGg0dr0/kljIiCOrxnETu6eH6+TDNFcAyzg36ybxKkrfJbTnEspxQgwrZGG
8RNUjTKF+alAiFhQ7rhYRSI8yGSGITHEQAzlUmWh3gQI0YGmdWA8g405vcMBl7Hz
QHWYhzSLi0jOJyErvkK53G0zJjo7m0dJeZqXKUuOBsDqXyUpgWeP89AmgrYqKFsR
BzHx4JidntUpKAq8xy1Gg8stiXJ3cdadrut2zYU7QrQh1e+Uc5w72/aMe98VxC+1
ljna48rvNpMcgGj2zA1mLUP1mtoSMUUx9sKHglUvSrkL7YJy6c56JmXORBp3amb7
wJhuesGHBweD7s2qEuM3eb5/sRG4X2AquCnXLZnfNqyk5c3QWy0k6eCD2D4B0TfG
9kqOeaHcRWRIq8wdsk1ntjiWpXgGguWB5tu0smJ5X3oAEFWYNQ2pgrprHAiW2VFG
/m3Fx5pmrKRuwf6YU8bujveB6QhBnZRs10JucLIu+XbUAuDij1yLbakGjBed7PLG
qWv/sez2Zdfb/7BAXRNB45pPymdyBRDhxS/AyxegUihYA7wUKIupCd3ysKftH5Gs
4gwW9WS1rzLwO5FHNTHEiw60RsuQH0kpC0umjbKO8oeJ/UJb6EJ2e2P/Jc91ebF6
TOMWV5aUA6QEfsu2NNjAq/f3lYAHyJfn+9Qpby+G1PDpU5PLYAAq7Lwnn0zAZWnD
MKWAMPkotjdIh/UQrOPN/c/ohedw9tijcuX/311hu+a5RZw268LRQdCShl0g+Qna
bpFz/Tq9JT5TlQ59S00DYnZn6i0XLNIUzew3eOJZGGa79w1+TiPdgJnRhb+NCw/Q
8pzfDw27yllGR8qOQjkkcway1ULLVhLbAur2bsHu8Xt0ufWqyyQRI+60G+nDPn7j
dVXJ44Din0TTp920kfDW/adwgvSrI/OWmA3ufCspn60MivxJ0S4Hkr3FcsFsZxHe
zPBr9Wwdu1b0d9VfVSdjDfrWoJGIiqSkbdJGuwSsiwJQNQ5jARvfHRh464/Oq5/A
mOyUYQVPCjXHaMGT/S74OzpNuCUIlNfiL95zKlPu9TWPgEtKGDdZi8uJ+xk9K09q
hFK5yoGxyXZIybD+Ah3Io8iQI/VCNosNO/X1QysbzSfp7P8kQH/FR4PfIjBUDb3E
mFcGee1y0/Coz+VUWtBfD/CtfUPh8JQWuuKQv38yo2wzg42ybGWece7ztNuiXWlM
6hid7pC1qHoFj2aKS2LVoOVhUsdkLOEuwnt5tM7tKwgjwqm+RXsf+6p0WNCg0n7e
7aQWBQhrcRZQxZSWI7AUDw17XGXcR2vBP0Vpv+ES4b2uI7jR5A8zMceZBD18vxPd
aIyua973ED0CHbdFjF19kmPLB7b38lOZWF7uz55S7JYVxePcTymKOoA9r0YPe9Ib
vg7iBbtnthiM88Wgwcjo7dL3MazHE3TY7Ej1CwIjuJKIPMLn8nVsTG34BK7JTSo6
81tO8P971z8XgwP32atDnXTeXZrAbxigxn3qKI1lDMr1PorZpwBaIDuzbBlUnF7D
HFqfxuEnREgbguwBd1SFQgAkOK0QrDNwDGkB9ykWA2N5Zg6SUeOYnE/sPHbkVwMG
qS8Kmom0fOHzN/8NMfCRvsXr948h36vhxMRwhLzlD1fCVArcj8te4gUXdXJ8dduH
9cYZ+VzPfHvG10T68LsaN07Ai7fx5REYFFjLa9EJR/2x2O8ZcNu6jVTx/Es3if7O
OnjLzZ+ZF+a4LCJPnihvHt10MNvsDP/oSBzpnQr2C3pSVKvZZu3cD9aSo7M0a9pb
p6DeL0XxLemFFhJ9tKO9oJbjxjrB2xlTYIpe+P5ElkJ6ZtnkhrpG7mF6Eeuq7eVc
uTse02b4PpPcYnojv+ey2nWRksOpCC08bOTbh/z1JmNpc/M9Ns1Vtv90Zcpzndkf
QjZjCLsSGlhUQMR1LE4r4F7UadES3nH8dyIq+Ee6fGD44CY/EG0JdXVadqwVE9O6
nJYimzpNeVQuCJGvzGDWZ+eqFrPvh6flDWtxAI0I4P87MCcU863KrhRWFgdKuGze
DqVvMoMzX93eMYNZ2JXjwVj+PWMBcTUVkv88JuSHHCSqLqVOIpEjKKQ6qtN/yU7A
qzaA/PMXLsd9wtSqa5yWJJw+RRv2gBk7JV7x7vBWuWrlHTI7L4rs19pbGYY+4R3Z
axSRajkyPdbzoeG8iPCWxHNiajZ+tk5TB1lMOMVhWuSOudkeCCo6f5WLVaOKWBOs
0cvpOjK5V1acthFXBtB/8gJD39T0TzJR2zoD0jT8LwEkvlbySob96rYEy6lMjL0o
l9GHVB65tAgd1QxdNlTcYFR9N0AVDExQxzNW//SmmrhtVF3kqsqnaMHzw3nXlUap
HtNyqPmKsoCdOHhIz6WqZoIohbZwXMGkdKQufrDUVi1G0mnlDKi3vKz5scByPAGK
APTx47L7yerYXzziyb+UCLKvTQWuiQNvqFr0nQMA+OKy5X0lJmttpkY+5E2d9GfY
KXli0VV7ACTbeJbFeCkGrJoaeL4UfGWIbTVpGuQF88SBfcgbxbG2aKrv4OSykqmn
7ILhW+qHNExQdRZ2DlaZdF7QV3mKyhSqpw3MAExlkFlQCORhH6IB/0PktK9uHXLX
53KdsJUjfqDiqsc6uGyA4L2JWrUkbMV0UV2Zu7kxJXzA7Ozni/RRKwtjJxlyMMju
3DrYXJFlq0CCMNKtcnywdmmN/BVzv3JgjVqzEbGVv1Z2vpNF0PtXdXDCTTrTODMZ
bA+PRkFf/c39sY13GuC1ffuWSyYSnacGv2gmck58a3UgigL6QIbbvv2cWqEvRJVn
tBrZ/2u0xwMDuvalXYcVjP/S2VKjX8XFrFT6wrRPTy7msFZB7WVaf2oDTTPcdfPK
ZFr7pUjN1934ccGFFSwWRdKU5u8Fa9NMHIcjQuZDzyWnABXDCmfr4IHroTbZ8sRq
cRdcDepDdbkXoLgGWSKQqfs9f9GCHz2IavOW39VxfcMWDQQYIFBhtjlRJXkTWBVf
gTh9os3osvN+iWZ8zJSjff/NBUicGjhPyKKyR56m3ElzcNaH3YKeJ6QAf8FtUaPn
8kcHidIESd20HnxNIvZIulktAALhxzGGDajNl/DpToxX4plg1HekXhF3E7lJsQc9
6TpJv3T7+JO+eg+VofyZVsfjRpAlgZ92tbXxZxuzSvPeCOmR1+4940pAYlu/8KK1
c7lyzibZGkSs3OjKeKKQIRzPUTk/3hsGutezRa+iPjnzTiPrV2oiBY/bhxLi93Nv
UPmDs+yg8qiW0UQCv71v1FqxdKZf5MmaHhxy8LRxnhFP5vJFatHSiM9SFPzfi1FE
W/jczWsaG+tbMQBiRdBgs+FuUyC1r17cS7LDX80ME1vfVNHzERVK+e4xt+AY388J
GweV8u7v7Tl3T3A1wJiAB/Cwy+9C7z6Xsulv9uinWG+bC+ZLBJ5KWYR2pDn8lQEe
Rq+NUZAk+FnekKIxQJ9zgUtGocxzVGK3/7S7q0TEVaj8WE2t/LT6XpmiXJ37ovsB
75AxxwZPDr+slUS14/+OmuqrfWnDeZPCThR305zAemY8iYDJBUfbQUv6UDIdt/J0
GF6j2y5Raqq2jBgXJP+D6M1kY9vK1WzWDSpwsYLLCS/+hJ39P7C542ZGR0zVOk0F
p/DtBWBMPF94p6U7cyvJQ+zBgJzDb4k5XqBX9JzK262e5ds0bBAFPSW/fNfMR94G
jHU8RgK6B+oXU7TouwA55FUnjgACuqZIZDhBLWecnv+NjLMVULNxqjRyPVDOfBtc
pKpBE+OYvZoFzJt6OE0YtD5Lq4+0aBoJgRiHi86wJNpd6K8NrcMi2A7g9MuJ/PE2
/WFN/a9t1PX4PPnJDh2SccB733NljGM3IBkoZ2ferR2t/pDvmdprLSgsdvmiQC18
S745vceRLoUgSBpXeXubHzKs5nKznrfpOXHQIleFthnpEfSGOHSk2eymVhxDFeih
OdsVjLoEU3MBDzRHQSFkFclDOwCRKnY5yfloTj/+5MdzDabbJbL4NxKKlGbUvyGV
PHtEawTTFqgGf1/w/rRxuYvKDuxanrhfuh+8N9FqFQZmg/Ujkf7ThwT+c8a+oBpE
79w6Wl5nom64g4wMRCYg/cLPH1Bxl+JukMfZfm3ifX01ibdktaXKLWhCS+OkT8D/
zZRN4SLb1sGLjLHo+CRJ32oA6at8gr5HbC1Yrg+LiW1mCT5mlmDiGB4CoKgWB/Qd
dRxzH0VY9qPlaHbQnAx8eU8McAdr0tIJ1+kghTk5cfCoaOk/IvQdxj4tkmJpl1Et
PT6ULIsM1cCk7UC5mm4kgk1i946bkiP8es0SRRRbk7uC5fAsa9GllYEXqiuunOj0
S6xKtJhmsoS6VnnUNszw4CIHiYUg5DFhITlI/EVFrKl4q+85z5kUnsR7RkQk2kjU
ffUUteagstClxTWy8GyPxsLGvYM43RSZ0mRGc85LG9nxOhuakf3YtXqYdJyG2+EO
vK8jzgyvh4s8nfzy7Pf05aAYmmPPPohnDNeWIJhWxdwQtp4Q6R6mby1Hy+X0yEMP
HyfKmJce8tuihfoA4L8vsBraVwSb2wxRyBLnQ3hwFX5HulG2XB0cqkQW53RRSYuI
Wi0QsmGxnrC8DwqGzwHNdxOGeKjLOqy0wc8eni794sVrkIo3WSShIbKS6e+zVTi9
S7P1XLvE8bZT0sWucOLVAz2/ljkkZdBxnbGdEscn+ptyWiOpBLjO96RXVMspU24W
mgwyrwM1GRGrsAk4r9viPO3U7+Zm69aPbfgk1R5LFP4rXwV+uP9jbtVQlX0fA3ka
m8nuDBUtRcGdO2p9qn2RW+f2rYiKersQrYtB1/W3mU/uTmh7vTva2YEHR8KA6LUy
9Mdxi0Jt4TzNNtchvZdl18q+x04eLr8SFC9qNF7Q4SLYZtgw/LPXsiaA6VeO+5Ej
SVt9jAxpjV5tZ8+CemIKzScpp7BrgMlGZlZ8+nqDPnKsa2TL7rzBoxCm9M36+3a9
hagjzGH8cjfhcskd/WyXSYFwttARqIEYIntpGUrSsBuJXy+GkmoyJ1GPKmFmXyga
GQFhOY7Z6xRyeeYC6ae6tzPR138KdEugQjy2iLm0lX0LZpVFizSWiJ+j+zEzvOH8
JtSb7hNcEWtbzJCjfuK09Lmj5/nbDn71IpfPJcinhDvr1LievSZ7BxJQyHObGX8O
Vjyf3Nzp0TIPsEo89qNp5pwOs+DIkrvM5+e6QFlo+V82OALPvIFy1W7YoM+Uxlbj
uL5HuSaoeIJtfobTmv7YXv/dBiXhqtTZK8CSto7zZeXWqEgI2KDfpVQu7QFeA+m7
jbllFMoL08VJVqt/gpxESgrF7mKdgs1OnzFt39HQDpMMsxUwO6mVu8eSuqdWxT9+
/djkdLzDUeMQyphKH94hWQgNNlEhHhvi1YP6ryGvtiRyDUGScjOiH7Fu9qJrlYPH
RsVM9WL331Zx393phMD9rdNwpjxumJoTFPaHH+wnYbVQw67qHyA1w0eQT3kkWno6
hLiYugx6WoQa4k3C7PLY3u/Oeh8kuhYJ7lU8NotDjJhNv44xzMNpk8FIQO8RS1SC
2WByx8SMBUsvOOSwuZN8Q2+XWUVDm8sP9xzYrmzV64bZyU2PuBMcVNKKa3m/G9Rg
LqGzEfiyoN0DV+u2jhHVH+F6b4pACo30lC9kq95sT1WaBrAx51DzNlUt20d8/16n
62wVpDHZg71ziMo3V64jQsLIeHaV82gZLoRq45Q86C27ElZb+FuBCADegX7B7hKf
uzXIIamNqRyRzSqj/CPw7IEFV8mvFwRnNYo1hD9YBD9LBTIEceWafcLyOOG+btXf
8RXROXxbRBx4X8O/Jz5uvZhuJIoudRPO7FHwGsaLNCFpAAbKh5FxbdwAU+2kjFbH
+/7RoWEw5iR4OHp9ieFuLv4nfjV+edZ2g3TjHQno0P9zPZrGYqTjJ4FQe+vxMzBu
hDpyExI1foHvFW5mSMG8NtAJ8mYcXezOLzCX3Leedgctau4y5Romv5GbwntchDBs
YmPVVEM8SyBaAKCQt2IvQG7TI2S2G01nSa0u1G48YFCL0ILPK/wS5H5sO6DLJEM0
xjDk0W+K1KPRFs6cjWy5+mLfYn2TN8FR7aek2CzAprM9X/pOLPkWfS5XWrSTCZdL
mR5ahC/uAvpbeviny7oPtq9N3cib4Ks3dNZtY1R486syFK8C5IhjKsVwjx+/lA2/
ya69vqioQ/uJsb8wFtaptYoxU5VEka9BbElwmkG0S3Kj1HxAm4UtoEmotosPseVB
Oon3AR9cc3p2aKYgZrYQYFdL9paZjExuBobab8aNSiAlhGfOU5HPx0iXJatcxDuD
LUztb3XXbCxcfuhrKNtO8eYnsGz0p+R2/bU4y91wq8NwHVE11ugH7uPkbJfNdjMi
66qZ6JsxkNNLVeVJFarW0cT+nsWGQXmMQ+5J5/GlYR0IEbVAc5Ug8koo/Vln0dzF
GY0Q1DkJjXZx/OX07NL2ZCuB74XpBZoPCm3VoGZqUBcFOWcXQGSd+flC1H/VSsAD
eXobTL84Pw9Foi11VC5BVIiXDUVzYafHz9dto9FKOJl94HKXpI8c3WBrz2n1j9I2
UOOCI6coM0hGQViIksEsU1Dnt6zBpN/1qkevmbdSxInLYkzArHT2aBwPBI1wAED+
iyzaV3nDbPGQMgNDemWsupW4s6gXSof7D0+TI2qw4AGG+eXtCenAWLb3s9RJ9MXU
DEXyAWHXCPtbQrSXDNBpBF0ilDmyjwflcLt+GViS9akhjerMbj0PUiVUHVunxW/r
M+Ew2efmMe1cJwOfeHMp8mezdw3iDTxdjkbteHPkXs1uELdWGwn5kk7Kc8lvuiLk
UdyM359E018UNVXVf36K8PM15zc6XdQHxOwaLvgPX7wqw+lBMg+WJpt2kUwsKbNJ
s5fxZReVT5jF7CsN7nsF+XcU8Y5fvaIQEXcIIBEMAxPiJHVJnJ32x7XtNVKn/e00
jbnxuJaQG22E4oQ5liwCHzKqP7FDGqX7BD0xmmlJ6s7SokWskt5UMgbLybsPVpiK
D/rGW+k0E24Ykcz5WFrQpdf6sT/MehSTGSy0uLPFbykI7hq9E2QBaItAupuxHjFS
oWm9StZJdyZv9KsKFEW8cFJYBZ/SXuX8lxq4LWPbe708G152L/Mc2iePzaooar/Q
E/q6c3hFHr2cNINdKH+pHWkhEvm117rmrwQUyqH4gZloeFq2Ewo9jom5xsoGz0kV
HgibxH3+2tK+9Cvvv/R+VP9uhXhizBJ7v+zNQfqclLq9cCqKDy6VcuAVAqAx/MT+
epi6dWpsItpGLlkMl25fu+45pnIB0Km/bJaShIW+fInjrkK4DgsBcPx+YaWWbN7/
Q9KLZLmLSnTVl8z9NQ2Rrrb1CBPyrNDbFfxAeArJesWYJiyLb1nw+6xHVrrH9oNq
faKbQ49dOVZOcanWOK9G7yJCC3MCp4qMvJjPy9QeABfx8v8zupU+z0jZ4jFeEFcq
VirujkzhXKoHB/JtKLC9RqTbukOH+0zdUx/zceRfD1Vy3OyJLueWlGirkCWUNL0L
kDRpb/OD5OFu9DyWitjShrF7+CO77rrDncrsQYNf9YGtrAklXGv0+x4o1Il3puG3
LbtedwwuqVPhlU42RePJ2ElfibyhHoIC+B9DtmHI/MG6Gnj21l7WDoVs2F/yDcX6
T+k/ZlGdmNltkngEkWI0VPw2A4JoG+lVHIMvxKrCpDUDQzKStZqa+7V0T25juuRq
znCl+cAxa4my1wOY5fX6xlQxMAbSXKW2MvTrFLG4+PKXIPxWxCsAtKkoyOxpMIIm
f+O8LSjv1icKzcEW1ivGO6WP+Wkk3Tv15phb+eVSl3ZjA+pydL+cTzmVALldwelH
2DiswIQtBQy0EIbRmYuq1VT4TWMSNuPq/B8AzQ3jEEm6scljF61IpMNa3Jtmv5gj
fE9qdbpDRWtisyDRlLi/XWKth+A9jtjbYQWcbIlAJS6LumEo+AUvg3PYXuKFOtfv
HHI6Hl04X3EYxh/sUX+gQmFcuLT/1bCkbxonTaYlPX8FJdENMitovS3R2Rm819/o
QPiF7vpVfJGdqk5E3KA8Xlp+Z9DTs8KHQXfLSviUjBKp9y9pkW7s/GXWaG92w6hd
avY6KFMkrwCyblUSuP0zEgDlyvz1ikncCdMyU9Cy2RjX+QxDSQRCrCeZKv1LcVnN
R5wJmDNgYNtS5Tf1kA3sgnYrLj0T8+ArprNVk58AQc2zF6ECem+jrQDYh98XVNO6
4/8fau+dq3muyoyhJtvBMPLhFqsIlQz1aNINSlU8nMt6gImlmwJS24ZjWiwc5kLL
U+uvxiGf4wu+RzR84xKtKekkLk3Kvzd+H6xcritIJ6Gg64j3Q6npHyow6cRIm4yV
ONOsIkYSeP1T8KnIs4qFpIRXbptZcKIMQWuk2Mo9nN9jlLYNVXeqVssNy7lnjYcB
wqrl+TuYejuC+yhYzfg6xl7FncOLuV6tzIC3C7zYgRby+MTM5A8cIZWS1QW5mcww
Y3NkXDroWu7I8tBBJhpThbafSMlCTjh4SXaCnTLJJt3zdB7hhaAdyCGuIdYNq7cC
AgfaeU39YjTAH0u0sDCy1zUPkPJdfqhkZifzkzisM711vzBzemJzM835cMAjOk3O
A4NHIZ9VEDcNvimE/EKKWV56QvJwYNkzvo7dAZEncd+Y1nE2vdoCpqOLUNiEUcEq
LeriNcJwkECFM85Bvc2ZpKgZFdia6vhB97D5SWCPWn0B7k0gWi54gqPkBT30BahE
wL4X1GL3+aU/xV8hOQPLN1af48nfckxDrjyEwytVv+7Q+sUj3DhtSke6SMBWmnge
dHRx0Bu03qN8Ebrf5Pl7W0s4IUxu2ODcU+CbL5/TBVXPzi0X2JKWbU0n6E/QXi1Z
jRoiY88G8YLyu9mWLodQQcyB/2R00juOPPJll2ae1gTch5GuZkjo9yc7reRhOIkv
+t2TCe0DBcU7NFFPlZ6r+zMEek/UFpz2wBSIqoVYhR1Hb15BvMgB+yVT1uCDSQs/
uO184CwmmcwA6nU1y3oryo4+65VMFPW25Xz9hmmJKByB/JcyI2Ung9LrXygc7o2X
KAWSg4UOlU2jXv0NP2OQFV2z0zIlNYUttEK4N1G+WSMLMacckGj7/Q04fOT1u8eB
3JJHjzMnM+lsg4JnmDBP5g3sNxi+ZjSKwxjVUkLEM4kStS2XJXhlzxuAwio6Vja8
1MndlFtJjJ3Ww7tSj2Db4/0BHhP8kVty4hMWpidmyQhEtGNG5SZk2CZEJg1H/XTV
8zXLln1RTNeYTHhn+9h1ZwoJBcz7K7Wfaj52d/2yTbrztBxdmMEpO/ixA7a5xQ1N
dvmZ4icTWyOIV89jIunuqR+SuQvUYr6MQ3uUrWbprLXqZ/r8FR/X+35NBmpfsXSR
ASKSMAVKgNoU5X66NpKOmRMyXZt1dZ5Gk3a5PCB15wx9WQOm1oJcOoNEGYcAIc0V
9WeO/aa3k4B1Q5TW72X4+DmRHVQPhhRepr+v7gH9dgjFhgMWhqZ+BXvFJCG2k65V
7XguP67XjMG7XmRroTpRDfxSDLXdpBGNhvlODr1nGJnkPOk/sj+GogT5+FLgt9gl
IpG/In1i/dZ4bX0e7o5JQ7ckJU4BwUdKHXPvdwRRNdgbiU57iuBMe8CsZw6kT4Tf
Am2VoCT25zKGUhz4vHdHOysZmGtriEQzTl91gJF7+fm7BvJWgBYDfzGabJGzYrKY
3FWoiaWi3OZb5iUSWKTlIAEfT0S8OmRGrI0wWEcx6+7b1tqJRF21n4jjnS0q+azs
s+1aknF6lmFlw+3rXDxxcMwkWbedkQXrQoGzkZKORrVYNuwHM0/iZQBVYcvE7/Lc
iGkJHg865dP1mPTcgAWPURdILwmS+FgmAE5MtEszPdnecV8cx0YYdFi2FG68tWe5
mTVdv97kAxzpMhL4ZMuLKMIl6VuBsgCp6ET8deVI+kU43WnKsmuM1K6t9b/UMV9G
8I5f3jTRLRil2+wjDDefYsCHUF7s/+n3vTlzwY9/5aMMz0+zgVct7CgVtZguZahV
OT8e8DpUfdbvjVV+xqBAKd74v2UMUKInfACZC0NhojMv8F8D87S52jhTjclPFPX4
+yT989+oBnFHxp3g6LoWrfkAib4wLZFCuLfUsd4ajgQfZY7RfumB+lA4AMV6V73R
/N/KavNQ066kKJZ80uIhdUh8UfWwjf4B4So7DWtB/RK/KXtx1YgmYVWQV4I8gpi/
MZAzmEAoT+jTG+N1Jt09kSGkAFD+OnTW7h7tnotfcXkGTBB0SPrr0i69YiakqDpj
GAqOjpqI+JjrHL2Gv9ApM3/AZDItNY+cWy/PqcgCaPpvC6hbsUvPETCMTCnBTDOe
bP/ELEnM9/GCaUwuxBxOuzDI3XwcZZDY/YINNnc9VBizYGEQYD2sAef5kpkekWmV
QWSZ0daYTCnoIxUBrDrdz7RSRA0SiuuD2apw72Zcj70WQDn8EmcaYA/fV4GAwnCS
uosUR1okuGyChgwpGfRn2UvTS6UgyclwAj9HKX+tv1xHUbQqCGLbzS7at9itobKd
QUEdr/W/kBKT6JNSVMigBoyaRZqTpihfGY/JgFSs3Qd8kScIFhd09QNxnaAtuqKH
3gOriHNaHxsGH2s4xRLS1P90tU9jRZhOXbbf2RZJOyvSEe1WziEpwiTmcInJQ17b
X7Z7NuGkA3Nr6yfSzTTLhfLhTF03Nr+SIjkSqP3pVz7VpuMRCJzlX4PWDLCZ1Ecx
znoYQsscdOiL3Fn8Udf6RY+rnoUiNWMSMa5EtKhXHhBMOeid4PbbotRVhQJ3Nd6/
oqtV0BqGr+eT19sOGYjI+Hr3+Z3FzU2KlwVFUD+D6xv3gdhH8GfYbjDu1qmmtx0n
RLLgqaZxu1W7oEHoX8YR5Dd5WaDFgB8MbvCHJDPsii6gsyXFEmK6Qc8Li2hqYdtk
ZWrhE1Su/BYdkhM3lvbu/W/HJliRIo+ceRAJTujl5vz26T4HPJ8F0HlLGXr+OZZi
TjaEn+5FPvhcm923D3pi7LKT6unfR9skQ3MZLq3m/A1bD7OOfKsUpMWgHJUAd36a
evlcrR41tpEWmAeHRxh3tSWkMKP1xCiar058yAaGlSbamAYyliAJtlYLZVvYABi2
daLXim5Wz/TfmgrSeSsIdbl4jmvwLFfdsOeLyCPeeLtzKDHqRpNCPb9nChnH3zvA
x/CwA6deVRbbHoBmMeRPH6SGmXtKwGRIc+B/UqAQk9UEF2L1BBGga9mTlzaY/KAW
fy6TnxHxgfg83yAAOOuGN+wATEtLBVxWxkmtlIODPg5r2VQMLgOewSM3hKcfoZ/u
7ic06kKSoX966X+r62QyfhYLGrRlT67mo9GBkNGdlEgm3LdxVHijjFVPrAquu9Jj
Eum3llR5oEswBeCyruA5ws3LkO5Q3M3T6ts4xrsWIq3hqPv7I2IfXUuBzSaE76Nq
E0yERbAio8CdACvG6ltN0d8iuTgdK5CuVvJ+doVtucYM21yHbwb3vXFEPN8mPEJW
KP2MHn4R6LOHtlqSArZ/dqt5X7Rm/na1lJefiYTn74L+CRqG+UWaJt+H5Yba3y1p
0+YeTlfnWsKbDIkF67CT1KL+3vgLFHzSrV8Ny0eUOQXWccJopQwDsQXf531tvZC6
avMt3JkHWtJnAt1vGDmbM2rwd2o0Ob0sUIY3dafUUkF93n+Z7bKhz1oQRXkDsemu
panX/HEwwPMV+Vdr/1pngzw0PVcEwAI/pE1q5/7so++aen2VkXd1OrVmHB+NawRt
DxwVcWulLDsK2Av3nfsbf3bIfmWFjrKCSL//yZzm+2Q+eYZRZZ+w7BGCfmVQSlRM
m/sHWeSrvpy2Uo8d26j+ZDVOolKxxhjrpInON0XII55YK7H6sbW77fQ0LsDhqEi9
0ttEoeV9SlBzM69pgzv6uOJElhDeyKjzoIpf2iq8vWUoSPh08rNfCLPS0HlpttLh
Z8i3vA4CwKEzlaMfmkhWHdXhxRdiFYcmDSKa/SLQcOZLcwrlrHk+476T23GkPZa/
hRzWpPMKFN/2pexuuHLtoGZo/8fUxs68yFDcEJGK1UQNHHXQ/KQ+PAqIQslT3RQc
OmZ/rLrmWDG74fU+Otb6BtwvRj52vxq3X1o1HJPsxSlt+PtObPuu3E6fsM2mEqnE
5qlfi2PcKigE//nx7VgJJczKdDSeTUaEKIwDFQ1iQIGx1ZLtaSMUjI/u57VbpGrp
qh3579syl4+G/KR4Buq1pmcj9uvShGYa6hB5I7JQhmKjbp7JCiHDM9iTBYJsQGiU
JEan4IJaZjpkdQ/t8waWZfECWHRCt7Q8a7CYJRonQomWfi6w1pGCRUcTYK5CdOuv
RppFUbsR//bqOMIH1pHi8zxlQOnkNqgQlmaRIfMBNEivkut4RHBEeBg7xVTTGRly
lBFZiwyW5c7FRX9wWcn6wlNWwa2usDXebSW03CAlbRAypgrc4G+oSYyZXTcINeHI
2rMSLn/RbSjFcnfnnNQdNh5IGhlFbTXoajfXKWuxaIRzsIb4ZP3X/FYFNro2FqEF
04cM1B/4X4fXpMF5SPhGq6cEpkx/upkffg0YxZDyW9wSuam3FGMcPrTMyad9OVsR
jfd8I7OxIGoZzFwo6SYsp0Ywa4+3gog1N2xcpbZMXbi1OES+SrbKOTJWt/SaeoDj
h+j3WNf6nfUqWzxY1WTjgV6WabR2orsofts8SPJXc2/9FrkCY7b5AxVKGz96ymV3
UU3j6843WnfWBSTQSRWZ9q80n4hxns2TbHMvlU9KGI/782JgWFAtLE+BkTvugji9
wfnRJCoiuhLLveAx2lj9tNuHRR3hkxJvXwzdrWaNYAxiAFIPiy4KVgAX4WmD4Hv0
al5UFsO/zAWzPl9tOWcsyUM+2sd9QiFu6b6SsJrVQAbpPPYJiuXy6rFeXNafx/FB
RC38I0AbjrHwo67acfG9DS0dlmybDz4DYB4Pjhp2nXZ/8OrvCURzkGsoEjADTCjh
wMcogLWrNbGIw3OFskG7vA9LTP8s+whOdizcs1g1GLvqDL4CH87j/w590asVvjTP
FB/37axOX3IORUIw3Q1xKM3yVUOQNuwuIZxfBqe6ZLPhODhzWL3HLINyNx/eVVhz
PBTKSpcDMrnWoL21TfC1jcYBewDMZnYRue+lzSQtNpSYJ48P7XmfCl+BlH/XFwz6
S1BZK3jrhKjtxXHLolNia+4FvUX76pAAiD7gkM5B9E9p54yf1PxMpjNIRi1qXhZR
0Raf0Ts06GYaJwkATTn3y/s5bkhP126TvTpIu4IYtuHPjbnf20gl49/wNuImDMj5
ebRh3xBBGksVunRQ1QHO+Hr8grNCeQ8N4YXECUSj2ClghGk4zRc5fmGztf3F3R+T
Vui2RwWANodcfLKdiQlnYTZee/OEJJXiQVxvUbNOvYAoCB5Kz3c/9gEytKxp0vR8
KIqJ1+1qa8gjG0l4ddco3Jr8oL0VSSrlhzoT+3RO9Dt+RXjGDtVFW9Aab/jOt9r8
JD1h4txlBrHyj50PobO50PXvrliGfpJThY4qyByhwChJ+/joFBp35oZWwZ+7q9nM
fUR0F+WGrSgfEwLXQCPp3F4Jn6OCzslNgnSN3IxFW3HLpTDgOJrxJRAEn6X8fT+F
EH6a0q+EbXRhyTHwwVkRQY+7MIkhVvjp75JKLeDCWMWT1PT3KnbVmcBWOV8vMjvT
1VxUciX+9ShD0CcrmEaJHMVoZovXCbUfdGn8PNqH+hh92Pqu2qXNyrF3mT0ZlGSf
35uUUzOy8pIlX6C+j4tJw4sj5ZeQhBtqZH50PZOTWzrteoBCZOl4CcJiVQ72ESsQ
/TylamQ2NIQls7gzpH5zBF1zpX9lE7+s1573frHJDApr7xVBuD85L7hI9TzBushA
BYA/2eSElaEkFaXrKQn+h0z6oUMNoEOGO/DiECrBf1QxiAWArwpF45SFN1/lnUzs
AwlI7MhAdcbTF6IpgiOPDZoXO34FCl0fhGjPoKZIC/bB77ULfkfiCEkFJWFb1nIU
KT91XnL4vy+OxHhEryzuBT1tl2iDQhn7auz9/g3OV4jRTeZ5h/6oYe7QKzwL5Tj1
JuyqtpunPTum9xgl7PycEreL0sI7HCN3U/I2VOtTctQFLDG+UcWUnReCOgbYgrlo
nQw2VZCU1tqCZZE6pFYPaLzHw2tT1kAj3s8Snz0+kNcBqig/7rW+zWyqzgEsQxcS
/qInwMP8MRmOulmm1lShPMRdm+v7hi2FxXPipS9jXZBG28vTlJEhXd1MkUQFFQMw
qUDjNR84uEULpTe6pw13x+GK9tV7XobaIaRxcmWTPOyOF/CyXkXdBstJRYaUJS0H
nw4K7SXDDK+WU4NDooKrviM5BFwmQLtuau+ZA0cqyzJETW1XKkqOPJ69JmEhPFj0
vlNAr1h2wRZz7aTFvgBHZ6py0e+NnRZt8zsJRGOHtH4c8aKNjZNiL2MWwrV3+bYU
Z5Iz+V9bgMerA5MAQxz4kPQ0uQiMkZoyxxODSaejZ/VEVXR7MA5RaTNSUBWZwIdR
B0hSX+Z71E9JQYCd+FMpJRYaop3ANQPBIXzQ20uL0OC+y63qYiblXeyDiu046QO6
MzDDu2geYoXOX0HKmO4F1YM0yW+b0gprkrM4hDI6Xsjh7IArlRqpT5k2P5UXJ4yU
0+8KHApTUatZuwM+bLm7Og8myFSGdIlLukFwphs6Sp7++6q2DEFbfLUXkBK7FORg
AOpgcCmzr8n92Vxsj0xiLI7jr71GdQewVGH2VI51mOP2fXYNaBxW4G62G4pn4p8W
yHAcPgqXi4JXM419zffuDnn15B51B+Zu7OkjDPXfbRDCInevuk9D4vyMQxq6GX3z
PLCZS5KldJZ/ALjU5sQYucCm+/7MAyOULLIF8u4YupZawTtist8nNu17M81Qw7vO
BkcqMoF9n9oAPM1fy1aLDb8mFUlhALXsvshEJsDaRybOFu5ASVy/RSWqygD8/SJR
RzhWyWoLb5sOcvRgNEEcnNuejQo2/1r8FNBsNaol/Vxjb1cewB1E5xhJsNCBB83S
vTeSF5uVu2bVR6NpGwKGElpx4DCjysAkCxIJ0xh+r8BP4jr+TZ0cOkaoQQ3Xptz2
K60x9qSU+WR01ptUONbZvfIZCPJGVklkS3SWDeXoOh5BqO+YYKk/MJ6oBZJ7yhx4
hiKpoAgLNjyGniacobid+8XUMg8EC5wOR9yEfQpHUnbj/6rzOkli1cfeLDbn0nO6
Fwubw669SMeN7Xx9xVjoxNNI5HQ9UwtRSKnH33DJFcnVOh3DbiTneCUQXH5C65wR
etK2Y6pg3hRLeO9Pmiqog7+AHACfjB/nM1skpzYAxuGdmK+aUt6ZgOpWiPMBMbBr
bJaQJMWkiNooCRVNzleAdTC2A6QgywE/zfaRAJ4ZieWo2anVZW8DfQBnsdehA/ti
FvBP+LWDE9rrw9xmhuOt0itR2cVu1oG19xbPWQ/idvA37oD3U1qvrS1TwKYoFRhU
VoHnJNMhavK5VN/3xz9UI69pn05hw2Tr4U1YqTQYh8bA+uvh2YRfBCIS++OWM+PH
UonwjdPaAM1wOt177m/+hIHny6QG99Pguck4YW5Bajq4klMGmNnm87V7OjBEI6AR
aZE57zskrXqGV0byKmT0U0VvlfHU9A6Xlq2iTpawb/cBOwJ/kgTWjQNmYDXO+SJL
dKCDMlc3I7dN6cb5a0eYZqvJVuHMAo+5d8RMb2m9GOMCTgurG3mPGnNFOj/QJ2Ut
jtplOQHqBnngrTo1ZcPcINmYns7RDI4nld06efQ09qbjCo3rODRBYxb473JND8pO
jogOH6xeSue/JfzIxfjzRemhTr5C9x/7RIw76pwqjmAMedxB54YSFewuWFfFj3Qz
xPoPfxIavQA5YMTNEZ5COhRmqkJrk8yVLmQzt1VwOcsjKGV56EoTGpH8Su+rKub/
5M1jFwzspsAETjMO99Zpkv3VSuETzB/7O9Pr8fIlm8RJYDjQNgIGZuJLtst7WBoh
siUTW1Gh2ljlYbojMHNqu5FDVcevq3ZWgWVdSr6VJyEAAUnJRBoPzJkgAVBHHOyU
llq3J3fIZ+XaTklG8jB2R1/Kqxno/SIGAR0WnOuIsPe4TzNe6kE6SQODUgsSwiY/
9u6TsV58RKJuu8crdJBItaUSuK6iivWW1+aL5XO0gs2ytneNMiamZCbtv+vwONJs
AJIZtORSdzpnWK4riC3X+4KG3+EHytcExY1ZAA94pRBghAsItea/eA+endYHX0EM
TlkNFQuzAcQR4xrKHYdS3CtSS9uuRourNeG6YtC7Bg0IzvPFnqFiO8lO+Kvj+E8q
zk4xoe+Osc3IwV9gsbdsU1Cc5G6YuZ1m7H1Z9CzL8f02n/dp264K3rjcgn7k9FaI
RqaqA3EzqmsXwPlDBJbHobJUlAdSiTdksQaUySKPQSiPX+nYUVEHGusvr9ZrHwRt
RMKdSSV+XjYAKnLk3Tf9RoVu9j26Z7GnJ+hsfZ9/qg9qfX3yOJDEj822EK0Z69ps
JkiZ4szJldOnR6SDHHdormTMxtoF90y0rrbl67rmk6b3ij4OaYEEpB73fsX03HVW
0fUvJv12a+BVw2+bOwVQH1P5hv9veoOuTLKd2iTCLKE+8Vuws/9hkRdH6sE8yuL3
IERIiNDa7jQxqv0v+64L3cNgDMddnPQIMzMbIIXVSUAksMSmha8ClVBpprbeIqiA
C1weVx6NccgsQEIB0QIdt3TzoYG2GLqzpWCEDok/YJtXTnq3CPnlRsntSwP/xmF/
KWtYp1BoPsGpS0cc//V3q7R99ByvgB8ZDD66+WER/PghL5iDuKvfAhb/X37uh5mn
E5GCZ7ddRMfIaPzXpTdcchJDu7WOPo8METZz2DB3MijT5imrjvnIT8k7m5lNVSrF
Ow4ndsKSoRTzJpKSfqQRBZywd8UvIxQkzQ/SMjBEMRTKWxbPm1xVWB37XteNoZXC
tugz8Hxsl59HniZ4KTjh3TfqacPZ9tH/9Bb92NWylXNc3oV7DKaDCSpeXA+d5xiS
Cf07pxegTx2rYHS7r2wJCTNp/IHiNBjWpXQuOcgtIFrNFlPX8Bm/HWCqXTO7b+Uh
+n3eS4ej/u7TG5YD5rGKE3mYoN6KcQFy8ubGUzpADcVYdd83aGTLTQ9uVKb3gKfQ
7bVv58Uzmwnupy2ZCfSFRkjjHh6RmC5IuxSfkY4HfY1smWQMHYwwWXdNX1VsDd+s
tfZSjw0dXVd1g7l8ESawsjoLScg3Ze2bEjyeW7DD1DoZvkyzzTEggeBvmOnqrqVL
i/jscpFoxMb2pTdRGimhNj3Z7MgAu/hm0miDJt4T1OFfkOsT1VHlYaRbLWmU4gUo
ctmBnIim4358dGLmQ1pgAhrCMql8At4CF/Mdjm7h0M6aE0AmDz6R+NX4TWDP21Z5
gUoz8udb7eDcVnVFBojBrabpG50cmZ4cZGxpKjNKsmd0RGlaTCnrXlYspN96CSgJ
KAqLSYNcLyqWwOpGT5MSUDNbC6fLTTKUBbs5ZbbRJhDPrrIPnkL+vmozh/I1kg50
eX47etBuV7+79sRM7C/BBSbrSii8sf+GquvIxobAJZ5kjkgEaF632GkCITIsI/uE
OI+EFSvMKWy9x0w88jJ1qvPkNbEy3JfzlLB2XcnVY8qexWovCuc4UgbE3uNvWplv
ceJrgEUYU8bPRojCqwSblqK5EsQ76hcEG5cjyKifhRcHWEr/pJqW+35paMAEOsKB
RbjRuMMZFKZ3kW36TcYrniBsEbmdiFN+n/BGH5CLiL25d2q+PoHfK2U80HGHRRui
oGDpJmpniGh4eiuZ1ofnMdHQMyzcPVtIq8udcqCJpMICevg4w8bYtPd1/Zbmjbyi
TCji/lYn2zQUryPOA0JDdCsO99KzIHxB7KpoP54Sf5/4vV7LxUYh471SI1Ytdn80
sFGGCkAIPKkhhgwh+t6EUrFlYhdPTGi8eh0Ol3Sh8IhNefFxtJ2GwFSc2HmNKUdc
ecMSDw8v0WgUDv48aEKMsDMmf9ltKHk0eOtrpkg4jrbDppAnl0Knx9s+A/sORlbK
vd1HxwWPOhgzEd66LnHNNzr8CN+OMpet1NFOiCjSH9hKHjH5uDY5xdK24opFRkDv
REO5PGb88VnqYtFBtSYkMP7SNNaHtdtS2c5vonHxv/VOmMfMZippqWmAQ/fJFDEX
wdpaUvmIIGXDG3aTC71di6QlBPjmmeGDpMS681JkDGG/WMqf8hfRU3qqMAX+WUem
m6mDrPzuzqPhonMR1tS5Lj52K2bSHytPfPWDQToiVCurrJ/xGMSv2+c+maMCsCW+
qLwLDhlQDLbu7Ci/k12kdLN+KFS9flyObfJP/RZ8kqS6pMxf0qs/s5NXa9gngRFN
nVGs6jv5TaTSp3cHgqx/JDoxhH7jexs+MvjeTv3NX5mpMo4vvBGLDN30nmsMEN+6
6+5bsPbmUv3xdiz9OVTv3XeJpSoxlsEEBY3maucDk8y1e6ewfsEQYhvo3HY+XBgS
sc9dM5pSMDu0hkG/edLzMDHx4WSuIIKMCFN1ns1Na0iZoqO+WkvUJC5cJKDNuov0
uVH0Ha7dAD+KimsEb32876DOM0smhWpcynA8fhjVgVtT2l2UoH06FPZ1VL524Xdr
BFRnSlu3rJ+eT0PLDsK13+46TDvwteFK/S0o/XssJaKIC07qHwyIm/srA8CO/FmC
tDQSk82PJf4EY5OuVCIfWxH2e6zLAuowJOYby6g7zMy8SYKQX+Dbt3PeR13tiq19
tvaIeoxxHGRhA4IvslnorpyRdYexDTVUYuHfczkgcgoBpTiPpaYCmVgAvel00AHN
xHJRIohJp89sip4l71k6U+THwaDqWgfHnK2P1EFc0ss6Ft+JZ1R3NAtrkXsUgfo/
Jdlvi9zU0ubAHa3//WryVn8zw9p59ZT5zaeQoSmoz3gVfkxdshD/Mql3aEwZHh9o
u1RBQGk6XxjwoB5Mh+C3JTuSUNXwQuDsc5UZq0OMojFAE8HLBEwKeBgqhyS2uRSd
KtnI14dmmCG8Rg9IkHYwRhFeiYHZR4LQUWQAS2KZbaA57Xs89KSE42vUCcYB+980
2jxPEvUjgQp85lVFp6nCwbMPHd14i06QbifKnrEJTVgFBoMmMYO/c40+yGkV+CSD
9xy61A21c99lNri0/EEfv1bREQXMpwG+YCeAsOH5X2UesC3IJqVroXpWdcRUAO+U
3ChfSYQBorlKnfNmhGBPuUZbW+K3oegqjA0TTAKQupp+W9ocl1vWckHcZa3SDDmC
wN0DblQXFf2LwPW1sGYYJmBnRw3nAAM3pYoBz+R+WY77UQSi0Y9aAdbV77BsmBBL
Od2avr1kA+mU+8zDkXLEevKwI+QPX6HjZMceY1ZXE6xuBOlW2tGv+BcEZbgXuvI0
xRuGTYzHnEJuuo/KPIzJZFnAX1ZUuMeymq/LRGqNe+KMrM5JUiZcemMce7wjxGN+
q+IaygOpTNnNQkN4/WiwBjefhkUaqWHY79oBDjIKWSux9E4ebPauVBnxn5qarVRK
n+wUp9IDMnNe63f2DpoGLsRm6S/hX5bycIJbOLDi0JAtCc8fJnJN3ocSnCA3XfT3
MZUQ5rWzoMmSRlYAinGVLqEzLn342UsuDc7yHcHLT9jJqxgl2h3urh54ylKVi8QC
9KO9pLRgi+BvRnF//bzbe8woAy6Er/B23XK6ANfxL1/vY7g2LtnypyvC/wEE70w8
W3DK6kX2UKOKNEFLmiBfkOtm3pLpXlarYTUSOrHyN1DMRxDglIFaug0HqrAPkB3t
+/g7Ts4B//FMNgnWm2O4a1RklHaa5FUcq0UTywot0rcQA5E6zrmGiHGhyCN4atuU
9wKWUTYO06/n1a/QX/pPqz8Ooqs24dQviaP+Sv5/TgrzSR5Kv17qFR8a3To3b1uw
gD5+XT2IjkF4fu0J1O6SufQpJnzYYVqSaBGr6+ajtVmMXk/a6g9jHw7tAQ8cYYLy
5WFxqOysveJYqSWtWe2mGSvsU0RO/Ejbf5udbNmnD8dtLvsEL94wDlA1z71sp/FL
p3Pi5Qqoy0LIhEvIEPISF4WJ1cwjt24H6e1fwf9U9VgHyM3gF62I8DRqTDymAYET
rpAaoe3BrVnMPq0h8jSmItq2vvKX1+PH4ZGZvpw+WHZTwnP7VTBFJXq5VlP0Sb4K
Sppf4r3j3+Ms31NdyHFu8sHMaQRGRxeEHyeVO8ZYHaqN/OUx0en9faYbBRciUcta
X7ShjLov7sRvwi5+sFGGLQeadZi0tF71q2n4BqxyXnaESOJfdrCkZ8xn++zl+6+W
PXULn7yDrttQ552xGLSG3jnrDmG793uNQ999nJLLLPdXZCkdUQu3hGpd2qFV1Ckz
kTGKjjs2YlnhImIjQD3o4opgAMkt7CXghOQFsQhTJbKd+QufTFjsXJp6PDGwcic/
5CGCH1N7/mZXdToEC2mULeuBRGzttO/v/L4rAMS05uGB88EPbnXmafbcf899U/93
RFvSSMoINKRK1cCiXLjmZRXJqE+epHi5jtxheD/bTG7NaIM7ddG3Y3f4yEk58Ssq
YvYNh5eLNu++oUYkMhG/0uutmWI5f2yZ3OmJGAZ3WFC1HWU1TXlNw3SmBTVtEks1
yK/ejfNAB0sEXuRMeNEg3o7QrraHXmtetVCAfTCz1P6b+R10rgiNmrYNwmx2SKqi
Zd3lguRn6jZhNJXKRHQEagkbvF6XV5MRbPd4Zy2Xd7/alfHxNKl5uFyLIuW72ZdU
aSuXNvev+iqwLCKs/SLLC4p4XCHBrgVdGmDvjEAtH4e+usmxWow6TEh+X20XTz+3
w9Da70AW068TeIpsYYzaYUAvo4zCCAprPvDb+TSD+E3Moitixlx+JmufW4/tLp4j
Qdzq3qBFHAhwbo3a3i0eW5Bj5Nbg7Vdv3/ORUSiZKDhBad9QZMVr8slcRFiZT/4H
rRPHZCKS3RjspOWO05TMCGs/48vBMQUQNtB0zR95OnGgByGNImIDzhn8DdksRhC2
9DpHC7ooVndpZhsmRoxywT+k4m84LFyCpyyONfOd7CYRecS+jr3+6ujg/IjcL0zH
YJZULpYLDgH6QHsI5mby20dqlFDIsAmHVXcbAAUjd9bJVvnpkD096Lzw93cK/ZC6
yX+kx94HNaZli+ZiuP3y+B4kwttkbSYNIqPGXdBQOkmBv1yiCB5lCAI+xzU7HaNW
7NIQVIs0tBbiXHcwhwofuiXfRzFYUKuE2M6OhUGfHk3bCZLh7rdayh5e3LWfhkW1
lP5s8uSRBRjD1O16xPlIgX16/DkZzeY8gMNUrgRK2Ffo/PhpvaWypdjEkea0cHAg
jgLXPxbAqtqwL36Qgjlll/oFzgF6hvM5msFUXX8dTg2XO6RzZu7CRdRbeg2UrvqV
t44EjVJwCuvDyUYayMgBqGyfTBpcJj0L8QlXHcbmFmDQOYz3kozTW+fAKJ7S3sg0
0lOOCXbUBGUQGYpAQF90YacrIzzqRUxKMs9IYVKzyPv8VptIANNGzSMCIV5hmTds
WY/K6Qx89RVXiFB91A/Nvmp7fICjiRO4TtTOkDiX9+k2Xg0CV2f8i8Q49CC+Cb2Z
HwAV27Z+Tu66tEWuC6U9B2BdJJF6dL1D7wBtpHGuvEFzZ8dzrrQ7RYkrr+C9xFiP
NHUYe+i6ViJolV53rbM9DFt4+c/4eFKSFsIG8rxiZa55JNlxscQdVNh5g4UQVHDi
7WvvNLMyXTAFj9Gy5gzKqu4EJycH/rG6R+OcN0hMErwwFYsSd8sVo25WMohEh08g
RCsxJIbFQedfE0amMAKG3DTv0yVJW3KnbeTG+tBwT1iAWrSbcanhcK278i4Yo3Cy
9UOoh96JcmOwy8GmQm+9F/ltEFiwcpwixYQvd2Bph87w3o/K7xvachR8OxHJ+rv4
2fvgqs06sm5N9UBUscdNWIFoGPLeM944/2mEP8r3qzyJzZLswxL/59tC5Af9WsRJ
rLwmE2AQ0aNE93HukkwvokP8L7ho5TqPRSQiIQPGmGAq/hnK7TCYZcJifVCp3ClQ
Z0oZJX1IAcN05we7dcMrWSIoC9gr2CcfeMv0uOThHFDd3lwcS8G6FjWMZfsquikG
Gd9aupBSP7lZXZegcfoProbqpCg2O/h6hhaSvwTzsMMj9WT8TmWFe4h/289+TN9c
VOlIMdobrq/w6LOIGeh1OAYu5kgTBkxFZtzObxU/ttmE0nz44fz24XAjR0iTz2vL
DX6W5FHM4R1q4BKyKzF4f0j0kZwVwT8tdKVBiPxfT8/tJ/GFHOvdA9OhOBzwrfTs
t4nQ2QCdxNntfgFLIpRkoCbq6SkKU3DL1e+kbr3z4VT9/I0bnDg3sb5BeaxAwqDH
hEaSgBUvgeOt1IgiWCCNxpP7ItR6k3HWlvSvgucJ9UvAC/RIoW7c3CKd1sNaxcq5
H4CMes3LLhvm7Dk9xxc11EsV+Xo2Kkj4jngFshc+lNKW5a5L+jQ9vq8pAtxYZjrY
pY9dXiA4g3Yv2Bp/MFayNzrF07ZeU2xjt2c92pYpZNyrTxaYFQvwOB2v4NMY6MKg
PDF7XQMgqOnDU7HSxKFAx1d9LOyDhO5kGyF1XkwdPjpD9iXGpiVSy0w8CTbTsY6w
2CtPlMNkAuQaqZsnyZDek+OYEGGpEYaic4jY7WzCXDXdE6n/5W8yz13rhjsEp7KQ
hhQ3GN+4ign+HyNW2bzlcMCiAcsSEPuZs44P8/nks+5ENXaeOD9GL/uD0/Gv70Wh
CFPXTrL7p/vZqggXE7TxLln6JJokOCAVsAjPze8fikOwO9KxBqnD0yzoDgoK1H4I
lpebRt1kocxdPjCQ/GZvt9r/fYL5PuPLgtkA/e63Z54H+lVX5oBlJxZc1iArge9v
+KOtdTRpConHWK/a3qqHmihB68CO5/DInVl/a5kTTytDjVE6yOsqymw411WruzFb
bIg1++kl6gkVSO7juygNmLIsQYHogKrwEpq1X80ZeZ71DfVs2kOnrEFKd/Bae0xT
IfrIAjSLigrp+YdwRqlnJfkwYMcrZ7EqzXZN4b+PgylvqQd03PpEtkYARhQkWrNA
eCqJxU+fHFUnZmvH/y5Vz6+7IzeGrTFxmmqfQxXAJfYdp/uv6RnS6BSVkmv7SkNR
C3anKLBBoHiU2/1yWFgbF8tRd4+u+gWarzDWkjYUOaBd1F5V7xPLYYyYwn/RkGKO
nS033dvHPc6wWc5lO58XjplnSnkG0y0BXenGKA9e69gGl8xIM4QG5Dchow2NDotU
7P/GnOObcvNbPJDHlILXFkMfU2InIvNDzW5/CpjNJgBrppPr3LdKjRZ8lSD351D3
JBc73c4aIFbZxY248MbQX2/S9InAUDGmygOHWZSpdMKfrsxYpuYWh/IGfOBL1NIU
UrR/bC1GknsLKJDgGtZcIvgR+bpiohN28CMftja/iUxY6d4+ksdDqMZEriFtcR9a
G4qW4+wIN25g2n8bjZ6v3yIsMpirPg/DUraOV2clv5VhvFnuu/Pergm3DyUW3vrw
YyWNo/eAME5uO19/pZjc6lZZE9DOSW7B75U6e7AMT4MCUb6gocQ48F968XNIcxM7
nQ1tgOdo1tcGjrz/jtnDXSi8FuaHPJOWf1bbZWJppRNQoDtgC1tejq6CCx79gbcp
cI04f5qAPlB73c3kxw8+KXWEeEfP85WKehDMHXaZdBaz7OtNJyPEKBD/b2S3aYsI
lYYQtmRFH8cIvgRjIJ6xGqMq9bwJOu7YmietSi5rkkCAzJlTeoGSFV/8KNP+LqQr
nkFaZb7VdtoT5EYwsorXQnRV0DSfu6MuTGP6nztEuCvFa0froF6nnfXpyie7NkDa
tNgwsA0NhosWIVqLWkOSabcUSX12HTJ+9UoTXmmU3WqGd33OAggx3YUS5w1kT3Pr
HPFBJ16InnFHSAljKzgne/+e+KkcuLAROtUHXqbpyZgNgd0qqHoNwdtp5hXNvLNA
2LdQKQFkrHTW7Hu8u48266taQVWlWSfDIyv4Ay2O7lEswg96SmF5DRYhhwMJJu2g
a6GAUiVTNrMp9bqtVu49Jna7mLlL7czcx5Rp+YlitxPLdAs0A4OAwi9FfU+VU4Cs
0NK4BLB6B0QjqjtTuwfY1HnTae9k286Q8D4RVY86EVV8pFG+osBtidfbPKfxmWpE
ah52wMvf4VHd16Pf+B715AxgvVmLOLe1h2iNWksseiylrZknlvrkocwh/I1TRZ8V
q8O22lqlm7ZjBgjCfcQUn9R5Q8jFoYukXE8Vy+TtE9j61JfWIVDJHooAPEcPtP9p
znD3bmH8pViTwFYi5+T79GCondVvboEvU6pdzwq5JL3yKx7z34xyUuOHt05k+084
t12ak/DrsgBF/E3926bea2YPCvwGkjq9MliiDnR/z7EH18/N0WVic/C0LiZDKFhs
Iexw1gsWnHKdgB+ufWrbi4MBsWLAhmW8k3lJ74hQYt3E6ijcjjKTnrsMRp2cKrNd
dXQatZGxkWyzCxFsxiX67MCysyJmwrh60cQdDaMOpI2XB/voUX2nHXNil9dM0WJI
yS354YvjgoapuHB1XOr5pkg9pCkS5CsYpsyC4BF6AtjkP+r69LgULTYYM/lszjxT
5fsXXUqr4bYClSywLxmoMhTVF5qgfxNtuMvyFWE9QEl0UCMbypZixR9MQ6yoVN6D
ciUXJzU7BsTOwwCxXPQzoLa7XpxEbYYhWbdPxdMHL6hRs1pF2okZWukal0ZMZn0j
AAikTfrzXt4d8eK/147sg+0KUJInZpz9/qRde3P/08nkoea05hffBlHrYwX1rs+r
roEqpK+nxOfxbxZutebJNqSlKq5zvYVGOMJTIbkVtjD4niPlVQ7bhmsm0qRSojpm
HjOs/gvxX+TlJm7JpBKgBh5gnYRbWsSDrw6OIIVPRXxLi3gUvpxrS/z8wVYh1F5C
VNyYv/qvqBkqxrriapvO0rcYgOoKgqVFSLOKzr4nURRRKoCsvcURjeVG6lWJYACe
f8GPCI33O3K/M/YF4oRm20JW64lNf9GEunzETvYaF+/GAIm17qDtBqrY5vF13sF+
A1f6IJpT3UYnjCo7HKUT+KLSN/hPTnywPqVok6+lxeIPp5qd138b4lPBkqNptf5h
4OvIa0LHdbf0/Kc8C+6mlRqXgca3ziMXq/BwmtCSwX0qfDWv7tF2SIzWWTHtTfdf
SwcO3uE6HY3v9FycIqA0Jo03FP9wY/9yiJyFWyXly2ZAaSXkF8xoj5SLFTPq+JEZ
C2v144pM5tS9B7z5Fw2Cvpupp4fXJg6gXmOzw5SA32VfJx8NmbdE+rD33UNPKhDn
g2YodG7KRhA4c+dGy+inldOmSHAFQC3IvZgPjutlI2+DDPJHhyoUQElFnV23x6RZ
ZdECJKZmAuIHv8DXndDNJKq6lKBHctKB/4/ut8ifO+LLha/GMgp5Elpa69DGLpe5
78TWDUibZoly/6WGfmiSMGdyN/bExzwYjnPb2ItqIC9uOruHdY9lVWPo5txMoVmk
xfDcG3avCxn3ofOm2HOvDNJ0qsP9bIAZXHgDzch72r3e4ZQryKtHSY8SQZYW2QuC
jlJNmAnS43gg20Gxn+c6qzLipD4teEBTjP5E24BOqZSHNzOhrVtgNSumpRJ6/6Fg
UMgLOeNmse+1e9oOgT6EMPTSCRmYKfeBc9MlS1uJ53geRNyJmlprEa8bnJxsz6uD
Lq9ZTDAJOBPlkUdJyy9U/kV3zmfEvX43Hl+wGCt5VzO4gRWhueovREAgJZ5kExFl
WCycBclgNlqplnSILiJVBgo2mckdGJ026k+oKrWI3i3f8le0oCiMIrBPrEaLaFy4
vUuPORVWtMZh9VQcpsads9ILeG31FVvwhWYH40CVmXUemGObia7yEmSX8QOoIath
CS3i61hklpwI12lfGTaA3wTw69zi7MGfjBmtA2Z1VKnslZvyx3usQsa5Lgu+kuvL
jrLcrVWPAfhcp1owPExBiBMhLSYm5t4SGVba5ShUqS6C+Z1l1Xd/fs0ZwS7O9Sw8
hI3/jF9UbLIrC+G1mp723kWhqo2WQSGCriIMIu0BGlNBkfWZmFasgEAN0eenvl+5
BapJ30CBHQAEeoX0uupU9j6Dm47DQ8pQ4DKtFbhPEAqdkNufHP4WQCgoqusoEXae
+BGyakQwswtuJzF/+xTIbacULa6+vF3f01nK5LK0RYFNfDSojivGYyoMVkY1v86v
6Gc55alzIcq2GkEVBqevpkNHrpOBKb2mB0WBNRaeVcx4QCdO2rKlHF/PkAGzVXj4
W2zac8J9Bgwxy8cgC0Vtju5zddVk91Yq0W2Py9q/w/rUZS/vGSDZqt2sXZs69QuZ
0mzk6oqJl7B4JrYt0x+fiXsxu7yltUsME7pBu2zV3cwz9TTV221soNnh0FwOyxjN
UvcIZjYUda2n/INNjFeph9Ss0xmqI4OUKJO7lZqX0qMLyBjAStQGYKEBQaT78sCQ
ynMmDN7V5oLBF0aTLpjD7UPWf1rpCmG4KhRxOl4ACeMSze4rfAwX/GA7/0y2kAD9
Qs1+yCYnIRlwNNpVqpy+UkPkhv5rntS0t+s767uqTKQHGQfAw0ivSAuf/tOrHKhk
DfkHP8gc44G5aEVhSTKyw6PNbVvN1KDxKYr/8qrleMG/DJ/QZ1VUR+dIZaq8RgjR
h5klOtjN2I50UPRtR24ycHunSDw8J/RsTjGykVdh10WPVMFwpEcTTGzsJSrdUNYY
aG4HtGcbpmCC8MIJniphcX3T0O9cuX2UVngWzhHFfHniq/7kAtMX+UcKa7nvpabw
GNq9/LUX9JErgRgbIqo7xJ0FuhC6TSOodhpSOthftdDxGgsGXj6BZz3LXlw5XkTQ
kOCXLVGeuIW6HFebG3gDzSjwTgmAyVinDqEddTu0YbfddJixHBPJns22JGlMTSpR
0sQ98ASsjMrAOswoh5xT3SV+88A+yVRczqU51SRrBOP77OiUbqf/P6HZ0RUGAt22
mUlLwAyDpyyFXI/Jr5rG5qn2hgZjGQk6bSCUiEkkGVqvkRYcfCQG8Ljhddzm+Yed
BNKb8rngiwtsg0tm9E4YdmRsb1lc98l9QZ3pZdX7s7GvXv7Nk8frq0Uy3ixIksU5
TuHxsTplDB4yvDvw6r7VrA6PpZIole5lrAKzwUWp286hxnnKpNfzdqVBgs1zER6o
OadVrue3tGap/Nc3LbqOZazRNsAFVqTgCRWuwhHoC/OWCG/IMhQVAhl5DRxIYf2X
LGLljJZ2564CLZNdj4Nd7a/VefLiJBMKG7WtZ97Iwu96IfyrHWrobq5zdpoLrqcc
QIlgd+CPLZ63ICUU/3Uf7A9/fCOtCN+DdZjqdD/+oFfXY5hA1NFc6aa8eTl0R0Mv
MYu6KJAhDG6jbVBxx66oBTXGpqcLHywzvWUU4zNwAO3JuF0DX4DeobQzfWOfuTy0
/K6kX/4wsVNt6dCSX7T4y7XyONrfn03GyFdUSCZXVDHN5NVO6UICXxdmKYu2moZh
gLptsrpywjrS9PZH1y0N4PXOLGTHbl2EaHHHMsyHcGW3I23pC9zCDPbin6xHM35v
mAdom7mQljUp3P+YXTyMPA6M2v3xDWpjNh4Yob/LWmZJfXUVD2uLV752k6sMeheH
a2R4J0EijkZEzZ+ZZkm7rCaP8m7j4qpsm9uevNm6Mqq4EANIhe6MzEvRNbH/Bmci
w9Vr8RRnpNgGfF0OPN7XucspB0e5rYHg/kf/AtevWuL9HwXjorelUvKbNJFvmtjT
QDoCZXZkPYZR8/xuniDhUwZpMNkqYJG6nSq9oPGteKZHqbYXud1fx5a/HDytLwDe
9QCb6nQx/Vlcf/bKYWJtMvJ8YrSUsdAPxXSkeZWnN1ZUzjDDLLPOrykRRkLM1QBZ
RDeE+YY/9Df8S9LJl7amzUeN6kU+XelAJNA8EgPwvZnQT1+IT0jZeOCCSTvWIrNT
rZizZZzwBJCDb4jALYTQWKxOhgD09d51ojJ8eapWMyTrHAlSs9sXb22/solGOHoE
3CK4I/WqbNB/H9ihIfjQkgWi3VKkkRoK3s1iCvJQ8qaafufNvMInrYE5Bks59xf/
6wa3Z0+ijt/qQ4WD/sTLtK+qLdc0XffSzPuRTe+pbNhq/mCeW362R0otVjp1wtzP
Hefj9wThP4kS57QVRjZzR1lmsXcxc+BWsjF6T7LW3Y+vDPcs5KkbdBrspMtT451O
81T4hzbjAQWJ49DX3GGaz/e13qyLTPjtcn4z+jDSkgP0Oo2l3w1txYTPhg9iyjUt
bBPr6GD5H+AHRd9VBRvACKdM46PQX/NjccpQvpGUtW6lX7xE09dBe9BEHG8Qloc6
dchccN++4KFdEIsA8yBjIOqoDx1lVSb10FQrg2Km48VHNytStN2+oXz3jHu9TPbS
pUH/w7Ju6vPeLK+InEKBLTpJRkKYo1o61y5Bar93HQ2+t92SNLZKqoTty5Id5gZA
Wj5MlYq8oqYSwVqza0D464mSymXPG0s/a/g4sj5xc/jVSGyuxrhw9YGCAbVe21GS
2ZpTTCxnWLXCmapE/ZNuMHMifgQ6naHG3UOME/kewp45F5QR2Mu0zwoU6oxpHbKw
1YJtJYpf/wT1zn2mDWoHa/GtDFYiYl/h7CM2eXMXE5TSljG5hMwOMzO7+tIrrcdH
wQZRMdp8uV1nTIbJxl23fdtEXz88A8b/KWqvY0FS/TnjUXqcg5vnKkS/VhirmO9j
3XD892lnY84N12U/NCBvE7K8taysZ/BjtoMazl4FIBvn9ZUoG3feR9ZPdprZWdZk
mazU9q4A/NWZUW7gToDVzulr6idyET+pFhOG9yp1txY9rowqteBryhb/fFst2J/m
Yo8+qcZ11urgge6Lv5DBAopqMunL5EAFlDYnlo4ahzwoQlRDB2R9WrvkaGWGy27p
HJlX2c1g3YegAWz0O4oHBnyNAj68/D44QjI0Ymmr+fyyUFrNcShirHG9m4FEkrKy
RTo4WMeChU9XPZnF7V50/y9UXuugilXUzjzyoFh4UvX8lgcpfTb8j4Ad0NRjeqIn
N5PsvydXFTn9bnsIdP4ihMSyA8CwzBHVV8zSzyYauF+Pg0fwHFGB+nmUyX1cIoJ5
lLN/KC+gkSfvOijgkw9X36/1Hcym5kMM5NSTQ4ipFB8ncLKeLTCIZMxoV790UCNh
s+i6ut4eraVuI6WAjxX+i2I98gSDi9zkVbaPgmlUYiJlZ3toxhfDNxzc+FvHEOgv
u0ear6Gn+IybD6FJwmFMObBfNf+TOeUXAINCSF44I/PHoc+ad7HA2XbwfeKk0ELR
Tm4F07tdoVGEFnYkK4oJimK2Dqa0TBMkc3m4NgqLUHsS5XP8bkm6xCHM3vf2OEB7
oLFArKIYgLYuIteHm7PWjHH0sCyHRuf4nPTheOpcUWeRmOi2EBC6O5WoMFwOaysR
YEjbG8hR1EHhvYZSBVGihLXoyuclfZ8OlQFNjXrP5oSBwLA27pJssOXMBrnkvIIw
Q+SVgTavNdqt8mdhmFUGDsnsmhZdjp8DTcloYC+c3FFbc35Nx6DN/P0fZB0IdHHr
4vMTSkzuNlEP7XtC1EFvNqjDGfqfziza0nUr9wKum4+RWEMe6r5xjMyweOLEcO6I
64LTrPVSFB/wNWnfRR7Jl2QO/+kESxgW/XMsadyX5gI+2TVoDmB1TwX5CuqoKsqd
+NtD5SVgu4Fhq2um4jqxs6eA1yLuiTFp6HmBpRgDp3O9c5hR7cpLXEfAFg6TGS9R
gQ2xvmgUya0kpZB44xsev77qJPxaHUqA/qkWCZW6Yq9EhPUHJFAdR4arjdPX34ok
fyJpDBNyoCGT9sbibJ1tqt1aSmYfK+lE1bvlkZVy7D+fZUdQL4xCAxI1OoXttQFD
FhAXS8zxIXVx3+7tsXW1t0mKja2AU1SyBasvqknbvZf7HxjWddwh35ilnfMSv0/4
XmmVbHvb9KXBGhZRm4HpjBnNbSk2PJhpA5gpjWFbLbp25VbqoFU7aAtDHP37g7+p
XUnRVNfqtEfoBCrH0n4GTVblbvWYKW9YBl/H5NQ4EraeasCK9xTxb0nbH4Cf6CRK
hZa7x1PYsmxQIDp7mMAftIxh1zNmczcEyqDVEQ1iS/VzK1/1BdHggeZTXdhulpJ3
DRy+Iu8ELjgg8fMK9G9wkxL/L2S3chmx1tj776VtLT7TRrbiczOMueq/sfuBh/yZ
EQTxKmfw1L9ouaGYrshTItWeMZ9laSjyNo+s1lNLz5HJooF3DSQ+EJz8MLfTsUba
4HFE79MZozRu7K0CBBKkkr0luOboUj5SPd5WIWQFIYiYFbIEnLnmyZ3ayhedGNmJ
IfNOKYT0aHFSI9QwpLSc92tTPKk2RtpDsbKtABMqfk9mXasRFipgLgVQvfHc/hXo
vdjUcUsfRDWnJOePNeL5C9JG64CORtzToxT+adsVlvEqhfrgEDVha7gb24ca5Iya
AfKfNSuRY6qjED9Hh7/i7RgdzVcbXaX2/rT9WYBUX+u79jQXibVd+fTiF6KOX9Sr
aVWzx727vw7dUi03o3/COeDwmOS6VGeEx8oAOurDrx6WrMKC75CTJV4j0yLfijQ0
krzwenfB0VY8HcrUjIot54Wy8DjNh3FrAZw45MNydZ5DwfokyZiJVTZZjpyD7NhZ
K/QMN/y8y8BuwUWzVMoFcSKdOBcIYfo8SXrbScIG0RysRNCfU+qnlttdVNNLxYS5
YXcca5X/ZzYqgK5M6hbJ4DvYMQDPgO9H12ckUHpTIrMNzit4h+wavX/7IP41QLyQ
MoOuYmMpGDEb3ZIySd8lzn7H0BQRVxw1zDpU3wtS2VrmdHtdJptGQmqn+sTXc/Ya
naYQD56TQg9JkCD0ojcEoQIXBhtIGfl13tOTRGkhpalpzwgsgjvh+U3zi9Ez1Ujo
0w5ThhuD3ww8plSQVHvNJPLOEmrIdN19dO7dUl7hOcDf1BNzcZ/+jIoRTD6PP6qX
RCLVR2L0mGaKQFVQeJocPUAjKlchZ66pq6CiJBLfnQjVV8R+IXIDVDPYNC4X5Pb+
1QP6ei955cvY5KGumnE6lHEFogq1QJPr+jImTx+S+9pNvEUPXh1r/ena/XMgvZbA
NvH7fVnOwWCaCZBckX0KI+TX8XfdDD5lkgfD68YS7cn73n9okLMhgMnYZf08bnlv
Ey82AlFvMzzW9/GTPqFkB1m2J/G/muEKHSRiwP05vSJ/XD+CWxuX+pTlL60gwLJe
+HciY7mJ7gDuYBQa133+USLdAnTYqN3kQkvzF0m7jLO9zZDIaT2pxJemWXGd4ozP
Ga2/MSplNpXgcXeVoPj1oKDfnnL4cRDPTEspanvEACnI5tnNikP7iVr9XujJKpZ0
ivniKFaxUN/T2biggF83DN+lGLWJBDcOcLP2niH+8DxNahZ+6GJk03sqpVC4hTnt
UsaMu9QlLq46Bt87knzjJTNEDoqC1McqPjESe1C3vJdCD41L+cyk6BweAOinUnJB
2Ouh7kOxaVULyV3XB+PB92R5v9tDg31kEYyEVnuJDFfVG/A3QOw3gurT0U0dLYBO
O7YCnpAFMdWFBl/dJlcAk5WYoZnafDRA3zJAtnkfhF2BMP6hpyOJqoqlMAadGbAC
wXa0CKXY1VLFi42qJP145h7lZgUcMTSzKx4IPquOSPjS4k8NGbaKGmoS32eG2pTX
dwpktUDvO8u9UjkELcT0CnSI4QAAXtnLLH4MZKjg/UJ9608k0+ENBMw3I5lxjgH/
6O374mvy+S3pncELAODB0NhzJv9KRe8lAutAjWo6v7JchpCViaqLY8KFA4HkmW5I
rtCRXYWDKWPjouKZJ803dS7xIexPzhwKmmGbPMa+Umnh87zmgv4IVbe0JkIawbdW
Z3I9y7EnjuSYeNMsyZezRKGkpFcDDaSCM533qYD3KqYL6uNliwoivkr6PoWI0hGP
xYaN9tLNJbb9+Se5m2BgWkoAmVGm0ZBNpUpfkDkYilkOl2+S1zxrKsAWgL7u4QL2
hcOnf20vM598yOX06AYL+F8znKU/G46KAuINUWtxs8tXORkTqHqxxKnC0Nols4lL
ab2hahbC6fGnC1sOrdDGXbSVJb197nJw4GR6LEgkAE9FgISUIgRxU6zPxlLeGiM0
GTOsvi916EV93hzZs/Yeocxo8hshCSrbydl8oPeXfJjZMgfwvaHeoCYDpAHcLIBw
0tbddCmmzq2pdCUotEbwqbtMsWGToW+sUCBFYVggwYU094CEOIyIsLq9NgAG9lsr
iy4bIA5SO98CT+bVGQZYW5YDP+BfVlMt2HAS6wo78w6MD6FmxjjFkS0gQsyCEcxy
Id9Ruj2wsPYjqm0t2g1OP7AJfCeDXE/gaDCBIv/W30HHB5VezSObQokX2HkxM/8z
LvEwW2JfCpXQ+e7SWlPhTTX8+xAIb/ULwFp5cD7IwSMR0+++2+JCLf1vgMFF+Dc7
BlfSNCMrIsX/qohMjYvfRp/QlpuYZz1Cc0AOBrSw7mvczXi5IiGvaLELzQcO0wJQ
mL/BU28CHEBBGqFPwIVbEMO9Y1nan+mwPotKyPTopPKWvmXDnLOjj4WaqHrIV8Ha
l5S3/tDfSxDOI1DkB6KSLClxs+Zph8HaDo3/zaDu9O6E1GQDFrKNz+ywUm+Fi/ZC
NUB9MXnCEemANM+MxUA9LoI4pYTcOPM6p3N8Pr+elKvOR+6lts2nrNfGb9gmsDvb
+t/CR5TduaBrrJ6XBTXTrtz7zJlava+U6KyU5EHHI8r5cT3J1gnO9C/OiFPNeaKb
k6P3DqKqehKGKKe6Jxjm7lLgBblK+dbwxlXxrsi/cebYPEqoV6lEXw3/xGeW1WHr
lB9d9CLjqKiD8UFSrFguvwRCheKoSAs3GlF1jzjk7OHneyF6hq4DGKc8zwZ/fJ5Y
PY/BKJJYhW7Heevai1qqBw9FADOdEw9qL0OIhFU86p7Q5S0jFbbPopWgnNMWmEdh
3P2GEWy2DyaQGz1cw2bdC+wY52EOfzxQ8fZg5+fvLFqcplKf6MU4V2KIC0hA5GLw
a4L/ft1DWZhN5L/AaqCCnscUH0w9W6WkvYHXUb9EC498EUzE5H0rFBu2i22ZYOy0
db9+9MHREa4xOKo64Ndg8gQf4Z/f7Pc2OVVkvtnCkHeccvGDgMU6YepCpEJpvu0L
ubwq/kDtO0buYT6AGedddUDmZm8apagdwoVnyO/xoSMKZAuKtDx/Nf2/i84jJQ4m
vsZ9L5bYG0zZz4+ffLxPtbD0VoJki/etYEXJH5Aio8TlDKlvXVao7LOuPNV4JLEV
jPUEtSkAL0XbgWJqDWc5RVY3h35mgNa5Oueh1z9V5xS29UB5vskBQDnXBgsa4EyZ
aKqZULDGLhIaQa9nOVCgH6hDov1dZfgB2nXH2UI6cJEtf69hpkcwxreBnSVhJauG
ntgNu0IlbXvbS0Z6Wbd2J7dW+uZ/hQWRQCKbudQb2ZH9Wwkh1t91e2pNiFSuN+S/
ePln7Q9oINKwQJEyTqOf++32z6wrq3QDGR/xyQHt7nfbAeDa8sCrur5ql0Ga2WZ/
YATA0jw7HBqc0QMb2GQYAR5/tyIkXALhyTSgPZ/pMP1QgxX+U5OPPRXSRUS838Ix
nwstgMKrsJicxepE8EkzP7otyqZm+brUDH4Jv0RwFrnCH3KIxYk3mEA4rz/4RT/B
IrnRgVhxTjXvx4aG11siBeKSjZjQQ8oImTqT281M5s1/OeuqcqZLORdcKuHENApU
m+ac1eBF2SMXEHQhcHk/9nQy+8IksZD1Ynbv+AtROfYU0MRo/ZW8tmwHdm30fbo2
5l079omQMsMTWCNEtzv/Vh8FPdLTRXDIFgN0+8vX0qyIF4D2eXchuMkAhQzRu5W6
NOQEjgSZIG7eNz5vzYqU0cfH09NZ5Jp15a9cPiDOHed6UPyVAGMC7LzIhc2IVScH
8dnhqCbEMmVvcQo/lETf8I4eYAEe12SKnOhEvEIWGGj41EPdvWx4DBJWVWaCYEG4
B6k79j92vtvuu+hbaiKmy8r8/QMpDyWEOHoFP1fpKD44XSQhOvsnF5Mi5c6es8v8
4KaDzRAJvBDq4e7g4z+X+fIA3GNH+zyYXOLmUiemho+LBDaXZZDML8YMuMwkx+Ub
xhEWhks4lXvi7IfO8p4MYC2Q7SN3kX+mSSOR5rX5I48VqlDDFsLIrk5xkReY2Qz3
D4rPJ1nsWIN66yzS/5CrLYd86K28DktayEt9kM4Vg9vRoHlpdpQJC//4OAo3TwHq
kgzh1qimq04m5goYllf8hAC6bmG+1zFBOx/0JWH8MCIHWQzzbWZepFjwwucGxjNs
j8xEcj+UpPfGG3tY53e1P0Lz7ffsN5SHKgK+ispK/w25myqwF2fihXvhPeFka5bw
BwBZ4xHIydGeJdEOsujh0weka787r/Jt/pgk6gTUW/yU3YabTzQuGDjjKkkbDdRB
Sh6oLXSMzZzZXnfRAs6iLWrySxswrHnWZsSB3WDqt+wkp42/OdJOb25rzay5RMRj
xI7GWHLGbKDTZMKMkBwsnHaBLC0ZE6u0Em2G6Ko2cQU3wqfGVfMqfTFr0U9BQm0G
NoySQt2A9rNFMAmc96q1jTEEHizXzVqKxQCwFfMnYD4Gcreq8NxM/yGErjGvPpzf
lov1WpoIAEOM6lCrlAAO1T2+TXKHfhIcexJaaZmszT5aq6X4FpPYXEpsPFXB2Map
sHJ06hzbW8Y3Jlb4Fz9IdmwJqE2RkUqE83XhH+FtxTwPcUA6Vg3sEpoD/nXFxvVV
dWVeTI4LKe+mnh7eWhDPSab1Bdz+j73Mbibb86/+rCaA42qA1ne8RpwBWZpgkbQ4
xpQZC08f8CwW10UEfKQO/Fi/ZhhCRMWcLegGTpd1qVgNFfVs4m9Fq3hUUi3w+1jK
2Z2JDuWYk7sJvalEn7gSr3+Fpw5AwtaczE4LxcKYaMTzKqXlnzap39CD4Ggim5vN
lrXmcQr2kprJZ/SyUhsl8YlCdlkdWmwr1x/+PgukxDZXxmV8oH5dN/kYQ9S9PVZn
1s1LZjkGS6jf+tILNEqzr9mwrnKUiGOrTcu826byRoPAcpV/mvph2WXFUeaclOBn
B0IPIfbmXNtZz6+x11vyY4cf9rRH+SwsuFIlarMUsOiR4JIWO8o2YqVVT75ScPBn
5frKPQOwbqKAVHibS999qLmvdLrFd+GoVv57baiCUFAQ+HkOtck1lsJbACYknPE5
H305WF+8ou5h037iUszUN5RSYaYzxldCysXu9d3kfY4OZAybLhb1eyE10JCrtGoL
lxG93y4Le50qNQNlEGJeRTi9phLrIbGiIqP2EWoTdVm/uHqfmMhnuLqESzLWn3C7
MXHQYl2cGqvJSFJQzpc434D//RMmtdHUuKbTJf5trRi+wnr7TGE7JyeLGILYcxy7
bUY9yNGJ9jLBqQPztBq5gVc5HEie0nkbVsc4jId3ob9XY7DfzRWuQ7Kuzs2+0ILM
0dvb18km5pCSCfI573oGRBomtVIsMTIwpWewenFugNad1ZKHrIeqilMYBlVqOkv7
/9Px3R/LgSroh16pGUoyqKR8dDcWEI1v7CiISywV0CJRf2wa7QasdudAwx9k55ED
yIeY54ootZtFkCPNTjV2ysM5RzJXaI0NarZeQ67JaWtyqwCxCKfbeOk6OQW+uRKd
BiEqsJ8xzN5Bf6UbA6Fjz/zL2bLbwuvTNcGaUF8TIygYWeU9oV/Hi6Yq8cEaf5fJ
cXsl/oMpbnJqkWRbSponPqEshTosX/IHML8Cmonmrux4QQMlz6MlJhFm65uUdQJI
+NPbliEIV2vTV16hN1oBMbMR2ThBU16xhlLFlp9E1pSUVQ/cUJT0VvuWp5qZNXeG
5WS7jv4+T5Ny2i4rF32/hyYPXYgkm4ET2A//8ZjcGneYvZlBuLQnk3m/emDaTcVh
GdAuffM3qesu9/lAJ5dZgJBRFI36Z990QOAn1X7weIXvH2UJJjXNn/gmPqqGx1K9
AX4qhaZscOHyKVm4KNGk3vcvf2m5yJ9xZkyiQaBojrjWvhbObLAddHb7W3zN3Cyr
FjWw/ZJo8AA7Xl+UQ7k/5ia1hJj34oichM9TI+hS7uPtzitcI1MBxL7HmuGHjNmB
42mQFN1LvisFtfQKLD26KONbnUOceyFKrKWajWjyiOV4Md/mB42sm1P+OShGSc0E
ikdm7qYb4VUAnbGFGybcOaYUBvq0+lVzC3Ym0NW707nLN3YdoH+8DKTyLQA0/kBg
qkmvubzKwqgNCLq0Vbgxy7+0+OQjxLDjp/kiaQRWFDrEkKWp0qqdqevz2F689w7m
Q4iJF467Ne5loeEYgUdJlOJAFHsYj0K4PPd/qpErGRmJ2W+EjLl1wF1rtAjVN1OS
Yt99+geTMu3Q+PwKFINivWsWO3grDl4BJtSh3VQUhpKQRMeNvvJJfCYEVZjnb3SR
pcOHPUx+NEB4SfIj98zWeFTsmZjEJMWaw8V90JBQbCRonjttY4s/PA01jVDUfMCK
Vb1Pm4eD6/0UDudns65iIq9/dM8RnkHOuZKTmQCElZnvmfCpcxQNm29w+Cqh62yb
Ca21lYMXctAo5lZnU39tv7jJNn+n8BcoYZx3higDZCzmyuCNcgUXEbw54DUSOcqM
CvXFn2gW/ZVFIQmthVC/80Goq34n2KpLazxwpl9kfYm7Hamd8Y3+4oaYvJgPAgLU
fXOX+ZomG/PnP9P4dZCXrZWKp02li85j9rJ3O/0KWLe06Hbkuwr4/RfZL/X50RXy
V+ANLtSBJhWdBEEq9Dc8EOwXkqDhVY8qCe/T8K/ylAXqXvfjgfPPlcLH4ibSbcte
FD5P8X5+Agnd/7xfBv/fKrUIitEFKcs0BLnvc9BLVDNLV9h8qH+dxxUH8OqiuPx7
9P9GfzAVs45aZo2zDpY0/xSYV3ND715X5XczEpJuj30bTWcUwtcWFHp9eVXQgrj9
ZfsEeTvw5CDzG/HH5c651mvGaCJMNFn53h/GIzr5bD2ueRUdoTWgZQaWbWueWKYK
WvUAWtgvQirVLI8w67W+ZtZBb7zfwCWORwAvkOu4hWpQscPhASiafX3HImy+7d8N
GSRYOBw7ShGKjozVdl/I+vs0HHf+TRRbfnMCZmw7XT3Zn9SGYN2y2kF/zpoGuGsK
4AAZO0l8rZk+Ej8jgH3wGm2qgZ6m/cIEcFMyqWqomcWGkYssVd49wpnJals9UOEW
HhO6asuXMFqgXtxmLOjRwrCKtDV+B2GU+gwio3H6Q3t3FK+UPiPiZLmwA4k82Rj8
30ZPVtd4YAbex498TmETBdfLQdiwCRMqyTJI9SDbwRFXO6w5qHfsTcdxm+6xtfH2
/dfJ7Ccwh/h4EZWMwx0P0EDGTDHnnGpjzxVFrUh/w0zxxX9MINomVrzV5gfImDDx
acXAycpGOIGHKSmsTHTPG8CHn6bnZPn1oZ+1ezje8/clIIVNH1Pr4tMB2TDjKKxW
Xmn6NnJwW1bhwImhn+SknDD+CPaXQZWkj+I5M4B0dqezmRp1npRQtRGGROYBNltt
hMUca3ZGhUDGFvKIr63gE8MKgXatFSg/o4xncy1mVv5Ac0p//lvFQWtYvC2jafsm
sFcnv5FqR9xNv94ZOBQ3y5BMNI5YHQg8A4glzKLQd67AIBnzYOzg4GkEbVX6NUa8
/ePvqOMXna5rTqYIO9Fe5RyJIsxYVcBXM0t8vr7u+/AgE+dBBPEtZX8CQ1YSLhG9
gzIhT0ZR2eyjXlI7+ypP40ayOCm6c5spRHXP4Gcoo2KYM3Is+T4i/+qbLZf0kGpy
sNB0zU3yu6qwKPGudL3lZMzfjQRGA/dt7EiksHUut6ZN+3mFL54+8x0wJ0nQIFGw
SuLtDyYqY774wNTpk9Ff5qthhm/owy3lcug1MxXTNAplyRBndTvyN7M3FY+VOTuz
KXB+gyplDuXNXrRnJs8Jo9rJ5rUI2lmBLwVstDg4RlR4Xpz7x2QERg+Y6WKUeEZw
AOIBEFUwDT/B7Bnoza+KznDyDqm6VC8ogUcRdB4vfiIfVa6aoZSlxa2bCfY1qEFP
yVFlwfYF4hlJcKx3ViukvT7Mul4IG5CsZYJXIDjrVkaQf+Ae6gFSy34bDW20yvrf
ROKuAEn1axfgfQzE/XqpBO2QWrF5jRcC9ZtOHinulmcuEWDadEErskXJ2/XJVZzL
UgaavxycmMG2r+upzTzY5Ev0HjqG6x+k99FrZvJsEPwI5OSWxp1ff1ee6uaECR3+
x1Hnu79O3ICtcR0SDgi0poIpCjk98sClK9nhbiO+XyLiYC80otRb6RUbdKT3VAy3
VHFNXwt7qRGzWoOVDR0doirEki01whAHIBg9sKJw9lhp45PcZfOOObl0eaWNtpV8
EHyBvj0iHej3OjA8Myh/hKJ8ou1F4o9f9om3AL6i3zpPnhVL6zzeoCKpUsV/8VbT
92y9GSjfklPsuTWy1gvxgZjp2DwfOEPhsMnORYvOgRzY3CrCgpsCzydp4rYMSyXO
CQiSudQLynNQKztm9djiPwfOKGnZY4hG9sg2h/seyOlPtseAi+Nb2V8vjUodcAK4
c4oa+zwB2XxWS1cV8S+Sl7p3CiJqdMMRx79J9cAnyUdosODN9s28PpEJP3iD9Fu7
xeDAJfuDcnDIjSXQzHspS1ojBd6xem9c1jCZslHiGB2T0rHJXzrkHMF40FNI4e2U
h9eKhkZAyJmvkYuVkZz3lgVxuNqCdhqDY4YKCObvmqiBAPKx2PFfod+q6rfu5PX+
xs+Xgoi9qWraUF8GKa9a1X2JVwOGkxD31JzLnwMe0dorttQY0/XpjGJf47Gvztv5
uygfvPrZyxqLXf+POzmwb9Uf/UXIQHOPx0uzO5wrO85UBkBYqT0zVURUALbjIXOi
7yy1483ZBhy1KZMVUvXS92zV3J0Uyfp4/3CJH4qt2k30XoNgWlCR7hCvi6FZuhUn
Q9Fl40PKIHPyzEUrj3fsxZvnNdDNo89j3/+gpmz4t3ohBx1EvF20FcuVfOcJx6xC
ihsyeJsoCfXhUNdinLRsq3v3fElhQ50zeoNI8gfxU0YyUJamvd2JpyBuCMyogYQ9
qD1eUNHwInlasVBzURLl0NBJJh3dvPi7oem7mfcYoYsoa/MrUye981Nt7i/2hr+p
Xzhi2ckYNKGdOSUFcCDzWjJaPFM1P2eGH6PxFUMySb0A7V4Cndijmli9urLsYQ3q
iToEYq+9sSt/sk/AjhtiUeQnVis4ea4WPQ9OkHF8GXtmkRRJVvIv0xvULKyxTwFK
JawCB6J2yEVaFOedCIqOm2mCTrHMoxIVyE7/PG+6oRrZCI+0HAI2+tXH8KUeYmit
qGsPBiU7Wew4Hp++w3SX8AfSF91xWvJcPh4o/gE9oDNAO8b5qs1+hZTJv+AL2HQF
QBKfUKO/xClTnbv19IFD3Q+MpXSya9m+ljybchH+yI7KBlcE9L81HmTAs+vi6H04
k0Hp1mKG1fmJcSbWH2QWBnyRIxELQhEwC3tcL3EUgJP3N4sXT//aa7gLP13K4YSj
jIL1gjneXnQCmQ7YH2EQoWrazv2J7AKKIttWlpoWALlEaATsYh960CbXrdkpr1Xg
MNw/0DvqNiUc+TuNoTamHROncDh+l2R5751f0hVkDVIdT8N8+U+1GtIUJakS9sg5
vZQFQMo7u0UQzwgCw+bEaJkVPyM7N8b/+VExs8UwN4LOzeHKemUg3Phb2i6Os1cZ
MSI34BbUDLJhTVSOj1kHo1A8P0aorrZyCeIQMwHE8kghmEqR7WHTdWcLVxK5qsqx
9GxYVOTmUfY+ObgoMxs2KfdKE0zXKbM7ogQ4Dkk5Gu3wtfGbjIlunxiMrncYlUSc
uq6ETgQdazgxj4t0t/2RUhM8cfQRR3gblOpYW4cBH7Cy0COqEm6wg/u2U2YGim/u
z87R12Xvs4SiQ6+HIA3xdrq6GtsFDDnRA6LliuN7b4mo8cE6cclKafej8JY3E79B
omCklCPRrpeu9D2gD4kFBp6c3AfQblaou7hKThn8R+b/IYKc4XuC7tbEO+CI+sgY
1jBp6JAqgdG3rDm3cCeD/QUtiK/Tdxop+DiVC89HDS11ak3YbGwewC5rrOrJ8arm
AoD+XQmRo6gbU62ZgbCYkYsYMIxUdn0Y0vym4eGY145NPI39u4LCuEnALTsvz8PY
oxjM1DvlO01N+Mr752luNrL4AnRVNxvjBjSxLRifUUtne2zdrND5N95tyt6M2XGl
GIDDaO4caRYXDds9O/MmM+6G+Dvax50UDfThSk+yoXUPDrbS1AnbxvYn0hm3RVt9
9ItK44Ntj3Lm7VbumciwpK1BCnws4IZKgAG7qO+2I89H382idTSi54CCoRZ1YERF
FybNRMHf0/KnhYHs+Yi2PTxHFuvaEfjVLM8UOEjOoHs7DUewNF8T52ZJleLzTGX6
GNJSNGNNZnbDoFdZ8QtMqGYEQ0S200mf/uAUgRyz2LcJnEqGgNFSd2xxx0IvdxEq
blWI7Ij2n1o7/cNjGUdTznWjZKKvH1S+r3lts1HdCdz8k86+LvuxIHHoGdBUfbvz
u4YHiuZJcbTP62Va+jH30ij4HCMI/E9SrBn6Wll5LmhRKpiADWrrpsythfpNx5+h
rCmeD29ueM/4XB0RZcYxzSx4XgByA5GDYNUwed5wT9vYSclp/3Zx8nP21Nc8Icvg
bSZyJ5oaH2urYvUwCwhRxP/QkxvNptppkemQOJ3VLQysp6uG9eKar/vNescRekUz
jU5FZpc3rIC1TmFS39bmBVtkr+noqSEL3EzTMkEFbmRdWMAEdfXDPd9bzQfgYVE4
89Pzbv+JxdxLKoLojc7dJFm8jRqy1xu6k3SdE7P1juZRdhfuH0N1EwLLbC2lJtHS
ppltUHogENYE4vhFVfc458bf5G05A+Jx4ylpejLUcCI+6pcnpdNEle9OqIWp7XiV
Thn4GPwdU9t1ozSx+5eGSHXYy7xHooS40aX0o6PuKk1q9X+pIkpUor3j/X/p3akT
7I1em+Ca8vwZqHPhpNOwCABFdzaeWxoIcpFRdOAUF90fQsA6EOanehVrMwVx692E
mZpJFZrzFld1Ordl4W4dPvwrjIb3Czdb0qj5rS/YJtu2XfxenZ85PIpKZL18hi1u
N4nChJBuP50JIcJc2EEVUbrHLuwHwAEDaIv//BfxTg2OzQkzYqeKiIWu/l+9NcVI
3YHKlOWiIqRcj7Lr6npQDZrEyY6uosku9uLldfJ3+Wq4AMwibINSvIu32QAbyQUg
L2meLOFV3xJz0A35Psq3tz1jufQD6SJf+2O6iIjiT1QGkoZ88T/3n4lGc0gvIOh4
XyHj501Nsodnr5LFjvapbHMIiEU+je1OcMSCN+rT6Jv5inKkULHzfBeI7yu3PnXN
f/YXihOl4Sy7cT5kBJG0HbgLCYB0gzMq/Gt8HPv/N4nLUQAlTDYtNRU3evXxghZB
4BEkEqVtF4GXdifipFSYZzgInZzD3z4A6tXOutIUXUJlnwN8ewvNf7/N77fE/LQ0
zGlW/eppH0Gyh85Sauvxo6T2cgIjYoqa1rT2O1qwR8u07NFIJJfXjBhCz20PWamp
dQMuNJ27cQ4fnEC+ES5+PCmm2nbwZXtydT8iJHM/8iwaYGjRsk3brbMYjVywFqIP
ScFOfMRY/BUVRKqYlteXRPmvwu7IgDYrQFKPggms5WxuzPUV4a12aB9xsCkoSAw4
LNnOoL3XDKK/7TcnA30pYPcLyBOSNcnlK3Qxep31dnF9y5eI7IOyCg5CNIIWkX5Q
2T4IfvyI+ZX0wBh/oWDOEJ3DzgyAA5wztgi/L91F4jlyY08JyYvV4K7eHzUZY+3+
cxOHX4PM3CFFHosJNk4B2jf3ovTEz6TC4/zgG+YwH3QDTI5HGPUptieKvpofFJR9
a6GoXHSFaWcRIoLEEiE1x17fnTfWEdNZPxNIIHx2WLVYhya/WKahDowjIPf0yW/I
DIdWpmMG0xJpXu0yhXzsoWcNAZtxbJuqLK2QqnK68x1g2vDGGJ5HqAZ+8V/CVUz7
fn3fdTNlXrAIRpfBNpwu7zPWMJCzPp5uzmHVZG5akWGj31QbeRga76BYgHWFu+ou
/nAwtdI60lRIsn9n3eWwELrVZ1eJInvRTxjaobnZvVr9Np7Hsuy2z+DPV2Yt+2QK
mwepf89D5texj1jrv37ZH8hqcc7uHpwrTm1Na20ozIViZA9jwz/QFLMNE+Zy0St2
7w3+MidSQC0/9tH7fHXY6smGA8iRg16YBYI7j4qvGqiUwfD8omfagMZJ4P4lKKjJ
Rs+uVEqbD7lzXejKUrCClM+sAvHDUX7OECQYEEj/ZPVWMcEaXPt2rFY06ZzHljII
ZTSz4KTVWz/zUSDEWVBNlmgowmcpVjeQilq7MuN3LHzDk5wPXhzYg48gi2SRbsXo
5br2xI1D3cEXu0TnFDBJyo5gIcRM20s7IqyC0hjhiPwlt7EaqWP2fuIwt/b/Z1AT
E2NVtsfgj4C4Ty8KCX3uYvc+O+hZih3Av8erGV4dnJYxIPwOU3ESMeqzauK5xazG
/VExHt5GpWbpjioDdzSI8Fvh3p0SYoyJtnTtrAcc/RqDf6rXD4YyZwp8QjPgcbkt
0EckkOLWMAZGQNLDa9D4m9ZWexH5vRixuosd2tQL8w38mmW9x9P4y12n9QdLeZHf
KUmoAN1JX0IujCfojXSd/vdkLjJa/s8gsSl5yNTurUDvBwIYmuOxQfnl7WHGXa+D
ukej5I/UXiuFv1IiYNqF1gXtvn0W9GJq9yTj4Ibx7yBTJ/dJNAzv1jcbj2Qj29ee
xAVsUZoSk3YlHP2wp6M9f3syVaHxBrr7XTiDqFNB3eiAPqppC4tUfBbc+yafYwR2
XZSYcJxe5GRsAsQYFfmmrv376cbptJmX9lRCz/3uwYBz0duFlZ87dwnU6Qnqt7AB
S0QTqaq8a40DMJbt2OD7V2beIe3gDwfcPQvUGIZqZ+fnIdoRcg3jg/AoZK2OrB8o
k3sBHGtUkxuZAW0y1HKuEQJPojWsIfzvYXFqJtPucLE9tzj+Y3lEYOJ7d22frYEl
DnF2LTJeWmrpcoEWJ18cB3cVQxPbU4ZxuU9S4t6/wmeVkSbEax08SIgBMQjh+JqG
Dl3liaqDimb3fkurZ8QVhU/4S8F51Ojxmpad+aINR+2pn0CMNzAzodVyXyrJyoSf
xc1Jflb5km+9jWYNxvZtG9HXZVrrZDp6jG4PJVA/MOm/7YeNY3GmCxES20KhmQKk
QTsywtgQCOoDjk4w4VKtPyj9+AfNiTYAu+NaDmVNIp/+tFPc35ecZY/4fl5D51mC
SRb344BEe04khJPb4Xso5aPXFlTGm+gWgM2fYQAjfSthfSgzamkzyMb7nwJNJUir
IHq11FbnK7y0VClb4La00pXu8HokMP2rKEI1v61E6j8GwH4CuzqEvrq3OYNHi9I3
tGqLXgJzosr90cPI12mn0Y2y3MDQMKIs5BcbyGgIxWRf+6BlyMFt0H5FZ8Kg6kYT
VAMvTw1lWc6y8zbqTU0hMB7t1h3aZDCqT0thDzkJVyo6sccuYKqP1YHD/C3jIIzg
8N4QwN5zgo3ZunbLeo61ksad9sVxyR+m7QemfZiwSsOAWZXYACOOl4nNLgqlDB+W
/CUWrE0q+gbMcMy10KPN8YvDSm2DcjvZ67ukA7lOzqAcRdNS/fLVbiuKFBHLs2A6
ImNXpHMIDkhQ7tmwlaTQnedS8HPCSVvMLjx0ZrJb9u4vS1sFDXPSAtYneFMu+Ih2
fi5rTBCKnN1a3wNwm7hjYZ3c40puB8pAIWtD12zBjUXx/c076UhWK4mh/J2G6IPi
ip1uerhfZTh83MfSQnRaTXcgvWY9o7nSluBgv2x5TP86zuZIDeCSqs3CHB74Qr9c
sLcZ+P9IHg+SB8/vO2xpMHM+PEutbq5MXRUOKYdCgSOvSgnZ5m4N+FOlWuHKkuwh
bD1ZusWp2YM5Xs182nYmUBgzYmVKgfS34kSN7y80HUBbeBCsV2e5JwUinXyxK6/J
PyBNJEpcYB73rdz4FXF5wbXC639PEKlf/n6UdukA/IFGg+n8HItwIPQpSOtO8dwv
mhSC4SqA+l1teCnW5t+7Xu/T+8LVtgzzFq/3Ya/nJIa9h+wdSxQxGD6VxrqPxSYC
vUFiioj6+uVbosD+beEwSrICPt7Ui96Ybg7rvn2bkHNgfuTU1SH74jFyn0btA5J7
QhWxg+pFrBDv/Eb3rCOvTdr4Hl3pa9G0j5iRkynObcSNhrI//tk729SEaeaemTla
M4y+jDlBuQdHe4qPzkzW6tX9fi6c1RTEA1t/GAiSEzw59K1ZTrEClRb6h73/naz5
J1X0aMMxDeFMNSpl/epNgE7SAmZYN9cMk4+L1QEwwQtoOGeiFbZ35OPpFfohmD41
jSTRd/KWjEBXNvHNbjNoiMmXfGt3IkW26vZoqiYgQyECHEOxiLcBbg8MmMdD9P/+
lTLdhIxaQf0cQifW2daggICy6pQm2EPyACbfd2JhelPdU2hRvPkyF6L7NxySVuZQ
H6P1oXrEcC3O48ERBbyl3FkNqZsWDJRH9lyOsj0KzQsPCYi+iYCh47Ys8fgePlal
Bj827P2Kdoj/pvBSsMffCk4tmealgavdv/XxbtADQqp/OGOPwsNNubdVh4X96/Ra
8oJ/3R06e9erySw642mpyVw4B/1leqt1CtMIhbs7l/qTcd8k41giz0KafWcmaYAN
3leu69AavCp8Uhh8s4eemLIYplz7Uhax7JaxhClg4p2B5ELszcN4cqoaGTSewG+J
oqCMwePsaW8N/wqSSBWIc5REZmFkfAx+89qAVmRVRXw3MPtWO4uAeXFNP/1mEaaC
xMVSUHFLmA0hlL8unJEzv4GtVpe+wtU7PIsT4uN7vd7TLk3z8cZsDihKXpi9D6wD
GGv77QZ8HEfeR8/PMo/Uq85fm8oPbbmQQqeLv+2R+kVB2hvKFLeqsvH8dEisy/EE
H3rfH+VulCQCU4ltGgTkjamS57w4ZI554svNLNi64bEgg0wSwHLAojc1P2SrlhEJ
pbgs+oQwAtXRCxmgPdb2EYIVvf9q6EwLs27FpWohqjF1pnYMt9AeqdBsAuwPe/tF
dlWzJq7bRhYwLNGsv8afj08kgKd5uLohL2y3J52q8J2kN082n8qAuFPYppz2dA1h
h8mw8JlaUk7wbTSz91SYKN+q2lgJf6ouq519fd+AGhC+4t6sVxowrTg5TbqG5vqJ
i3x3km7QWNWwiSLaGGzDyHL2EZZtAGW9kFoHKV7JFC1yaO4mOnEPb7XQVQUjGHtn
4HLcUsXuctGim33S1xg6w32MoyWg+l2gf8Rpz4OP31Yg3dr9/wbePDAptWQJnCfX
j2DWfPSMFOwmi+AHzEnXefAq0F/I/faLELx5IWJZCUdVHL0tsOvhb0w7m1N7wkoU
V0sMPb7kVq4C0jkiLdWdErcH1Zx8/utZ0joopi/gnH7Oo8KF7AjI0ENvCLrSjRC7
xfSpsiPS7sCSEKzlhcuEbvUzn2i5S9LgK2upsaCa3daGqy/5TkSeMxfoarY7lsOP
7+1jObcfUc+28bWoB6gys8krUHiUkQa40+kXjAMkBeI8C2hk2QrpkYKI7IAYu/ah
Mq2fpO4aYdxjxIUw5Sa+vhfBpWYGgTJAacMVMCG38DvjWcC6l9PA0tjy6ED1lje2
2H/KbJAfv8NqygsJzIZwdgTp/qj4Xj9wBFvbdqT+HqzgJdUi0Kd/Tac3p2AcmI+E
FXf1/AwaJCAJ+1DhvWePSqM43fIO4lcb74YcFsUwUoJH9nCECTNi1MvuGXcdqu5q
p46xBOQdKtA4hAzgDykpxvROq2Gvs7OXxW4ba3rcexGEyoQHZI6v93XB2zCg89EL
Zk6opHjxx98VoMooBORYpB5EsvtYYgKNoM4cC1ubLzwvvF4s6DMfV+7yD3w+4kkN
FYPpTfSxEfyYze46KLrDtZCzSotqgxhpJjebJ6f8lxecA2eAlkc26lmUOwfmFqaS
8gHgkf3TV6CEtspN0Oyy4OZCpsdnm4Qz8qFr6GjZR1zTB1sdVxEkmZAe7xbkyv6F
1D4YtUZavAaAmmFjk8SDCM8eIbsZ/Pogz9PyT5BSyrIPAnotQdCTk8SlK3YOivqX
MTYkY5+R+AQyOatrbH5K3aBN1od/320X4Mcmii7HAHnE0Vf61wU7ZJOIZqfE75ZT
rASR99FVWnIT4pfASnvN30HOir95ZQo2J7i32WAj0JMhoYF+ifU22gRNgPSrqOAE
RSnqd9PqLdciy/+nozSvcDC0f5G3EYepH+SWjqZynPBV17zYLxg53eBLvvU2zHfg
RbgrVTrDkNp0jzjX5r4eAPA75JCAWJGHpMLove00b8bjUUJXrE8oQ8jjEgf3dnFI
7E3hdM8EM+dzZjmWW8XlsYvJ/iYxsz6HfyRLGyX0jxJLHgWpy6s7jIl/TDJZomLl
KfdD433QxXUmbd5fFYIkxnVW95vPuA+JEqtj6BGjwSdKiLnKFPSBea5kGt+7b/Jn
fhNq9F0miEDh1Rrve5Bw1EcBSVqYNJmmTEjKBtViTaY+FRDIleszENyvaJ9lloK3
MLFs5Qlsnd9oucEUQYhtTVTUtJZHsOkZDD2p18XppM+pAnbV5zDn4AD3AgXHIKU8
jkMZyt01JJknLWyQdbOS+5YEA3fAAmqnxBnfR86neM3OYitqSvtsnVdEqIHpvMNk
43JdKx630orBTF+Ep0Doi0p8/i5zwV5eVjwZc2qCxBlLCq7sGLYa5Ketcm2BMf0b
vcjzNQBfFItmD9nDgeEovdLPgMUErXGYKLOQTFE06hAcu7wxqOXT3MQrvMTtGN2e
jgNxymyMlHj8qzT6sUHkPx8gXqQUn/NIS2QQhbJOu6TefOeQ0KciClggSrhzItAQ
eKwXI9inH0drXo2Md1WDky89xaAoGSlpg4IeF3IPfSFMCXdc5285IUSERS7Tu3wq
gVO5xkfrDkYtE+byFE0XdlfagkUda8o+2R4txAmCwfGPdhdHcPBENhNyZOorO6sq
wEpr4vpfOP7Vho8ObkHhmFqwfuMdkZIw+uGzH196ulpHpP2YdJaEIgDTRbsDBx5N
FrNZsu9fZLdYJQ+ZQR811z+jMx9L+MMmiPLyYZaHlsld9+0HuXAK2kHzOTnfYSoe
BnJanCzM623Gm3CGpOSET1XSox25q39kdIPgoaz7RVj6jULQVQkcRN9O59iRmKMD
W+xR4FgiBrPKEKPlztYuhRX6JN0pbzt/c+JNemrNu/LYsz6MbLaSUy+4E2i2eZ7b
9cTinQqCP5b7wOLLddMbDL4lbg72yK6zJKBP7+NHwnYMg25G4Pow6G9QKQvUwGeY
UZct+FS6Vs4b4Xik0efDjSs1h06bcVNFjLcytQ6hhukSYD3L/TFEwlDf4Bs0kXBc
Wt62qqPyrHtiC8iBq8+wK2YBWUOSlm1+d+qSQTz5Pg3Ywt1X38ZvdZwNO8QagdZL
UcX4BBahCrWi7aqRKl0XJGFU5JoOIJ3M2vtThX/+85bGfVMbX0bx7nQXj7QNM9i0
N1B/iw6M/s3acA6DZVoqcqi5E7CwBsQQAVvz2KMAst9PMxGc1rU9CnTK7JTio52g
l25A6XAhQyKHvtAdneIei6X0DWwtpHSz2uUC1Bs6L3HiskBXmzoyM+EEG3mkV7Px
4+4j2LSPMSofPXBFPlV2Bvyx8UNl23hGH2xQ9SR/Vs/DNwXw8MI6twwvg9aTIVRt
hELK+UxPAnQhTuRNC3xXncVfEs6wm4NOOanvhfsWV1ruAtGB8K83jtILUzWUGxLt
MgieSM7BBJep6l77mlTYNjmO0XvvUrjmxmDx8jUyE31d2/fLcLQ47ev+kVVD7NJT
E2AEon3NtpZMgLusHU4jt+19OklIxJFfPbt16iltjW98ZGd+Bwb7OulkLCP0jhKi
aAdKavIoD6xTmtHV1KTgD3ED/tZb1bYzyNX098KTzuKVl17TX3IhLL2CalLX2zCK
vf3tmcjtXmp52EDHbbBUVSkO6X8uOZ0USO27dW/JmUkWF/T+1Qv1Rp+M1wwbXAlN
A30uQi+k/5nfXVW/9cgws+7unG+ZUC0uzRfprwUwff4PXAO0m4whigvRVaBJQK14
Hnl51QXrn0uzttd1BSMKMH9Nb9OiTaOf2uDhiDM6sJeGAnjlIi75MN3+p7Shs5MF
JQK12saBmJQV/V3J2yeWq2GrLxYhNcsNqQtO2hca3sC+OgqBP4VpzK1oSzkR6wQ4
3DwMjy8jzy9RAlwRNCgZqnMM6gx9TiAfFXqA2akOY5aiF2E9hS6obzBcLfsMZd7X
gyPZ6LabXQjszf8sIeNuIbJG9aUbyA6XFFU+3IbDVqyfvNaWCDbxb9FX775KlICB
dmMb70m8H/UOCWmHjg9jvgQWIzHuw421hELeyfpX9NxBbU0yPT9Kx0RX3O8yqYOR
40qw3nHs9bEY+tx65wfNik48y6HgIpTjXlXN7jJgnOfIGQos7TLE9t833OzcB5As
Iak1fyqtBYGaJt424j3GMU5auX++8rUsop3q4x1JMn4BSMU4CxzKE64KDRihpgOg
5IzapDq7BW0wLonG796eMQvO/Y7nW3OJ5KplEyyzLgZ1B1lgWpn/sRvXg/5R1fwO
GtzYzCbDQrTed/8JauFQ8AriNwY2JTe35OoUOtL0tm0uGqbaOJR/OwskZkHzhNXm
jC37ruRpoXeXpQAvyNh9kW3blv4zdL+MobiF4ECyGOJDLkOSplA/fnOGpxZyDc3d
+7vlfa4vIFWq6cb1FRMMo/mlqDfw1X7K10AdwkLCqdQ40X19E0uiTooEsPR2A4Lg
8qBYJWVSXlOUBg7KWE8049z5DWeXj8eThKiks7ezIeahhED2UNXzsaMAasVIooKS
/ljAEjOLqsSRFbjHpfeuVqf2VPD24YjEajPa27xL9k6b/s4SWRsN2Y49sF7FsEA0
+U6EWMQLlvyoBoy1LCCze4OjKXMT+ihf0jYMUbZvkCNEuMZU822M+aHP8gSD61a4
CB4UjhmadjpdR5bc5Y2Ps1+iJ2mFZ0rCtCddiFkIe5vzfgWnxxOXVCUHeoe06Y2J
/oX7OoQV3WMZNk1kr3o1aDZBW8OB01/uHnEBeu+okgssvmD8FOBgKxIMMsbyuDTE
LouwZGYqLaiFrMd40OcyOKsADKT27G+5RtFqYVe4z9rZq/Wc3jMkfauUf4v2O3k8
g4O5Q/2QWzKWNJbwpDhsQkyNk4nR7a5vM3c5YeNEeplqtPW8ed/CM79v0EBcs/lj
rBXYzc677HHPXXrmpD+aRek77iEyYIR4sPnTbvwufkh6Y8/X7HpTV3waa3KZhO+Y
kaEn97uOR1ZESsXhWxXiPIFP6roqWeKJ+mxshgD8M6UbRo6v9m5sik+luk9ZNx/E
5p1lD6b4dCfCmO3YfsNRlpWMo04pKAjzJsDCoIktP9Y7Xl64yAt8MZECU1AC7zbB
jjEDykPas7fPNlCbOCbSBKCOBeeAV3zsaQF6UkyAPGjuoVCJl9+JS4F3aal6PA5D
S15qFjD0VM0nOMd6UFvi8oMRW2zg+4vJ3lQq9sXcTutyruSsR//GLFseI3EHYwbs
DZfhE0oKGw1wu/mZ6AgsrLIryp0KZ9HX+b37it465du14C/eZi5Lj/k39Ol12n5J
wYQlUt2BAjZrNG1vGN+NVUUY8cGDNmV5pc/atVfmjaY1jVgaaKiyfgz2DU6iNNgn
LLzz6qdSIPOEjpqGCCrkSTiMvvlRS7vOLCBfz7lnrd5JfNW/aMRIwSgMY5ti28C5
Jbn2NrwQvpUOD/+x80WZwFl1cWg0mQKJHpuoKy4qa+bzWNExc1NLtcSNHLRdX2Wx
WlGup2rnIrC3HcTraBiyJ8NbMM2bOFsmms69tbL94sAn/AhTgs460qnd5UQIlIw0
UDsImUD34CdyAFbf4c54Xn+5Pi+Xaz/TacR9sSPb02W5bO7b0xHM0Az6jW5M88qA
OHSB4NT/oMURj9Rfw+j7WfRDs7EOOebcqqWn1h3ow849xuAf6emrPrkfLgRtCLxL
P3ULNvHfsOwWHZEhXcGGjqvZjxdgh4kmuY8I2vscOKdFhEw8t9DbCsrv/s28swzM
BpM/WwleyRPERh4VxGZv8OD/G8NN87rbiTSfrZ7w/0VuRpjiAqXtt8PEonCz6HyQ
H+Qwxl8DMI5drPQXWes7ImkWh11D8yRjziivZ0HbFx0rlTl8/wgDta2YRC2cbStr
qCqOYXjvOo3b68aXBWiVdIBijvb1iwOjvnTGdX+L9L99g2rtkR9tMH0qj6PTxzN2
cWeZKwWKomh4sdef2R4ki23K74zehNv4zBVNqa+YHz9+fSl8P6+u12RcjN/zL7WS
a9xrLxpiaiLD6YFkdvg3NW4YoIK+C7KWEl720KPM6WqgsHNTBfOatkEnFto18rCx
hmTnYu05K0ow7335Lltiuf75l6Jc2n1rFAZrs9Iwd1TVNpIO3ezq01a6dhT3U8iy
bXD5BmH8chesrOOoZajSY/vWLWzRbrh0hvGjMp1cI5Qft/wg/o1Pljle1ZwQo/FL
tIKvAdxBmUdTsUg/kDTOEPtAIUpC/n++PjFC4QOEi19fOm5lT8xksRDev6n/JASD
focXGMRs5MaU026mLmU5dftqDCyNvoO/cX0E2roGPcjsCyHlnSEywg6++Mq3Zk9R
K1344MHD+4SnNx1pRtmBem1lkXMpZzXt2VkRKGCRtcR2U3uPIe8mQif6e2TwJwGT
64976FrReFKOQISgebxWzYGsNS96k6uwF4bY+TR471oa2SCdW3tyHurVDntpashS
Tdo1XwBjbMhAsmy9YdtyR1uF8seV9LQev3NLmCJL2tR2II9tg0P0nk/7n2Vnxc6u
KyhJRKZml/5gdQVG7q4Lo/lil0TUmNmec2UCXmxQ0Wh4B9MIX3LBidwSnynFldEi
Ym1Bk5CGGZXD+7H4Ky0Y2XfODflSAqaoQIS9UCa40D4MA4s7r7Xzy+Y/SzHRK6FC
0nH3ruZgYdu98mdotw7cEj891+UWJT7lplJgsgdbQq+oWWsCOWv9GGZBMw83soIU
jWnrjf9rgzdXyjCD5Ex5L7Znb13sKxfgtIaWRWMajdTuoGZV7ACCqumq230wLhW7
wAF8sAv6Xnuaka3z6TOpiz988NqnwNwgfP5bm2+6OEVNJzuyp8rqy7Fj8RcRYUsc
fvOKxIxJAYWWdBlAultixivwGES8wdvXxfmDyCcVMrZrsKmxkyXORqG+FOVshJbo
myH7IEzdSEsRgX6IhxKJLEp1TvcABsxV8RaX0o+AZbUaWCWXIz+K9QBGAjbEYrOy
0Hxo+KYeeSEdsU2nrjNywXZo+z7ABSB4YXY0mxEvBlFbkavhRTMKRtlIcCnveFGo
e5AtMEEI0urFpdcxZpRhl1tmTKUugh9qNlDZllvJV4bz6DgirrUHNWZASx3MM5cG
o8EHz2nWAv1M7X/URaX8/HC2N0CvZTwe0h+SJXJufcxeCsMZF2bJ8H6iO2KtUWuW
jqi65tgjDtwC2JOuguRr1GHeOZpQEDNnSV2tIpDptuNRLgBesfARb4Rg6qndahUq
wzzIhxUOYy/OJfXBTkjPbgOlSnYPNsyqWY1Q3LZ66l8lfAUYlNalEnu9YGzyG3Rj
hIaFtZupIHv6DwpNfxhvpD6Dfo3AWNRYEiL5TTPFxeha4zU91jO9EP1qzamAzJCC
DpAg4J+IkeX+NaVC5A4PzN7vRALjVuI4dOF3OiMzHjLMKpWbtAW7sVp0SY/6cfcO
SfV6G0qJCaVG9qwjBmPVBGs+v3gR2slLH5RDVlbe1p38I7W0kmZjQKReA4AWZDAD
8pf+sA55nIhFcQyx4d+u5gh4aAF8B1p6aMMPjgmBhcvjUBDvpMsjq1zAr64vNqz+
9YpyBATF7inxXU+EyujvN8bHyMubPH5+uXHOuf53Krq9ukifKeYCWL8Q2U5bIcQa
XACRFJxeki747qXZZl+KENS188GYhprf6Py29Z3x8fsEffpdpQNrDHkIZ98VCpqY
vJhkDZEIMWaQxAMAMrrF1ZR82QrwJEsgZSbxY8/T8KtKFXDZMQenZClvcJW9m3eQ
SJX4XUHHb2cZ8hd8wx2BLYWH+XaVISTwQ5LOwVSG66uoWn3o6qpI7mAQzA3VF3Qx
rNmLx7mA/eUdlYl/MdOsPGB7nh5ytRfV+wwDHLd4jvzyc/SYg0xNNIVwjD+r/fRo
QrwTVEc4STMorLz9Gof/b03hnh9NblwnhuPbdL/pUsSPOh1XPZd4n/+4l3YSy0py
qUfpcAcmE0bL1QzUElBa2MG7x3AmU9WDQ+ylVlUTTBuLEt2j40veNp7cb48owDzL
WlboqyvRHOSuA5g2ghFn+cJm8P0iEs86icio5VT4w0D34eOsMk866HXv5rNqdIMB
p1jm1veZ3ZMGnFFoRAVkIN/2bsSFu828O/5H215u8Q+Guh8YB7Yr6H4Y8q4ahYRv
YoJJxKYuca9DDHgo0NbkpLJgPI+MVr3Z9Ax+wuemW+1XcOSGNwTgsTeA3nAhM4WG
P8Hw/6YI6DB0oCj2fDCmwcyCHnQjjdPaNi6Yu1WJldoIRIWEJdOE2VAMANb1WE5I
zPdDfuS3Ij0PkdMtyjsF++wdGK4GyWr9rO+0zjIP2ltEmHg6/wQ6buzndVf9V6QQ
H0/iKcBBPuuNZXkN02xtCHpVLgiT0Nq8QkOLfufadWxrTmWzITrQLTEdgYEp+zx8
4/0FBuoM11mU4J6+rlUC+hAPP1FPbmVaXiB6MaaQ+ql6naBkQIDKGyKfG9GVvV23
YxlzsgzWO/RDm81oEkWgs6MCkpyySleSGEiOjw04vCkP+RU3RpEHCQypW3uBGRli
4ckZiaC/tw49h7/R6cu/7eoLVVfjrvnRPhP7ARtKyiUcIKibYRIzItkDC4kNOLM4
OxPDfM/scnJCRwW2PyPWnAu5bLih2JAMmzI5lB+F97vNOvDI0mvwx9vzwuY1xqii
eALMC7vQ/cUMrbTHaoEwIDejlKwGjyvU3f7ibjxCu16wjmpSCOxMnaq92Kc/4bZU
UGQEq1cEAIdFq7pIrgypvF5vuv2E7ArgXCeO2M/fFodDALrK6H7V5unhGbSrPWzP
csJXeqnyw/U6aokR0Xl0A1fWtAxw30MDN/kMEwtGO/n+eJuMnQ3LcFlBqrExWsYX
sGsl3plYAq2uP4ikelD6DYoXKBSofb5ivjEjUEXmawhoSOkZA5xe7hmv0/mykP1M
q1oEbkBDuMou9+GMcPg7Q+PFHLQkCL0AlQjLaAYjGvr4srid75hJJZLG3Kgv2uyC
rX67fSnFhlNM+uN8Dk4/0v9Gb5aR2rKdNCZpTSl1AjBsoGT3JITXw1A6/FRTOyN0
1/7ssaB7T/wSZn/lkgBXKJlHb0khnDUWPOggzyWCHd1U9iONV+im8Pk96uxHR74L
QTBIdnlMJ7Ajvi5TVCGl8apajWOPCeAd72wHcu+k5KtBqsv8qyq5svN1ASNKu9xk
YI33cWsCnTB3EkUF8fJWsjswcZ8PYAcGBqVl9WdDEkiC29NR75mGPKU95qwH7MGl
//4XMn9cT2OfvkeIlFwv4p4jsBloldofAV6VUz/oyEzi1chZb+PmoRzvV6p/sQyc
WgDzJHkLrkQK8ZTUHORE2uR3UMKl+iCdphHUkmLixFwRme1yk/PXc59db0EZlnGc
w4JgrI2gz1CiiP6ytSIfj9wMyYzsKUEYTDtar+8GMuBLUV04YCWt/wulpwzoVC/a
xdXRTYBKklt9vGW/qzGZ2/NLB5skb7dCswP/M3PuF5S7oTW0mBmaBF9UHp0wTySY
J3gYmPQQtw3MD8sdQOVr7RNh4MOSBZJEuXNWH/XTrXAK3xc7bNL5FOqr7IYbj4dr
JhQ8HYuzHYNuMb65mQUqu3fnjGwBxcb4oAgFnH1Qp73UE1YwqW68PKa+Nb3g1XBF
oUc2Wojdw8I19F12T/OQXs5OPYUEraw1th1aPLktJut5cjN/plqSBoUDyWu0cHuk
0lZNeThptSwO2leLZpm7nq1j2iiwAPsOBjzwJm4OOnEi8qkSHHz8G79YB8eKdgAO
av6H2LeJ6yHO4RTG2PSbhT/C7l/LynXNLwuCjecuMZ208yi8BFx4l0hbKF5sfM+Z
izk6MIy9Igrg+q3wCXsIyLgjZx8TC3VhK6rkUqdz/hHJiZZ7K0zqoxt0Tv/X5bWj
H52n0wpy2hlvQWFx+Y/B4W9KR201o7091H2LccmtpgPFqX2t3x3G/FkVrrdolNzN
vxaPX+SaT9IHVLQaX4yFf+QzgSj7KMIMq7r8OcS+ug1buK4LqCgrjszq/1JwcBX1
O+UB4DnOCQxm/OInQAnnTdFIpsN5ITx2LrA4yZEbCEswrLe61whKoQvWSo96RR2N
SlC6em84lQZyDoOn2Nos5gShW2Pq/x6xYZYWwEQwnLW6Q9/o2C6YbaWtxcHRVpOH
6UwCCOAAip12xdS3LMCj5uGnurwYGbAheXAAkKZGIFCgviWBt3lZD3haMPc8Qvnn
To0s9wnhAf2KlOo13GYdpUW7EWLGu3raguJUyrG2vFjk43elMMwlhHFUIN6Xg+ia
1wO8BkOWEidMyGXU//Y09AdvMv9CjTeocB/DiuHvrWf7pu+cLlg3B0ey3dkJXGrX
lOj0nSxhVcnDj7nAdcp/wJZy3YqM2xozngKt0PxhBIbvVdaZb30JzCTD22NjDXpR
VWpH3sUyPeLVrBFh6e++7UKOcsPXX1pslrpyZe+h+eg319W/pIfaD4FgorE0zpWv
NmbtsiKdWjmxAR/l1y5kk1K3UYJNUryNlzY3OsQiaG6OLCdgq0DVwC/iEJPjdXOn
KuuzpFOrfZI2ylH4cKDNdoxu6gN3gD9moRNKpKtPJOUTLfAEGk9ITutormOzqJz6
i9VZIwz+lnYewPRGM08cS/eIPZJz1U/MitIwFH54VNn7ymy6KnRqOSwxX01Xo7XY
DVBLcPMXlZfEN0XkWuYTn3BgYrawNqsiMjWUMEwRYZ9BLtEE43iRXE1i1+LfjDkQ
f/G1LdjG7CueCaAREvva2UMBz7zeFeFKNVTHXG04wiNBR26c4Tzr36gG0pdVWMr6
HEH52+dTF6Jx676n0sxEnham8E0pTs+ezTwlsSCZvfJPZpa8URmswbob0vRTWqye
s6mFS1QMcpiy6pb6zHbk492zNLTESNVTcp/BWvgy66JlsMkjjBP7MCGOtitB0+EJ
x5/SznHXsj9yP25+vlErGM7OyrmJ0GsIV+C+jqNCCiO2tGHmEKqWnUN5ra/t0JJA
uchwOSQAiTfMReVfqOYyWkMzxscYg3MoxA/0eTnKPuWaa3+kyuppDCDFQ+X2qaoA
O8fku+NmBtI+v2/JdAdP9WTp5TfK3gA/RfTWZ0+lm0PSOz8RlADyIgTECQxcC6cB
zLkmLTWjc42C2KDVrPoTamGSKd1n9D9TWzxxoOI4mKQlqPohOkifFJSNHs/oNzhd
dKn33kfJm1uVbrrs7psFSHMPulzNF6Te40vRPgVfoEmyLesaZaCVmdnmU5b71jLy
boLNwsD/boAUtvi1DM3mWOzsQegqDosW5MIOaj9aEso9YMyEINU/kV+iVzzpBiAe
+4/YqjKYo36rZXI6scvdWVPDPN5MtUOiOwvCm1EtEGGNwXimH+6irlS8CJqSoVVR
n4VHrxxMgo9ncfcRCJBw4PZmiWcxAidFkGPseXt3N0TFgbBP565efplwHSpHVbd+
MeMcxhylymsurOfT5slsoIggVGOrG41aeaFg9e1uJWPQBNTWqVq4OJlOnvCEUzWK
3YwL5D7rdI7c+9hyEXudpirQVcX5Ui3O8LBiwepf0npPPtDuRHXvxL6BSmtSgV0p
TcN0i3rq5mS8XxyhdwsyAa3LyBk7zhuaF1WeyEoljTmbF0wZHkjyFCi2j11NC4qd
iwiU5QOSwxPN9b6nOqB4i3UnuOLuILpNAuvbnyNLBUns3Yk2Gy9Az4I8PfBkgfSg
GrBcIt9NNETIve15Mnn1qAC5nFBCSrE43V4dbiln5F4TKWWwCUD7OhAJiWTkaraw
BSb4mqOzt6szmrbQSArCPI0jwQe1AMjmISYKdaOGSR+fDEkcIHsWJopuXscwB1Yw
6MilX2T1+Eh9MX5S5UCjXxdFeKwk/dPMbD29sdez7/quLHIjT1ZOGjhoMor4U8V1
FV3yF+yCsQg3j7oPvP7SETQA6FTloZzDjlcj6S+u5BV+Sq2hhjZR4PzRUlrpMdGw
UMyPvGLA0tWRVS5h29rav2CnuuyhmC5ZaXCez5O+DCDHDkp9WqCbZ7fv5xwitckY
4hpk6j1EWXJYAyj3x+QoRisw08mVHrQgM8X6mebfcVc72PjtBXYQZ/CFM35Pn2C7
s31E++zqc1cfDE2XZ+Ckkfj5EjVLS2VdKoAubvlYMm0z+dKznZMqWSVCJ62AfoLc
jc/Jrx36ikTNf0IU0bEbYOVA8eBV46inpMIso8wTCTMhr11FgyZJw9nfv8am81tf
CGj4ZYykGaDoKmO/ylRt7ixbMjqO4TN/jU+5M7KhOekgNaEMeg0RHJEA3FbyYfZI
CPvFE+IFPzvg2uXUdG+VQD4gPapWgZuJRVo9/VbCp7sydXlD2U8didq7ejlGFke9
ewRchWUwFveKok3niNErWvYv3jKvAo1lMnCKxPRJ0Yo2YRq1HXlpZ5UNZFEiAiAx
vzTtZFkTALnNCmeivW3v7ToM1NhKVmS0SldIoplve807slzlc0EQ3PADgy0pkb6f
PYEOW/5411B/e8bIfqBWus5edE5FDLkf4eLUrwheI5lUuJ+9T37zVBIKEDnL0xMV
f0g84MWwv6b5/uEXrug599Ryj2DV4lmRkvnEN/n/J0Eq5qNwz/wSFyDyjZ7UtqQV
Y+njdyzyfnQagmSxzkw+LPH+OZdfLk/kANXu3pa29bdKCpg5lbzDFtmpSoV8VyTA
YuxT0fxQLLaxJdbEqNc/ylb3cuFNk9MMyWvOsdEBmso1Z4IcoBAGFYBj//RRdQFr
+XjY1F2V0pkY3scix1CXx8Gv1gkloh6zcz+TzaekoTOBbhUxVzfD1eN6i5DYCnS/
EscgFUrvrkL+s7470TaOTWtaNM3hnhB98pm/NbsxUTTIxL5QaNtTX7BOD0NT82ym
ShzRsWw+VWawHUpGFWe0Sjs3vaWyyF+slgy4qBiFMiVLKskeP6YkG2ETG2Iv/hfa
LiPMuC24W0unqtdlsaPWuPddkPTolfQeJ4hMd9QbmXA/J+0yVFOOcVEmXaz9PM8U
941lgtasic2dcFFQTmznBIMp9QlPuFqt2Zrp4e25sUoEpW2rzIF4ajN4gm7HFQUf
p5XrOhdpz3pSUFToThIZlJrzMLtfDqF/j0iGNhf/I+hvlUb5bYohlgyl/wIqJpFX
mL6Ys5t/4N6B7dwPbJVPyGnXPMSwod02TMpZXe0IAYgh+dITJ5xeWwEunrfbU87U
S2wrBZdOBkLS4Z1E0B201+BCiTtsi4KT+3/NphHmR5MdYm34g3XeDxT5GJ7iqzTI
lMmz5qvMcefOrYIY45cvFTUKSdOhghFoTgtZW/AN22Dz5IsTnSek3CdkQN23VKtE
rBmb2TTs5Ok8+2WmmY2X2cbf/CvvoJ0isvcYj5Foen7G3Zp+D6V5bcRAdnnPsLUX
brWLJUncbLNlBz8d0wdtw5y1Ezv4+HWG8PezG+l+q+RiwXQhrFwLOH8/sNTOZSUm
u7FK0JLCrQSSdIr7zzU6psqwBGbKDG4KU+u8QrSkT1BsXFDMuhkHMmv9FYib4wfO
lb9HeM1/da7cUgSw6BGh8NyJblPhPjZosYurCwwIcEp0FpPgdyNVDD0nTpIl1wBH
asYqQTT5u862ATtUqXdztl/j0N3Tel05cI2eux+qVlBxr4TILjeb/rgbP9oumhEi
7FMiCq96gYp7YBWefvkSdmP8p2TrTRwfu4dFZo0+v7HZRDViMnVXE+vFQGX/azcA
A3PU4lW4A6PW18V9fBHpbHmiDaM9HNzt78d1wyH0g31BVgpuOI9VdqCM1Nl+MSJM
41kS2UPnJe5db9fP+zGCW0XtenblqHHlbR/BMivqvtYAwZBXNqJ2Jtx1/pAigcG7
9PySbB7Crc3V9Rmek5Hn5ME3Kvy07sDrGLA4ruv55d2tC8U68F4dPL2krjVOSN8E
zMG8nhGbH6tDIxt+nWublc9ma+qi9khzTClOcGnTH8CrkcrRPAbQJYd4DCBbqzjD
ZeW9TjFXtFNuWSBo/OcFeNIHp97KgGA1MgGU/lsdAiHH5+ClUPhKzQS4CY8Asrsv
X7856ODiKxRTZLE8wtp7kUpGI08gqosyXm8g8jL/z76rB7MDDnx5DG/S0c6FFg/e
rTPR3dJA/Py2EDIleYKhkLjGFiQ0zW5NBmfTOJSnbC4Pj637PCzK2b/52fYDwEEq
BY6CMJd8Y+Ci+zlaIaIj8vJ4FSaqpa/YQCyHImR+qnKrrpOAjORUwLC0vcocHTax
iSooykFXZNR+L795OXkkjAs2V7L+Ip2ONFokJjkOP/nvMW14MiGxO+pNMCbrx2NP
L00uKaYG0es7ux3GG9HAVbBd5A5lLY1/Bl+cMNAZOZ7Um4sQalkmJ703JCiwGTxG
f+jr+ALg1F0SQMbcEJPYXo3Gca7CJn7Ec26WCJYKx/HMETwqeFBR37Rcntx+/swD
uEhaiYk20mWpWCbY9vFMIYlBigngDL0F352BnoNERlhyceK2eaRiFEF/TJUWxMm3
1OhM6X2YVbL2SOsiL9N1iG6tvQysSYMYqr1+4Uk38sd92fRgeG9uKRIpb72FEsC9
msCpy/CY4Nq114bo1My+tGPEgQzffc6bWZA2gEjd9HmQt32df0hkK5AU8rys83oq
4g+1aszdKUmyEGttYt16v83gAvHI4h8n/WQ7kSVK+dCtZo7SBX3li33hvxuz25Kp
mEPRXCBvqKYwf8jJqm2z/gaF8536ibvuEQvso7r8cSZy09O0C3tVSro6TwKf/g8M
SviWZ2ohlfv7EqhkKOq/V3NTE10wT+Ghz0lg2sO9CWSFvZzvtMqEggyYuO+BWK8C
VjbdpcsPIdM0aCYAdMlzdxOW7ctJeg0ml0f5VPdLbK/VNV+JAQuZAz+xVRC/Aso6
zKQF1MPqeYLyynissE2MyOPvc6c5akPPZSlVKZ/VkK9nxVYohxv7j4NDbY00spL/
7Lrk/sJES5I04UrA/Fd9XwCY7semc90hrevRDGGbAUtcyttbiJUYJ85rd8T8s7hl
5glsEI8yPuEzdDKQa3p9NzyOVKEs+l+vsQrYBysxBtAsB3yzMB8vehSqFdxSAQy4
Y94a3vGsE9DtKaJX6xzsD20CmVKw1kBdu6ITHse2Inka+xR3I+BSf4+4Eex5urRB
1PljPAsNbBoFTYI3poJ4pA3/xKVDkXnKU5l4JvASY5E0EYcnOF9ZmWvcD2eFd79N
byhgAcVEn/hmsNlI22L/ADniyUJgCTnuizSWD19DnQ3LNMzRybrGbtSRrXXlj0YQ
i9/e7RBRgWCuJzU/aw1D0KpnludNgtBWTVJNZWGGY32LY9mMA3YvWxoXWJtKoS+k
xQQR4fOI/af4A2yfGx3q7zJNjZ94R/1M/gVteQJkteezBglTsfkhRGDKPQYN3zgj
AxYnvSHw9GNAD7Nx2QA4XKGObvfs6V1VUH5ieSxgAtogCCdc3o0DfvrR2n3DbNT+
ilzK0bCabjDnv8+6UXW5s2PcqKB4x3uPrY033ug+wWgkGmhPyn2yY1sU6vzWpAqK
jupzjTOB8fzBYJZKOnXmXy4z1XyMK57Zt1T6JaZ8ZEOH1ECibYzRPwjH//l5yQ/c
OKgGEaswZ0HTSa1Vp74zhysEciNu9JXedTNZqz8XmaplS9eUKl0miZRuwGre82mo
T1aHOSG4w8vj3ttweKYPvtgYE6ouVAqZVn5ltlra/7+wq0GQg1gyr0uZysDvQo3h
U5PR6SPK1Vnq96PHWvFUVnH4ptZ3n7knIhySljjAq/OgnPtly/pJkuQhDL3Up6ta
khD62lKWLO63lQw9edP6C0mxBGSh7geqJXlKsAaLG7WMe6hM+ocG0yFI0gCIp/Lz
uvln43q6am0bZpdcZBJnH6GGpcBmqwucyx14QTTrDmYRKOznJGbZn2kKEwuRayex
VVq7HFQTg7n/m3tiieUjo0sFWgERsIwU6cjU5pwjqPCiuoVn9qWzw0r93i9zls/M
++nIfSZjKoKnK0FxnXYO2zLZsbYpqRznWIgRv0hBy4Up5RIzBubexfnl5cwuAXsN
B3egdPUQoOhYfImTfWFPH/ZdsQYVt2QZWGNR+ysP1Nj6WsHW3MisM3v9ET4YtI7F
yyFPeuKO87ql62ppd/ySEfO+uYTdl1BVLSEk5Wbb63IFbo8EjBDLks9NrBA8cxbV
/+f9zZR6BG6bmYjIMNq3LrYdnQmodd/AOAatvPfdTz44ERBsJYCpS/QjN3ax5Ql6
ZZHwe+ga0y1s7PkyEJR1AJoo2AlJwgR31nyxGEO7+Tf+tb8ucp+UvA42dLABMYm7
TjdpYbDAPm+5IWD7rL+zLpC85LDJY0oMaNTm4Hm6PLRn+bcZGZ4euGc8184Ifooh
r3wwdgaS8AMLddnwp9gLyO14U3dyJ2NY4f9tPMm2C/kQPTM2Fgx7JhO+Xw1qFsiI
WhvKo0vJ/au5JdFEy6UiLF6OC1m0lGEFZJtzTTWRAcO2x3i7E3UyInOcc68xKGKe
4pEvDnqt/zpIl2tWK5xwEJc4rBC8lEZrqH+tjJzuln54pETBH3MeqIj2oZvDGpyp
mW5T+sTkwMSl/drt03D86nbAMJKdOVTwIrEJZDzheJB4ab64iCgFLHL79tYvYGHS
yt3mxwW/zMBVY6cIQ2MWt2G5/d5CXL/LpBXArcqyGdBk5//0MkL3TNKnM3Qym6VG
GT06/10LwAaQpA4+kVk+T68OQtrkkkEz87zxVQab2fWpOFsk0nZyYDt67T9A73a0
74YBJz390D/jH5VQmzManVQdLWoz75exZCrYkJx2KtYLjcsOecIq8octuaWZNW4G
9NFoiJIzvobdO4CSu8ezWyGPjB4m7+TRxeqIjXt2JGsmHz11tY7jsBZ88oV5pCGH
dUny60ncrXr6mGXauUfOFHgEFmJ7Q2pbuI6OWs+A4+AiPBVtgNe80ng8cIlb2+KC
aZbqV38ODHY56kKysFldf7js4D/iWgv8q7xcezB7BMWt3hEG0lcQ91cEBgQTQod9
GayQTL7jqI5544eNilssjojiAT+TmC/OW4GuQB7HOMGe3vYz+7De9TC3XUInOvqf
8CsNyODJnrMtFJBZ3+3RhV0hvuOOR6x3ACupEa20Jz9kqTnj/tmJzNV//Or5tReG
5raSf+CCJ5W4PwdClwNwOfWm+1yAOepCt41pVvF3h6GHTkzcRgVg975JF3MYdUPC
m5mk6CyHtjE7W0zB88tqruls83nTEv/Y/aHXrcK1u0Pi3mnV0Pa4JR0Z+armSUxh
SQjS2sSZx67P4AD5oHXTE8JEjed7Lv/z6bpbu8kPLVV0jEKWTX9+Y4ZEsyLali50
+uo54WzDKypaxFdYnty2EObR9omW4SMMLpMkqZ/nL5zgpWNp8ypifOP/+qFOREGO
WoI+ys//Qt7VtINvzsHmzjXF4QyCxZ6eMfzxyaFvl88bpJHE/E9rdu6qIQUYc4Dq
atw5GoT8qRy7W2w+XnBkwdL7nVxlKD/voosVXnHcLiAWZYFO8WGEs98cGkmmB6I+
DdVJxYXpn7nnVJJGye0j2h65T3sYzaHd4yk0ZilYWAZQ/adxJBuuaigZOIlkqCw/
g1KsXVXHDuUp9BIx/FYpKFrXx7cFvEAxh/VHBr0LnbVi+j/ITFUEddYL/a22gDeI
x4FsIt1IHqpY7gIXBz45lsdiOH+dYfxN+as9wAo4xRGJaQVHJFyfUvDduRXDQkWC
EwA/gGLFw4bpWJKTj0OyDhcMH2+hXOCBZRJt/fDxl0BRaE1sDlys8B/9/mpee6kP
1eGUmfR+/wyzxBo1TgXqCrrUnIxyOcv/pabJtca27/H+d7N973vLOOAGUs8aIWek
KdTMC0/ugbaMgPpYC07lIT1h/BmgAfLb9qhQjbWNsQs7TDcTWLFqTVZOF5ulbrf5
zFl8NGouTs0e4JyMythL5PqiTbhOuNw35hWnnlxUh+PTxUQewpYO0bMO/XLG0v9/
Ugt+R752+VZz/R3SoKt/5gXIV1thLf0isyxPgmWEnw+qXRzJdcr30+UwRjqxb+HX
EPBZT5fYo6RM/JCjjL/wcXydWUDrDo9iAKqR+uqh2dXoA23Wsxmi0eWhqCuRPUnP
VklNHqFVjDO0ezHpbSU5dQNNgXnP5dZgAvwc/lR4lAW8kyC364pEhI2tadALUzK5
iyAW9EpkthKvtXo0KOgkrLy+pKNwLTDS04R/78zKvLJIBOvMKueqrf/mf8GAlCu0
+C+FkYVDzBmpfy1XCGyx6SOvoUwPBp5Zh2E4VIioU4PYy9yugrETaqscm4YNelhM
znAoMYkZoHcPt6XIAR04wUxlSRjfxQmiJ2d4OqTfxdUnQC2dyJFc+jYV3i7PPmlb
H0sH0WfPlckn3bULgD/alp3BuVQWHgVhoBEchWgCTQxGiTJTwE89nf7OMuFSUu1Q
jTvQS1tE3dz6Zjv+wTgqo7ykk+M7dy4OX9TUls3BCYOBI+vf//qkDGl0fqFsyKX6
M2nphWOkU0WYBxCoq05QdwYPhErKbFUxzj8Yj6KCZoaYozjbkeOqfpwhCkO5i5u7
YuiOp51DhuKPT4go6/B8VwkBTZQKqT+rJyzjkpeqNCPOoE4fpoMRzQxmHr2ULouf
ATZNw/PibStYV5Vu1RvfC1Asree6PedNYxbviySxnNKlZVodRTwrIQ2WHE00wKFO
ujWlsTcA/3mZ+atZ/5+ovBiD9eVg6QwuktW+obQUD4+r+DCGOUBjvIHFf+48I8ya
xZpBwiGl9ZRYEA4DXP6dBmC1AzQKFhTJbpCs25U7MyoASuK/cPt3bvT9yL8tjM2O
d87V+4YRM2BJHDJfszyF8LjMtyvUaUpZXgCmQrOKTvwghr5m0IP98KvICid11jsF
1YdDhQEmMQfftoAsyL/C2Hzt/2YOdRIt6Oi7/VFoSZA1zMdvjr8fS1ad2VAJoOve
hqN3RtR7GPcAx3kxrRBPWHOrJHeOygJBIlN4IyU5D9NzXoTanb0eIvuxYTwdxQax
aWiCFD796uJfgtShABCPCZxS8IomAWY+n9kREw6rEXtq3z+EuGGQSnYrUaxNu6Y2
F8d4Wqx+wp2sNvsXQyMTzpp8YDUvK/vMOEfenKGGe4ZwXcBjH4s7fdRiNZu3fHpv
dpjUe/LioAS0pGSh3sP8ioNW93389X2h7Bgb6XRajcbas0za7CLqrngxd2o6aTtH
YCk3/o/IA6IDh3PLQavwQighlVsGDUdsxCTAzjUUMjcqF2P1z3xsbMY+6Kyxr0lL
QH7LC2XQS5MErR4RfJjwLsSLay54PScedpqJCbsa8nmROZpdg9MvipH7BHKK6aGp
Ar+/+/u9Jf9bdluRxw0J7BbxcRQJlnss6Kl4NJMKLAscqWmFC5MiPOSTNWgeGcol
yGFA4WOpIQvRMWpZmIivG2Wr1QebMuoJD5xhBzY84/ydNK5DT+4JxW9kIpCQOV3p
XXToWOQNiVlNLw/yZ/wXRcovlnaaFhDhmmKoKzF7tunw844hsRvHTP5rgPspGJ85
VZF4vwtxd78zVV+a8GJMxoLDRGpEgC4GGU9EYbo8i+3zHRY4T1cnj22u3K/qKHuC
RPM+HI0ZHNsHLIUEExIcZIgUctJKAMK9PPlI+9V7jtWw/wquZO1wgCffqQ83hIsR
uGN++dw+p+HXQh2iilOzzLk4f0EtNsj6ju9yfmAlUrWG9Dzvdd8LAh6BlY3BQx2S
H2m1CSTVk7NL1Aqhxq1DWlVscykk4zrvA8BYO75hlMLdSbtcSXBMJvItuvy+in5z
L5IgEEa5XxlmLvbiKNhi7aMD4/vUO6CZknIu5pV3qXmRKn6ev0bcRE3TzAY4ORXz
uFESNweOpWZ+PN6jjpHTVi3eATFP+LE1IvANS//053AMM8JtDDp4OgWNuBlQKFeR
pE9AtdHbbVSwzjzqct8Cnge6r7kJUe+11pxecZlrn2zxhkxGohdUIgUnJQ5vXYb0
k5yqWn/eF3ietIGKKQnuDXjoqiqFTpFVerzKwLAvgG0XRjzyeMel2c9DDZZWFmOC
VIuTkmlUgIBuVfIZ6kr6abJPTiaWRfFKvlQOCiNhBqGVNDyXtRS8N2EpGGLNlxwU
l0EBl+2Q5SMyShtMv0f4j1QqWIaqJjkSRzse89Ce/jSCildj/hvt2r38ungWpeBQ
cjPRqtNvcYYX1NUBMM1uC/eq6EYrn2erFhcxuNNmVMfUPZqQyxkfJrKca6AYm+Rd
CEH+ZOQKVGgg0LrsDvdTPTYFqfZ1Cv3DazXwmNeiXunpFRmkY4eMZUTivNnwgJ3/
KXn2ZY+m0WaqTUCG6oPQhnKBTFZH6+UDKGy6vLL2MGTtiuW0HXloU4CT5DuBjQ4J
A+lfL/V8IIYeSFbtRMDUSdBRbd5HhuxRhUI1Tdkgj/XloRLogeehn5JxOCxSky0u
aPWhvICU2zh1BJpb0heAdfRLp2bGgezzeAnpy+ZyOoeN3rGOI48XKuN7dq7Iad8w
9PnxLIuZDTDuHufq8rRN+LwNlCG7p2LC6sDV71mda0xpF06rSaWr5e5xfFopcCec
X3pJ3y1Bu2Yx4o0/wDqN98QVJFQaTmNZ+1vI5ixY7mRrbGne6sJj8+gwSJ4gSntN
xOvqGh1A7+R4i6425K20Fer21R86f5ll5dWIwIoR2mKPExVMr5V+TH5StpJQUKKV
HeOEBWiRUWn8jfBYih64Wa1C9JYsm/sIv3SGzI7b4eB1VkEM5vSwodoIyrG5sPwT
Sn5dJ/5cysyiyzMolqgalXazPQQUjG8YSbd4JaNmLka5qGZ+3SA2gI5uPt0SwCDE
tjLAwUpWide/5qmUAldCcATINCwrlLRJ12Jb0sbJBSoCj0941ucykpEkYwpBiJoH
vhxDWdHsjLYun2bD/QaKVApNRAuXb9gPALnqYyxxI1mm0YOCrFExkXEnYH+aQCkn
yo6GitRY6LgfpRsVuqYCXOP6MEGdKX2ozmwJugwhSB7I5/bA6iM2WUIRKf19T5WI
RL8iCZtJSk6Pd8ybRmmceZpz0nOvuPbALJxWa4rZeodqtnT3kU8mld8kYCKtRJ8q
BMcSVjtPHZzLLRwL3BcnjVineQXZD2nO7EfL7+Tf0RVJgw6DGwQ0pWNFGKw+l3af
7q5yD3OxtG5U8x+TmyFJBUdjzkzUTKqL1BrxZgZ5a13t9vQTVAo4BucLAmDUKsXy
w/4p28fIs6/u33SPKm9vDRVGEyBwDuAuv4sB2j50IE5Vye1Au4sUnh0P0YuwhzHU
dJ6ruI8W2fDYYOe3tIwPQTxlNomwLt9fNXIxnqzdEJfBT5U97MejDjG5CAJaHFpA
rxI9zFG0rCyv7tJx9m1AlnpTgeombE+sTgoRc3zcX+bt/X8Fh4x6znhk3wwmi6OY
GArYjd+ukNRU7DLKWRUeiOwIwJdJxKc9lQv+0u7ogcFrgKq9Qe6WRQRi4CRjFihQ
+fIc3D02iTM4c5YH5Oxug9jB6j1oN3c3Qyp1t4rzohzzZ6F5Ywu7U2XJEoAusscm
Y+KE2GWqsz3LDCbOpNy3xONqODRSX71kd7lj53r4O0krrplI8LRmn0EDfzZImOxU
YvYJo5MPlfAI/GuCu8ZwhaQ8sIGVhF3yj1bqUtKm6EsA5Z58uEgcijxZdIfAK4ld
OU98aa/F+Qr6Wusa0rFX6iOuT+mYUQELp/SAJ1wN69NWDekzyiyLYGNQGw9BEWpL
Xt2xPgKjeNUf8rbfbyzTM1hVyoc7zVkgAha5jvYjRUz1KpiUEVp7E7V1FHegQW07
Bu6+145xHFAluK1k1GMYOPooEv0SI+bzKMmLn90mkEoj2pD1Gov9M/8BRPrbMPfe
hte3zk9CYQnrcYL2wuYedbGSxO5OE1zf7kQn/EgsJhdUWJwXyyO3ZblUSkLw0gAs
ZZHb/WqtDprrItIgE/cPLDoohNFV9QLNO9+08651rZUbpWUStWp3Q1XX9pMhU4kK
H27J4m1U7QuLwoKjl+6Yg9LJLpk7eYH+MSdaB/QABQf3bFRNibHAIgQ/Hx/81YbD
08M31pYLKbatfhhKuw1uLCP47gHcE3SH2Y+BSL+Y3szlPMHke8BQFpspWVl2J+1E
LO0/jy8WFpOMzh0+19sEKMZ3kaoWyhIKIZKTSiCZS2jAgov8YE+PU68Er5mP12Qt
pKAb51U2Z4ndEOEiFUnfSbcvsK1Z1jQSyvjgTyl6epuTeVUmJg10PrHtqhhuKZN4
RSqmfaxYpr8hgzrsy4Ie1PxVCNUFJuR3Ir2Am8YL09moGsQtKwDKp/+63a++kNOi
rTw0jyoO9wMM8unI7v+sgdz2GVExpKri5Aw7LO9NpcSjWCaJhdr/azHme/6hV14L
EFC+HVy4NGWGC6X7+rkrD095BvcIXBCrVu2rg9kYEuX1C0PAOtLmr9DaavHj2VHx
uhmIhrAnIqFHpsrUELHVs1+DvJ278yvICWMfK/tvv/O792G4hkhyql0/3EwshhFb
H3t+5+9C7r/CvH5HXFsvg6F9jC9GO5uTBnPpY2Q67PJ98Q35ZVshRZYR89IZA+2Z
7AQQH+NOFqdgUlpkWpjw+NeIhBf0j3dt0Eic8tb+MQRxhM4nqrNJA2GO6K4eWCZx
eFkYNQ737Kiy+4WmBoZFFsCNTeM1iA0cJW66Rv/XNalnNS01dpgpkWgX35mat33z
K1xtuyVyTZTQRWf4zLg+7CoGoZl+4E337q8/Mob0mTStW0VI6BZyJYUF1Wv23rjp
86w9Yp25pvDgYS9pCsmn08rsxFVFmhPein47Phhudnz+6QsapfTryyZjqKKRg6Eh
FcnCj9VQ5ZjYFhPctHXAUnNUiZXAg89NgLerPSGkaLQ4IUkxPgWZQP5+FxmBtw9G
IFbP+6px6LYMwjUvvUfe5sEFWHrPRvXGuJ4WIkbjl3V3P5RHcKw1jwwbuG68PZZ1
qFaRPdO4nuDt13xOk7lIX0Gs57QUDttRuNgqbx7Xq6R/rKTP1kG813KYewP5GJHY
6yRbcyCUlAlnPo6R9qltdDW8XLtVhmbo1wD55+4xfD9bz0Iv0YEzugmZlXo6ursq
IkvY161DOJsLUOrFIWjrQYL1kvJYYSRAsJhoJFdqhsMKQpExl8HnyLYL9KLgk3v9
vWQWNircFMsuuSHq4yBFFwY6q7mIAbRYFAXwObb4YHBtBtozvm28FL2qx90wM628
p2jJgDg5n2qEef83rcIgzRGvJZ7YQ8ivxATiblSuJp3PauyysnVGRYCSDcBMXe6c
vhe0RBHEwUzlwUVmS/He/eEY0KdbPuQxGjuMPeiK+vSyDsHQeXkH07lHkqzpGK+Y
12jBKS1tOJeNqYzHBms3m8JQc7EHAh2DVejL/Bu/EhekppVLPqAWr9FZmwWLtf0Z
8kMQVGDxYuMOpHEP3iIDl0MyuEH3+Olh5+564ggMyUOuKpKRhWz4vmMS+wUG87tJ
b63dA7+8qEVVL1IdRxvrRdn23L3q3/pOaLv+sm/1byweuDkG0BnjFuqIy4+NZeFq
Y9RKjXm5FIeOuJOZl4ci9lUbQLwV3NSTDLXwpG1Qnh6CN73t0hvWHtYMHAsufS4/
2JRX280RQMu/CLaiu7GMoU4r0BC/Jb4lMx+G9h5c2us4O3xY1q0SEmu1CJN/tpeu
K2kbT9nBgF2t5J9QCsq5vbUa0Ut+HZ/6R+mj8YSVDQerONsZgpX/G5GlHw9OVg0h
PNy4Ae9mK9ujgfJogUApRyE7bffmtSJWyHL6bFpFxsUXYCNeCXv3nJthGuMaPHfa
xTWMF3A598lC9Uc0wO+v7WdgK177puqVWSQNVhi4DpCvFtd0tD8dCzTPQtKBfQay
9pvXhSAoBOx0rsbNKtDti1bwMPr4tSaGCXI79Xwt5RHuB4GpcX6UMrR9Nry1sDd4
NAqvhL7Y0/1Inelg0lPSV5Kp4M2W5nqzki91bYTLM0NTxbRCd7jt4KHpNOhsGoRm
p7X2UZ0ZP5k0ibmb5KeCni9JBZfOrtEvBVdqNxIt4DDD2tlecF0WBJVJgCr9jFNq
D3etARMG1GWvzZ8xEW4VXRoxoYsBIBtMoOjFfZQ2irVOT11A0slmxximpUILVxE8
Lmc4s3OMmqKsnRX5TpTHQIx9aijZEuHkbT+t1Sb4m9dFyTMhDEqaoeGnqCCeFSXT
IfHaAP58rX4rkRtbrDMNmZz+a6Lqtc5rq/fGsVXfW1yEVePIuxfyb3HuIxkZsGmc
Y6Xge32o9qg9Gy+66zCk0p2WoynsukN92fXhJMZZlKn3m3UZIeHMsE5rfQbDMjd9
lZUITeeuXTy8olkWS63baZ5qFcugmmQa723LChZ2gj7in5EdgyyUkc/N2Epq4kJv
o2FvNfck1D1qfRdWRaAcasPIz4rNd9mzwUB74e2fw1l9EKLiOBEMl0c+Ehy1gzac
Dez280Jp3LMfcHbS+e3BxDYC+m/D/RukeIPGWwcbVcL2Afj1INbo8bTYJudPtcDi
oY5fhkd9fyut0B/LEAhRZ6R3v0uy0I+uYzjGrHAlTZQJkRLzRtfGr2unFRrrREG5
qGr1n9K1MLK75NWC3rn3hHcjTSYsQZq0chZpqqzTzuT4b1P0kEb/479yU3Ce6fv4
NL9eK2wn7pVo5crofOKulnBeX7VIWz6C57ulDinorU8T/er32Qem2zpDP3OS17ZS
0ZY43V69BgrTybiQsQBE3NIBGAUoSGi+ThxasF84/juES9e72KTl8hBzywT98JSj
HpO7UUsLes0oiOkXFtvdLZgvtHS0182ai5A0W5/LR6kZ2D1pGrS5P6bsgtge9m3I
yHXbqOThUEXk83saCB2mi1yCeZRtpl9UX4ecvSGfAvegRaup+XJuGxpKzmWfGxeW
1pMNpTF0l0A7Lcfh00xoIRjR8e+M4hP7EtU18TWPuUwcb2JR4BYE2fZBZvvPBKOd
Ov5ApGMnFpWOQT58URADGfBfHq9qeigArwbxzeMw80t5hp1iWBulNmT4uYzfMIgi
JRkhSaix94XW2PAFzHa05UwdcdpzRwVWtSHr5A+iF+DuRg6iGdC/JAIcf5tKDiTl
fzXP3G0xbTt+ZtJqDq7kUQfn4pWwTJDVXWKxU50XkhsB29gxz6ATWFS8j6fyMLv/
REEwHIslw0+NFCWAbOlr/yMGw0eAUS75Moke3oiuTa2etCYaqzmXYk9FA5Xkb8Pk
Xaxh3lA8pM524QmCHcBytFOWTdpWFcxEv3j+m9i34DJMcXlQQW0V8kvfa/TF2G1U
vEe6LvkDKxt8XXziX8Tg36pQ4ak66XeMdxI6OP3TOvigz0KyHeJDVOCOC6oTl3jW
f1pyzxtEDDyMTL/W6rpB0ht2D0bUlwFaNqUiLl5Mn1dtYR4OPEcamsyZRtb1JA35
TmMQFJGsLNoxjTKL+bIaZiE3z5O29uHMXH5GHUjm/s7t2jrE4JDGTZ1NSNfvJtvq
2uuvwOxU9B1lg82402fhuMgDy/lvTrXQZZLkJrPUx/tQDu6p1zq/gS8qKjaGbf1+
FIhpWtfKQ21nOuvGHQpY05AhGUSlPOmTVDygjO77TfbQeXDEa9OiAHmKEOOlMja+
ZzslQ5xrzJHc0Zj3wQr8gX8fN34v4bmTmoJB++vp829FnERJZ+Gen3WldGmLrHSW
YE8SbLb2N8/lU3YCS/N5X/7TqwkXogKcrH5jJyspvsdOoE5BxiVa+Om2MYPgq75s
aaZUbWX6DZc/07FAc39UGHcZFGlK0ADKnxe2IRu0lGcG6sgWIr6PkJ/++kpuLdsS
PTCGy1TwmKPMecNClt4eL1k6FvBZblLoVD13SemxwkrU1Y5ha0rNogVQjHDZvXqe
0Icxz+TUPM4iiIWxs3cj7k5F7K7x7GtrIQGBEC9RAJekQAKYesM9oKRzQw1oKkXM
Iavp837DKtBGLVsyMog95TWGAzqu+xxR2eBnLt58vsBMXEVal3y5owO5Qd55PJPc
yAXMpAmAJ966V4b4WsED8oMwztTockxsf/T3uq+bzRecBs7yy6W9uwvvvgI5b1Xj
qq/+uQY1RHK7IUGFCN9ohPae5yyfk+M/V7yfuVGPQIFhOGc6Plib3sitWuY739pu
wSygE/33TxGxeUsJLLBXGFV8jzPyNN1JcqC9hQQ85DRiqkyZIDRoNUoiupy/s4KK
qb5fhWHANpIwCXnmquoTU28Kswh/clVv8SIiZ33iAh1GXDaXaMt4gbblaI0cNC9w
0bvfmES6pTycTCtma7DXaMvvEwQ7PyN+55wPjuHOGZBURE2JHuJ04BRqF7DI4wxy
XupDzcdLcn4jiMh0mri89NgR3qF9kDjQ3sY7eujB9X3N0K6J1lQZ0gHm4CdQCkNp
hGGvndoDJlJ2RY63nwPuaRbtCM/bkPGgKlPNJpHfImB/KbeAKewbW/N8b3uAkj14
qRWQUzR4y/sdDvzm7LNVgyfP/YuF518NpW7kOA730wb49CL3RBazpvcBdbCYYthg
46yvy6H51Taejf98fhx3n+/EgsfXCKFaHWJSD/xJh8qAVZjc1WR0QeOcBUaeNn86
iNdi5WLZYhh+ejuL1Y1MVvAL0T2Ik6rHxqQNjabN39G6+Ogfil+Ib0PBcQ4blocV
KYw6gCs/C9wiyHXj1iyDrLs3gWKF/ryZjROOvbfjcbqnnmWGs4KlsIqbTNx5AfJw
OdNcWnHLvlASWUje9yMbd/I07ryWLfHfFCkMD1mpPq7vAWlksoXrtyHqBjPMw0rn
G1WFO2O4SrakimFY+D5IPVjiZh9hAcf01ieE/f1MDknnFUNKdctJNKeonnmS0HHe
+SdgMPj6Tezb+yT80Uzlpqjrm034aELmyedUmg04NRdGsVM35yJmNDTDl6IjBVjM
eDiQo5pgTDVWf+nNn3PAb/ikyZSyrPoOQw6oXsoMPH+B3CDSP7D05gAZ0zkzjCAr
9jJJgf2Cd7f4yesi86iUA/XS+5Wy7DhR3PlwUuSnIJ6AbcedE6M166aEUaFgAhgx
jgum8mq/pkdYTAzCybfQYWmoBMnEGgZJev8xZ0sH4KvspL2PdFLhCU/0wgj0gQ38
+eYjwhIcm69txANGLCVZXE4pe+YP7QvOUTr9Pj7PESildSK12vy2J1hJh0DSkjNc
lU0ovKdaCejLbQkk6uRCp0AmZiQ42XZw0578WJBgjbEYRuI0/UXvB4DOQc2DuN0J
NGLtmAdcoW+f3/60/6PPZT8zuWB99oM1cDCTON+BaCwbn5pB7f0UT37etbSSa3XC
EZX1xbDfcx+T1BTMCTBML61ZGd3YHqeUwc7oSh7DgWpj+AhII106N998Nyo2hMMx
Znke8xzNDDtHu9eWhHTu/CRU0wUd2c5tCl+Xl6eSS667NxIeCuUsEnM0TFjg3G0m
RD0mcrcQbPUvTNKwwit43uJXBL0fo2TaRAPo4j61WjhJ9wDha5PRpyRtaITP7oe8
6weIzdkfCglCVkOwfNSY/1l3+SexfRdZ+0ZmYKvO63x7P1nqJzB0WytPPelkL5wo
k+GlGVZZDamkMkYweY+//ul9mAhD90tC9dsy1jBkwJ/cARGsO6Mr+VIFnmwGklRi
apMNSP+oFwYibnRzc2n7iiHCl63hAkPKTslZji/qitZaQqCMm0FGn2HnYlnuOJY9
kz7VEuuY/6YZqJ9AVTpSlgffjCEJMKBo5nrEGbzjjsII37x1UR270F9w20jOsri3
Qgp/gWN4fvn4KiHRHUuK231CZ0Fx9yQh526/57joFMDNxv/fgxT03cvoVTBa5nTN
2pz5zKGG8PeUaZcPA59xCzyUBZv5KJeLm5ipFKq6UhgVbl1gXb3a2IsvH5wk2Y4k
tfJvDG5eSZu/FMa9ik4kJN2bTjsiWMIXsi2BTnd241cOnXs2hUFt3LL+KkPhkK6b
0SlSjMv+zedBiiSPxsbhXWrtlNzOULkUJNCh1qQM4zknbgEpMWBD38G8TqpFg16v
zgWzF9r+n+3GOb3jbMW0Tl53y+A4hBUJ0jkncv8AQeFdwru9KfudgyV1F8EjX0eS
gzIdbjpllBnoxST/1L9i/yj6JQ8+kN7AwP4fiBHyzN6450+s59fwcm1mDosxzOCY
DHbj4QswgZ+bqnv01+vc06BHOUpeFBJOVFIg8mnnprRukB6aNOyxzmdHXQm+JBqp
2DDTQgphmw+S79+oKBsNtsLP4JlS3AOjNUhN3iDdKjS4+71MpupllZRcM0hG0l5b
ydXSfEm8aRJVZKCYEC6dWg9No7TrFE+AiTL06edgetZRokGU3QpAhJosSgWUD5tr
XVhNBYyQPF9N6Idab0IiNohugeTuc+BGhZkKl3LbKQsqow0pxRVgM1PJTBF2Nff3
TlSLoYyH0pBt+wXf/9Ko0ic9XsfEkMp5FL+Ixs1O2HuK4PJTqfXpaIePKWEiZJpp
rIQeL0jf6gmUt0d80TF6L6Zek3u0faFEFpJO66qzJMXimgcSldUCGgV3lyZ8PXbK
T+3RG4ZhTRWBXY2yUCK6XjENw+MxJ3p8qzn+MdDTF0bkrF8SuEO91B1x3hsGpv5O
wjqtWZ6boXhG1e0AxYc2T2KIBGQqhpMBXqJxvCEC+IIZVMyN3gXZvvCv++7+XtJy
r6qKREqriduiSHKWC1erBIwfXCv7taaVZyMTq5ng9StzbmEKnWikcTR9h9TZctMK
F7Hj1M0bNGfBK+iciuxXVmgJiM1K7h5BEuxC4aAO73ZFdIv130SiJ4lBsHC5Im5+
XSl824sfcRpgbBKKm5rt0oXZqtiQb30o48I33rtwNDjxqXYGphdM7b3ykbhwhEpH
FVi/Bx0cAW2dnr9YGPK1OenADygx8VCc9BxtsmyfXOl6+sWZg4pK6uxUnoiEe4aa
ATRZeC6wd0/77jYtC4BR84T/m2FhoDmFtYlmxI/7Zna6G4mxsDrXZDY1AfpcUJ9V
WUNrYD5QFvQxqd1Ar56+Adn8NAvq53Ny0/k8uL8R2qgK+JX9JQsBORN/M8YhzmpX
Y/07Io0Dtl5HhnanpXf1+LHOoJugf/Bbj9IXc9R2H+kUKXuUZJD3H9ccA8WrXxmz
w3XLBXL8uG6e//2A+wvWguHONYn3ZtGLfb8rZbUryNhFZFTg237yfuIzLhoCsjds
ROCGRdjvBYvWU+dcsxATp0Kp7EI5FDDtfKHwSvH/AhcWLIO/xrAKQBsPFpQ0iKy8
h+0qbKIfuEd7QZmWWhEuWx5a21ZGLJmVhxN4fESK0fZCAViV9OEAun/JvCAq3iUj
paGl/E/h00bsYfL6x15fxDI9N1/GvH6N3/K7M+qLbODvZF4Lv+2d/jIvUjUG9ib2
01m1U982zbmbu4QT5/HgoruQVh8NMT/abuZmppu/Ngjk0krnlPxEFuq/Jm6/dbsq
hPhjSIUGth+Yk/8WAJTAKXcMRdMnirsN8YRQfQH97vvLadYAG8kMKdatcMI0G0Mz
wYpuXGzLALqG/WdyNk8OPqNiXV+SQ3sN4gkHgSebATaK62XaYYFL6QYs1v2eHAF3
XWcWpnDfJlD6v52NyAhJs0ojHmhQVD+xqR3xIdehRCHbIO4Yb0zsPUYE0zYfpF+E
aSyJIHoa0a2PprowqRLe7zcge0bIDjT9Y86jb6Gt89OWCVKRLbzfWmTzSpO9w6s6
CarU83EQSWcpuAYVgdjOApTtF7WEMkBb2n39JoNpWkm+Vwhk1DiRr/EKyUDdkThH
tAT/P+HniAgcxNpYwtsBXYLw4x/5L9g/Q42xo17OZzGmXpACzGt2Ds4w55dEkKat
UeMXxSWSDu3Tr+ga4FL5h6fTx6s4QYXDNe5vCN/NZPrRgUA5SaN7f7iLDUrQwLL1
GCLdv9qpQfMsF5Niw3acOIEM/L7pVC38+nc33DO9XlffEpcVotFkqjDV0kn10W3k
2QFmw8HeXMffltu5RbCHkSwm/OS5+4Ka89XJM0xcj1bDrjwx5csdUaPYMDQUs+LK
ul8B6Pv4KRsaqFaFYZGs9koO6N0BN0z5alYZYnI+Or2qYZJj+fmCy94BlzxPNBe2
vASjqetz2aR0+tZlVRbhl9uT16hXOPQJITmJibkzXQICzKqxZWybrvLpEte0Z09k
S/brL8KQKr5tayU/+5ZqM0TB4G4YOsgmzvKezSsnWOwLWq+mJFLtkTB3L4ew8AeT
jX/P8BiL5B6NaALDTdRhFfDKHoeyKG5n0+AkxD6mWwju8zlJtvQXAkd5FYEs0K7G
V2XyR8d/4sxyR1qpOEu3/wuAqMqvWVrqasFJ9a9cuV/PE6nzjUO/PLdLMxSn/Pp5
PDhwdW3DOdoSe4qvoPM1UIOb5eKtUmLqk5LGjLIi2cqoNR8PUt4rxurEkgf8krHh
3W+9zYWtk+aDZd/0ViggGXTmEZTrPTwnft3Z2itYlokIBkuq1QAP1J0JWSI0dydm
Fh81NuuSsIP2tnNYATG+a4ZYIXZMWrQQZFUmTv0xeupCOxWurr+ohSD4JFHD8His
HHfBDsQMIHKg/6jiWCfGV2vW0dk5rV4WU4ZR3ySYilgT1xl3Nc4/2bEFlDyr1bKc
D8Zn0L7tZ2devVt8biyQPzeuE2b+20L19F0/BqPrDPhGB3HdMhC+ikF2wBqnvct4
sLWAcigHgpqr08sLf+fxoi9UFqDx9PPeqK6AgQKQwkW1LfuEehry6og63xaoH1xL
Of5+Flms2z9nFkMp+wH7UGtaGCHsqwJaFknnTTOJkAuzf4Cy1jEjtd1SzAzMLM/h
85xF8lW9JAD6vkCbGosuQTdt/58KJndWfLyh9Vyrgc5eRjs70AY/L/RgepFZcQTq
U9cWtOGSqQ/YYuskdRyJK4BYWXdhvyLlxFh+V5UPlKo96CYlhns91yu0wNopwjpg
MhX4MKbu2tXb1HMaRR+0nDc50PDQiGAYKoEfoUDUDXjP4EMvr7+e0j63fyAg5mPU
eJmHsy2qeHq28jn55smNN+jO4IOK/VwbRCeetZKCezwaPizkFpT5navkzoamVf8n
NuqTSMD9O3hWcvw4qIm/IW7yx/wACCJvCMRGq8I+9fq5qSpL24y4TmUSDI/foxwB
9TahmzDDjlP6MMwWkbHsTrMSKnyakRg85iLewg7xAzHOlwBWwUqjMSiWX5g0qhqu
0CBlBqBsXgijDSPI6vL9wFJ32WeeMiFklFdyvHJpc2pxmcs8voQ2rtqYdYVTDeKD
9+9nyHx1jAfEr3rwFEaGMLfmFgPvN2PJEluCOMXRh3EYNZtyHkSo49GEOIfT0Vb5
AiTgXdgv2LvyC2bvWIzVNCCC4qW0pW5fR3YPpKzmCoZ1nW5M+9yMAKWrnHXLWSrx
DaJO2n6rmXM6Miu1ZYt/c+pO8kd3GT3UuchqpXMABQJL/WEWRk83S03sx1reRKCQ
1h9o8NpqQ0WjzjQ0zhONQ5N6uCsjXIaOxG0gu8TXiZE0GJ0NqfxC/78JzmBPWZ7W
Mj1KugH+2pATHI25stL/jaQDqpM4qeq+Fxwt0JKVLhaKlSsZH6XYexPu4mkdXfmE
mJvNlHH2Wbm/tjxPghsRNjt5BYRRSgBP+w7nEnVQE52VXumtStng1vtBjw10OAh9
URpuvyQS5n5COcRSQYAhFvxScFU7w7sM6iBpkh5BsPbSR+ApYVKjmeO4y41ipLCV
qrMP4QqrGkqkBoYvsBGxdUGpwiEMi77YhWk02A/PCCdAxWDmNJPl6rSjKrhrRppS
R4/Sn02Xk/vpTiF0Ncf97RywoztEu19/g2ZpKSlGSRHdrAyN/yZAv+4+umwMtZH2
LgNpT36Xf1nRLRKvRb65B6r0QiMq/E+MKhSaC4eb5LEdff0mFOikNPK9pO2oGYj0
lKnmUXknO09kezaHD6pV+dDhXsj9iDMos9hQgkTl2SETp10fda1duoaS9BbWyuIf
MouKCTTAUXURxEvQn8+pnanxaPGPbjpbOeyegYRa1p6FBItjCBLLPQowh74DGaPU
4nusbrOAaWLzvKd8BVQ8IiLSc2UZKN9rRxnp3p42/9nYq//Y1jmS+vlkYHl8NTrQ
g7PYsTf+3ljpuBVjqbM7SnEn92lsTQNiitc+xRmMSBozRB+NdeLITN4lPm8EgYk/
26DeRBTOIRKmhbFusuz956WicBvmDy6su054x1nMZkQBLixFeOWYjz68gGyyFWtG
U/Mbh3fY4/As6E+LS+zW1S211jogna6u4r7peGrMizeBvaWsaox48NKQf80HVMB3
nuy98G5Stss9VRkAEgo/FxVhr2tzHUQiM8TfIqpizAJu/HWoNc8Ghskyk3AuLMmg
zHzjpS2zK8ZYAsHnjLKS8WR+ZONF3CRhC1C1nkFY0J3dgbAl9kHYPE509La6i5T3
Tv453DuSWTOHbYr5MzvMUb40yuy7RlePrvjfvFQt5EKcXUrS1HLI+udggqXyYKV4
TiyN3M1g0YGcpRtE/ctS9//UCGnH8FtsrISzhCm59/hJIbrEbkXN5NqZgBwoejVx
C0PY2c7YlHPzW4Y4NNjV50ZIH50rXpTJ2WO/6qPWKY2MkuW88DkeTJl3Mm4KfwXm
fmTbXOkDIcDV5Qqp7MYKhd7vVR934TJTMZy4XH3eTdwdw0wsIl8R9FuPDRoqXOeF
etRP9vR3FnXKf/0Rito3fFZJO+vNMk8gJiquaWXIylhjoFcbc94w0EPaaikbimgJ
XCPWAEWtvsNZ+I3Y9ppuzqHdTpBaURvpTRVOOKtetIZMTBgDwQWkUE4SeOHdqqIn
+Ohxf+ebnRVl6buzqrL7Z6qKxEUt8pJPYT1r6hQPWJOoE8ACv6NHp82yvIiO9XvZ
vYgro+s7kZnDq53SODl9g/TVvFFG4UL6i7d7FCGZI0cJ/+/nLBIbscPIoDIDvwCd
ggKvQ8JxbnUSohF0Uy1f47/WQGsX3q5C7m7WPV0Mtsqslvd0q9UgbtDgkZenlny4
vI305M1lDB0IrAUQ5X8E0iPOFbVmWX4dwZ4JBdtKQeG7X8taXz0LVJYiQcV5bE01
CXA+DeDAHdzz87nT8KlBKQAUrtr/b4dVPn3ciiPH1M6oLoFE+/u+RVwUSMrlHaaH
OUEsMIWYw/8T7nMPMF7eXW+D9v3oQJYG5XBNtM8P+4FH3qhASbze0n6uYWGiD0he
K2gMNmVZatRCXgRYDKB7jY2wnJHSdiPC4lsGfvvJznhPUd4uxFwUXKj+klWieFHh
9GUD8/xjBVXfuvOKk06+0dMSV0LOtf86wEIly2CLfsnAw0k8rSFm1hH7QO3vMJvT
Lu3lSOVMvN1SHDZcWirECWujXe6agGcz4ehmyc/DDto6qMoes04qbiwePfSKpyPU
qSM28Kx5j6DIMcnOy2LgKMOqBZHJG5lhqx7kPJ5OGJPOG03APTywxQGNizwdCQBu
ah8m+ZZn0qc79rKExTGYo0G6NAl0CXpwOL3T/Zu7O1uww+96J+PlK+K/tOIOogW2
czpw7bMj8tihthR9XiUY+St+oSPlXs8B7jV2Qlj4ScIAZOeb97nHfvqg+bvrmnUE
DtYzc1uuysW++f5QSN/saOsF9f58axrTF9R9TuRCUJ5Bi1x9Eby3OatMJdAlcbAe
wJNQYT56yBTgn/V6WuzGGMKwuHxJfphHalva20Ala7FhfZV1wJysp64PqII84frp
yYwCQ/r1/NdfsD0zVLbET7v4uxb37jlYwudYKytmHYVhWOsptESh+HSha6h7F3tq
YyB/kwXLBNbLqpqTnUrzt5Lx1/ogdohUpsAijzaMje+oOYUJVS4aAPOjRAboIC2u
J1Bq6nWIEcLfs4sNNWtaBAR5jQkUqoz7E2R+ygXOROx1rVBHzTvlb0ekItC8KeOX
3imAhn+nbvEBUrng18KRXyWWMBmyIrSpyC3L0VTSLAbFRLw6/oG7AgRm4FiF+vhp
qb6YAKDNF744iVmWxGSOz+R486gpvpgOjd8fpUEm1mii92z4DL1CnsFm9Etp5WyP
tBINSK04im/PLVu0OOoA/2ZyoyG0at6HKVZ+k6GCDtGT90RXTOO+jl+3fZQiDv3g
HDJ4gRklSOUO6ZtNwtvvmj/wF0xV3Fx+ANc9Rpz/S5ipdpTmnO3kCwQSyWMvfOKd
1TYszbOFCOJqo6RWmVpT2dvQepcJlGhzyXi7O2f2wmxJP/9o4BPH9i/OkGxx87lI
H0vh3DRSx2MyUva8EVsacZDwmElxEmhUY733Q2+/JPchFYNCqo26P+764N1Yqkis
agu1R9NoMj2YiJTQ0B9u1i8NIBseBxnKzs51Dm7D+SJH//MKjttxJPWFvpW2UwH7
hUIjv+7+bd2dWDR79BH0lnJWGx+PHQO863tP4OvmLEvEXm90K9c3+EHlgDcAvLmW
vzw99wf1cyQXnbm1Tf9rcexp65ieB22UduWC1ttn0UM1zkw21EWm3szm0jHK0wsF
Sec07usFSzqGHDsw9/3suZ6uyEJL2WueIC4mJYsb0jUwaNZsaItHeOn+pbVmPKT/
ZluzgICZ/2MDKrMZF7MHYvd2H259hyxVTnWrHYZSEo0OBl8Cj7KGnZb4pKK5CiLP
PvafCSQDCN+2RsAJMp3JtK7yN2AJYu2GdjmkDxwfhISt6eQvsnJL3azbfHqOnvwr
Eh0Bask0oa5VdL9sHCAYbPNOiGEQluUFFMwrW7vWL7+iQ9qtbn+L0U7CsJOvBuUQ
S8RRGgpuS5M5T9XYRKg4/Jbw4nlqXtbZV0ILUUkNSOSw2UTuTiDiyC4IPPGoHH1v
6aTKKJ06bOhA5cXsx2V4g1CQUJ7wknK1Z7syUwoHGGdpAV5jCDpg39jTI9FmWKHv
+tdEOe9wKNYJ/iZLP1hBeKREfF0ezLUfu9PJvNdMrhYP7tHIoGy4YG7WEDtoHb1i
/w9tt95O6kB9P6xUhKrA17zvOfJT/ia4oziDXGlrZAl7Stbsz85IHuhEC3Qyeg6B
+mzIBjRjI9AOXIuDvRE44C/HrP7XSNBt8Hnt1Zw3K4TIef9Q4Ipi8e19jy8tJAUu
v+W7tEUvAKXA0ih8GiAtWXBpQPNn21aBsoTjFx/ggr9iNHzKZOUXsyNkX0k+12cA
+BgiAMyLG2+wX5QUathDbr/A8KDnMJnCjaxtAUWEuDVoBY9plBokoWERvjWJl3BM
0P8Z4I5QySNoFvsWyuPB/uMK9Bf2b0bsBVgGFvur6s2UTjbItvgVzJiOEYKwIX9p
zWzwWDJ54dfcSQBCMVWSDnEpJbMM8KybE+I1jMSn+hor1rJDDEblVjo6B/pHh0Ke
SGWJrdFlUS4hDiNEjXDnyoT8LmwvXVTWbZLWxe6tkLRsHZuwa09uJrE19jko3y58
oky49e6oi4PFrdHzT07y5y0pl/mDWh2xMtCv1XaR9P+fRkpaBJ78Xzsq6zHZl+ZY
2OX0YqTOC6YdN+kXgrHBiIUstKCbv08wtHJQlPnA3J0jubOzndxO/1nyDEG2LRvw
X7W2uRNGNeJ+syIGmSAWHCIVf+hOWPU3mEH+x3bDIuY03zfb38gVYDZAkBe+agzf
sfWOFNK/0dn4Jz5We5cZxhEKZGXQ1xBxIJZq4azb0UoPfggf770dcj55M6K03P1H
lteEbm++NmWhYGfMzfP4oC589eGSKWAHEQgYo248ZQcQbpnrjIWUUt1c0g6v0ar+
t/ap5IsviX8zsdwWmJJWvvkrrxwkXkEhMJ9p2ugXgAP1FoLUQyP/G9noTBiBYdho
b/jGqv8p6usvWQzonCz7JY21Mc/XVh6VdrDvILrLBf8WKgz3A+g+pBGYPfrquF9h
OFunSxDlDgDYrGJbSUv3ANjLHi6dP/OmXMQhO77/oMlQtEVyqkghvrGfojmRRWcT
PJcXnXDYhplcEtl9mhIrpXUlm7GbastoEt8h5nzLNf0/IfOLl8LD9KNJwy/RYD3e
4vU20NBXeFgM7OF+I86cJySNj0HJlBxMm54cSZOatFb3g7tIvSCO+h5Vhvm8IDro
WRLUVVhVS9z4ilKVnHXkpzmeeXNawSqSOJjqVBOYtOfKL8bNOd0xFDQuWbZn24Wz
aj+Xssu6kDBkIktnKPGp8eCvuQaJBdGVYnk6XnvZeuWtiSQLeWmNOdHK+F6A0TZo
LLEjcy9/1x4DL3FYpByb7eq7y1faM328mORwG9yuTndaZoUh+SpkdgFL+2BJ97V4
2/8Wa23qzp8BxyRPOqJmA98YaXmKLTt6txkdSqZAuzONUu3cxJ46Hb+d1pa77Gko
x1Eps0EIHClFcw1ynFhxz5o+0hZg+xlSYv63QacpeQiov8AXE/DV4H8UszwqkaKK
WIv16US+bMBgW5nIiGloWwN3vbBVkI3s4dxLMhB0RRVozbgYFU3zWKlIk+XHNXDJ
X7ExlhkwjC6yL78fTFvnmZXjjvdBLrdk6Q+OeiqjmRWOsThLRMHr9swaZNH3HMm/
iknlPm7rs0XGsLVbaqpXdgS2DDP2Jb8T5Ys+wNCKrlNX3xEWG1kCu3t08QxnINQ4
qCqjUy541w0LkYWTyqsCJYe0iwLqgSDZ3KsCDOG3dRsN2MzDmcRiVDZHHfgbg/AV
MDVLFMnRHC4e4+sMMJli0inEl8ZpzG3qbsGcKRJ7lbpvD/mFtBj8z34veHmGSsE8
1LLG1kpqqTEdFXF1DlTpivdUpx63+JgGGjlZu+3EBOrhd6z46fiZhgDiXc7Y/dNZ
bG3wj7of/nEc8Ax+Awons3AAp+61IUWVhg8veNJFU/20qYe9CPMQjSQ4tFFEk+6w
fnEKP9AjD0VmIMi2MVx0fR+kgDeSou51ZKZRkS0pzTs4uxMFz5G5GQ46U4ZJ39pE
vdhqT1L1ot1Ln52wJoM7Yms7JlRUhLBewukV0o0Arwj9EXEw0VP9Pkn/NQU5KyG+
iA/hXZ3GKr/OO6g0RwWBTDiMVOWLbKTbmhJCmY9RHPd6Zwn6Gpo3tus5X5doaoRR
EUIce1vPIOLPEP/BvSKx8pPETq5b1u50DrPfuEjUX+vhGXg5SxKTE5vCeRgAqQTt
dJ/vwR0geXcJuvmXflOwn1x38VH134IkcdqFXRUPIxY55z4DCMrw24BnpYPICV7n
vMSkl4PyxR5TzaL+hP+96O9fXUBRQvim4dG/U3yY5XqX+C4fgGhYyNSSz9tT9S9I
mAW0qb0sMfF0VF0fb0Sr5Ixu2ccMzfGl3GolU5vadPiMeQUPiEx1LEjCRG7VMtiF
cROlBPRmOoMxVrKz1jauRL9Qzp/AvwaAOAFHjmwO0DNXs5mXTLkPOZNFbsxgXjEy
EPXZWXx8Lfl7wxIYu6ocQM/StyTycMrA1GvE+r1qL/vbsFho01iEJ7rTSTjoSfMb
HmzYjd7poKexh6gGddci4ROEZE3ZjLJcwfP78Ac4d8Qq0KYbLtrtjwSLQk0jXFaF
c6QdF2F5DbOp2oQmt9R2u1lgWZ0Oaj8PFbQir3Tbr08AboAQ2wXI8+haSuUB+eIj
gHV+iMvRX6qy6w3dDYgwSkxsLXVB4sxoZCPpDZGdl5gHEV1NdFMJp7Es6sQ1q2wA
nRZycNQTsyZbqOK7wkRVui7fW+ptd3do+NP9ajs51E5BuPC4vXg92koGeLSUihze
CKLXg0pOJrfAdvJQfgi+pNN1XjEb1dmtnJejDN75f0IbX1UtQgMN8dsPXB1rkwiA
geMuMr8Z/7VUw7JcVskW3UWw7HJC07mAqTK/Hat2fH5SC92rIpli6H6UZtfVkAPr
zVxDttjqasMZrelv+vcsqR7bD6iKpILvmpzaXCKENDTRrYsftUeHPWfgG3mdxm/l
YWjXk3Vl1LJhi2QSBk5BvmBzzEM+gCYOAo4Z79g4VB+Li5Vy6pRlxQTtfKOXOYaq
MvjFp9eW1XBQK5IubwhYJLnQ32ol5D/mwcj6oyOkPT1IQq/O1T5Ov1pi/PqJtBSI
jIfqhjhurAR1lxffnryk8B5s+gNP41mPqeqHUU9MfIiaCNbNmLC2/9eNykImLU/y
jUFBur5C1av1Sfum/mRcpzYAzoP0ZadbKmQGQ4KyY+O5kk/r9thekah4hecLcw1m
m+5OkU6oMdX6ZG+9Mc4dKgbbcHk1WqX/358TtZDhOiPqzRIkwvwHfxQKDHHq6E7h
RHGfFG39S4CCJVA7feWHVKGtb6jqpsmPBJdH8oZ/aZEIpKp0lZL7dyIb8veT8ro0
mxh6ca17QSw5SrDB+VlVKxWvU1LdKBlqlxzTsB7oSOYSy9ElhD9KPg9XaxMNhXwK
wQKPWSe1WsUI7HqLC0MvO+N4HXPCJCU3zfCDMJeevpMHHvHKI78rtYLS6Kwx8E26
xKIbsKU5t4lyhLDGuoUR+CJ/McgpCJDkkqklrqSXzfza86NAcDi0/yljL8lzlKB9
gUBrrajew0SykChOSlmiPOTuoM7LuydXsFEXYkTPgb3xtAIqjAR67QH2uRjror5n
jG7S60+0TxgN9hCumLPDchB4j9f7n5hBNpqVdiF8YVcuBts/qt/0Ehgu7/WT5WrO
0hs/kBXIUnIeLCCERgajev+fiz8AJplYVmcrtcpKSwbw5+YiZGXuzt8CcBCS9k+z
g1wf++hVmGMnuVxewUOOaMOJg9xQMc3JYQ7SwFgZjavXD1qi0eT5SuuCBgvQZGht
dhrnuTK2RyP91F9WgcairuqaEnw388mAXqactJ4OjAjZHcNPmOFKjy5VCGRs/vYz
PhcKAk1iivNAX1csl3gFGS5wGneXroGr399UY1fxcJ2z/Vwz9SQKwOx6tIGmOkNZ
y4uAHzDPlssr6fXEthE/eIzyuJT5hEwPQWfUPwsiyVFAMeUWEPg/8cP9jTZclP94
2Ua/zFAyYp6eutRfCadG/3Jp6/thl6E0locw0D6gFIQbnQT/Pnv+SbAk3+q0Gm/C
L5IIanN+E+C/Z5g7Hjv6YlWT1oauD8tqIs2lJ5IJ0M4/rcv63J8gDb9LnLDm73d8
fj69OJe/GxD6drq6UZsYGrXqOizm8nJldFdPJgbMfUB3Bn20IMWAlB9cuiF7E0dq
RNhvLnFr5qqUu0Xhq6qdGlsvtvemul3XmsTl5q+RiZQpUnBay7hHEzQmqfP3BBNp
jCoe8sKb9ZgT3ARyXxagmAvaagbifRJg+0mgK0Fi48dwIovMWXwWCVulMoPh/oWi
QjHke9fHQBt6+VLXjxX1iz7T5bepzvk8AqzTEGIswddMFnW5CjaklSCANny0VQod
y/mJzoY2YY7Ec8Lu3PCSiVbGw1Vpb65DO4FpI2Ol/L2fd0eGO5Ln2UM6q+Jqm7hh
EvPatq1qGKJazg1OHvve6L+rasYF5ljEG//Jonfhl7Rb966kz8etD3jEjNI19FlL
IIcveeNjalpnkwYPErrqHNO5vb5iGWonzpGUzOb5PiWSzSskt5CewfbqDf5BO3cj
Y3ez7RYw8G1PU+/GJ5q845BmKiNTn0h69Sr6uG9WTrCeuexIDYaaSy9LSVgqCu32
0mWDhRYM0qPgDQQ07jmqUAuyuZlyE4TNfhxXesr+ComEIKTab2OSvdeXWI+4kclv
9U9oSAGwnrvQycZihpAvFubkSs/22GEFKWP3b+u8MjYNCb0FOqnB7pIr9RkLyVyr
BthFolg7goS3zEFwc7NXClWLG8DvIBiI2dtofoncFkvFM7sv68rdKCEKYyWSczqC
zneWR+d7n4f1NzHUWEI4JvpiAlPxr9J2JCVlHMjecEK58qxlXKMWEG5M4D0aQCS9
tsbNSDt3cMGOVjHLarJGeFu7BZWh/Ck7o94G8oehBzPZlLLcryIpdpNAAa54Axyt
E7Z2trUSSP/FiYLbT4hLhMXWqnMrta6q2WXRvzy8p3MFkl1nKIFdL2Pbsk84rY5c
q/udx0rR0eIw1QXJnylWySjMno9zRzYuQsaOIoP8JS0ZhPYdlmuDguY7R6KGIbcj
XS6SpLoJJuMdWnh2WV9y2c6CuufI2iX9AYdp2rHXAbbSRYpGoGK8V8Wj5Zn3Spr5
Zm4WwMGc9Gy/TbbckTxPwQPKA2yvEJdzbZur1CLs9J0BWi6EW684l2ah0a2XiVJv
xzV7tD6fdeLY9r6X+uweKYIM2Kzv+gzoq/cg6coek8Wdgv3tTsjWwWkY2gQSneGm
MTVhq++hI7Pv5WHaiLZayWU8A43fE4Zi50VDDWUz3Ny0SJNAxtwN6N5o9sPyiNnO
68+3xccmceg0bNMkeQXn17Bvy6bIu7GFAMYhXRJXbODKz1a6aULdJZJSl8YsVURz
IoWocWT799OHDWidGbvDPV8ebHmHgz+7IW/buspJWWjny8DzQ8BNKKhmtgSnaiah
RqfVAI3z1NXlp+IwSSpW3/1NbGWes0xS2iwTonhBvTXpw9EiARtwVItM1MsX79sd
4NrEm6Th9QDz6QOGZBeijZyDULPELX4DJ2SuDoSIO3klUYHxtHlGC3r8h5FDzqKn
/HQST9jDOhv5XmkUOd8avXh57xbYOm1uY1ibcuGX/d9VpyIsMPhpnauLQtTqpIbd
TJl4OS2EGlRRacDNyBpQumZiJrgQJE/oUllz48g67o5O78JbSjTupZjtA2EVUCnv
jWKHNTemTkoLcZ6vbfvOSonE8l8o8V4QAPxOeO6H+pcMzQDFyeJNRQOqjXfI1UJB
NyVtnQugaACYGOs4ZyRiotL+KNuGXjH2be+dUil1VU0zicTE7wReK7MQqU4RznLS
CJWL5Nci5WRd6IyT++s0cPBa/WKj4jIjKY1756tXJjdcIOaYl/E6oi994MllHGBk
1VYjD3hTGcAPxxuUwaul2P3iTGl8hf568YdrsGX/A4moPGo/OPD49i3VNJe91zgG
/msThX8hJdPoS22cAAZjRBVgou0uCpvRsQMTpkS8q3vXpjaSTe68SXFCB126mEIe
HSlqt+zsJuqIIZ0OqXjUjpb7/tdk/XqKh/BI28cfF+ZyxWahYAE0wuOB4nU7NxoH
oPyxqE/KHVGqdRKIQ6Qhpt6JMm8NXTNUC3dDzGHLYnq3UDK++mbGPbW00GuCgm5c
v5Y1x0OC9uOsuAPFagrhOdk8kBdOOnPp4/UKsuP3i39AxuzW9nOUgg5dV8Tx94Rs
YpHCi67eydn500TBcmUBKACum87p94CIEwFVFv5KlsDxNOo3UpCh0MKSOP1QITfK
s78ocP215M1cDlsT552GyJk0lrMWrcaleIJmPNq9puBp+mhgdHFYRI2rLPYRHKth
iL0YEvK7vlE2YNG9wfdfcHg2+qWpFBg1gtJJkKbvyzq4FWoJrlrj8DPVYunH16Qf
6jgziCgNjANxRcY/KT3yxB7wM2xWJxX3Lq0QA7x50kbxCFmrFvJe2xalJbnFz0hB
RuQjq8HD4Rig6Aehgb2Fm0w6e7dnqMFPwMSIrrj1Wloq0kZloCnnUAWXNnL24GYs
K4He1Zm5AMUqQ32rSHg0rvDrkFyYxHjIcEszF9XnBhTJsnSoJ9wxEpGa/gBBkxzJ
Ixl+kxfpXXInPQIWLJLtSZ6sKqTGfcXJfa85jeuFdsiwAI6NCf5cUS7lALAlP/gx
P0xtbkfnUG2E4M8a4djneQlVMVRR5pC6xXee5r40Eugonv5wjslvZIXZP2/yA6tY
f4Ahydy+wy5FV0AYqJ5+moQRcMPGuK2gGDfgYNCCTPt/+Q3cSuwXbBlczI+ijZZt
jie6i3JY7E0xaAS1qIvx/RpvSSXRlghRQaWxvjFDs9cs5Cl7IsJUVa5CgdT7tQKZ
Bc1BApySwsq3kl7ZBkZxMH0KPlJ2fAN1L69/iAkcX5Um8ctqkIlg1RQ92Ek98Yx7
3m7nIxiVc4t0Zu3kjAy/xp2jofw2b0zF7NZCqAvQA01nSSEFy3FncXDKYuElcxuU
CMTyZoBL4jKxk9bxxfQb6yjlAXft2bmljH6FHfXpYQGJ3/VG70YahXY9GqZrHoQW
kL0CpH7MkEfIUwI+t6kG9Wmp3SOLDBItk9HzcxelZZYYLiLuk/2/+ebttYoCnDG7
EJJMCV7l0iSIP7vDwou38suniIXuULLyCN8hqt7G+rrIvTO/mnoE0ZoKL0bgTXOZ
tB9ZbhE6zf0zNtcVoW0kQZtyQ7ug0UzXe4h8HkhIFkMvHk/Sp/c9rJt11x9ibuqT
PaK0rJrcZDOQIHrP5KuVK5lk8jc7CYZE/5ZHnwkdqy4fAAV9x6HXOPBf9hjCyeCc
ma1m3FWbs3Ly+GLBVX4+gEioAqLplzuXQdncMqqzm9EF/iFvSRTX8UFybuyspGl/
yzT6Vcu54l9acc7ddBfKw8KFjKwlMBGBCMbz/tcz49kC+YGcQaYMj/PaZzPNg9fc
0cTmXhnA5OeCSSUALFOmLu5GaNU2LNbnB8PB4YgpUoHzkeLaylKa8s7yWt8oiH7n
PQKHA2xj+F9xIN4jxdvqF6dnpF5kwKDRtrf6hEgx6VvS7zgIFZ+P/9nRgf46IekI
s5TOEYQUQsGl5OkVNxtLcXMFYe5C+kqqLBj/pGBe0JdGxRXoNdAuzJVZtWRTnfqy
FvwN4e42eif9UmdaWkphGAYeEmd88s1xGm5FYW/r4klqrLTMn1bLeGGacjPEPgUA
9ELF7qj5b1Ou0wwb/H6K5KlLDqukFwVesFWHV5vMuK7Wysw+wZbUb0xX9Os29tPg
feMbrN6Gw+dGkun6ZDAIVDktphsmVloOPdqxIBfF52WCRE8zyiYE1G3RTX5oJo4f
s4ARy0sDfQvPfK5aY4A9PexHfJpFwGgh2H+7EGn53betybQBwdqA05LeEtmlK+12
k17oDMqPHEvh46N9pfQP62g0X+9eh0iXijaakZFgwiCWBGJ8Cfg8tUNvb6TxSImK
i/7P6sNhWqItUHkO3RFf0YAmSpVSkcDDr47cV8UETa/M8SHFDIkQDaPr6fJoodfQ
JjLTiE3eCL5gjYK5ml+JUFNPDM3yRQmiUuRJzchWG0WMWrPrCfwn/Y9Q4xzWPTA7
qIJaKHUcnyTpTN/Kodb3URxNOwzUoo2fY3pX1Gs2Z3nUM84WzNpZh7pHG2TZoZCE
neN5Gvpq+jhTmFXDPAcs5Yn2BbmWowA0DmIkU612euq2TbYheGu1T0Kiz3m6n8OL
dyIaL6QiNuivfjWLc43TEAZRBL9+iXrQIhjXP08O3iy/i8JeFB2ieChZ/QFO0CVh
ZG3KdU5l9WCl6aD/3mlJF4bqFFoQv8HraSRzDu2nSbhjnciqSIl9QvOz/NjjXh+n
PFORdkquIPf//mGzDiMVWc+G0SlJ0ZOdQ9G8FEqTmurL01uQpd9LgSUj+SXPLaxh
XA5Hr7QM4XCHayRqN8/JdUuezUned4i8w3OY8pD1DTRcIa9q1B3HAXy1x2LyhDcb
FjsWrCMNOSbmqb934Txqc9EaZOfhxMyNRu4sIhmA1aHryNIUIpELw7RIANW+8EtU
QR1pWFrwjeEuY6SbtWqvnCqMeHDdPwNS64vOJr0rwmeauNzCgNAHm3RKc4bePy53
zb/EEUvd+AfCE1kc6CXXzCkWlpXel116ejMKODhs+tTZWneu0i7h/1WWL/ILilO5
fvkxQf1kQqsbFpB3td9x46OsgX1h26dV2MlK2KSe0UntR2Dot+UxeI7A7nlwxMZQ
UsLz6TwHvAdGxsXMrAEq7Pd220zuDa9XapOPiY9HfvHZFROrSR0U2Zu9hyXHzGjq
9KyUrHDr6jQ8EO14TBbDzH0/0HjVzATrCCE8+B9fIclPfcQEc0nBHgYPaUcmDpD0
zHQDr6YI8l1RYRt5aea+RxOyLe2cpTW/2T+eZE6HdEGwKIEMxVFeQBNmUtK1oNYh
Fe7OXsG3lfDszac68tQ7Ob/FAa3mapLufyohE0mnjohOGCBiTAUn1rcAtAe2yZtP
oBPPfcHIatToc9WQUVha6a418QoztMKPgebZOb8nEpLOEG39qkwGixT8JsdVyq88
KMbPVF4woyoNZgphIDEnsjg/qc1/eIO8+fx0rq5oNbYR87qCYQP5ke6orxvn9LcV
x1uXFfmAAhN79fFb0Ivo619+TR8+gE7rTwIZt+OheK4twonwxn6R3ERsMMbaauuU
AM8H6vEI4+iyC1ydK0E00kEULBn+3xDT/L4UOk39wIUQOR+ZutRv/h8Nx5nKeFt0
qkctcUo0HxD+BYu6a18oo26ZRH2vyH0mybU2Xt4YgKN1XWViyNGhgGh7KilO+Pi1
yZtTGPQRpxk0ZfIFvqgGdnoG4kJ6QnyySgybOKjbCAfgyNAcJ2+ug795oj/KKo4Y
O/ph/KMTCPFxr+fO0VnuNHGIhpzmmwpiwQiUre+cCJeyCdtlrR34LBaIBMN6yoBu
Bhnk0++WAy59dKVryTRhfWXB6kDwKhJ1X7roP5NkL9DzETbnO3/4p7BnEUPrmxr2
daTJv+CvV0iF25yhNm/tvXA/IUabAEHVfpzPQL5Dcfvez+2Nb1PsXdBY5i8u2l3+
wvILM0D7JrviyvIemhkt/LOAy4R4b3bA5o67Bt+/MsY1TBb4QrAenBJjEZ6zOSRQ
oaomxDj1lPOqoGcjBeLGfTNDCd9C8cU8lLCxU0oFmqibVL8EUCiBg0GsVNwy4yQ/
jpnUANovz1IczWkHzwqswanfo1DooJdlPZ4K3qK7I45Lzv5A3rpb2A9a0LbMcaW6
DyEB4BHQSvLzCRFJnP7MC3ExM4TVwaUtzZ2d6+0lllm3iLxyPrRNtK0gFx4/mlEp
mOCZh4IFWhBZNnqgHu5GFj65fXWdLuhN9wDgQcJlMFZXsSTEXWN8kSXIiyIenGNE
BrQ3hMmgjPcNy0wcIsAXu/U1L0opdsIMmvg4fEEMP0RPt7QvNL+xLVFHLekVCvlM
A/85/3HsT03RdMxwNplThJKMMdXLsK14AuYsjZtLF27LNj5kdgYHmS/CQIFlQEZH
XpbppwS4v7wGh/xOXfHWijFbhXNNNIe96kKvsMTs5ZapTBG9Knyx55w6OghZfEBE
KaMr925ROHkoarFpLfwZ3ref51d7q2gP7SG3gSqpWgoB4jsrX54oLST7O9Bqy8QJ
VTsIo3PDciYwelCL2EQOJ5hopFjHu0dmprVPrOQPrGr3H+SCUvFnuTaoBIuBR++b
2BhcfpqC2b0B87TuR9GkiX095Ipw7oviPvOZkeUlNIEYSAqoL7ozvfrSwZQhNohT
fYHT7VMqtMDUsjBpujlToQfcBxAEVzEDqhCL/M5t+wD6enf18Swbnim/wQpcCq9g
R0pi64PF++0mZKr00z18lkhadB0BCg7IUp7tWV4PnCRo68R+QHyk3I2LNSJEl8Ao
/giYVzdvspJkN1qSQIHPl0eFpy6k5DMVQbveanJYTGCnYNA16+//YQB4clH3XLYS
bD1AaswIs230kUigRznu/4epj0vB1EnXPphTdv+P8tvU3nirumIiGOXaNAe8V/tK
MFZh1oKr+zWcw/UWuR8gWCnmBGABNKqDWSx5vbp6nd/gFw/ogcvQ24hrapSVzUC/
T1hRHRZpJKLRHDPnLYxM+fRH65BFwUrNyhcaaLb91XgYdYVJVq/rnvxwvKA5LNXU
IbFMo7vJs7fM+gvuHG36Gpm7nNn47cp0yx6Pp1gLLOs697bu4PIBcdLm/c66UXbW
BU0AYLXcYZ/IuFp/wACWZKJoGxXS3pCfk/Vt9cmr812+Ck6BIbqnLuNvdPW9vO+b
X8JVLDATyI7RzO4dpRRru4GRvkQlQrNYly1gQoVuqmvpWNXWNyZ7hxsi1j2MAc9V
S0NlglqjyTDVniTZVTJXkSx452I+gwMQh6vq4DwD6lQtT9D5lgZRYuyYWG/puEug
6UTiAnlekqroOMFeU/731tjgC3nV0Gzx7aaDqtyyIQ0tqn8AjZ5LWCk0VgFNIq+r
cf4N/CCjop+jL61gUrqyW6XbYarD4+NoymV3r6Rxtc4O/PiJQ0X48LwDqxz8/5sc
oy1G6WcKlRnE1jLss+KTc32yMdInHCWpgq7nyOCODM0+GaWZzwmnbb2RhwgFVMec
RpDy8sTuZ1w08rO+VzhM0VYr9k0jkpkUopr4WvkVyDllVBeN+eBKJBeNp/uGdLxn
h6g7NntZ9Gy6u2rHrtrlY+CL544BYSpvFe5JAsL77D8RmR7qbrF/SS7KgZeE5X1U
NpfHe+dqwXbGw5Ha8Z0fbyaLT2/5dYKaCksybpG6rTXuAjPrf//6e0T0zOrVO1Mq
Z6zEGDdnSRHlnbXpToJEjcYstgefjOz0Hr3yihm4KpGxu/bTfV68CZFgB41y2CsF
7/ooJxfiDYQzazcR4VGqZUIOaOdoalycdXvG2teMz4cAavRBXtfPN7m4OuZkYBBb
pVAVCMAYPtfXnCSaWT4PU1YclvlIFa5MxUbDvMf7rbFaUtL1dcK49VM/am5MudvR
2YKniNIM348Lbc3mhHdwO1S8Re99ZGkL3RCpHwkLorkJfy9++vfuiEowJg9oYKDm
q1f5bANketCHVPfT7dK1HvuIDbnYhnRHgv/srY7w1dYfVtxIRxOFgs7m0UqZvqr/
P++KTLJcUfDjWQkdlzufbMqVCAPxoZ0AkjRytfh/6vKSXJEQ0ZeO0fCepuR4GM2Q
uxGnabKxL5b+6hpQ4hXbscAI1mqYCW+k4GR/fQQwmyOLOLL7meKYaVklFFrHkdpY
wNHMgcVd2Yg1C7AfHoZHqpAlsJyLGzzlqcO2RkVnLgrvLQCE4mbHADuOj6AZAYzD
6gxK9Cy+boZHKjc7J6T82WKQaZpTdGguJW9cs1uVGiONs0BB6tpapFZDtMosCRFq
QPKrMDL1zgrDeC765pmlC5Zn01UK+//OjHCUi0CwEpQyD9Se/PWyFAPA7sOQ59cI
/+lDOehxLtnmsmW7piFLLvOBYJfPE0o5QMTk4FFsND58fk3s1or/BUujoRbZxAiK
nvcyGeViMVeVJomOEMlWeOqpdCLAiy1A+HrxlKuN3VUVFVZD3CVSu9StprLlWSIV
0SuVfNWT+OcmpegGuMP60XE+1VkNX+YmdZrXjnwGRnG6Hr4SoN+QNAyxhWDSuUQf
+PxqcQ7XuZX6YyDB4qz2WnECyfkrxYKLQ2T/jJg0tH3YuiZUwGHLVkucrJeNumqz
kPZWrCLP4oonoyoKx2zH4YlUougDGufhQFJiHoaBsPu4cWXiNzVojl1YGyKHf3Es
vMeJdxhzjCzvS1k8mRPTa5MI9IeZYUaMfEbv6+wlXBLO6c+IqR2aR7q21k4IEc2/
mYEvtv63PR9fU2pkxAjv+saVVsLX/KuEXYHZjmk6otb/pk897jyil6629YxIpDLk
bIGOIynlO8OB6jxXcpdvwQgcBNki2G5pEzVRjGOHJu0HeAaSNrc/jY6PoC1nTem0
XTRCDomZPtbWRpYKXpzRXNwGVXoG/nIpD4kVfizhRgSSk3air8x0ygZ/BYhupLGu
QLWmT0r9bFxhPeRte4mO3Ox7mIOYRsHwHrqRoqNt6lhAbIZ7rgJrNljKj3/Cn6wi
m9cNm8fNc4Pm9Djv3I4kn7BBoXoRLG2Q9qFDqweFaGaDrmItnl4aOaoXO21Tsl0r
rtW53ol/Ql7s7pe+YX2PL6t4Iczb7KVOZIBvfzkk8BcY46vQTfUM5QODRfmBZWcE
6pxyWVdNzSxmkMrMtZcmTvtiL7XpiIydt/Wmu3rjha7pZN+iZu45u7zUN2+spWRY
mRLREL/Ih8DsdcTIiszSD4y730wu+0jOtKiUQmK0G5Hfwn9Nzpx/YgM9Dq98Cc5Q
G22K6Xe92kb8UuOI74Ydyn0UU0VhS8zFJHNMeanfyK831oaMVhFzecQq12Ovjcow
fIQb94xcHkIjF0fmL66NFWhTvrM+mUVI5Vv9OtSFxEi3v3Pn2pNO89VTUdgm+klr
mFzt7HV6JGAEaihHZuKRUng4wmCBZ+9Np8A8Xny4jsgEeghe0jukzWoPzDD8quoZ
fE2SAh7WBFEUVjvMIeAzNI2kEfdTSp/VsAp9xWjRyeaBNcz9Efr0B+blpMZV6MpN
e3kwlN7e2qcoZ2erRnYtsNu7PXsQxukd56/vt/G9//CsCWkkk+1xhBevn9cTYu+K
iwGYAyzph8GRyHEElztcQ4nQk/3BN+MDX2EEZAFThsavMx7clH2wiBccKnwHpycA
y8P26JiCt+L9AgfFeDyUs8U/lY0fabAI3nfhN/iuHp0k8Z72re1ZNfb/7r/4FPET
QPht2q8AdjWkcvt1d/TXyMVYQwtJtE8yhQ3zXAA9IODYInwVh1sPMPpvs8z6gsvw
c8pENy6kGdT88qcnhBsgus07+oTHPi85cwIeFg6nD9uqWSTlobbm+AHBmICk5Y3r
p91fd1DzLSnZgMCXI/iMFTfMLfr5TWbiuqn45qSQVdwlyXSV+TiETbBuOo/cK04T
y51hEPzyawYEmLzAsePvvt53XWJDmP9wpYGe/UZeVZ20NaBaqtd9tCX1D6EWsG3V
Al7klrnb2rA8D+SrEmyFfkaRlnbwZsMWYGmv5ezYx1+JqYZ9lAe1WWq/q80YhWaU
QwWMU1PAZTlVv0cvAwrgoMppBtzHetjlgO2vv5up+Z7cNt4NZmb4h82ZXYdtvkn1
ACgEpjlEhQ213XhYTCrtexmktmWNSKlffUoBD+ORV1+DR10OoeqtmEuDat+oZNUh
+W1DkKw7RoMwA7pEJxBtNf93bcFLyAPizmqMJo17aWhq6qAjn8aEE30WLaU49sxj
O6EQCs5g3UWSxX2YsFp6f/gP0VBVArNFWN/GEeOT3/l+GP+3Li5aAHpVCkLRmsCY
cd+FeOjXnwSsqVpaLuIX5t7e8Tm+OYOgI0dZ3J4AzsuNI8FvRssM5/yDuKZyOjo7
PUEIlhTI8JobbdPsZax/qy1Fdf6E2vFsPLGx0UO4UO7Dl1tFFgnPfFQFhdN0DSWk
qmCyDEq5Fy9/jGW7qypSL+DiiKY0E0X/ocGiVB5az8NYoYFDsGf5aJBdNS7gn4+t
gPwtVLBLJecgsM8NrkFbcOZ/qMFWPOkEh7IX1wXI/Z0kKaO3GRTDdhPrcJ6G6/8w
d7O2Di7DCHe94ItXhdAvMGSy2YOETA0NMjzIzqi1zgWC05VdE7OT2mh4KORvjT+X
D4nx7OjbPAcvNbEDpQV1t8/5TYMFQASLKQ7V+MGuj4Fdh5JvzEUQ+6HObhwZBJHP
nFib1Ax4thZ2vKks6BFW0rNonNzPXOUE9cVGbHCgHSHssdYDkCxxQasT6Q0SzPTz
GYm5hmffGIkZXisRspuaeSsPC4RuGj2H2R3Sx/4yQiKs/npEs2sw1PqW6NEhaK2I
KFnavjMTrwtfNOBg67oxA9B5/5eCCqvCpEQsNTh+cas+fEpscS0j4m1AV5UnfEnr
hdDZk0cUqpC+vbqs7oBnVvuCLigewLCVo58nkiT6ONtUyiLZPBj+EVrL5qPA715t
Yk9NYdE0f2Y6b56jurmbXbn/vJiGN7YlJEyYGdiYmYGxVLvRseoSlS4l+a+mXxIP
eVcvvHTrhuxtkqKIWUSw1o3zBNpPdJxHcc5i4TjIJy+XokI/cWl/KyeVzeHUIPIV
UYANtdqZ/26x7wVbrXzZfjMd8HeJS4Pt/Ua4rPCND5qShp0cJBDY2crBwCHOO+Wy
aAMOTdLdKLUE7OeYXzYX2qutE1tE09hwdJwn9H206F4mU0/eMfujVW7OIezpddPD
Wfhma9Z4+E1PjBusJjlHp4oZF11WtXdczoEFkCh9R2eaDTuz8lMsYTFb+4mHX9Ty
AK4ELO/YMTYZDcDx+3zjcldH6+cm2fYJvEUeKFjwg2xbBx9kJk8dpm7CyJ2annTZ
TlUpZOG9cLq49xka+HV4R8Nn+bE2Nf6EGf6gsRhIMiMLMRWSQlt5BIMo3NtNKwKY
UMVuH6BEuVKYnoa2YDdBaktaaK/4GLTAiYPYiRmVhba2gQmVTVJhJsrWky/UljrB
0llfnP3X3//Sq/vvqhK3QCXcTKtffNEkeebTWoV8G8RGjcEZK3zRP16MUVlUMTCv
HL73Q/ukIysCiokl9PdUsspgjuakfBOMnrzGdn1RocBbDsxvHZckRvEmzJapCEvm
muMlw/mSjLoRJAlM6XyEKznJRYmjSfM/3R6aUF8i80wT+j+2stWc7arQLwhYWifg
XSJT9yMK4qfdP/OEi/ImZ3Na2m9mQr+rR+o3jK98e1Nv+/pcJpRIQMRsulmWvI2K
MPeqay7GiZhk3sCjcxjE7O2k/xh3ZTbPkVHxfSN3BgqpkViB+TZYPPAfciElGgQQ
XeR8M1Dy7JnT71xeUQd2EPYziYJMVn5P08z8HgVK/suROwksZHkQBAlJ48PX5LYj
LQFqO0Ei5fsqvPglAUHk3nMo1as7RHBHXrcz7BngZFnZANX/KMBRMU40ebMiyR/D
BMg+y+F5Qml2/Lvfgpjt1OTi7qjPHzwE/yPR/Kf9p4PhH+kurNXHRUIUevD3YgvG
QVB35MeJkteUqCbAEjkVpIhZr45QrtGNW8ZEQltQSAsHzXwwC/mRXDnxUEtQzcLE
uVogyQI6mVVK65a2Avuhsw/R32J0Iit2tzj8WGL0UOJivMENUDo3mqhqECbPVqUd
QB/vFn9wiTjN80RrlvHpOkohbIqZ+KQveZctvJelpj2tOWb88+6lCUUuZUJiUFSu
YH4KKXGTH6/bgaQXHRdpug72COyM6WIN8OWJjGZo6KkFG0RguGLFMw1RHYnzUon/
OMGt3dY0LBrEAm0f/ay9KgyJWJNg11t4dyx8C/Q4q7ZuGA9jLmer/J4WF6QgyJ1F
uVe4Gqq+PkDDbvuup8bpbCyxHc4Ago6t9nOKvFLLfT/srKT2TLYd/N06+ScCTjv4
vZdUM0rzR/zFup26+GPRvNsCsBkXQ1KsM0bUbI3Nabyj6NcX710CoTgVn/lfDZIF
7Skz+uxL98XeGeHLkSR/4r//2xLercLo3PYYPR2KmRoOhwM4bjtHWjUtoam6aqEX
nBWFEL3yziH1uJVMGptXCtfMpDxBDWESGrlGoxkzJk7vaHaNo8FEzquP5wtI95Bg
30R8mP3D+WHMk4O92HNI4cn9UPxUez6wPAVfY89lO7f/bVFEunOG/OwlCu/vCSau
m0PFOn7nPB0a2vsn+JKHSk+t3gDWWAlDFyo6Sf4YAUV+4K1Uvo25poMYu4w9Xj/m
YoJQTkQH5I5zXRxOshDUZLFXjX/FlzAT6UhP3S/Ae2rPIHtp4hHxiCPb5w8Zmxc2
xwTLilAkrq8zEnY8QWh8HDFwGjf7DHB9JiyIke/Tv3I6tpqDWdUM2ehS32k8ltYc
OYjAdyD8LmFwBcpJkIHfyvJr/d4g3ooZAWgiFjgpk3FtNYLgR+xyO2cVBXkyRu2S
3pRi7AB/+ehPtqtsa80UT+QFT7WZTpFvhljzfLEBhqO3mtqcwWpX2DhVzSJOEeW0
ryi4hE8/4CLxfgo0vWwTbX5JlG36J3Dbz9j3jXlCX7dRxffy2b18wYHqfdM//3j2
J3aBqYoJg7ztLBIYiqzmU4RxlkDkULUr9tapi2PLdTukCMU5ka0BwaefFguQwcNy
/viM+BPVQSHmfFaqHPEfOyIGSA7D9EPIfoeh5SoZ67lQesmYhtHDpLJvf/eBCN1Y
pQlZ/8CBT21YcwJSON12CTDP0Uk7ub+GHQknpOtycrkLYcNpSk+BceKRiiI98ld+
DQhN1fHJlZRBlHhQj7Kry0iylFST9DD+7y63Gt27FNa03owzXOEDNBwWltiynFq8
Rs9kjgGS2+G5pBulpyQgl8rR1XpDZg3jOt9T7sgBeuEzRwvCFduW1qwH47Yn/vwv
HPiiUz+1Yh+rrgzShYAXZPZAPCNiY8dnFHQ5wCdE7h7oQhRNmggeIID7FiDmxUf7
SxQroxD6GploedxBagOOJ2W25tKJQDntg0+CIz/Rox7/ODxo1aVtms16aLetpJ/z
ScyxcDgxfXAL1WZxo+wdPDnPHRv72CDfkPBg4CjLKFi03Y1KvbHXsHs8jSXPK586
LxcGBoMsx8IgNCpzfWH601KMpSXwZSZVi3ccMJg4SEPBYCRkGmRNNbovncmaf6yq
W9+aaTF5JYEYpDtCPOBjDOSfoL364mI4DBSJ3A1S47rPi8lDEunKmdR47CFQCsOW
xw1EdHwT/QEJzgWFEzLicAwi7/lRMWd/Saqzl2GyEZV8I7U26L+JoHRENcIMUzx3
1QSlv+VksySY2Kq2amUzEL70XApDWvL6S/54Tvg6J6dHsz7ndWFsxQnDhUTE9rFR
Nud9Z0/6UlJDZaIpU0fClPz/rDgxn6CAqOW+9ngPcMMya8P6AtigB7epCd8As7z7
PUTld5kSSdPCaoSaS013S2dzLuDb2p7PjBzPFcxQwgRhDnrDEiL7Z4nwsyytKNkh
aRwhhQwlqs1Mgp3ztyg3vZsolK2hTzzyK0l7bPBgzssJ17kY8XHCVBR9dfRJOLp6
mhnV1bpoyaNcqXysUgwtp4XE3dcij9FCcNAWydq2MGx/tvnFLtFBbwtp698Md6+u
gkji/Q2nptleu8pwRkkrdKjyHOk4wpyqcRzYQTqTZP0K+5Nz3ENva35F/b0ltIs8
s93v9NGFxxGqOQDZ3Z4whS2xPYykuR6SuB65Iy4SzS0HnDa1p+qHhWqW0VOeZ+o/
x94GMnpFyNapG+4KLWjAXT22fcZfJnqPepfbyNw2fRLPQhjyuJlo4tRF1xNs0knH
43qv24eEB0n9yLJkdGtbawXGI804K9IJ3K0/X4AkdvC8+PHCWNuCRhUS8wQdruFP
CbcGFnIk2B2bdhUHz6xIbkpocNo2L0T0q99cqx0zrDjS/E8IecU4xmpp8CsnWHe+
XKd86vecXWqp1CtiE3u95MuGaBeOXRRnbmNtezz3JDQyBKJXXa06v3fpMz83wTlq
oANDkuOhNLVTNH/4OHSQIRpNQtgLCvceqEE3TWLf5WVz4HrDmIffKIwtw+tVZvyN
N0l4tCym+kbqe2/dkF/aXbxUJrBIXgEJXGH0a+tThjZRBz2Kp1vQRqbR0DqWDCWR
761Tld3I3yuyz/xPIAN9kf+c3TCwiDKh5Jr17aprB6jWDFNoygx8YJGP08BWPPZa
WaNcso/nupjmqrd6y07J3vN5B+sH4uDlpm/kylW8K6IHkeEMSxetahdOkXyXq1sU
1iE5ixqc9TVto+K2NYAvzFpn4NR8pSm22WqIxcHfAtDIVgFixl2DG6Rd9CLZgGXF
yDx0QRl4lruyLIQFwZqoqQS20PEmcZ0PwnQx6kEtpYsUmxFZVfN2joxZYJmqgXsR
d3qnzJPzrsFQNGG9rYWpxo5XA5ZaZB9RkuSzTDtPDnCX+2xkkbfzZXBv2E4Y0iWp
rqvswa4qSGYOgutjg38V0UK9sRK50Elzcqd1V/exo7kSuSfCDigSrvAPXMqkNaWq
jxiM7UZY13Puu9nIkZtsjAKBs09xAw1LxmJOtSBEWujCDVm0ffGdY7QXyHDjLiMs
nrAFcDzNxeVbL2Moi9AQ5PZz+gcwsFjAue9Kt0e6Kt+d7WcGijZqBlfqO9tbHzic
Y/k/TWqu5qFYFSIFbgvV0u+N9zPguJIiGYJCbB6cJdFT5AdLFp8QMKuR3pmjz2B6
RbFtEnLGd0sCVawZJdB4UtOyWK1QzQui9hyWreyIs8qW234PdGhKwgXm5CMLaF/0
UZr3o4BZdzpoQyCtYCdlKMCBqiqAWqX0I3MUKafD5AWFi7sJhi1kN6CA3ouNhV+u
l9Tp3kSSLBA7DyQd6PUjc6tf8Ro2QPOfpeOQDIjNS4cDJvIYqPsmMYTILAqx3Q8R
tpvHgfCkkKBExFsxMBav1r3XvGLQLESy4TkwINyPMa7QgUOEeqQaz+t0yIBYyfDP
vC0dUIvU+lvP4vsmqBvhX7lDUVL1bHE2pNy6/C/MNc33Yj18yjrv/E+ezS2bynFy
XF3OLo+VFlh5F2zDx2Ps2FqRaet0WuxZTOtNakhfNHPgp4er7EHuIUDzXwaqilM3
Zk5uvvL00r3n2nefY3N9Tjvf6+eh2c2T5hRV56Fb9LT+FNiBZM/Uxluuj8Vw4ajW
AP6Fb7dlHgXXX3TZYbs8AO1hxFGhhrsAPW3pSAuJ49g3a7qteJrXLsca6YxAYImS
sh1CWFIxrA9CQWK//QyLx2HUvN1V7psLseW0pBpmhOchKo2rKNm4qNAEjx+m1hyf
YxmrDlfbIBl5DBw4sncsmeWsUT1RNOg1bLcmunmLRkQJEKhOxa3j6IcTSpcmN6A1
63lunZfH8wMOSut5QXTdtJ9ICa6WeXKZELDWkR2VIZDgji3J3uUxZmS8+9BNmnu3
WmoLIaU7RmiuSlmoV2vIMODG3IEbtfC1n7fLgvnXWmijQMbaUVydA4DpJiF8jiTt
GqUeeo5Xxl6nKB2D/PNjhFT3HrmrfKksJ7MHZLJ+g5f1jOTKl112qVk2vUjurN/r
Ke/9PNuByehUBzBBz5KiGtlgKqrncWZNY3q0I+QCvE06rcyLp8C5LSzZaSqoN5Wi
9HCfsvyzk4i8ziZ0FjngM/Za6THnJu3FEcxYFCJnm6sAEqy1zk3igMG8S+8UA5Dg
+XgmLMdt+fmIjLAdPAfccq/cGHrDX2ZGLBYiW87IdNt0KCtm/Z5v037tYV6k2FRp
aN41F3n35m6Jf0LVGltSpWWpaPo/JtD5nY2gv/9YgNcbouB8umtj2GtxltN3xuAd
TbGFTz1D19o2mrz1RHhKaBJXfN1mYgecJ7omI/9VavKthXvKPvsMwo3tvd/OiE91
1qoAdZZksKnfrHDd/tkpIhCrpF0KECvzyWOE9E7KZkWVVNBOzs9W60OCWHzEVTAT
k+Vo+ted7EZ4S6OmdUkOaSUawFe0FDESBkda5CDSHySqBdbkvoyPi75XdaaHT9Ly
nnjyXW5MWGQVhUYT39vh65uzweuUEZRh+AoBHogf2bBRq68/Y+EIo3LzdCMSCssD
3wL+FCqnu7bGqTSwBOrRvEH/AL9QSBTwrH+orNGZCqJzsNEs6KTPyKiz62KI0liR
zfOUB9ifmJNnSbNa4nj+hUXFlXj3mURilRFm7pPE+RzM1vsCFzmta4Awh7WP5GWX
06mhayNfERFUrQGADEXW+DwE/2FUtr9O51hSFGTEjO/d3Mji0V/yisqiet2sRCTO
d9Xz4zuIncUzxekfbqzN0rLeWaamDoTqS1EH7PGbIUTfP/spguP18xQWdGkNB5Ck
DG56LCr+SiecL+y1OvlwjOy6eZ14yQyO2rcduahGk7mnJJxvGrKNbEIXt+6RZBBV
JWMd0p/enUMQRWAXhV2FYAjEJAPYL+8F9OsemdPGGakVQMgJsnGUoNFhjv3+BLpq
jnBTaYlkCOdmmk2EfJ+deOBPzEjPIluGNlyAaZ+AySXYEC3MJLdbjGNYQUwXeoqV
0hZjOf0ylVZ7iLBfPCYSRvmou4KsY04F6E5b+kY84GVgD8oUMVoMXVEcVcRqdH6+
O/tD1eYfVHof5RBpeqiODR9FFrW/hdh84TNqYqAHai5Vdb610h89ZDdrV48dIQf0
ZNNdMT8JggyMaxlx8zsKkOouwdBFL66c5anxX67Hp79n9kaeUGmsN/CMS4Qbrp2a
7qRA2H4YVLHZtHa7Q5XSAY2Q1RM3miu19A+ywSYe8wBTW2lFC6/b1pqdv23TkpZT
rwQupKeDShmxRRNApb3JJzdHb5MZiBMIcV1uarKOAKzr+2iL0IP/Ou/ep2jY2gmH
t7bx+9UjlMKWojlhocQTwKnKfwBWNZgk6z6HgEXAaHwHqaFodgjD5Sav56PFLirI
lWOD7C42vUDy+meTHmnnm9nIVKrSvh4iDGlEPU/77QeMjf/TVFmwaTzE7Mq9Gb4e
m/6Ta3cSYvGsHrF7HlzW3Z0nmjyNglsOngOrOzgU/kHRxTcVpaaaLljaU15PtJp3
ad6Z2GlCsol6dysae0p89qI/11CGAqPS0jILlZH5UM8QAjsE7YqToQwKkAlnfB+V
QK5icIobcXa7Vg5ybiveSMJKgE3eaLWZHdZ6j7lxGueZ6sRj+2OEfERuT72xy3gL
m01qqOihihH8oXeVHklS/VYM3TkCMqsXuKpkMr79gHIGvUVlJxNGbVFlyjF2+kYS
fu4e0DA6f+vQguKtpd42GpWiho4qGo0on8fsFvGW12VlwQ0nx2OdM9UzTnMLkrtF
AKX4fPWhiDN+mDnB7Ik1Xn4R3pzFVUJYLuY5SWoAuXke5hGkEAV7GtoXASxVAzcU
IqBDm+Dizmou+erKSxH7k9uCacz790dB6SWJL0VcBl7qlpYqZJazVisnyoovGr00
wsDTuP4WGabeaV/W4WPLe/dipXSNHsUMOsCrlYDlRS8xp2L8yRzX4RuSM58xjpKR
vh265RATiB/0sLRLVnh263YRAFmuS6Y41RUUIMdvBpYJdboGQBQbzvdJuzL7Lh2N
jKcliMvQ/I+k+AxKL7zOPOG2hnZab9Y8vUkogc+cS+Yj2ZYpANulDbY85R2hG2Ny
Lj2ZxSKTZO4vnNche68rSnHgkcCFc8TQTjyNbBu84KXrulfGbcYdRzNN0lB0wVSJ
Ayrouk/Cf4ngfiHBn+dMdRr8SZP+sE0erawhCYcUuuwYNU1W8v/oqnmtXdue202V
zo6PFohuVK3a76PYa02CaxeuEfBoZVBteuCXc2HZNwIoauJ8r+0mt7p8Sk9/WC4D
xAUVal4PvOGycbatoMsfaYlinakoTdIgTZbl+dY/0MyM9jtAuJgcly7JaI8Lsk5T
iRMxb784ct0L+Eqpm3dZQu1W6zsWIImTK7OJo6u+mimAR+dKYUz1qkzcsM5Bea75
wD5lvrJ7ns0paxEIoZHhAP80/nwiId2902MjQQ83O6e4UYe0Dqg47uHjAU/ZuYA/
IXixWpdHyDdfVMLhxRYSkFXsIMSKfDEvgLm7QjGRmnsS6eSDw8VT5hCDwfdJ0///
FAvq1fe+LoBh6H3HhuqHG2mYxzcno1MGu5Zg+Lq0GlgCl9tjnHA48nNGqagBfZKC
i0QYbNbLl5qMi2xiqPTQDHFDXRu45NnYIsz00uLwoLL1C6D/te8NQpSTfK8gvkFw
ayfO8c7DjseX0yHuc0hPPNIkuqx2hZuxFzU0gP+vcRpqbInPUykr6WRo2HPLijpy
tfv5/Hj30HwgafjmtAhsEbJGdrf9GizzVPzs6hAE9MaQZEz/AGE5Wead+QzswYJ+
Vi+DvGn0l1mC9IDvrtwWvLzQVcTgSz+le9bAstGMVTaN7/5UY8h5xo4A9Nz0hIN+
2P6nAW1xV3NRAFgd7/3RoWdPfA8sfPSWXKQeE+363eTQlLu8X1TgjmrLbzetcE/Y
YvAel8jI4Iu/Hz2TvzoCKLOdIpUHZ90mTZ783mAMBI4SLAwRQVYYycmVXArkPze6
xRXH7uRHFYibnrwWdOAFIWCxMAcQ1xh8llRfjxzqfLd7M0E8PMC8y1mqsQyXnNjf
vtWmzTibmzj6dwN43buc1TzWdHz8V+b8EYu7yPfDEzA6nwwx+MFVDTheDPtM83TF
Tfn/cK1d5ynOQr6m1jxE+rGsmtm9wInLhd1sHDhVtyYz0rAE3fALY7DB1/aorsBa
tb4arMr6qWvGks9nXSySCLrbn03LfPO41r7+jxBtY0cD69b3NFbr7nhKxOMchrHu
j44Wr9h023x5Xj5y9O0GUoez0sgS4YW8EMGALPJ0/EmmGcTmAXx24bWF0MDsMOr6
fmc07VgVdb46BfGi3tDUlYAywY6zMmRIp8gsg8thyJxdBX9Ug5GKlB8D0Is5NMg2
D4qKlccTDEcyuRpIzsdqGDriF6eRnvab/kUYv/n/EFCh6VoxN0cieVyHIuVAACy2
e0UMEGWJ/UndHH7DYneoh6Nvxyq2PWFkp/h4itwAQQojSPg8hsn0UhrLScM1hooX
JL057dOjV97HujvW6qW0ycRb/S2OnnXDMJTujIEAo59EOfV/810Crgl3izX04IOQ
fLIDXKeL72/TIFrN/cnG2o3o7U904r3QeglHmsttNYhv8cej8dGZarD3h+PIi79g
6MHQgtn0DahRaFmesCIbD7V5V+HLQ22R9mvLzWB22b/BI3C7XBHX0RTKkKw5aX9v
Icyae3sE2NvlyCRO6cU2oej1+ZPogjeNyGSgC3veIIobDM7nQ753d+WvdmUSGxD5
4U3F1sksFEsQ/ncmCSnVsEkXkug6xVtgaJ61/ufN8YtOPi3hwfuW4RP7K3eYokQX
sRXexykfLfrwfQlnVdvo0U25vawu8ZDDG7t58oe5FNqi/2BaRTgOqEe2jjqLXRYp
UVNYqQyWHEMN/6a2F8HNlFvonfMBXU9OKOZSCALbkObJMQra3tounZB9pL+DTkA8
ETfzIPuR987FhK/JmYwAKOQel761MZpOblSmP4iK418S8cWgi69b98QR/XQyrDIe
RcmWWw78riNoenApKqa2YTD5W3lkBQL+AcyO/K8cb0fQzGKw0QSsauZDVGM23qK4
91J19uZINVnlK4i2BSUysOW1NizIXNz3/4bGDIGUANtr0Xukrv/c+LKuL/Y0aMcn
Yvrvvsl4EsQTrUxPtA7XS8bPdWIShrikyuNQfOUhXawoMHLjibpSBmk3MSw/Apmm
Y5sQ7PwFRbqTSzfW6fSsfc/t/PoVsGOjyIUEVL906h4RLbK/Zjg6EtfaLhmG/5Qe
aXFxGrZjr1fdWI82kGyKB5umgxUtRsKq5AIIyWp3TE1Ie0tCsWMPWrDa/XIN/SBk
wcbw2TyFjE5/eq5/ellBNRiQWUZ5G4zOpkzaPFBlNt4291EFMnCk+gv7BQ5Ek4IR
3Z9adRZDvu9pszeYWqZUIdS7M2cVLTuPxbhA7r1/NADb+byogXFeRrYN9oZ5rzdq
vSTgVBCS+SIjUJfkRLhfU9PHUKyQVtYDwSvhrLNZyfRuInVniSIRXRDwpsgqb3Ie
pxICT7sgmen7b3B1AmDlhYXcgvCBCJWqWHeY+RKJVbHsJEvgmWO9evMF1fi4KRZT
z0faWHM5t0Jxhx66NZSi/Q0APYq72vlFHdOd59y0Tq76InCQF9BcNltBHpSw6IOf
+iRaZ0+autM1Y1EHyE0Yyeq8K9BnT9zF9q2S8On1+Va4H39wx/6iWCjZOMp7RVOU
x7MMbyfoBLH2dtHr0K7+wL7SrFmqB3X+BbMVQaVf0ygi51I5nYr/ndoP8Umo2DTf
mH/DC1ERcPpXyc9Eyf2aNCZkTaMdfJVPFfhMFTNNYMXi8/5tTRWZIyFaSgaxmapq
2/FfiOJj+5FbL7orXFCWdwIEQ6NKxlDFSjmGejgajrkJ41ufzIi5do1N5CILU6Us
/fLpmIvrMhaMEgmWJGCfnmAmu/KazXPQjvwZcv2pKfAn7n4HzWyBCYh9v3ZQPpD2
ZbjCjhIa5gKPOiszGfBg5+cbEwvQgs9MxyjPeuVH5V0b6MelaX5pLg4ZrWE+BFG5
kqNK4enzYsppdibQyuGFeZbBRf4LiAXCdSdPUiz4bPvQS0C9e6WC4NrCTWxNrJco
u9fZDgy01NwjXVhtllnnKHGj0E4wklznhdTAFxdksERW10PKZNhSe1L36QfARVx6
TPXmOTqH1dkv4yrqvjMWoU4FIr83ppYtBDULLY0HAkiIQdfaAQcl85kJq1n9C/Di
ET4iYk0zC9eJFPCTREts18Q9dlclOjdbrONKOiSOQQ2X6hz0NHqWKCLxOX7ZNy9Q
rDGJfjjYR77DwrBS2Vqi0GutgWElY7h86qorYn2r8x7F4jQnVgHxR0i5hfp2I3Tm
oGtwBUaZLGcg70wvj8/yRFWJLZKudWo8Hi7kV2xwHx2nuMznVv562DwlMv2OnUdk
9TpqpbnNAckCZ5KDTl5ru2erxlkJB00uy58QVoWLE+efEuxk8SmjOvbd3X4kUB1T
ccs86TByu9IrJIlv1QVZKim1P25/H8X5v9eqYjQG4yTmpJYXb2Yd4nJqiYPGtZa9
54H4aBKUcoEMTBE2V1eitTK1+j6SE7XrYNh1EQK6UU7GZia2+79Qv0n3cMxiR2vO
5YIrZ/mFp2kb2TTsVy9GRLaOEPnZF8JArXJrxqL0MGXQzvM0DIq37dStax9QuoLH
uz9m/x7gMOpgnszDDXTwt2iRQWIdFZ9gOoY1LOfT/g6CFybYQsaBV/rTEes+iJp7
VnK9ufTlMYC/96VvFOFNgL9dnqZqG2hjnrgNR5gVZl0prJzKDyW4geG6RDJllfvY
iHsjIgSvdnFbiseu8u3B4aWqx1MDEfdDXVCp5QC1bpV0PRFjb2GQWmyzVMxHilY4
41G3F8K4tYlvtTK1bu3St1exbgHm4T97915Ml3aq7j4MXChrVrcbdp7wA9ly3HZp
8oThuh8inZ/20m8ENy65aTR6ZMEuIDG+31hjNLjCb2rxBURirqpGJF4XjOI7A2rO
gMDxyXuTScPZXeC/TTTNFb0y/mfb6o3w0GzzAMk1qwZlcYRUdsUAEuNR9zngWsLF
JsNTbVaUseDOkWxXTSWdw38YXcHY4ae+ISNtjza5rAQhSH5aAp5C1YAjQeU/5y6a
Nh0EptT4zOIqZrTon8vxvFs0RrxUCG+CVVjQeziouzi3FkVTsfs6K39KCHblHM16
OOdiaTTZUoNGDL5b4rygfVT0Lr1ZYwNFk83dbFoL4T9c788/IZTId8abt4z6Qdwp
BYppuEKTX4T5a79aM3tEycE/j+woGUMocGdHJwgkSyFdkQYARTGR9YYRWyWJmfTR
gvc5PHeIrZWA+l+ET6rfgqKDElCYJ+FiXi2qTmzOsjzDAh737QpJThHeaoDHm/Xp
9UYq7vSiOBF2NIsL7B60nx3a9cX268eT+ODAstLL0QJQWTlWnmItl0fwpuEt0Kem
+MCZokqyNw8I/VGNcXD8EGqLIhzJyTpwiDBnjfuT51DvN5Fuv/bkVg/VrC43VWKO
kFzyyB77G41W2DYXuWAaScG2//IKmcaCtMLQoR0e1WDm3Ls3qXefw5XzvlBkdp5+
3CoUtpmJUB5PG8lAlI/QEyXnyHK8i5K2r0G3gI6mzh50JqxUK6DKN4+E9R7FCHbM
c2bVM4rQiL0ZJ+4zp1TvlrcPLdHHcmLnAp4rJT5K9T7X0y7WpWO7PCqvIInzhFjO
mGmPi6V+rAv8c643aZxUvPwM8YDT0zh2cmtkXrKS9BZ+V4Sn+nM30wWo53K+RY6H
oGEViSeFsGH3z6Vvj0ib4TOzdbb4yyj0EotjMi59BYdGqKUmZOmajZqX3fTUxgw5
bWnkfAWBJJKG4FqeejJJChT+yi0DjqYoGIKWYnTOSBe83FR57qObtshOoJLOGvoJ
XE3VdY4O3eUVv9ZZRaAOVUHf6vvnPg5+2Yf9oqq8ejVCU4L1/2DeNoLMT0XXEhtP
4Va5dTPsCrvk0x5ZixiamaAQYPWxFWlOAXKHY81/CYucqoy33TPeykdJp/vrZzUo
19OENCgep5KxWOlJdctk9+X6HxK/f1I5swbz5EcXlohil0I1iR1KhWWBHOkN31tx
Xh7pWJyonjAsoQESeuN4eQMsoU4jWoCD7VlPtwuL8rkKxSnDvCkCecGn6V5T/ZRc
cQkQaj8ex3X0CvNqm6bDKDJydELOI7lgLHYABr4n4ATN6+ivNPcjqRL1+LNW6Q4l
ZDzUObjwjfNrgduEcJ/e8KILTg5vfuzL01NFOQlFpAt7rCLYf6xLQ1/dOj3X2OBF
I8KuHIHkgXbykbpbyaBUruhHdj0oHXDB5mDOe56ZYbZj8Kas8wRi7NdK+8BOOdlO
TeTpohRBpj29XmkFRH/S2uU7RGbALOF6jgyKZxnfpDwWuUTg5zX3SgqOP1o2ppbc
UB6jloCce6mbe8C3l4N6MxgwD519OkzhfAC2YifOeY6NHX6/WrjY3ONVtjzKv72P
z+5zn+n3vNTyxjW+ZPRJ57G9PRmnnwcI/njw2X3K46QjUQCToEB5vod1e/V0djxP
iJ5bYSCjs0PcGwSmF2zG0KNAR0lRHP/HKkSbhoOJIEeJQmvlSZcfo6ZsHP/BntmL
WirYvBfgPrwlU7UdMwym/cD074pypEKJhFpONtHq4pVlAQf2QxzU8g2HlvJDNqpY
lG1xz2YLxRg9fweDLiyKVbORXXZzg3geAhS8lxHva4amC3vvJiLB/jweLMN8QauS
EeIsupEGmHHzXSsr1NOqhFcve3C2OVH9fS9a1jtBUXKAaLcHOPwp1GMZMgBPHENA
Ekr+bz7zXHqMfeGI/a+80SLEmLmY7rGrNEcmIWWdWD07TILFrdZka1Ihe9h8r8DC
faSwIWA3GZudyhw+Bfyp6uJz9JqYDlbDMdMomo/rEDSsDKn6JF62Y5bAIgUoS9gR
M2pTCDCc7MCqHxbdY2LvfPYDA5ekZYI8ZJDMszKioA5U+A3uNLPP2/6k6M7InaAJ
931ATdLJoeeYT9YPybYsejqsI402FojHj/nJVJMt+B+lrVIpjF239Q+VQ/TBjh9m
/ldlJ7F6Fj8gxNneGXEtHR5bikKCMuQqIIsXhChuroNSXMQIArjQ6NjBnOi+oozN
/CN8kieRu6rl08Q+3B5hx0+nOpgenB9WH7/QXnZcRNpCyfFetkJfD8tc351ELbHh
UULRdXIW2NUgFvYelOZg26ZYwelRWTdiV+KhFUJzZXEAKIA3+pQRl0tA8OFQJcV7
yFWt3ZwqrPNZi5UMOO/fVbgNEQohku8zNhZn8Cff4VWS+uX4UmmvjYEPJxTOt7J9
RQh0xoNVN9790buwA7kXJKl0GnaHaWFJj2G5IN4dj5UjPpqGTULfK546+n1ygiqr
T0jtDh78Ku7r6h/wQE4/zVYsjxnGzh9Wg+a6Ief7S/bhW8A0N5SU05sHGiSlr/tS
jlNI9ALQ2Jj8tvtpBZ5Sl8nQ1M8nIn0KPc7fUVBjSlNqPXm6VxN3hFGMM0w7VUOo
7rXMlgldZ0XHh4ab4ONpMQtLtMz4AN+wzw8ga60TZRWXZJAx+/VMGOpBrlgUbwXx
7D8uO51OPng3fM1DKs4Bc/O7QCNtyEc1/y2KDqr3jVkXKl/C4zSNktvH4VGSf1vU
hR0dCnxO9MJF9wESE4/EvGcrrBIgS/BFmY4cPJWEvCU/htAKDM9beb72aDMKr2fu
oY8fGEajhMLC2m3wQqYARYYhvdlS/8AYdC1vuRL7366Pn7HIKCn2Ykq8gKP+EFKy
HYCE3hrtLybZ77bmeMqRuExrB/wY12dSDUQwiEvK6e0lolnADvmGrCoCgLpJlLGj
Iorrvozswcns/IgaV2Ve7DwQCq34BC/8OmlGfKCN+o8BpoFSIRF9+RJ1PWWbzKJ3
Dp2JqYdBK3fyC8vN8ojTGrrv9FNIcSYUMwBNoodsj0Oh24dHtJqGYUAqiDXtbkvO
S262WBrxpL2vfMmbLjODTFMcgZW8mgcJ783v5Xvk6US0t8Q4Wj1LmD0rfBH/slwN
i/+R0qR9sM57DFhKjuJGrEb8OFMaSitzSM3d7/FRdcjWOmqrHV2v0ctX4uoJqG4l
lFRxidfs0Ku+fCsQVczs1eim8Spgh+RV+iRk2d8+iMTaVemgniL0d+3wHBRvS2kF
Z63dX/a7jL6nP0zspbTO8IbM2+CckQYVfBUau7xsqY+PnLoVoweV/ERD+pkwDuRP
pNUCE7B6TE0fSZwPGg3GdzY/Dqva9G9EglDR4LiUDkXzmhOiOLGpLG+QWIl3Uj2O
yPOTcwTwbs3oIGNokPxIXmCMqkFXU/FnIva769MNUfIYtrcOPtLeDvTj1tn9ry6Z
Ev4PbVFo9VpzBcQ12xPOp+0rIqyh1xuVwoyx2Vw41xGA6mUXZnmLCskgiqId+Qcc
LCL+TAF1ng1YI0gLy0KL0aML/ZQYWiKS9JrIy1Qyu2hW2hdT8P44laGAAtOLIgRe
NA6XHvkJn8dL8wridv1MuoO3wh0wCjUh1md/4dMGv1Xt8YwyYOp4ge89xCIJoxY+
snPvBkWQm0lUxm82yNyNwF26OKFdnzjlOWzLeiwItQfVx4WUtM8ndxx86yt9UFE7
iOARVBNW93IlzAVq1xLMzoFLJTRyQSCWot72+5zD1uxHnhen+thEcRbRyh0zfLMv
CWUroi5S3cypBTPDmK1zckn4JQdWaAlikIJ4J2DVzXBlJsL1+iVcwjdtZFOxMfoI
jwMLqaaEKO9ikDijbRgbK49/7xLA48iKE4tBCPMkO8+1jUh5Sguz0nBAo+aUSJPi
tgY9cSZjfNmAV/uxMFNzCPYefq9h4O9LY8i/FMY7oUIdK/1Q42r3hVwwBmGdWTq7
wZeb9um26YV6pjnqCha2tiInRNo9eMmPjT4wKxOjVR8o934VC+bxkOGhDIJIvSIP
ENuRLBq5fotO3B/VtIJbTlW81iYUcbBCe+RFBQj3/Lt/lZfPcawP6R0JOUHYpDX/
OJT1YZ8XjfcA7fS5UP001NS9TAkGzL9h9LugECelUktgFpVXYpM8J8vMnxRLQhe4
Jpve60ZMJK1PWq7t4UZeBHYizRs8nvjqqkExP48VxCChOtoSNh1wKSLczCDiO9OP
T85jcTAfksYtoWe8GT39yT7dZIzfTn3zYbwJ/hIXFFqYsjjJpcwcEWJ/eXITnbwu
KO2+guw9OzZY83iyNUHc8q8UeKeIV8Lp9aRAUCbiPVMBsYyAM/kqfHcs+b2cbrqv
xi0yrUWxlh42MeZb8gXnKDk45ny9eW+BlG5UD9bDzO6k6NhAcoPD7mztquzV+G96
HvOk/IWkZw4VO2iblhD1ErS39iJIabZ2mViv6jjBrFvX4LQah74A1l/LFbMYgIlS
2sfWdB+sDLGktT/8C4TRz86AIUiJBhxv271gceMGkJulf/IqVcCFB0dzN3zbDs9W
QF/VI+Tf5z45LtvgBXM8Gt5KQy5rvGLptqchOLUpr7vFwNdQfAT4Jv33ycBXr6W8
pb/5HTep70nJG0krilfiTtUpGe8Q1iZIHXSDLClCL0VlKmGcus9+8CfHqSFP0SW5
glJNLpSmWMtU88AcMhN6Q/VAMk8BY1d0cEJ2W9cCutjx0x53xtKxD4n2HrStVj5P
L0M/lTJ7p+0HD9BiSg26XgZYoHRHWQtcGGot3kCw0gbLpoLkkDgXNYLvSq1Adf5C
JPOPf8iWd2tuufvEg2YgKLAJbyUtUiSXFESjqxfv1cre8yHQsv9SCJiyo/zNY/iu
9E+jWEmhLwtFfYfIRRp/d9Oy/a6LgYA5vgT6hachwNcvr8tVpJNYX40ZEFHmGx7i
r1fml4LAmajiCfYPiWQGKk4w3uO+WA1bd9EKD9Ryg91pelBnZJlQur9ubnccZiU4
zTwE3aqlS4iH5sXUk1U05KqV7+amNIs/gUcfmvprZxNgALHyL70GAJGRGZGH+QxI
3/aWCdnmcTzqvefO9a/nrbCxUrkcl78m5EOOapZUaFLHXyBW4obtBFV4tXeyE7t2
CSpu3KrCIntxtPx6UWOe/k1NQ2QlY8qU2d5SCCH05TC0MvflbVEwz0qODJ8NwkrQ
r7pYyx+Dok/OMqF8jfUo5VCAdm0jR4q9ttpjZPvxLqcRHcVC3LbkMOZRg6dPX8xl
+Qri/lEkYgq+TScTF+D6JZqC9nqE90QwYozihJiIJybPS5gac3ijRRsO9un8NZdq
CYmuATKW7HswXuFEauNE2Aa4NucAUuIsEy+hR0Sjgs5aIF7jAdb4iQ+5IX/OLhAy
sP90Ss46CbO/6+cjN+1pmq6SlaZx0cHgpY604z23fNRUAqgNVFA5IPyv2Lw7KHE0
M/+bUYcFpXOL8FJIKMkQjfhs34pLnmX9LJeuxq+FflO/PBnZOaz+q2pFZcoRD4fn
vSEjzHjPaSQk/mu9rfLQgdtg6/Rtd7Up/V7sWM2ws4hjAoMl7+y+ipbVdj+aw7xQ
NNN8+av6KSEWuO8GvGyND+09POvteeiDJuPTwimUVP6TJvXc3entbwmp4bDOqyuU
NcNGpde7e7rcRWv/hdVLtmCu/OMgcmzNK1DR3WHiug1iBNQ1lhgPckSagy2HX5Yg
SoPyBPT7ILCbFh7HSSwRgNZfUDAYjSuq5E9DZNDwfIGiibdQFlMyGebrLXDYzkux
ytYI05P4d49HxhgsAEa6a2RTLoHPKNOR4fFh+eNqBfhHSiH06SLfHnWvqQ1cL81p
XmNnoaPuW8ZsTlk8U3egkN46IEYu70x+DYMi/wMMPxjqjAOeV/XG2ukQgH1hvi6R
9C0IaF2a4iL9iJPkJoN1qdMuzliQxO4DaXmLDYiTz0YNIXgkgLbNo3slMl5hW2PM
IJXFO4/IKFM9voDyaR6wdWBKuAnlgAAtLQmg5cN2Sa5Kc61JLhmW/iwrVrkoG9wq
AD4YglDT9bRXsMA36VHuQy+cxbqNm7iHhtDRxbH3WFXTgNp0YLI92+dHQyjyDzQA
ggbrTYctYJuvE5mmTefIYwnaMhWnDnPt1OuDaXTM6uEqmlwlBJuK6Y3v4EnvrtMo
+I8JXOSVx4qV/NAch+IkGyfsPjtR4sPFE1XMhaQhmSNnJ9Gb+KSUl1+w35oigbxk
FtfKREOTWdhOLLnPuvLdjoI+yHOTWEjcGUh2RV+ENqAWReigDGpmBhzb9Qu/WiMC
0ItXALZ4M3QZWw8FGim8n6YmstfA/wVp8iIzhgDZUlvlO2uZ73Scvnqbl6cXWj8r
xd4Dfd0fzD1QwSWkII/JvdhooeaXXC7VGgHmW0uVrR1+iPmXA23Uyb13hVfNtoLE
M8hkR3Q9DGsGlTkEtSuYgX8Vq34k5QqdZAFceJ9Yeez+y3LvqATNvDOHPArGKxz3
h2ZeIaLvHR9Kh4qbyeFW8uerUuQxbyWZqI4oqLRLOrmBdrEykzfrdWvBxRGUfORr
ka+81ZA8dLG+28Fh5gmGecsvmaC6SkKn5Rwdp4OBymgKqTKEchm6+7H9CcOG2hNJ
QEA0kC++8wDslPSNs+AXqKWOl99+UOUBcoc5Uvg9jaRSKSR/JPpA/cDW57gaJn0g
Fw3YTLutPUzqxznR+/0lctExOE5jo4QdgGY+DZLYBGs/PhXJ9LMwYRLADLGcIFho
Rm2wsxb7e3lerYSk9vIuCwFJpmvn8zfKotpqx1igioCZmoWWsuVsYyb+T8V69fgD
RV5Cbesgc0QfmQ870DYwHV3y7MCmDJwNgiR5OT9d8UZEsMuT85OD+FxSKAbyXsFI
yTxAYTUSoGwN6eZ06RSsBsiInK31IcAIqPbUk73b9GY2X1ZLaySPLqBgGjy1/hHs
jnOArXfcxw9RUnmdZYSlt5aa+DFFZTHya55wkU5OijsLWLgh/xa2qAlB0d5M2H0E
lAP+iNCnPY2azKPOjkGSGN95b8/3O/pNjtJ6jb1Dovkz3N2Y6Wi809hkxGQcWcuw
kJCK4o+BJzCaZIwP+kl0CxBpifEY9YhE/RTWkzvFYafPmyV6Y8KDtI1mjGLGqRYX
Z/t2Hvg8a7MwPb0ogIUiNwksnPw7fyq3D1XePRguhqWqT6VZAoypYt10MlWXvRBu
RQu7EL5uLP77CyXr5nZq/JpRulFf2U6M9x1ar/ADaNZypGFd9V0gzH1xBTIW/1uq
SooPCQXdftJVEE/pN6qAWMsyk1zACounKxTDiZq1xafgVPprUZrSodQr0rv2UgDY
EiOFygYIB8RVeBBzV+peBzeHSgn66MnG+vJBzY5/zFF68drhaQCtD83LrARKka4I
a0AoMyumAlmuPIZKl1yfez4VAEHkVbh9SrNWXSOwaMNV9LaLVMdHbf54mvi4ZdRR
8z3S+uPNAtmgJs732tTBktraEYlviq0/KY1lM/zYfNvqYYUSDw/pOfOqdxUkIhdI
LouqnSte430QZ1gX6EwnaBeuHOVFrG3lgPy158nb+rFMPQp+Eau1+Mc6N8Blap4E
U5Xxo+1J7d0Vu+8BJVUyvoDd0qIRBuVeFfcxjrAzZlEKgJAuLjiJnV3hoUGLtjZq
hWtRr+keI13jr/Xrw8Z4S4mnNjDZCcy1gJFl2Vd7MTF8z7Dx8ev4fuEz/wR/GDPL
6utI/dZP82B0OwdNlEECo6CKOKajTp03hCefQbjmY/IIxnc3ZOKQ0Ui2X6U44Sty
xohkkE4QJb41Ysdvr5NsRKjfQwuDoS3mk5e24W9bLwYjhPHeUJfU9ZiBPFutYwRt
M52+Bo+BT93gI1+6bQOHQUcC3wRIuy3n+EV+NKoG5GO3GqvkoaqGTF/KOmwSPSPq
Q6p9jYRitDUgOwruZhfwnZeo34ZOsLlX6SahMVj0+iLgrBC7ynFVrd0bIW2dvdMv
hBHayUjPO9s9CkodLmzXJ5EPf4RjH4XvVXm4UMaQO54nfNYuVjArttNw+49fnJY4
FR69FGsqcpixKm2wDbGf32/pVa5RRKr+7O9p6Goxfl0T6hc66IiN4OhZB+hh9alQ
5FqcTguVccNCzmSI+yM5zdTrBLtYA6Akmr8HP5pu9j2CGDZQEVXa2J0B7NKFXKOq
UtuUTlWbLJ2bMPZvdilVNSl6nOtCUHrrkMXbu3D9w+Kw2x9k7+YxxU44vxA4IoJ/
3yLjxkd+Gwrm+YI/ty5HtsCmQZvSvO+/q7TvRRqM7C3r0ES0Em1O3xc0qgeQiDbd
1q92y8KrgnzBbSAhh9OCM1nKrPCJEeA4elOJ7kFv3QJToM0IptVIu7y65jcTeYXF
U0LhFuS9B5Q29UyogAKdm7JtI2P+VzuCaROK7EmErEIFx2rDp64a8GjS85Sy0yA6
2vFjFmVyNfp7eoDEGLd76KkLJcd0UzB0xtgwFCSEdnfQTkF+hNOt4ZP4cqlCF5/L
X262ImzMZG4WcLa0WFzYK9W12KsH88RMi/CEe8z1u0yy3O8a+URATWc4zHOcQoAh
O7tOTkhPAj3oylowFpfh0HqFXK1k1HLWfUip5pjv267RuQr7bFvBSEShrxKjglgY
BTZFV5YEg3ArV0J66aDnzdx0Yw26gIdDT8AC37ltvFckM8IIOdyTs9GOGa80bYaS
ZUfAGcoC5baF08+kbUG/0JS6L3zFH8VclaroiAu+rdcFb4uy5iRpVh2tQzlDxZ6u
m9pc6fNyPDQjpTmUMbeWDGJki4BLeP0l8z5fgq1JmtOrV0/F6MZ+xt/MWh928TSO
3ISVeaRZSSqz8Dx0UqI+ydT1TBlU90oGofsh+qKILaDr3OtgY1EDgpZjqx/cSlo9
MBWB25C8ajJkyVvf+2cWj5gqN1xE8zLtABto/K5in8BTp6WG+b6oQPpp5tWNEkHa
anzogXaj8ecesbPLLGKpYO6nGeS6eT3CQ+a9GwrkFvTR7kKimjjgeSvLPKfg90WF
KFmrx/D5Lh8caUekrRcV+qqKepsqGvigiNDU52Jg+ycKhZJ85bxquerOxRaYXGgz
HelnGmU2Ky8cUF9bRYrf35u4EaYgML6jEBUL4Cb+OxmIVL1El4pfwlEZJIQUzWja
fsUgw/o6JTniyfM537JQxPFN3EVDT1KvYpp2ZUSFHFU/tw2CyKtM7Fwsq4B7Jus8
N7BauxGLo24LfjkKhtUJJBLGzjnH0XIKn5V6Jgf8ZZZgvczxqOPkacIKRdwMdGK1
KbD4L0Q3Q2efMV0UucJyxL5aMpgB+L37VBEIsIh3iLgEQW0NXvkmwFOAv/RJ8KH3
/CkRVrB+E3qxfpC6cmluB9auxJ+/NYJaH3BT4Y8u9atktKzGBY0U46Y7HuqDMH7w
b16Gnq708w5aLOCVH6QnGGEpljJWMaADE/RNC6nQBbP4/YPcWeDGAC1hDz6nXMZN
jH6fe3JXnsL7g3KLsKnoqaBxxtih88BgFfdC3Pb21z987t4gYFdxrDmakhwRbfBQ
G8scC1ryV6Hj/49Bknh9CsNAvt83xL1QXvhifvnRmnHqaoWY41JpMl8hBwbJg0ge
wj33QMQ5L9nq9e0PUR1U/x05+k2C0DUU08ep/RJAHHG1ESF8Oia/HoBcTwvIv1E7
hu8sVcwhSXb1BuvmOtXs6BYIIuEfSz3LOwKua3bpeNtuznealakabrZC3PsCIkiY
fqSg1Z261XeXVoLdHLGH0WJnNHR2jAbgYRO/b2bTsM6ANV4N1dBpCE5QvAWfELLV
f3XF2cFr9te8LdaQZikIZ5K1G4gM1LGQCCYiVyLzmzOcFwL8WT0dbJDRhs2u039r
/iqFs/N/hxl7fsIriSsCW2shdJLr/IWGLAPdix1kg1afw0KjZ2gP5137NE2SpRa4
XQFYi3gQwWqxBf3ws3Q8k7YaeMW6XDxTe3ZS+mkxXdyOFqdwj0JuYcHRhtLeSi7+
u3ARboU/vhQNIkSESkUne8QoYY7otZfBK23jugf6ztRKQU3fhVSh+t0ms86YVPG3
GZ2W2ijFPBdZBm+vK0gevSJ4WLmf4tUVpEdHaCqo7sLpDg2fyuJlekBCw8puLE4q
fLRTcj7ThfvaX27kWBVnOc0QptJX6Mx1Bqmynz3tthEplHgsPflg8iUIMUJZS8IJ
46fFAudjbldUSgUnp1y4ItUDtCYa2e9P9aAxpWWGKvOpFKumevSHqSUMzz4w3obr
6zZinKNJqDxXbytZAw9LsEis/qIPwC8b1yBvh9Eol0fywlR1s/x/iuZMjaK0VkLC
lv3E4yz6gEQRs4FcidHGGR48DPXGGuWEnegWGioHC/eaHnpNubTTpIHjpamgrHru
oh/ofslZ7mpyC87Mi33smEdEJ0pth8pdkqzmTFSQQ/qtIqTwNb9t0GOeAzb0G3rT
XR2ckdyqXsY/maJIUUQZp2OA/h0CSStVrgggbfl4dHgZUhTyLsIn2h04I0LSVkWd
VYLQdi7d6OGIppqrDyUqryONi4/X/OX8rjgsz7mgUk6YpO8bBDYuR6hlkrM48CG4
BnMdA/YMGTPt4Lx/t5D5/ITs7S5mfQaqp3QxeriZPj31Ff0Ayahfoc64uw1KMGuR
C75Ja6gAVXPDDSDoEXxAMad+lGoYq3/mTA0LddePevGXrcDr2bFrz34CE+Q3q/2k
GOqTir4KfvCH2uEdUTfTA0FonW+tiqwPZJgxa/fmpj76QldVzpvXhVQGDx0BP/UH
Nx11+Fi84oJwra6Qabao3HChZmcKwi2l3aCpR1I3DzfCTWX3nfEmVKegl2adnUPM
kQ4lbHVjMfnhTV9gz3zba+zG1pX2c9xurX4gR6PI4Lzm+Iarwm1TocoFszbGi+6w
9OGmnPKYxFGIjIarLn4G9HGyvG8Z2Dn4s6bmH4+tbj0mwRbDMPDhfOfJUC1HJzrR
SZI39TjX9APLVMpP/BAXFJy+PaqcZb2CmHyQMJ3VXvEZaIlqzCeeJ8ZtJdcNFq7b
hHaYitUlHQIu3Op22DQSKl5/K62/ilbdLxMyi5gaTPtoZP+XqNwp+mOuqSThPxRq
HfpQb3+r9/Ugs3boksq2tBBe2lh692q5yOwww4QmbUbDmlqYGkYcziJYIKzUt3rW
rqUFZXJpBcxafa5Cw9o4s/J+mYj2r8LyjdlnBNWab31tXsJDFv2y9VZY8eyWvviX
1qXMrQvSYTqZFO5i7PtoSCeNDuf/1I/CDrvudvHUWELU4I71bbnsU2k9z+Mncwdy
FeHQjJSXewGm8NNHPiFWFYo+mLoeIcJUrSl9NeOWAGg3NUUCLBcPINUD0nFk53s2
VOxBd4XjJ1yodVZ4XrYcQ9+huA8BPkCAaIv5NBSoI4kEEBY+NnnKeaqmp9yW2eph
MSFCoDtKjdAzRDnYv7RTDM3ml+r0Y79r1CLLBDyaOVaHLYxGUOiUeFvytpYppjj6
v34MXSON1qeQhw5w7fu0OTe88lB36ImHywpAgo2+lp5yVs4qm+3Sni6jA3DiMgna
B5CsKK5ZkOdG0TtdY9/p65wZbNajMXqjBi2zzcStbV3HDTbdZQkS1isJdiPB1Foi
217cB5GQ38+KDo9lsb0R4FO/R4Xq4T54nxsnTTvLGtmQEuhs1MHtDgmt2UXU5NcY
t/rVhyqQoEth3w9Lp0yN7YuA5zokAUEqIjiqakfg82JCwJvGsyFxkvH2j7nGlYGR
gIQ7pJrm5Jx6fk01PhsmHFyIZ5z7lGe8UMIIQoPiaSCmHRorR6I98ZfJglN8Qdli
gQzbIUS6251YH8T12qKN9kfrxCzouS8jac3eTh6tTQElNEYo7owau9NdptPvpO5Z
Znbfm9UYZBP03uuIo62g2I+K2ymoNdJUaHs/kfynhiCXjEbAKmvH/0qlTyd+ZeIF
I6RtSdaHj6imuNjNoOWfiwR9XVnAVD/DGLjAHKg/YfppZbAM5qY/CQNXMJhS4wCD
bpxrs77s4UO9UhCGNpGGpzgTukLUbj9cqcf+0VgMOUgIjKAXLarZwcojb3qmpYoy
QMnN1EvStIzQmlrw/pQdWZTePDw6k+8etsqxBr7G132RrYlCCppyzz/eKhB0A/ow
xabP6fzrfCLK1q6WwQA1cWf2vPaBm5CAeSaeKbCqjeM9wSz1vQI/UrtkGA7B8EPd
rukQkcWmvJTJ0FXbY0HNYA0U8ZW/YTZ4S/zEjpGGLTsLXQjQ+4uSveEcu1zZdTOz
sQzR+dh2hgL2pB/fQ1Khbuo9a91zMBUK7os1chP3OKMILKzYGmecgJcQFArAlFSh
4jwRVeHXjcbx2sVMWsoVfrDA+7bGEFYxsSlInJc0089oeE7jyRM00DFT3+Y+qFii
EG0hI3OhjDVkts4yzChsMLgeDUmBXAox7Nv2N/2DEAGH20XsRGNC2LefRu2BKKVw
WlH0edaRvoMVXUJ7gR1bVIyYHv0G9MQkpxuxJuUbYBb6kY9RRBDb5k45sbDIHFHI
Ew/KTzl0ARN9L9/peAcYSlqL4+VnPQj6vo7Ev4JGzeyxNd06oLctS1adKVg0mzkA
AHJqfEawR8jvmUi999PkQ3fbvPkxXVaQxiGbwcRJpzTYnbnCirDTBgBRxUteeXvr
X20mGp9nFdpzaS4tINxpswo+laNAD71dHo5n3APf4g0EyKGJHUQ9njZw4Yy97n29
1iLjkhDk7r+GvmO0barO+ee0gFfAXJcBwtIJ3e02kcYRmrVpuAELobfq54E3Mb2G
3JRIc6rL0MKFi+VZluj/wB4MhpZt4U3NRund05jqBjZkLkfDRadFyox5g7icQ4jk
ZET2Yc2l27kzFhUi9sIhkGF2klv6rgNtKBihpO1z3sdwG88YY5RtingdMrwYgOeS
XcE8q9Dbjd5NDeR+w1uBdPIf+GX2zSji/nRdez99KKnG7FpP7oXbwNxZALDt6TcD
KWOam8dNsS3wr6LPYCKpDKlNs8KNfpQk3uPX6J1Ra2dWy3A02iYU3jNYCocpT7KI
fK/NC31GVeRxj/U6K8l9L2TXaKgj5KfWwwBG+cwfd3QRniSxbBwgj/loojQiIhIM
mxZLHzfEBXkswrcYuUBdAZKKXIbEVX5bwQR+hAztCYn5CqoGi+YLf6weuZ+eYmI6
+XGmv93fIG24zAHALrioKwcXoCtlmrrGlRLDuuBY0CUtIHTIkGD6lMXgEvyYJj7a
7zTl+L5QH/dn332yvrvd34nRIUsxznWAjso8icoPNUfHewarPGLod6k6l7Rb4Hqr
rTtJTqbGlOcAg42TQLFiGNSP6/tU7NPFdso+CNhLBgpx8VA/qajcuNbUoVloENDq
WLTHPN1ZfeDiGH/b04uKKuWyDQlcV95T927BsGsUTUZA4xu75mgsn6T5TsG7LD6C
t8IclPiohmHxzJLzD2X8pLesFpmVYD+GjWomxYW70dRp+eY/S4be+kTjGk5vz0WR
aL+gqu0+vfUVdAAZtmsKbHLySnOcBYWlOiARrpepkbeXedTLzqSw9jO1OINWBtdN
g3sp61IaYk39F8KGPkBqFErzcCieSKN6tMw0m1hDVPfKcfmxl8OEnfKB2sDGVeZ7
jAoxa+566o60x599Alx1Ou3cSAQvjSA8+pDKPlsiXemHr+Icldr1NZHnzr6VW09e
hF8uLZBsfhQEOZCeSn1klkdrrzCIw3wXMR6R4JJjywNyrK2NuWWYROb8TSyElXpP
n2qQZG8jSFwcPpozY8iv1d9mQDQLGe8mBaDZ11IlpnbVZDP4wGuLTys+0x3LnnWW
kgphUbzGpumO1eRChoQyM4YTcx5QE3ZHAohMyKwH7mkssPBTQRy7lhlvXHyFCIR5
nS6di57AjOKi5taa+Xeaac5gPDIdNk0DYfeOPj+UTE4yPcEMt4Ig2pjY1YzzFDtx
iLIIdUK4932KnS7VSWY1k6s4SL49C6f5tUkQfzQUQ4wSso9IL4SuaoRGD7QXbTln
Fkz5jtX7Eelnv2Ap854tdk7NiPrsBOXo463e8hRXgSMJ1rW5LyYh3nPFqucvnFFD
czKhyeqJ5mhbcFN5RrqBoyGDq5dKv5xaoGP5dtgECBKeWx2xqt0a8/2NFeSI33Yr
TdyNvulBQa9eRT7ookSUBjPYPhc5uJksef0Y9Ei8OvgrFjIiELwyli69pt1xOWgj
nyo+01nzaZBdGGhrS7M/TSdsZpS42h9tGuGo+Y83Vk44tJE8b2VszjedjaBcZtEL
tOCzhMJZWLQV5+7uf4E8GIa2krI8Gj72zt+sH6eJQ0U/HgozFrVeZd0JKsYCo49i
9TFzOImnQ2XL/t8NaYPDkUCtwHR447fQ4XlOvXULsI2x48wx6/7POmeQRxIMkL7i
TDSaA+RBS/V83JQLCK1eMl/Y1l2LW4IKf4prxLI1hmMLbWmC83NfFgAfcn6UUq6L
P2KnhfBLiKkhbHw2j2GBdkNTpNJxHFMhFVU82DYWfEfWPdUddY1lXpfeWpuIKdYF
ih2pAXjJ4u1h8Wa4RDTEchP2olIZvt2KIX47eFYOWBM9w9XhodQH+6B27rZRG0Ht
mR9V7O7hyUfc5OrOeJ6rP/lgaJreNK9SNr5uqabJsxG7gDpAA5V/MvH60EybAPgI
Yknl7QtLShUea+tSXiUrsPdyTN2jCOKdAFk8D9KAOkWxPnrCOWN9dJudrKKmUNxb
gim9CQwotQa5pQr07VVMTCFMWBkIN4UNUy3Ing6gDka05IU6duZT3m+a7K3jAB1a
X8GGVR7Fg3m0FA9HKtN27qp4Lfb4tE9ztEbOeQTLdqYWQnryvph52OVK2+gZq0Ey
+IYy06hcCL6dW2orQywVSXEEjQeh/uvecrT3V38TJHljIUq8pl64z4aXvNvk7OPs
cOvV18yYWYUSenhhlzVWtqkFZb19SG9VHteljTUegXX9CJ0TkbGfT8nadhDAxMYe
6qCL826els5GXy9ZddakyWDpBrtG0GE4270ksKvwbW/Y+tv3q2ZgVemPCN6f3zzA
jK0DHswnyscRjhGLfGU99MX3G2Cg20cLKawP1l/Jz2+l1vltOVILbNmig501tbUN
HKVzKAK+yNBjCghMT2s51BeqEyKEgUgQdc6rkoPkJV+ugQ9zo2aS8/YCfb1zlsw+
wCZ4T3txYU4ni7yoM24/4CWMjYFg57qqoXWXzkmd/xqknKJX9gc4b8O/XrayO9nh
JS+O3KvcV4Ez9RbgmsrYbGdmysdL2yaG1YipYth7X3TR/xmMnkLKefaG5aL8jEW8
eoLFop+VGHiAPgFad5lh1KsTGV4ifRjXweIpfru79TnuGZklmWDrvRWEyKhnY0pE
ms+YzJBXDh3iiFr9bp+9QY9Adr2eDRxma5JLEQOjkzGGfsJDBu9/a1ku1dh90jrB
y/JqcL1jYSvwac3dDY1TmJGWniwWnjUUkjjklHlStiRXyIIZXqo2oAfAyN0ezpIh
KErDUCmAMh+bpYsGeM2Dw4hA6vyDsUt3F8WTjyg2UqcJ3KfSVY0KhNfXTT5OqV15
bRgKt7iny8lzb3NDhU+Gkm0mzMqP1MzPAu+fkUxMn12OaQHO3jnqDlSO3sQZRqq5
9lJNgFq3JkGEOmSLBBsuseCzVyADuVJtZo0FCWxlWQOQcel5k0dF0bWAkU1yCgqg
myDGHM21wsR7/0Q56175Iozr+jxJT9mIOVWbLcfRxGh8z0oLDLwAaMAE6y2EKuFZ
dIxyprihA62d/+APCupQvErmgDOF0n1q5zVkpWdHDvpugM3xdTFQcZZswn2nZFKl
yGwgIGzRua3MOhmfQdDkT/mRNxOCBFBMI0jYUTTx4dcDdTKGzUpG0Lt3kx/xgi1N
xOLacxRWfA4/MwNB/oprldCIUC9Na3V75gcJhwA7SADeXSfyAouMRxOpRz7zSRc1
lf9pEOurCh1aeJ9c5lHfBF0pILRsBapNkFkV2pA99f/wshX3xzuZaxvhhsJQYB7W
QbGWKTdwC1zedyqw4YIJM2aJJ8zMMUePkKpi7meJAx9MUnq68qdAp9aSYkM5SWYY
wnG7iMLR7JYVEfhPtQKYqesahQEH+stJFvAPaIW3LXqve7OY73e5/pRMN58IosZH
etCeHBSlPrqbJJ9VnkAdiipOJsefAzcw+NQ3BsXHmBPb/eOV3KKWM397ZLFqqp5P
+1RwUzRHQrgKhEj4cqwhlra3NAeFvlyhe5Y1SOcMhUjK1YE01eV95ZOooHknO/6w
VSn/f2Ab8mAYmZZuRfGwW1hNstoOx7DjlhvWa7rNWFCrtXA+YDq4OfdvvViqby/n
0k7hy2StYeFgWyS5cy3XYFD7LEVFOHPjbXpkqwl9L1EUG5bMamhdWLyw4MdRrj35
jxHHOgPOhdrQcC2Qi3B+zQzXiwwLAKc7oP2jvKTZG+T6SUaarPul9134n9FxSXmY
fcTsBRuzPVXtKyQ8Nhy4lAKXlHAyxUxBWaBiNk5pn0BchDIH9eIMaVSQBIBqIUWL
Z9BEcz+gueBxtPU6+iEjwNbIxDxeheyN8To1moRKOxdBmVMQGffoa/bfOXX+AwDE
c25U2wikEVoUAsgDoM7yGNbkqWK8Y9YwZXdgkaeu8CbLBjic6VuZJs6QSMcRVHso
TD6JKKQsQdr04eOSwXapefjzsMR1glm4UHKcIWPYMLxKRhxwUXSLEnPsh4ElSROk
XcLVI1+Mo+/y7PMbN4zjT5HqNABRMuB+odbpulV40C4D7BDYRR4jRF8fOTsgyw58
uO2rU42k+2mRurQRoQawsTMkv7BxJOQWJ37eYQyED8oKr2Xhb2AfglCK5DPATbmR
ROjYDz40EmOfunsUv+0BoI0QlEZXBiTOXWW8WaGYATnNqjjwrZAMTbSGkiL9jmKK
4MSButjXVb2yRCw/VvHHjJFHYYcCJ0I7thryBGDjOMA9IT3NcjuU/n8q/DV9TZKH
6wXb/+Fh/+hbdyg668WZYQz3T/R/bLuFuY9HJktVt2FWJr8rpMNt6C8zEuRJH03t
DT5AW5D/m6/VGgjLSQAbR0LVT4yQJOYuNZ/aW9ORsCKKW8mhJ56yx7JOd6j+bPs8
1KGLCnGr7BX6W8CEkjX4qxnZRvG+/rSu1JLOcEXjN+xFD1p77/KBfGaEGZCrmxRf
vvomrPIlVPbgE5wSkfAWoDmKaa7EP/HEpad75WfW7QIgeSsBLEsgtMb3Ng5hTk8l
9nKzOdsg3OdB7NR5sd4vsKhQEdoKhGmj79J4eeomzvbUHlpyNMKekA5eXr7c72JI
DmW38Pcnp3ToNUX38cLBHk40dCE9oYkfQUddMCTsOewQ81SaK3eOPThqFR7kRWrR
K8PnH5aiDWcLcC0txugrat4cfA2PgRnjDqo1kKihA/YBF/kcCPsrxdO1f9WfAswT
TjQKboCxJ+/vO3VOnXGyciY7taafKTw5fRF6vi9zFXCq4UPQmE2+m6WYfaensXUf
R+QpG/k7XKTTd4BXiOl/oKhFZau7s95bo03WgWj7BIkNc6TlcPm3Xut4wDAfRX84
iJ1dv7ErBGE1oePK3dnRG0Eyz5dUnbECf6mZ4R0qGWv2R7tZqQgYnvboN8LI7Ve5
cQB8h+qKBe45HwyXi5XGl1TCzKioXw+VNjGjHfa50o7WPzqvm+cRbs6GeK4C0XIt
pd5Xy3AXnQxplg8nZQHRmqcWUsBymXeElS9Hb09Mb15E5fAF3YiYPn1aWldO3rJ0
0i3CAk5xVRNkIjvgzqhLX5EkVeuU3FrzBRH2CC+zuLtBbmZrUZjB468Yim591jjG
4NJeSIDYs3qmjAC/NddmCZd8RhW7wWi8jKdYtiO7FIce9OtO6pIVtzLfdiI8da/5
o/D568RM8GbU/qgatynn1pd+Y+dTyyyzAoUA2Q69Y3Zot4Bzyg1FQbpldF6DJjgc
97h+DKfiW9Eu0h8kOslJNf7pAZucW7T6IsSMJpz7ukmmtxo2kqtl/r6OIuOsGKAy
FoZ3o7jdXY4C62bD6WDuJzSXg5SkPs+ZxKVPsGlB81eA3/jVSt6rhVkJeYmzGN7J
n8ZoKIrk5U69+ULUGQ5yYQN5X54YvEjk0OpCTJ6HE3Fz2qT1Mi2QS34enISFofxv
L7PGxkDHLRyKw2uB0HWF64buqDxQ3F2kdWc4w2gLYOEFt9Oz6djzWO7uIt4MNR1o
tWvQlq1IA7UF4Br88lVf4PFhvpNpvE9eNCGHVA2fQt+TVc2S2zmqxEZm7qSGWqyZ
vLzPzxN8YXBKt//p3NnSu66/TPjLr/Ly/yj47QY8kX2cgwO3RxMyPtk+wnkAdsWC
x0RUmU0mhkicgrXOnqanLsLC4QItI3rsQeYQMbrlG4dutyYbnaRgPPtaLWsh83/8
CZGv+2zf0Dn9Txdk3IQ4HSiXiamJpjVmVWt5BItrxAWjdNw1AirIcHS94QUuH3jV
5hAz6eUjtxzomHp/SU3RP6JIGb3qQnXZrJvSkjMk4Tc63FE5WbuCn6TTbq2EWK+s
nRmjz4voLhqCikwFn094JCjDYHj8IbVmN4na6wnTmdU/WBNW1PxvHP9GkakRd/8E
I5a8ih4QcCZFdGttws0lxnOXNU62o1gRu0sypiE6FBl4e+vAwTuqOHm3XHNq2mAR
D6znUGS5TXLkMmrF/mvGFyTQ+KRK/G8orB6S+OvfJMt8xWgzFdR75ghnaK2S/yR2
CX1cvV1jWtD045VP0vN3Ytkn2CkI4e+d/CLzv48DwvdefpKOWbWFL55ZG8sBIcgC
ozAdyo820oZiP4wsvMiZfv9e+rWMDSE5t5PokUyr88DNAKhKOrFn3kirr17HqJF6
IqGk69ghFbGyigG/cV1hlW3OjHAxk9C+UqDUppJq/TmZjAjH6TtR4bX5ynr93fX+
BD6yAjAbuGErcCyIe/Fu0CEuXHlogU1vk7ENnxXkXwuDgI/wy6BrlhPMgnZ582KJ
W+RTd6eXIbugyTNE2SsKpkqypMvgByfQjgL45qoPC+xosHw2/3BnWM1iSBDKrGCm
dZnrZqIu8sWHJzPLgZQN3jBkzsFlVquJ/f/gi/9edU5NpnEHYQMs4GY3EYXCs7Y4
zsgxAkEtI9QbXxDJpqWY3L7lAnWQqki96GBVDo8TScjsDntFD3Bax727Tuwmifam
zadHbnck0YFbO34eE9RooNtVOjUHxbRt9EFrKypo7RvA7B8j+Rxp/YhzQFJqNlLA
6GqBDEBC5VMaK5wM45YHEiKt0gdlKivrIK3pPr8qoKuNFUxXG50L25K33o/qJhgj
rBe3hS2LpqqKzr353/z5a950XfbTT6l4arWwKhV45cSwcC5rLUyl8HrBLYln7A9U
2s/4urrGX11O9fr3jA3QRZMhSOAkiARAoym3FwAZGvEqdm0rtgzdDEBvQt2e4+2q
9I0za18L4JCiSiVj8WspKIUTLz10IGmxCO6INRZ1Sk+jGxSCB2+Ly/LGSI13+5dp
N6qXuBZacW3ZlTfTFxjta2wk0v9t25uLAvxh97vzaWbo117mrfE03tys0fX6KPQM
zGwnOpZHuXCwkMMwc3o83seoZLhMABHKaDiRJhwtnrqvc3878VMPY3xAbgBryRrH
uVW2oS65f0JioAwsaDmzzz1FwSHgolubpjXjfwhqmWFLDxqzyUvy5Iqn475c1EF0
hU/n33j7Z3Zk3HfP+lErnLlRWe5IKBeBALuq/a2PJcu2ziqnpT1vJMEyJUf6C9PJ
/mn/ItHYbmJU93NLexKakueBa+/Uk/nbNYDfKMCh8yqIFmLshzqSWXGXp2PHknh0
o6C3OOCggMe7Noku7Mjl3IKDTm2zcMSpw2APilNITAm8CHJEX4qDiyoLsjnSk5pQ
1hg7K8+Pw0SErBP5+D5o3Lahz8hpYsc2zXBpe5/rS0+SSum8RjPZYSecHMZkcoPl
41ts9nxQUTWhHvuEzks6xEIM2zzWtX3dbBd5B5mT1TAtbW5m89mbaQ4+uURutFQc
0kydrTg092Ix3WYDJ3buA9cXgSJnUhef/GKP/TkFX+HbXwsxDMLeEXZhB65OuLWk
pNfePFaDlD0p6X2g774fP9fmqMPBibbyuPxcDbLz93phE1z2L/3yry3KnY0ByHaF
lgd267nCzsRQmpdLY9bCaMRsu7F+pdBePKLHS2JhgLIN7ViXdR4W+xLu81VncuoD
H2x8f6ky0qvwbXuM2Yr+Jee/9qZbyLHLCU8Be/SNiIBAiK0MUrx/lsX9Qi/kabFS
qvSprthFuw71kEWx0Jyxkzz7jho8I/VyusoCfTrQoXivh4JeKPMV0+D4DxR3bos7
PBWImX1FnfitIkhp6mS6S9ZTmXXQaNgmXp0RtFKf5LcOELub7gSd8rSC6s8mkxVz
aMKXxBLxtlZ9e6xWK51carmz8hBOsfLnXJw+aR7YiCpxEMdxo/nEwikOg1GEdBwt
z0SZofkodPEE5oIjTVmn2whAPRYIcobsUrCAU33FKdKu6hUNLLme69JKt2ebAubu
VESmV/eWf3QBSgxTZlwX3E1fszRxZ757mwvH6EbE69P4nM6kti0Ql2Pp8Fw1X6rx
NY+QSFT4IKXt9vllQmZ65apLFRBhKBE24zwnNPyfKHgvhQx2RSih4JwvydZ60a9B
hUiBHTrMIPiBybbt+VoRD0QRVt2SqIQQ/6y4bOR7GfMEWeJmh7oARdu1li1P7UYe
MdrYWrRb8RXv5XeA8784ri4ZoCN/CxGmbwRhAUDD6VsN4NRMDCljlGl7EuLTo6OU
r780pEpCKZyJjBS6qqPGLu9qEdvMDMDK5zObJUBIOxESX6/7LtdA9UxkWBR4XAQC
WfCUdciXjOJ4/xGjIJtEuxOWMmr3YeV34l8PVZVuCWyDhL+ULPKb2SXK+A2SSjs/
T/B1xrEODeCRk6j0+PP0Q1+n4M6PvRDzPTHYOK/6lAEfSOXunzxu59w+OPjH3Vux
JCNhKLQOaK5Xb65pla58B8BCr9HnrJZ4FRZFKnNJ4Lpbxk9PdU70t7hSPuGJJ+vS
4F8chxnbjWXJh5q5rtKmjmOIGf34UPBhntvhdIAHo4Io6qGGupu3FTh11xO8TNiP
iFVosBd8KgtW4VZaZgxfJD26tQko/cbquaXIeYmoqG7eFKGAsYUtadDSNPzU4atO
dD4wPBHqVWPRnmnKej0Eify4YaRr8LEiOkqLsG5bu1Xnzj8QVELhNvM1V2S1gp4U
9YwHLMBkd78JezPovluSV4vxvpgr82ch108Em0yyAi0Isk52nosaMqCxY2Y2JhiT
XKq5YEvutvlKn5qCdtxR7q/9G2TeWyMXo4u5NLbB6FmZzGtTiqfU0ljxKjhr+kvy
bZwCp6MXpPDTbSqC45Xxb/rVY32akdAERtmKXhICozwxVyqEAv3RNK8IlIpUiAel
lRZBBz4zgJOOOAujPK79IYb0Gm3ITq58xdOAWwHIHufS6sBpCL/QU0IsjCLoO9lJ
sJSMd+bFx/GY/UuQ/9HAS8bCg0k2jOvgvZYRHtaqFrzTWXqFlvUiGff6n2QQmYR1
WedTJ3KYfyi3xe6Bz+q/luZPcutIPWlbFQmTHsIbYkRc2DGTllSEZQwNVN9svhwy
Rl6VVYfNCLOMPH+Eer0xp2FN501FaegLWo/9tC8rEbnpbwFwkYd9SFpVPoWJvcfi
2wA5RfqUMncap9J5flVs0Fc+1aFdil2g2UxTVYGeuOyhx6ZTv8rcFRma+oceukvT
MbmKY5utPZCwWD6p0km47uRa3LXyWItlUXbXSzxgboCl8aQIk8rbITuwYPJak3Wv
rzICsa+1EE+Rvn6gBkYUC+yLptDzMTkmCh8qKxNnS7li4ZDHkLRpb03yQ0QFAuda
u3dRSnhaqemLe+KU94SPkH2bPIalCgwCerwotjpwEzWuLrtAEDz8Addta4G5q3yV
ATElNNs8HSOWEM3JVf6DshCwVcwdNJmVyuhWb0FyWnVdM75z0eNK2fBhBxLwpAaN
OHNfvfA5oRoYk23ocX3rZ6d9Tdv8lPCzXJcmtXgHZljjYcj+FGZQljG6tu/tzLJk
Q8Z7h24JZH7J7dniGLPmudch1KNoZg1leF7/D/eoCBgEZwcRIfa+Mc7ALfA7ZNow
SoJG3yrv94+nqKRynsT2wQa3qsl4h9c2A1xp+RiZfkxckcZrx6Zw7k80dBrooNQ5
jfXEPFe4PpA53xF8dj23CSvkAGrSi4d19jSCsw7S6Dl1Y7hj34vtHBOf69+hs4gH
RxcQPrYZMe8Y97y0YaeXEdL+reHSHYNEdgBe+2KlXlsgUl6WPh/o5q3yv+rhpaOi
M6C+4JRCz2TPH9OMBavSVLckK5U8zHjDPYMinWT0Hjqbt28pPRqsjBs/5JddIf7V
Ij6y31PzouMPPdoEsDa4ryouX80Ne+FRW3gx6EtiOCHUB8JRSfWiyw7a7Xxj2kPc
QPs+NF14YWDc+K2UXVTBvc8x7jTloxFBr81LNy4aIha+cKlFZZ23exKZHPThnIby
ADIw8lo3YG+LUIpGzInf0W1eFWL6cWQ5I8oZFLRsOgw0zPb3+IcQ9zttQ32LNEUj
+TxKgwiuwIb6aX8KpnVvD/z8D3poResP/Z91cWQoY69RCi2pmNxqRuigItRN99Zn
Y2hL6RAANxg1mA7Q0RLH49QXGzrJRW70XXsAUDC54Z+lZXMbHXTDvLBMY469hV12
dSWNALlUMtPyoNMLpwxfbcfHD4p/Af2gxuYJfNKvxHczodyFl97IPfvBPOJ61THX
uqiKKTLIYwJlo42jpApNKn0agZzjJNvWqRThzc+gZwEIyP234QDBmYVcPhNgwTd/
BB3i4qTlO/LgnjIPoY7k7OEp3vfgWOjRZcpm32EQiwSNBUcQt6p9WXad+xR5Qmel
YEqQ8RHEUafu1hjHogTMlIUmL+oo3TR6gPVUOGAuctYjqv+PbBMZwEIwN/vnXg2g
u6SzDc40ccT4dpfAkzVAJWt6wgdjtzjgWSIznM7Jl1CeaM4UpV7//V+VfdzSVygV
c3TOqiqYN8cdZ4rWgvZKtCHH5nk8iTuE5tMuX5joOcFO6rHfnH5NPHQ+MxNLaZLU
iFlv1nZGTjtXWDl6wf5b5RLouVSxQmDoeifomcWWEiPnydl+pjmPz3FFfHElTXv8
uuUtoYCnJaiC3UOjZVZZEQ+k6jNmo/uLyL6Jo8sFx8tYMlzLAzzINEE+VfEXfSN/
4ID4ObbE3K6JiWQwSP9jZGFAVw+9rCd+eHk0zbGubbLoeRfjPOshSDku5/N6lq9r
HEiDZdhuZ78MDO+0pdikEnwnwbXEC+QgoVTYaZ7i+hvQkh6ZFGqZopwzVYKIJQGw
P0PTnVHBXYD3Ql933XR9Y2MSatbP7ErDmZIm1Db3eYf4omY8pquYSQysJtg3d8ku
buKV2b8+N4Icpy6eOK5QcUhr31SSPScAs1iKik1iAkM707Eda9TtG8WZm6w2T8vf
SRiuzNhh6t/jXI/Nx4VPpAMKZGopgys7sRcZOPxPnrOU8Yeq5XcbmvlO5AEGsPYf
MLIatM5hJh0syejqt7JRsmccNCfynG+yMLSgvj4vzbx/T34gwwoCM+daYyBvEtun
izI+JZiphncnYzkx1JFi1luQMNNpFbQaNEt02aWrT5R3FNwdKvlSqsh4neLaFvsV
64ev+R0S4tcsQ/3uo/fQpuCCig+Ds0AfPd1yQSPa/DBl5NJ/MjFCoehmpqPCiMxC
LojbkhlU/4a7K46uTzt3mkVaKnc/FiU5zQvFItx142UFhaWoVPa0N0v/QnbkQdKg
jTckXMrCXjuXcNQ/CAqkDt6FwdHQIPDdyKPjmwUihXB/CGFhV2LH5XSxAdeGOFOk
F5ek5pmlFQCQrht3IeAdJFBRBdyDuFcUCh3W0yAnPaMOpp59+76M+jNc1blLNU3F
7Kduib+hSVY0XXsfQFeAYxwbWgZqmBZ2qBwR/PleYeJPfw5UiEtsact3rTeJyhZ7
7Oa1xR5UAkBWnWBEUO6Y9juzWrTEZI48YH8fgrzVe5d1Qht2fM/qQkRl7n724/+G
mmAEhk0LO9yaxVnR162uKMsXnKDOiLJWK9BT22dh4THCL5LlDIjqhn/Q5UdiLlcq
gwZwsLU2U2qhj3DIuwfqxuEO3XCiyvTk/BVnbDpgfAP95E6a1LnZqmGK+8mEnu8A
MkPcUztcSXrjvp9i3HqZ8HvuFgD6v722Auv7oOAqQXxTfWajf98h2TfMFF/g4Bu1
ybAQWMcIE09jc0pzLi3jnNa5XvyDo/45wjHvUwDByMRw4PrRmHUkC3qiqagSoGTn
YerENJTy9hnIcqO+ciwwNVGVRd/KYiUan2JDEsqzKckzIuvh/rDBBwOtVGse9oif
raW+LjvnrDYf5Aec2082NjEUN+OMHU6yHUj6jr7KAVRM4XRt3H1S5n0kPv9H2glB
qGZr5XJvPVVlpOuusmykRjU8AE4R747faCFM1tXPWUSnm6/n+ZMePrJmbMOCQikK
2A01H4yfTyELn/p9atALCJNDqMU+ZXA5cSajtJf1yxOI+aZzVTFTQgLHxIbEwT5A
LpVJzOU/xuU64iBmVL2Nnubi9vTpneqcrNbzzK72ggXMih2K4+eeFwcpScC7P6Yg
DcL+AmcKgteABP+zqMX687S2tcgISs0aWVwt8GAIAyy8RhygGPdpDpHEAr15m6yE
t5hsJq6ees1vFE2SZ75bnW9FNUi0/Vvfl5HZKl0Fcsy8R7+tVwe9o93ywR0/pKxN
5r2fwDDG79KgARC8nP5+qtsexXlEvKVISDBp5VbFH0emhcKlq4w0IKQtASPr25y/
4yMjDahhaIyGaz9yDiDxJsSinHnQgK3Dxyr5SmLRVY1fycCYlhhz8QB2hsbzo5k+
Ug7hfsmNayqCUgfFRejQz+oMoV3HRN13WwB3MH6WleBLBE90gHJP98Qv3BDcC0P5
aq/YwuliIAukYov9rBNhzHaoLPS7jtkfNYRSwF4N76nu0p48+Pf5TFatewF5REZK
NB1lnJae3HnVVylL04eind0OQmBos0dJV34gVcJg7Z+d601IWPqftUaa51muGIcD
OnvuRL92+2GNNKG3hIC5Tv7ku0MH6Njiy08kaouVfpcz9j0I5g/SP/tQfPYL/kgt
nEXx99KucEnUn8MaEbJ6J8P+OOqTmSDAtqo2W+Z9jccSFIX0kxce42Peq05jusCv
cFMg+T7byXI/Wf8w4WKVkDlpQi94XYkqorNu4NTpfF7WQ9WXQqLTcz1KbxtqGPDb
yQU1ICy3V48TGYosyAyk+2uKphURle/FB+/mx/Sj89IC441qs1TWKFxtWzTv5izw
ez9MpbDBLrSfkwAsE7UM+MEMnk2MgmZ2fFEXwn8sNg40Ub+7WbchhJ8Q8xOujMP+
18IbD07khW+V/GF1lSCrt9A57b43UwY5Thas5RBbrHdHr8xMVq+vpfx4p9N03AxU
T1zKSCtMnBj6cbQ3icBWnZ+youIepdiXBAFYHzKrNSkvhz8KoBMLcJ/ZAg1hYQA5
iB2uPUtqRlPXcoVWuZgc9BdUf8eLSQYYJavHxGIdhLxFVX8yeocr6LJ21StjRTES
c+xY79JtAD4VBRnZID3x5ST/KcpUB1B4lDuRAom8hYx/3nJkqIY0vt9+16D+hti8
DdUyI3GTZH8ZDxMCCn1ZqElt5FIXjzGARudlwFd4t6265RYRcO6XIcsgpqDI0UL8
ZfBi0oNkb8t21uZhA1xuNcTStLMANV+5o7/S4jP9kA/8D+jeC69S7m5TkLJMSXwY
F+CIoXSOFMYE85kM85+AMYDToOzdN2FdcOlrsxsis3fSkgBhoS0HBLSBwuSLWpK3
M5LqgdOuGQVIZoav1YG5yKNuohmI1Mj8b3jTXOrfWkdk2LDCcJELEgj7Y3aENMvf
kYXGgoUDBgdgW8kH9+HXeANMT34/Ep8Ex2PvPi0IMJ6uTN9sALdBhI6aNSjDqR3J
tLC8BtxFUInJCwLhEbQV9NATW7H2JNvjCrEjfM9T4a/1gYesyXkk9CrkXzka70rV
CTVqER8SFDet79L6ZjatGgTf6yq51d4Itb9tSvHL5oRanQtAfKgi4o2MM3MJEQQT
CywnykrBQRoetCISXhPvoF+083CPLX7jS+TS6zLWDYg1Slw4vN1KMo8X6MJl7uQw
mGREQIWOANuwQfFusfSr/SYLmynIYr6+LLIvIukH3cPOS0oCeEaIK+kMJ8jcbRiT
mSvKr1UVVCnQ71XnlAPw33iH8BO7ZeBuYUUjQJLGEE/5dw3TZDSYZ1k0GH2Ta91q
Hi1VwQZFKWXv9KLyJsaH7NpG91C7EBWw2Q6FBa2I4kJExa3whuPeCCtHzqPq4yjD
R+WK47h15AYKgs3IT264xtS4yNdvb18sIKGGoti3o/gvrv8fokdNMpacPptXTAkG
V7x7yRVEeSo8IO/oRKTv+eGl5gmhGIW3T994n9FZnAOChbvh0F7HqjxO74kcV+mL
bSwLpgHOfDZgauew4EQ4OdhGJHaEQ2aC81o/GCFcqjTdK77x3pkePmv0qUn5LS/Y
WShil3FAsuoeFhi82QpQm5fKHQf9nxPEcmQ6AELMf1bdNws8ILlndXQg0AlRe4P0
Qx8+2H+7vIaOg0Y7J6PlysHbdXt49+ShgXEr0IBfqmMJE0n6E8gVnDBmM2Ntx2Wl
Cq/G46ayGCrteU5tRZQqgZvCU374l71jCTAIWuBB4wlzTBbuSKx2bOFXtTQUE+/b
XF4+sdrlQJWLIN1OjcJUvD1vucPDHFTXZPyu+YaU1sE5ftr9wyS6JsKHJVJLstow
OP+GU1jodncxN9ZFSoBauQbp/qCrKqvyfJ2I/C1A3vRnstP5Cxr6aDmSScq52X5S
/LW2xH9nFgrkgyxxrx5untWqbAWGwdtYktZ2MEE2WYqexS6PLp1jTYJkMkpxdBvk
YdGDjDAp8dZK7M3QvF1Gotfg7s71tI0jtUs604PodVufLjiA3M5mV9mZquINUdCy
TFRaz4lrmHPMVTW53882hulpwLrgKduk6n7WZ3pWETwdjsV/ShCILHZYk4+Os2pm
SK2XpOggrxXrGnOIZ40Y0lQ1YzgYeVXoInIatnbWKvNhimcDcOojUb4eZ48I16+h
NSgOlMa0CXzBwTziT46UPRDjhslJrIJFr2qpZ44tba7tPy2t9MPBjaePWwLM+xdX
rtc3qlBQ7XDyFmSc67DhLiu2UXsmvIcdCoZNq6zBcKUnuYvCMDMvJqcPK2x4oXsG
zVSVOyoVBy8ywa41Dmbl7dcKsLcUsLsbLJ4HA4ZUKq689XkCR4WitWgHLqLFfb4o
6QbtyH61KFV+hYk3BkmIUeoss9V7GmJDuvdmP0BVMWr6Kci8WQoQATglh6w7ztqX
tcNV1elW++f4Ft6MjcZccWkoD10u8v1v4mnnA9jXm2OohW75Gg+rMILzqdR1RCEG
KSiOHZIVnWXCP2ev0Lzxtbnmx0e4jf5FwPMFo/mwlmOQrtS38PbP/GtI9EdMmEZt
+WVPsdU/jk90y1XxI9q8Nz6p1VwiF0pvmuEA0o8ii/5RGWInat7noy8in3tqDn9c
oFdIgK3Shfw3JMQmrdysQb34tp/hwrV7qC4jBGuSEZDiAxFYAxLdn7z+sIfdcCyR
/phbQFRyla7lawIqiEZsj+bZL5t9TzgDxmPLESR2BghPZ1m89iOV2cQfohgXcQuB
m3jlv47KVeoKtluMX7x2ed4v4xUivV2WR6ikWxzV6UChPt2Im/98LyT6sVZkXOSM
A7KZ7sRG86hf3MEyl7AOT4dSovpta4b0JTI23U/DxMyeAvqQuq5TBSJTeZz03R08
BFLD6jeJbKlKh0uatbgdJQReXls6Yw4YCzjcdBoztwPvKZD3jn0m8G4PeVZZkAAT
2AvnAHP/Qx+BKQgsoi3d3s04Geieh7jYqvlq3+L1TcMiNcevSa0liHrUR8WbaOAx
+ofCqzQUrrEUqCWX6MoVtXEzxJCyp+Xv+UtAnFMl2E6MoqF7YSmXfBLrGx42H0Nx
FGQSELmNLO9R3ZE3ZlFQAtFIxEvykJIB/tOGesdvqK21mPBN+cg5b1UiF7F4XThb
9hxTixUq6A3C1RRX9SZpRoVqmszP0xI7bbyfirk6jlKiiFJY+wSKTiN96mnK5Jqj
KSNx9D51Wi+sDbM528VesshomUiyyOxbSgFlG7G3AnGMfvLQ7DGn5NuvQ4Tx7SrR
Pz3dezX0Za+bHt3CK3I2PAEpLn21xG95wn+oVf0nsJX1rMDUewIr3n1TZwey6Gv2
E/XJ/6gmFJ99krYCM9CraXZ5TppN2/MoKTEnQopdpDBPHkoNMElvWEmThG2+U4DH
kfTW+1mPuk3bd8XltbebAbiX5nxDeMPzUy/IcOLhBCcWT1wMWbB6dCezpvC4o2Ch
qzlIV3RhRkZWgvCOtW1OZVhXXdDo6i4JmO0uLo9vtPG5VBH6jpcioDGjse7CndCZ
Ber5fHGaBvhdw7xmwXwAUFZsl0jjnogC4dE9Le0+WftOE8P556Oeigz9dYPgVMJg
gvG1FCqtp2D7nG9lUMYnJBOkH9QbST+MrNxGuI9CEybURvhZ4Qi+X3nyV2/sow6g
O1zSv7jdJSZEA50rNMn+dwwqDmHvwJrUvHl/Mda0IefRDry95CZfWxZje1B5taxX
S3aH+fGQ+r/c7TVfictS9Ng0XWBWRsjzkBxbzYhmURISjcxQKt0nlyhd3iaWFsZA
g5OPTe51U5vU52QrG5shw4C9RlNirAGazLPXGOjzS2nRnrA0qiyz1XyqlHrArhUH
8WXtgGvHRytYWld14DFtUQOthlxDT0ksbzrBKzf6yIIokLs/hasZlFRBZoB7Lbug
2b7SQ1MykJwojISbWxQiqNNRigi9iRPIKC6Ooph/hXWMPjvPvM4qvdzD/T+YsjT4
sWVSJ0dF2klKl54qS5JLIFkC+PxDmH2VMiEzfCFt0MQsH4PH5kydp89W+um/QODV
HU8IjH2NgIJhnn9i/UI+8I+dFmsxHAViwa9JyKBC+ZdU9R5cY6WTAuh5SuVGz69t
LsJh7bO6PwHWDjR0+9cQSsJ2hskNp9iC/LjF7xYU684EZaSzg866/qoopG/5gqnP
xcPaa72drfHQ5cRH0q3lGMEG+1/+TcKHQtesCAf2stZ1M2uUjsc6XOTfdTAJFYwq
oGI0IG7hegdfgUpT+09y9OJYKM+TlAbUHZ/nvaTzMb44Lj89Qe4i1kTlas+e5eZf
3TAZBAV9ottIUN3wCOj5v4NlWhtR4Rpx1MUdIyhCUEwoemwz6pxVIrlBARs5ytly
9CsBpLh8DwP0OlmzpK8Cyg86N2sfYN3IS8saLcZzmCBvJD1U7ycdzDC+gLI8BKLh
CTHuejX8kqr41Q3xcKCi7oq46Y8yHJJK4Q8wQAEDspM9OgfiCrvBBGek0Xw6bEkL
7NryPqjabbDx0HKvXyp6cJfkAIxyRDsnGKLZkVq/0S2k6zAgv5AYqObHH6EA010v
r9tCQtG1k+E5v9tmI8BJf7GmJl5TuQwCgb/Lwwmx7Cx75Foe9grLsk19KXUIXN1Z
lpI+QmqU5hkYgQygmpcRIByoRW9mgvUaxjZ4aC+aKwX3WWYGDJ40u/oWKMhvvubb
vEh6evatuJen4cN2QuiM8pa/MuAqpXGmtTN+7ACNrqX9QepE5MzskkOlx6tEQ6Wc
rt+AlIJDkG5Ty/8vRHlGwgsO8C/G79f43gu/VUc45r64W4xR8EOJeV80uXs1XqPB
eXvRbJJkHWIzzuaWXfu5LNghkf8Tf/n4N0v4qDs0bjPkC7fWlAYVmeamy5gCFCd3
0sdlVf0mOg+Eju0f/A3rlp0Sst2nw+NhOwXFaFPVEVkA2kXKVfmQu/KDuROFX1qJ
KICO9hr9wWKa2ow3868eIFtPKRlJYzXVfgYHVDrvWS5N1fn26u/dZaACIpKflt66
xDCnbvut+QqvDHsEKedzTipEEaZlLSd1TBYr41YTJN1MRTkDfQggLfOzFE5DFHRA
PHTiPl4ETi89OLQu9j4ONp3meRo1ydl7U1NGWIMqY29fJXlZ2oXuwkJE1+1kUj0v
WohM5PrOD7RX5FZa7/NrtSJMwiAYcVTBumu25RJ83V9MtOXlgdAQZa+HNI5DPxRC
U+9Dp783Lrjts4Wa1u8HZ9aigc52oTpC+jwXltud/vawGgZYP00q18cJjtU/kqBA
OjCDTPWKB/jVB63+2ig0ajCgUYgJqSbd/lBVEdyat/0wJcAZMSLuCU2fUlHdhVOp
YSzB3EMAVAtOmTnk10lgjR2dg+7GSb7IoVj2sqM54ZAGx2akSj4sq9n16eK2KFIP
bLjf04xx7IoMornF9ZDPIF9qiKC4XUXOpRePPBUL56V2jXJMXrAyPFU8PIPfuxwU
xkMit6tMBd4nmcVUphGihvsy5YfET6Wrn5TqYC0pHX2o34wc/y2VisqR3hWkPznq
80ROTh1eeUBKS7FAqIqgbusdYH+QkyjiDcgq79X50+9RPCawD6ujV4kmeT98y0Je
py/PHlhAxYvlDNhbgXPg/SY8DqkLbFxxIA48pL8EQn6s1tVNSA3Y5hyen/sLZiWN
Azg6xvzN/bKDnpFPFEsOdfvbmBGoRoExIkrg18KL239BXx4aM+3IfXETuQkwBCaK
4ucxNsGUqJ9UP/+reCiiLz4qW4SOcMrQNWHUEBTh/GSipZv1JL43i0WZb/OwobQw
mPkU35QMoWWx/0qEM1tlEjC2+8y7aVi0sFo/IT5ZHuM/EBJjfDkCyYm7qMIIJ/YY
fcg6GD9sP2T2sxkqWGjO6EmneOyAWKU/lxD89ff1lRPAbMvZKCbp2m/cW39milWH
WmbB8Pa8uFPHdTR6HoIwntzAJ7sH0D7a60VIIwKCX+DsBh+4IQ4FmkqpEdi0Tyjx
ASgRgoqLz2Mzn6sw2pMbmRGGX8hsIwiQ65RPkvOUWCm00EIFxlKXuSb+n6pEYVDF
mU/JrqhT7u0zTKsDdHWNkS/oAhH2yFYUuis9/BrcgpeUITOOGeK9v4ctKITtDHEw
twVokPrHJQKeqIpTBKaMLrXWsfx6CmujdiWAmayubeoKOwLQs5WjH7OUueXWoyfk
uOeJrwdEWDyrJAkroQuwpC31r5xc5xS7sV0zA7h9+Txqzvzrv9lvxFd5bIaLxXhh
z03sW0MDEpo0uVm26F6TcuYmXY16H0RhLiWYCAEsDzT6xPYJhllVDTPCCH/Yzi8f
lkXYvh4UuKOXXm6DkFMknO5VpfhhHVyKdLs/cPuHCRhUCGwtcAgnK2hHQGUF1CSq
agdaXEdGLTPblXzzy9jWvCZsDzm/ZXncIWl+kc6t9HTpGo3FhGaP355G2Cij7hAJ
GcXIh8EQrVKiKgkK0zQVY98ydPdirL7PaL3/lLvBCdz3GVgASCHYEN5JQ8VTXOGc
5vA2Oj2wioT8V+13QBIXOsmSbuO/NUEKIpBb4iVQLM7Bjz/06Yx3DOV4wCTYOBQx
PvZ2f3ttlRtaFrLwZcAnMOAxbOlCqLygQI7ZvCwXIfDliNfHZAKWEJ1yv9kIQHhE
tqHhzGrEiMPqfLKI2Lhb8NvaYcxnBLTwNHO8GCERSmTRSU2yU/BPgMYoz8LZZLZG
29huDKsROZmYfEssOYwGLoBqLAqOFvrmb2+w6DL+L81TbyfJvIX8Dy1EZVdheMzV
5yiGasr4QFJ9NoP+CSBNcQ8bGmd0SmuSWUB5C3vH5Jk0BATpRXgwLc5NTzMK5JRV
gNuWeNjVj495sYAghJtPWyGpRtuRqrgCURXMiRzirjY93usLZq+AeQnqQdKXsx+d
ZrTIoqnZnIJ2pyhbdBYyD+Fa4YKa81fO+8S0wDMpybCWG727N1B21Sal7iX1bD0y
DRVx3aN+uwd8qFjofmrQWNKhvqAcTtIDan2M4ECY3EBIl0pSqG/CtCiDjkqUs1F5
TNOuZ97EW5jJztELbNBo5lFSUbTBjryfGq0SiyItMhJGGcAG/GxuAtwK1itWEg+i
XU2yH/vwZ5cirdKdS+G+zZCoUETPP2sWlFTR10T9Tu06kODCcKVFvDO+HDlFoUL0
tESd80H9EqhnIUwVLc6T9IFoQpziTzM7g95bsvb+yTwulN7nBgOxuOc/bhcgVMJl
VEvXDlXtc7VUcm0AnUKA38lSvB35zzZ1LDvITQT7cS9Elfsc4E8jMZw6agu0+3vG
L4Y60B31l64hXFbVeayjFfhckSN00NjF3+QPg+hdWlm6IFVPAQshn59zgAz2qla5
3VMgrDSsih/sSCfqjEZUbpeHEveX0SjfhoLakxsLA992iOP8HV8zVfPXazsHtYXk
AtRWfOV2YFxpmWdOmlN5XmBMSXXPzk9K+Y2LN5zrbJbsgdkRg9Rpc3T/fi6fg72k
UXKBHh8/+UWshAEpgJPuxNZNpGvERHpSkkRmqEWLYE+SpCU0VrYkE7H4OT2APy1P
YbWxT+zpgzOzwloCcP6KHfgR38MSgpHgwic00sgm/8nF605OzEYsrurgmZj9qIMo
5EashidCkCljnuj2xxXZexNwYqCepo39v7Zrdwsa/PCwqwVGJgpTzawF/GoCOthx
ZgUSHjQGzqF5VBXEcjpV1AJyWAFZrlS4ZB/gbo784kHfnxfcKyZ1Btwq/FJnvbl4
UE5x0rzE5tGJVMkp/7tNFFRMz7przjaTaZoq9KapJQOvJVe7wU3ZiNtoLt26zeOC
WoUwhh3YBEFlFJ5rQKRhjtbZzUDYZNCtm+54MZN995AVYrsG84t7Ec/A2eLySY+R
RiZF0cqWOyNovhFxgoYb0z29LP0xLOxryy7cERr1Yta2FaTWV7yow53nNM40wR7s
Y/XlWiEfqHfSCd8pVqnIu0a/HJ1J3JZGGBQiqP240HdNVSAbQrEIY4X3jA4Et8dX
qqhGilabJmU2+MIwyrgDI473QOJoCDE5q1t0O1MMZOCRLvuIXVQBKiw8oOwr6hwy
8I/3pl91NoZPCBEmLBk1U3+KOqQhGMmD6W9NZ80WcQV8p6T5heR6sFF9Bewux71S
pmFBtggtUyTu19dOwmgvJYr0YV6eu3euvY4CucU8MIoNsZxYvLnQ/5uHEJqgWLuY
Bj+lkguFKJ8/WiKnqAeJouWgxR5gAdFUqSsdM9OuxR67I4b2dBOW4Y23hljBTZnK
XXA10nMrJARQLdXrzY01i0ZPT9cyjh3BSqyhj8tfVEltimTbPPopLXHY9leOghAd
oqh73i0Ce7/bETfQh6+R6LqoCOEJbRxL7/Ynou18P3GeTv6UFL8+0jotziuXUMB3
vOXVyDdoK1oPw7auz1a9ECvRnHB1SF/RbGnoV/ytFXdMkja3SdpUK6u+DZcvny0F
bk1Nhbu7wi9F1UakeZM+gn+zX51efut1HSgc0nhquqgX+rdXhTIeHSAoQA1iYV2X
wWYNvPclxyEQ//BV08nbk/hdB9lEs6PgxGeNJ1idPaKiIcZWN4ec1hb/1ffJ7E8j
3fOxqYdFm+7FMSCVBOPxGYx3n4lkcl+lfNZxHF0bB7zny2fY46jQmmEwD50+2n0d
4QlUat9qpfv+OmRFWoU5PybcNayUVAPLyyWjMLj0EnYgZvhJ8QEUYjm8DvwG3alZ
0IgU259/kqv+hqzfEx64GnvihlurwHPTDe/zgW0uKoWUSx5UiIW1YpnOcgGavbXr
scgPN/G4dUIZmspYr6tSUsglWGbZfvkc2oTYVvTgVIuaNYXADpWYYjl6cgWX48Hc
dbpo81o0v+CnQWMiln78WHfuB9QyMnvw9JLOFKV2ED/YtKcSaCUC7+nb28y5tTPB
fGUwzNu+I7W3SCyxmn0Bc5tJv6U6ABWjWav7Mz87AKPRK24B14/kCW8w36vdiMJA
in27pzcPRmtDCPH32uTyWFw0FY2Yo0+vLKfdKe8w8h09GBaRYvAtIxMpevWzpbMn
Z3E32VYlojn9wVnwNHuOEO6AB2Vjd1RmsXZoIWqb1oVEt8biiUxRgHg6pkf6m2G7
S0BPlFWuGR5PqTaNvNepiEOWsPTC0sAYSxRDepePnT0+xx0swvMSGZTPZizUqS71
2ZemEvIOMSF7179MQkvuyBCqOiqA42w0aS7C+Yb1C9Rp/rewLuEjQD8hHc2kNITH
n6TClflfyIDcB+Le1Yut73/ImYUipFTos8xI0YlPHHSxgukg84MgKQnXaM1uhKaW
vDuwZu4TLP9Un2MgjKyG349iB9X4zTm9/QpI5rNvo5yFZrmQhNebnnZoY+lZzHN8
c0bvmjlRGtGa6pIocrx+pF7que/IQI6SHvh2/ocTdb/aqErXmQj60SKXx0ne+/Ky
u+UYf/8eSZMQI98O66JsmpwdodRXJGUfncG5lYk8wdNHPuPnSf3lgy2/uR5An+y6
omz2IatbKTXAd2cUFh6fxs/yhydr9i+NAquJzmrA+qofoV3kpZNxUBprDht5SMiF
6INZmx2l0I68R/i+IEW8+DlBe0ZpR/tO2m2SyFp129b8w1gQRkOhltLpfGj6AdXi
HszsUfX/F8x86CevgfjDyKVaTWZxnrz4hCf1YBmm+axUtwInRcf3u6hrJyTYLrIw
s64fOQ/7N3XXYcsjlFBlTYl/MEGnEqICREFmTTxfYj9e6nM6dKrW9KcCoibqyymZ
5TpuCRi4bMC7aVl0JLwMg+XL8VrljYHTiN59GA7YEJaYdTcrc0vV1dFbBSntm9zA
NWWvPZeKyp9KrqUIgZP+AMhyejkiswaaYdH3Pi5Pj1MJ/s5DTDrUAaO6i61JXm+E
trMtKOuQdEHb59/m9pnxASUjFukQQJjXhOIaxRKUoUpZpTokMp5po97mES7f2Tao
z+C4CWdt43AMCKDDWWoT8HJ1l2Vm5XAP8rv9bfs98JieccmmBCoBXogPyEPm9sE4
LUKD5VP2zIicWm9VlSjBBMnrMUMq4Q8NRDAvqGFnlbP/bbHmSyr60TdnWNSLIGdR
RZ/RrFcCm3adux3AeKOCTieePlLzz5jAnAcoNXJ1q0QHiIHF4Ys/s4RIv7GB+cwp
7tA8ExMsXK7VlFx6aIanWcsu5Bn4g9Ep1bjpW9KoJ63PqIRuMNKWmHa34a5n0zQq
77uO6dgpPYa9wQygJ/UUKx+kPcgP4wdouVvLzowQBsOBhThLX+mR6rly12eH6OyJ
A23gIphFKas6Xvw0US7UAUcXd1qRM1Hwj1yAnCrg2vGLuoVkNKNm49PyQD5kL1IL
8SHaYIxBJkgwRgLwuPScikbbQmmIRWMu58s7P2GoclDD/6l7XIIGVcmN5kC9aRfu
6SSu7DTH0SJCw/fgOJH//BEhM+T+nl3JdPO6n5obU+h1If9TqgXQQpt+xt2A66Ur
9OiYhwtZxXX2PYn0zMVC278PaZaasOb3YGJHSIwBzMX35T03xjzw1E2cT3cUOnNn
ME8uqEWQCqeKqxBdh9AReUpnVSYSdvkb5mDALpnW+LOJ156X39st4GKODSL/k+v7
60J70dBk8UrDaYcqaiHPySichuO5FGS1xc9pIdTSYYKt2l0dhLqiGIUK3fHB3XfS
gRuAoXL29L7N4JxSehHUrP7qYb5RA5vimn6U3lRF8lb9RUlRNlxCUsvNRu6l9fEc
kFVuofibsLE9iGWSnBf36qz0g6xNou7rvafeMDioXRMggXrAocPfrhxkr/vZGNIV
JL8ji2qUqgjvevCb/6jEOvUdNQzViSgGQ3oPC6jXJ8KjRyw4utfgGLj8m5GpPwmA
v4EgxTfino3HC/ds0VBNz/bpAjF8CUtHAITcux6jUCcXQBh2Xnk2Dc3t3cAGjrRA
fqy18LfQPfIm5Kq0AAEs4Wb+m4mCkbuOgB8Cr29t6mzTfnqxoGSFNM9xzNwtHn5d
l/PGksnBSPvfRCMyoiwiHFPdKh1qYXY+kOyV+B6mNsj1/v2Vnf2+LEkKHLY2mPo9
J1L4hN2tCeGvAsU1LPImCTy23iYzj8ep0QEJImpWw+xI18FimnlYYhP0b6EbrVwn
pxZr6Lk4BVvliHCayjTyCRuYCS7l+PX98QqTM/91jpFs2nHUOZik0+tc4nL2GuQG
E4mXifd7Sotjt4Xoag+SRmoyLrbC66W53AlCVRVN+UHczTKmIqf0hslVXPI4SHke
jmQRBG9zEXnW4PyIsHteNXi5sQ+9b6XEvHCUx2R+97hnxxBgIZGxqkW3vGkVUFPQ
tgOOGXn31dPVxiHHBE8Zuk576VrMICcMgWngpc9xrOkAG8cjkzmo0YQx87ZK1fdn
DOzoW4kPL/V3q+0HJi0lgrDgsVPt1Xs0JuP14uZKlEEMHnkS/Sq7DkBFsX/ELJDv
5Q1osFcbx3MuvhRMu5BP7XD2YOuthAae4o9mfZAYC8+gz0iMrmNlMnYCq/FjZKgZ
QQ6ob9+/NBIFT0DprVddGGkrixx+8MtKile6OlMyDdcU6wP8xWb9Qd92kGFQ3L18
cdEDM+SFJ+bsIF+/uv+K8OfneAI1MxjkJhzHollJxF7N8mH0vrldGM0dfF6no4TS
DroDss8PTgAM6k7atMjYocFLRii9g3AOlCi48a9Y7hiJUfmC++7N+OLYZMD//sxx
3AhZTY75eRMh7zcbKQfqLQymFR2S7yxYHkVVqeQslc8SHwCm/vvq2o+z/f0RVV/f
xuDSXzOcGU9ocs3pMRNsa7uj/kOoE3G/g/GzJinIt1cdFeoLXQ99sJGGJ1rV+xEl
cRG5YD/5beSI79xhBDu3FMWpLiompbC6hUH0KAoAML7dHHCZJr8fhAJZsX/dIaux
1z35S5oYr79MV8mVEsdxz3idZ2f94k1h3lecguSrH2TXvbufXhB+C7jDQ/shHF9t
Ge/27n86GqGIXV/RzI1JbNJe4gK/Mv0EuuoQm2KYTkXtOcSx2Itly6mwUwo6XeYa
xxc+GskzXR4QZ2jidO+rVKOkJxIyh761NZ06P79+No/IBJPSbtESKzfPGfnxzi8c
t8U8vcHy8iU9IUXWprxjCFuRuaZN9FNRNPjC0ywt94F9zLtbfCotx3IfWpdYnpto
ooseXHHiLGvC8o9sSj2pJib92uH5AYCkwp/qr6uMZM9d3JX08YRYZmvXK37dIzIB
Odt6cFT0OnDerBkaJcFJhmYg2syplLZMGvjiUARTcIcWbysMxiZ52P4SEYLmnPwT
bcANAlF3fC4xkHjxaSlSFN2SvUsW22iTilbtnl7qAVk/ES73XanQzH9Ft1vKYsLA
1AlSFll/Dtgf+9qFyDirDHEmxTWCyf+Tan92tes4auaHaDQ3Xnt+ooW6l3Xu2v15
+rBLVIvL24yNEPIbbbk/X4UzD29vn112LT8yEdEmDYqssH/NAt8GxTOFWnvfaJnm
CO5Sob4Cgj8S8/p/d+4dBBMGsSGvcLmhbJ+o+vXFrXrFGF4Did8kAwc3fzOxbnFZ
dJtO2KCi7CBorn+YrOxpoAVZfbagz84aCaT232J/I3EuF8AojEzhySycZ4ZRA6bB
xurFEq27Tt+caOGiPxGTlDAZZTsGERQHFNfh05Y8gh2+D3WmRtsoCVeseFcPOyRR
V2GrEZvcPas3unPalk9RXOzp3Kaz0muVNxkkasKe4dA6uTomMYM85Cdgyf1GzpLJ
Y+1t60WaO4eY/w2ysXsSxCZQylp0Z5oUgcE4cT++cnG5qk3nwDRgV83u0nL9c2k9
Bge8TYrtIKk7jk/PF2gdNoxHfsLyqCd0fDeMQgevkzJsUfyz4eIRkuD1uOF3mh/5
WVtB4MCwF6MFXcnqITf7yg5n/xCEcL9B0kAUvJ2QlUGTEZgty32kSxafByU8TUzk
NgCu6aGpws6zYEYcIwn+NzfEDo8TP1fnfD4VxGoXnO3P8T8ZR0Wr4euw6fPkeQIh
6dsfae+oSl0K+0zuM/vaQcSC15evh9DthZeKTHgafJnUgmKF+nbJFOfN3BR/C8l7
yqCj1dL5uOaeQVgHeE80L4cMYW6ayPGHa6Pc/1hsLzyHFkiD43XKsl86LGQzR5Tl
athvKKW33wQJh7fk3bMwb5u41r8wgiATYnajX4a00FFHKF8KcuydlKTFvj/P+1Y3
wDkGx2DtEIXuPWSHDVVljwqSrdy1syA9yrThIPJPo7U4Bmujyv1/694t7MF4i6RE
Na2l8XROnh4uPz8PlWWO1Aehl1cQOT90PU0i2s1YM10fiat4Q5sPK66AJhMRGmgd
luCtoimdrbKMD4RWeR5irWUjgG9q+xhtoKJBKphVZQh5KvsYGl69DBpRenFk1A8S
uo1p6k6faQk5RQzJmu2UyRP3/4QYXJqe/Ph2dp/WdF5eZfllw7TUYa9HbKXlG3W7
54Maq8LnDhqRHCuHrWPfPdBn4Ltq1FLyhmvWBcdm29DrvoJ21+LGJrOqLEfq0iJH
7OgeuOZZLFppIWvNF+NO1Qr9299zJwzD2Kv5mCaRzgoDNUJLOwfvAPVP+BQGNA9l
GWzHuAoPDQBj6BuNyeoS9xYMolipb7l16NzTm3m6i6Z/DeBQ8m7Qufmy9u2w9tsv
bLM9h3ZwOL9Xajpf52k/WZ7W5a6eLTHHjvPB73jLCkEa1zitbEAZUZLfdkL7Vzmq
kc/xw7dRtJyQlAbviCj3elr/D4nvhyW7jP79S4P4vrtWEXDDBfd1YqeCOJlRrzmz
MZQwWnkCmIJHHTdMIznx9kAq1wrtybioARb9CSPjz5G4fc28Fc/NGuVZFeRprU2E
xRXgOnO5+DB/wX7SAPeFzrNs4ZojRS6AWSWtYnjofem2SH4YIR8tFd2IrLC3GqAU
Gqx14j/2V9TchpPI6i9dlww/PdOFqENy3GPTSDa2GeZ1dg58LkOysvPTqhLCYPnJ
6CjD8B5Jk1X2ldYJOk+NmP01ygEuQ0/pyTNSgiCAza8aUQW9D9cbwbvcmX63d60s
R6y6TzOEnhJ8IjqWaGSGuj+QwvLv9LN2Q/mKe0Pt9qj0CTfdbD257t1zAqHuHm+V
x51et7WDWH9PmnUeExHV/dLp8YFsgPjjh5/Pcv79qCkxdVqt3FfFg0btZ93T+DD0
uhaLheyWsrcqpJnWomE+owGXNkF9BtP9jjH/8da3GKBeF5YmDoDkGqKMH0OJdjl1
l5Wrue99pU3CYd0EMZ/JEnkLqtra/yo/mERAXivJnyHAetnfKKe6dSjSmptrXiQa
icRrpiW7Ce5vGqIV7Uh8C4CSpnfarmt4W1og1QCzkbgngo/YNx0YjzPT5OXOfbp1
texTnXnxtqHc5NLbtEX3wU+G8hIwXfwhMY8K/TcnaN5GQV3uhg33XOJ5qciCU4B4
Wr787b85cpfBdSCptzIDPjM4P4okyhbZwHh8598kxyVkDZTsxfY6GVsx5MqvpLGA
sezoCe20zs2rpbZ+1HZ/dhVJxTE1X6o9G6zlxurDY4hPEPPwrvfF/4/+ZLm3JWnk
GGrXcq1itb1CENlO5pHgeLm9GzAjAOSrYNzxvzAlYF8+yvAetmqA4wbLKR1dVqT3
g/GONOx6Mln+0oHiBTrm7MBv5CBGRn6qxnhbszobzM9hcgfdziQRKtcVfMy/BRcF
GNeqiIE8KhNemZly6K3GRuW0tDnOy7Ix9wumxpDC+PtCpz+g7czSElPsdxjIDpGt
oJQOkUDcFYrqQmah/mU0ASCzHLEtJpcc8KeQvAQmmEnjMvMWwtgGDiJtcYnXmxtJ
DVFxTlmHmGDXee2Z0Bk1OzkD++CRRkoLCG3OO+UWgpSk7mRgyNmF/1az1jrqjuyx
wvW98quVJ+xcOJLdyY/EB/A05fPo9LVmqbVHeP/Koz9OAU4Sx1+Nmp3ESsHlBQ72
uP5bmWEPqHXYC7UzeATPxt/GLwr/KPFThYsOSoPA4rurV4UTrVu/5q+yHhmaLY+4
r64lNAbiUW7YfkiQo3q5nHu3KoIWeK8/0uCw3lwty+0+GRt99wxKFcJMDJjIBg8v
ZTVzpQ9pMikTvq+owtTwjLGyNIT2HDi+skLtTkhiU0CJ5QELVLglyz40dfE1/mwP
Xhi0jcIQB5NMqRCXhzQ5wTwxJZqDy35rmUJeFwCTPl++z8QPij3cp0J9wVhUI0Ae
XcBcIlfYv1FZoDyrxtq/Qy8TBCkVKwSI+c4gpUVM0ZHWmJtWr+U0tiRxnXhPv/uu
KJnSHBN5InzYuOElUpfmFKxSALL/nhPeNo4Lx27HgcJizeM032Lp86B/Fp1EJRDD
5Vk+VfQ/X4dcDy/PwIg6a18LG9+/B+dz/mHFZbVo9LSnaCaaC34H5QJqT5DVBcM6
xQ1chxV5QMl0V7Vb7wcbhgkNTqejacq15eLsGumKwukcAzkl1+8f2iHa/SgK8DrJ
iO1XrgqrQJg8kcBa4TQVJHDTQglZLkfx1uYbMHzHzkB2gCQgZm4J6jICVB+3m2eq
k7T4euNnxh/gB9HqfuNgTrp7GyEteQ6vhYW7JnA7XKXNBnXAH/MlTw4r0BTelHtK
rufHxW400NGyQLJ1l5W8fHF8rq7wZd7cGt35ds5tKNgpbLIqnw2vzTrpuHvjBiEj
mgSpmuryBSfteNydC9oHJyyI73zyW8AU2RyeHFitMcVkSAB+kMWAnn+DxWOn8ulF
5gjVxxuRIE0Tj22jvr//tQrHM4oqlV9Zuiw8R+QYkIfOGgdteplJN7NNDO5QpnTz
a/yITlU0d5K3VFZYl/vUyNow+c073y0kC3pMyqs1mKqPXfMJ/+2jY3NxFpK9ege2
xZKh+oTJO2qpft/io+1HYlIeZOG8SpORNquMh7/e15CrJxygCHEFMhED3+/n/mFJ
hsQV8kEF1YBZj+hoYpEJjPMwilYJ6iOS92L7mk9j34l6U8RPXgcgKd6eOSsSglbB
ZoH0LAOHexm4dpXaIemeUTR+Y2yZMcDEN5yXK//X3XRycXqmw8RTNu1LMgWic3b6
BvPCFDFuPII6ZvL6Brl78Rk/iSlW4hmbFwoz41fMAz4c9pFWfZesU08sJq4urit0
z/XLOi49uDe0Ch5IcVgBEOZDYroFMOgeQbN6HeVMrN3fDxKkF7vA55LDy3eWIGWD
N0Zxrt0gRXehi3tgUma0ycTqtMKhEAjUXYdw2D2mc6ZCTs4dfBeXO3EjKcxsyHlM
dTP1JIcPPn6UdhmrfVybCaaC7Ewr659PBLkdDNQYizSw2n8mnkX38+6W4nrp+Md7
tjbk13EiR8xCBS/S3r9LcumlhnW+OzueHJ9U903FCeN2BgTG3SQgAvD8nJ28js8B
ViFueCharHvWKQpBLsJ1oWzQQWyjnCKW3N2Dr/xqd/jyXYuYeWn4a3yDJzN7J5De
FU/q3wpM/+UG9nxJDcm9RcMerguSKstsWngSikaBP51a83hBb/V8AvIxzRe2GKIL
0L3JaD7mVDvrsBbOUzLceT0EWTmatRbJxfQhul6GOOXfRlUgZkeSOr9SKXxVaEJL
ahq2Uc2WUhkGjwrbz9Izax8d7sSOXa8sqkhA3XXIx1qUsZehnQzNylDYPl8APIv0
GiMEEYXOh+LyYctdk01nJsfdOpMJ8bbCQmVoBKDK0TW9lqM4qDDAkjUcF5K500q4
twr8sJ0bT1OqxX34i2pGJTuE8k97X0PvM2eQKJ6sIJ19PY6Cltei0jcShXzm0YAt
ZsVncXVmzXAGNrLFCflqbH1YLcZxmvcyr4MwzkyEUfgWcsbh2rq/cszBV6vYa05j
B6AYQv49OkLZG6isZFRJdelKz87WjEHfY6hd1chw/d+vdFgAcZyqGTo/cJuzTQNt
xN4JRBu6rVUGIdk9zx7ToLNu3CFvPqrb5+Scsj+jKEGISeK+Y3ZfV/5QO/JqkZP6
qelNEZO4mXWkzXtDWNpBCYONcq0nvCDQl9YOE9BqJF9lqBcqK1RPm5zMB2li3cTX
XHirnxUTjBbA2k53C+Tq/C5THzjnhZUxE25CCXZj7zqGSgjFglUw7wDQc/irBUd5
sKA0QN9/ufIMVe+ACrrdfWqgmbIab5t8/T/VUpNYsKgoF3/8fZNgCBsVqUFTghQ2
N/do7OojjKQ4738iROltkZUf0/Rlix2lVila64PtMxQaaDTPpMb3wSDpdw/AV5WL
ack4YkGQ9iuO2QQwVQRbuSD+OfR/fMjZoe8SKZvRsGCIQHhs0Ict/BbF83nZi/Zg
Ns+Kor8saTRRmc7k3phkWCmY7l3YQ95jQ4Cr2Ecoon95rdIAvA5SGjAvwhqT/GzY
vvF8PdkpBw65aqoXCCVmdkwiNkoaaBgmpEmsJ2l1vGCdNNoISoEyiJFhuibLzP/p
Grb5KbmBEc72aL9d61/+z2QqQCOzUvee+yMkLPHtnuzJyeJ1lwr2ASZ1yvBLdimY
lw4mTRhHgEFRtZ7+hksp/ncltmrEZWICjy5ZTlefvCQjjHPoolkGdIz8vFviSbkw
vMXTZNi+F8FZdwb7R4OwfIh9lly54DAry671ScewCfrT3YYVuvx+YtRQpMhEtKZH
zQSY4b/AlHT7zD9XkB1vtZKQBaET/LRDLqT1TBXbYuqcLxhMXvj7dho7CR8WfKuZ
EtYUICm4vSyKwbevBmPQVoLE2gbCXlTt2FCe48uqGco4evNc1TZT065+6+18KvCZ
mV00DUeNvUi/xXLq8fRunzPma4Y9xLkRx6eeP0W8rI/ecc4SYUGpEag4Mo1zUpB3
RDAOjrmPqfkl4oicN2ycJ0FXtzoBPekQLtvaqQoU0DpSvIo4SkDnZTHiLL/8B4aE
VqTuuMkf6rU70jnRhcfjNMqp5xoqX1AnqghZPuaumewkzxN5VAohnLpTXthXKSlS
cFhN3vaLDTZXc65iUcHwgilIkvKvA32683He9LmIbEhxg41u3aUx56OobWdPyhru
r5qztWaUQpgJQzk2DughUCCBqKMOUKViuJ0hsZMDwvndsj69X2QgKSfLt86PYv4r
QAS5T8lsYYJUqVod7UdCbgbIVtZPKcyWNZtQofC61atO5Wh8Pp7iYM6V1Xtcs9B+
lTG5BOpspWN42pivEEKGpZfy1allzUI2rMsAa6QwWpqg1ih/dfv2u4Y1IYno+kM6
eaEGU62DNUhnFKLxFJh/RZjmbrmsiDSw7hP3BIZClMmVgGiriDwDiORTPxFYGX7x
VCetvyjE3UZlzmr9ihnmETBy40jxjkEPOI7fMQUBU0yWfYNnpcljwveEGp1aicpx
zFFWe5VLVEd7CYqlLHG1uwD1aDLAKJj4orOfAjZbK9sAKth96fOLON8Ok37v8/IW
bWFrfQmsuSRySRkq6gVA0i8Oi7P3B3HGonP2i75jApyLwz+JCYW6NSBALPUsu0uK
0u7Zv3cFcDUYgVDAyHjxPfZqFYP4lTi8FRo4PBRdMCO1UWBsl6w8/TZHwBv2c+j5
vOF38l1jtCBSukEyG5/pW2w1Utc5+9Ds0a3tAyGZco/xxTbqsChx9e3+b1ZUC3Mk
Bs+JkGryijL9gFfd4zsPSgtD06cSxa586TQ8JH8oRKjp86hXasw/qDmTY+3S+uSz
VV+rH5dypee3Emw9SU1x6Kdptoc5B3oEXjLu+23IftuI4+S83F5UQRcuwAqpttvK
ZfvAkWOEtXvuEuLBqmBq6vCF31FzSBWgJDW4Ojm7sLmtX7W0sxRKRc2NZyHY791K
8ruGbvJ0/SaCb8GE0EK+I022hjqrfA+vU0V4RllYJ7cQycFxpQUltvZ6djCQ4M9F
3P/0u20sx6i49JEwASyvRxTG5ZM54iQJ6RI6dK4B3UER9/pA+Otq0Er8tBFMgPAY
yOX6VgPFiMU329D0bkbJGjD+mXjO7z51ftp9L3OsIPWbEALpuxqpQDYGIobND6Nt
qOBPvwjhO9Q7lAiQQ6VOqhzcKatK83C4WltuxgXzc6HK2pcq4CrxjDWTHn51H/kS
E6dUaulIY6Z5Vl2fD3m9Zvo/JWryca7CnLGpKQRLOinnpi1fasXbtf4yaGYz1/TI
pxdYTAPfa0TrN6w198XWWs/OXn95rswYDtkYLPdY4Ijr3XCyCMeGue2V8iuZRD78
b6AAU+ey9yFXBPJg6huHoGgF/QkXqNovoMxur0bSzZWPjglOpFx6wUO8fDutRc83
+fspvgMQgOHAK1JAhck1/G4pVHCMTd4+IbeiTeD694SAQloo4htB4qS6S5BHkH4R
5iByVMhx+n//BHTCx9EnNM7qpP6IVphqvDb8qJYlKDpPPsjha8Mo4Ms80sJvNgR6
OemxZqqYC1Pr8Pn0fnabxYsKqxqXhUyuK9pP7XS/PmnIgjRJ0/aga/rTjkg9V+vx
gVHwhbXwtwd02njHGMPEBRSe0bDakq1KkTcJUx9/s7Z70+Cnz8rCWmaPgVJd69MV
kKnP3ssHLIXSfZDg/NpmMkLGO++8n2ZHF9Tkmguln5EkYSZmxck0+FZNm9EtPMSs
FA03DFhPVQux8VSd9X6KhI0s+2TacPPZEuHNgrY85e8AgYNtxio0cWPscLASj54f
FUJELP8vyH3X/ogtDGvpKUbH/R9tiZutIYUJlBFGpOb9z1sQG1H4stpzQ61ur/Tj
UILRMcn8bYONusRXvBWsUvi2ipJ+8rxmX7UA5MldfSBVBjEOR2I46CbB5IloY6JZ
cyoDnqWU3FwOkInL4Fn8pRZcGc6A3e0vboMmzHx/I2v4PnO5G70R/ojwPvdRryHZ
k92ucwXuvvXCP8zgenRciSMG/+6RfHFiT717NfBHjKVQ8Uc+vPgQiM5XWImnPGhS
A8iu+7Tpe6HbpIB0VIbBpB88Z9VVJ7L4ydlzNp79b6Kpi8+pajOdPXkL+wkzU8Za
2u4CkQ4bkmI65gcWHXAorJLngCq03nfcb0Na0D+mbY1DXuYSWGM6G1PgSkawqSRO
zW+kYbS82gxL2vw0hOrWReMcgZOPdHoBUWU1rakUuLJMltEl+RFWmKmQ85+sSH73
cRKfKaAV5l9syNRRsVM3Uatohs7ah/z4fdL2J1bCJd9eP0owlCIkP6MYXEYwkUdH
xTcTcPKRN0LlmRu8ICZyWVdsM7cCj8uzj/ffYitodO/piWqFeGZb7ngASxd5ITv6
fO13FJwKVHxtwnw1iQqaPKFr2izPQJ7I0k58Z/v5NASeHZDRf2WkKvwGmQMjvlkK
kA3rEv1BD4cUJ9MPyyX273xcU+gXKNOBLyo/A8v/MibOHcfgrfvK+9/xoAVzSx/m
ANqF/3NvTRqpm0jcGbYvowd1RkZ+xsFMye9RTmthT64yR8ToJkTYRZDq5G7iu24y
e6Typ46CyDlpM9KOF7Htw/HsS3BOER5AEelhKKqzbeKh0mkDkQ8DCum6WLiuPLHg
8fjc17JHanm9XzeUWJdyJNGa/liJ4NfJ17uarTA4NwQWzo00DIqUJX6buiI8XZHZ
Gdn1Q7j82LdnvGcm3tagfLz5/IhfC3h2XSE8Y00jXWTLlElHWND0aLHTO2A1z2af
qpYo3hOK4dm+CULYSyhBYRJMPWD+n8dJrx9ib86bxBlWQl1cA8TEPpOFpquNSt2O
nZOpRa1at9hUeFQwltyUm8RbToYVgMcwUSbP8dEAQH8yWQ0F5URAup334paOz+Es
QemuvMbA7Q6OzayDp1FcTiG3wUBVRkGzsme55eV7cxhAZMrXfj5wR/1Wq7jNCGom
gb8KS1KEp40GhtbG3vrplTWytPfBITPapAp2S2f21il0PUpN001mQcYJMiBAr0y+
fvTmXcz36fG1XlAmAAfQmPYXAFz171R7z9jGEyBqfgx5T/Nn74MX4rSbBgatT40I
vktsdAp27DotQYGH9oeIAECRWLPMEQ/uy9ETKT8OYjFEiNpsejY4vppWAC2W7Zq7
PQXlLesvjtSupQeWpXiTjWb1glyHS3cwxXIndm9BY9GbZ0MkBUSvOX29inez2Q8c
Zq4tg3Irwo+n6un+63E8cHBiy82gLVDjaH4cxXeaFDHG/aAXN4roTqbvcJvILZVx
szRGYAP657x5Qt+oTpHJCrOsC24tej24Kqo70lHXtS4aJqo5J9tWJ6CwPFruGIts
4WCTxuI/0DJSVjr+V9siOX5Vl4arErU6I0SQ+YkZDtxq+9yLVzkniqQLPdjX61Sy
8wZN8BGyZ7D1oPzSnq9txa3bpgQYgNTddNNDIiPwK18KGipS1bQkx5qTY9lBa0Cz
hMrE8RpbXY0ZwZjilcfyFrm5mB/8AKH+yQRxR1jVL7l2Pwd0JAYMHP6GvBmnZmDl
0RYpaCQGrIqon4DXh0hAaCArQGnEYUQt0gNdU7VSUNhMt78trqVjAHHXiZCPNiia
WZ3V42llJa118NGYTcJ8jeE+Vf8Pl/GcVl6maHBZ4BxtGKQwKdy8GBiULR2UqEYp
wFacELUDTlbgz7GZWFiAQMntPPk5ts3QOwneSJfm1AHpswEM9lBz4Sf4z1YOSpEn
FllqSgze2NjXX49m8TuPD/xrjw1Y05p8RDIkUb7uMUHX+r5aVAKg0f+dErGDnENO
613yL6mUqwi/COxCJhX/C0N54VR6mQtet0Rah0oErKnMtoJodvsZzEy70H/sxseA
wscWVa4nfq1DztGB39G3Pq0Yos6i8g5jhpip1rXr8X7kTje+8uJsk1OM38Jux+2x
frU4MHuvxNN6FQrTE8qTUXZxUi4RW7c4tZ1/5gLk6Ej5+kPM35WXQ70ZS49RjphF
8JDCorPea3JJaJex7OHTY9xRdkjYFfo9ufZ/vCSxozBpZBZcHKWwmKLtarCa2WQN
yejQZLaM/sJBssOlYGktl/IyN3T8XQqztXziJI1VRmsDpEdgZkupbjotkadeRZKU
mKjsclj8OzkqZVUCrrhOfO7rAcgm42XseNT8Ee/H90btZ6HM4KnP2nJnevHeHJZy
em/GSWgSTkglaWRWR/FPAf1RFU/41LIp+aN2Vg2Hjwl39aQZ4aUOAfX/cftgM1kx
QS2lI1+W8WDqdF+z3g59runBP5mEKc/9/Nbldugxa6o0bqWQADrMutBnCFDMJ+JR
Fe7O8KjPbFbOiIkeKS01FItPWd3Vrqnp9+Hr7Q/lUuvES6CaKe8IvvpYRhenrH/p
TabSD7aqcMQutW0LVZCi//1KDReFSn3d3BlCRauTQp65a1AaghAs7U1+s0Z+SwaP
uq0IFgvCLPXQ0jdkOXX18sDAt0CU297+FG5jIbqqLYzBaWe9PPORY9krxtnMLtg/
1G3mqUyjJsmVp5FhhMtDmh3jIaaGVXyNFmH9+J/xlWU/yvK51rhpn0ERCS+hR5NI
cBThnVzU9qO8F8Tc0rzC0/ijVBsP1l54SFrRUMFe2UAb08G97U0aGuYIqWHkM8ik
dpxB6xj+SFRIikWcVesN0nMraDifhwnbbtm+TRlXRRg/o4VGrLjaLO7cyMjtGHSr
WWTUqVYpRVvCX39Zw+7zgHFkO9AtGJBvrolFH4Sx0gbFOtHWBoJ4nMjHXkac9Uxo
sptLzQVuJ+Fv4ivxiKsbPEsB2WXfskV4Mq/AovwEfoxS9tTb4rqHvJU6HNkFYG6l
B6Uh/jWN9EtTKBKkWgGQdrswUlduULhwQmTlreY9DIuaOKILfoxbDTxJkQEcvqai
l89A3KliBE5JyujxueAGsnUmfnO3fHmrhUbJas0krzc95F7dbkUg5FydxY9+oTq7
dHhOhffM3jFnzLSG0lJgSmietaGbe5EXvGgt/MPuSIsWrJ6tM91NWW3vnFNWlptd
ehq04o/faUqPT6+9rNwXtOze4Me/y0sPDUHamNjtx3lmmXLZVOksfIAiqVwMeWfl
tY/Bb87Oc6dWcNUP8nxolfyydd+fRfY4EyRJiTbeW75kiZ8AT5LwCnpC64+9yLhI
LmNYO7Qg2bJsMgtXaNXXOquwISTYgckEaCJZxbTB2ywjYSKp98Wj+zvlqug8GbdO
A0GgfXfr/3KHqjPyk7yLGTurjvdShWI1yOboV6/VwDe+gG3yi6vLIf+As6f4UF7R
Qg0JXPJETrcXqhRNPtQ/NbNEkdNd7xAmJs7IUdNfWZyKl2HTXecJdzEVOoVfeasY
6CopHkuLYvSUB6pIg1RS4iql7ygOkFp8mxei/mULStwppHq9x7/md9tsOiTWhaxG
cztwWlpixoAKyiWCA0R5tMxhIm1rOTk+6Ldnh0mswL+FGVno7vg4FPG50OYTKWDj
GI51p2Rcou7FJtyprEdvLm6hT2ZkczIbZI2yReOrMLqJNvCNpeBlTI8CDcQzVBCr
cgrH3cdlc0vbkNuI35bU2wr4DBTKaj3aEIdZEryEZmJRdwb4SW8PZJlt5K8OpD5w
Wc9v3DhyWkhAECk+i18gfleG5YavsYrPZ7KgKpnptiw5tFDQvIdWWWLnjyxN7Z01
l1AZprX5R+6gHxuekkLpyohvleUGEDzg4ITzFXM2iF7gnYvhJ7915n+oELc6KL+a
L2PoQEhYCVgPT7+BEQpjnep5v3g4w+ZFlPGIc8u89sgBy2d2KIAbiKy+JHkvoMYm
pWE6R27W29tytRZdNsu7fkQInCjchUw30DPL/zlUNLAldSkz6cOxdu90EKDNUycM
HwzfzRczk3VjksMq4w5vvqL3yGw9b+FhQJyQoUxWTyxaPWHo50dDKxEWi4DIuE9U
ZJkHHc3ZeBxtfw+Ud+TYSt0IZli31G7yPv0PzLNrZADdZKEFe5ENToFUjLZnfY3b
XxXFgMOxfMhzLOO93ekfEjvHvlzeQluf5U2fEMd2tE+BKoOhLfTvEkzBreWGPeiy
/cWTJ1fwH1hZS80IIJ+arhHgWIKozNMKMelyMBFSdKH7UySSbJGZs64qRUoSHU4V
x8KhtaXNPCuiV2Kd8i8h4UiivI1J9V/O2IjUJ7uje/fQ1c/WSh4UesZ4r/CkhsMP
wzFQn98m6qCMmxfwMls+8yy9WqBm6T7gTZ7gFlfx6t7nuIi5nAxufFOrjCp84yFx
vZk1rjeCZMZBWvmAtRFpIiArCNjLetch85Rm9y1nEPqrJQd471GTDI1dHGa5klj4
GqW4Dk+B/teV9SNDkxOF/c/72O81AoTA9IKTWlNMdR8AiGrQzFoy5cjF4Xl5YOXW
8RbzGZ7qfK0uE6MfUqi24c7Sj2aKr1Vk3NdxvUnfkVZzdKCuFwsg6WNMLzckokpi
cViZS9eUyZm7W3OWYq7gdA54hlmiCtFHvIsHT2aIiUI8yfMX70lkev+cKNf/8Ct8
ibmNWgV/8/o6p1L++uRWw7Djr3qK7Mas0Lj1f5dQ8qbnX+gko9tqEEr7MbV1enQ0
AhOrJpeVl3KC0BbexyvFTBC6Z3pvYMuxeRlpeAh3/HWi9jP5QpP/sQ4JP9HpVTzV
ixRKvtF0pWm/+TvROMT367JpRTg8tB4Vh99bYBVkNLi1kmiXZ+CoGugqOoMIe9tN
TsXKikCVnD6FKeNsZ5UtI2DBeD6bZro4MKCjvJJ11SLSNsXozClS4RKAw8aHnNI2
i7DYpR6P5j375E60ZsMsd7qFWNDj9M7jxhflWkCWGQnkF77wo9Uom0a0pB065E+J
NxOiXZYquUeCrqu+Dlx3NSg31PiRJFgSQY8MhYuq7lkT3TGCrHjtzQ7qZA/xlW/U
pSqMwr/p31+pv+CM+lgpaUa7rCmmjZBLR+4LXdEHxIsa1qHiFTrbzNNwjSBWobx9
e7TeT17ftiuk0YrxcQ+ySYvwY2LBCl2oiIcufh0QGENiaPQKNZIayXHQyUqfKCq/
ScOUqF73C8Lp/YYD5+dF7RzJoluy35tRdd0ikCKWnWZ3MnriUAuuwf3c/NJ52y9h
gKFHnQwyqOk0tJOLLV+9P5/oMXrNZht6XMy5bCEFQZ6Lae+ajerMd80RSXFdKmdX
Y33hYs1tBkYbXlatUlLQDNMh2em9wFn/vfx6dLB7f5J734WBK0IlR1OzngypxA6u
9pB/CGtNxrvyHBLjwqBX7VIoj63gP5jO3KiZxU8JKrQeHHkG1dg7C6BGI2J2Id4G
ZrJ9Uqhvn/Zler3AUsIHzRIxsKFFsft9T6lxqwnP8mkeJNhFtd08JAJId3a2qQ3e
fyyfcSDAGCz6S99WaxiLD49LTKfbrNMBf6Ly8bQT05IhkobgNxWHQtBxn877wKLr
T0mubZ/A+xkDyD1AD11XEteiQK/yhjCIBQ0F3uIvZa5BA/8CQoQjFJjTbBzpLyKp
rz5A5wNh2u5/b0IkrB34ZBScHBB15ZMWlhfFe5bJDUOU1KJv46AB0d/JNUTc+v/W
Uqobb+8Qr9J1odRwgUjowD28NSyoj/vfUzkYlLskinN87R5KoKB1k+VU0NKB8wE2
eyDRWXbbfZjZdA5Em2xDHdC/2GPWGcRl0r9T0CLJsThWQaaFFhiWBM6ZcVZl9Kz/
3PAm1gHPhTdiSL+rKnTfcKjVgf4lWCQpSdum1AVVNLXjR+GZDXguH76uY0OHhXGS
dena589Vo5/MXh5Wnim1BntJNSJfE/Q1kRROL5McbRse1S4A12JLOi7pgMGU+BrN
z33KQLYZ6hpyaUnqiF+lHyAPz1M0K4YQ6qMAljKuBzwY48+AHWeginoS1B4a4N73
OwrrAuy6ycIp6HbZZFV2IqVrhZvb65kgOCWLZK0xuABbZFAlES7VyM9LgPRMZI0f
n22Up86dSBi76L19e9UUfcdYPD5TQv6rwmbp+SRd25UrOX0yb5iz+oVpK4rPfBOj
Y9VdfzsGmqw7uUKFmfydciDwfe8cSG83na3yik5jeud8LhNZnuhJwtIhOUtj/uCJ
i413ss0q83aGYddJCySGCWg3LUHe+I0igy+khX8+3goBFTKZw5ldf1lvzuiGY/6c
WCWF8ga6zHOApLWZWyaEPh9PNw6tQgn9xiLh6NYRb4vCu4+v2222ERlat0p1eZ4t
Ey+9Ue6nf7KIoU4Vqr4URSIlys3C/3NQk+qBBr3Q9367zLTdVCPSv/ohbvqiebdC
aXVBrrWPSD0RxHXVTwJvRqDrCDkif8WQFMshCP+7/ptU2rwpq5QZYEaA/BWQUzkl
Fm2f81Ey3AIb8amS2nVfJimj/KKlNPWWGKwKU4jFAxvAmlDyDNDm0QR9LurMPF5x
gmllxQOysdmVShxsbs27HNLTXz+EqEL0jhQUY0FXw0+z7eRTtcdgcuFu2gELGpWz
iKjPS6PC/iwhpFmAvcADW4mu/vl62O+ed5jMbcHfDgCgkIt13RoM5k7Es9DvMziQ
5cDKlFSq6HHe2kaVkzkBV60sivJ1Rr09+TZ2vKOMV/Hdiqhpzh001zTNQqXcR/vi
wz2mS+uoJeuhe8y5BDBjGLZ/zcwC6Noh+9g5PtjRQy2jEzIMha5ctPvVuI+a41tM
IQRfqVzQ+vZ3em3RQjpVlX1XUoXRlLbDqNjkgrfu29VVRQpAZl31t3H/MF8HX73X
h8AlPg3RcuUagOpfDTBiVm5TuGRiEnHmMldcd92gMMmP8ZdxmxGfwPP1LxYsQjuJ
K4nZ+HTu2SrXBSU5fookT/WWAJI8Iiy2ofpHaEY7+wNM256zUHnYmRWVpdKoiGk1
1Kf4gixbAxTOrbgluduNL7IxnG1l2tKxzCr9ASi5co3WhkA40/3GBB46I3pGv476
i8Ig20gdF42Bj59HVFZvHXGpyCOs2ztuz/6dNYt9iHjEFD+Z6o6Ly8zJdyo7Wr3Z
P5APxbYK1NIuxg0DzO4HnhaHpSx77N5illJFSvKZK9wuxin2QGtO31+DICu05Bfc
bnw2rSxWMdPuO0g275fRfqYixVytfC7aPlBI7e8BZ9gqFTO97zzSI9xI0uLPqAa4
PeDI0b7Wy9CBU+G3d1506gmrUM5Jm8C6qiVUZlAdQ8Dw1BXIi0j6VXLGPGKnRDkm
xfn53p68afS8Pepvu8JQXtArnJqI5sg9g63zucQfdlmO/e21Tj8Qkm0/FN01qjo7
Tw/F2Ln30U1rWgXdLVIBGZtsYyJa2jJ+wf/qjNV4D1brjkRTrQEaNCYw0PbnljR+
U4NlqU5G5tYt9XdIgMxiGQQVnM9O+Wvqb8afDCXV3cTvLP9+n/eHsiECdBfH8dBy
nOQljQXq86ZTjrS5WBz+pzigSM2M33JcSwi5+1K7qZk9XREfafpVkrk2VMPfSpm5
zKCcStJr+NGtq9M7pix+8cmVgslCyfqnjmXbPvpHzf5TY6MwOWLz4J66hDveFrYR
5D8MmeiYtzeur+At1LE9S65lPPkRVrXteGAl2PiMFr/4GoL8Eh7Ouru6h7hVH7Yk
KGT3u/2T4FJWhNnBqHk5qvUYL37qLTe02ORvSj2VeETzkGSDPd0kkDCSpaL3NU8R
0s86eoxDOna47mBlpvXd8UWzQggJnzV42Wd8E4Hy8VXJEEhNSpnXbwkCws4z160p
jsR3fUXduXNRY4RlEBWmWm16OJxniv1BPP2zYJykbqaPlTc9n/r5fPebMTAKrZKn
g9dtp9cMBG7WtQy/TD8Q4PjELWQ7RWNAtPLnyzLEvrUJSS118euGUs+VQZZMkUsB
/uRPanhK0HEf9+5T4DBgc62D+LL/XRMZ6IC9IgcxGFQh9aQa+Bnh+b47vs1pWXTT
WXRuTITNYRkJAcFb/kXiDThS2yl4FOMVDMukuks6qc7nkg5bgyihB8jAT7568Dl7
OSmBJT7LI1Z7mWJ+o4K1CNaQNPn4y5JDWCmzWRHIctSCXaoHyyXFLHGnCQOhVmVX
0PnOvaHLJyGw/Xu6J9wn80mK735WAtEbRi96ynzllsd8wKNDKD/PAqKPfkbvgvIr
bOsSIVVCcb4YA/td4bPk0KcCz2bUeaDvT3pV7oFy/fiTk3mXcbQUy1ZggrW+1OmW
tzM4bOkR65ebTzaKEHtu7PBHtDWVZM9+1mZl4Ss59k8geEq75cB9cKKIVIzeYkWN
FVTMl1r0fI7l2j+HZMv/adUmEJXl8hxBM0CGOxxzk6skZyfdLpc6GRWTb7LrboVL
M4jvxMcxiupIw8aYPH7cbechvT6ip26yxaYQcFFLjWmCBRN7d8HhPYb9MzJOeRfz
/3TGDjzZg+CLEWnl1H2y1AN0gGRhCRzHEAgGDDFF2TjbupGYqDvquI5CNEbiPLZy
KHw19KCjV+qogkgAfN/mFIr7XNqFq0KiJHZ/TPDJZV5HNr1pr7geXOJ1hYHW2Y8f
THh7+lqA9aTgwuYkSrH2+1DPoPNE9nY+H8v9Pu9wWMg25NJqGc95Nd5N3JkEVHiq
MW9Nup3l8LGUhYBBttIF9Q1FKIfN+Yx59mhlTaG87ODXSjfgOEfzZrEhWptsv0LP
H4BqtoGLfZYv4AmWfecYPPw9D0J3LF0I56oqeanFlpf22K9rbAw6wltyY2xs6Ogq
w0G9i7fINVHXg+qbGhBBkBVScXnPVB+t+50/4z/AknNl3NdBFKzasCW6kR8TYooX
/wOA81+QXtwHFRuIdNGVmqYKOo5Qd/eqw3mfjpVaj2HahcMRV2k4PHC3+SVFu64J
lRqD2KB3qsdXtAhe6gHUckyBWBntJHFRsIQKVs6ucGINRfU96Khx4BdyMima7/TY
g3NnHgM+FwGDRxI3ps5ng1f8xghy7khmig1v9z1OMIUZZHA0qYCneMG9GVUYaWkd
SIEROx0/cjbfh3+/Gx/y8mPFP3Us0X/wRfu9mracKhofoc6SokyjaJVPCwnMcjnZ
Y4CYVjeu5/aBaY4I1znbEISgByW0oMnozwrFisjuPzbSi/UQ+ICpmBxoBQZFo8n5
t0IuHf6CJqcNPyPfe5i0Yq+0qliC90ato4eggeg07rOPcosc7EQ4P41SXwA9IS5z
3MWApgeavLn0rHKukmYBtfrghkfnMieDKXpl2dzPl08+XomS6LTVD3IsJs0vX6Pz
KwAPGNRDR7VayXbQw1Q/AGXD7qFGDsmxKuP2X2lxknMAdCMWcx58GmnzA7RL5MDc
TPFHmL9PsUciTFF8GVAi7LHAN1bn4rZlKcOgx1onf1VyyE3eAnvoeufdSKkQCPab
9f9Q+qxTexvb5fAPSAKZVeA5rGtUozjJssMlhq83NFqAKKJ4gdFtmoQ6vTwGTXwc
hiv/QG/8viHpzEGCg8Gtr8DTTc+n2KJl56ZMAlZYTUQZJEB3Jxvqat68+cimhnvd
0nAuArsHF7nBzlsfdln48v4vdgsA+wu0jXQpAh0k3FNgzV1aM3a6ZoPp1dQxVcnj
7eRozBZxDdRgVkwr6W+v3lMCnovjIJEEhtbfnodzPckwnDppJ3hYMoX0a7lRHJbH
VetwZ5PP3HefKLB5lJTZgWQqfBSZ2cvoct/R2XJT4dNeEVOsOODth+hbdqQ2NKxd
V/41FoXusk/8uQVzgolaVtzp0yBinZ7to0Mo4539M7A+vTjCxksDn3sh6SniGTXS
NUV6Gz4SSUFbDmKW3McSaZ4Lz83vr62DE2PqsU5cqzl33iRFv1F6FWJdlFoKdNmz
7guHGg8zbZNX8ytorSxP3sUAgWqk1/fGuqp0R1QvN4DUztKnkwJAc1/tYmMDPUER
9SfqTv33IAjy8GnbBkHjklXESHHEbPHwGW0svMbgNCdkjjalgiEKUsBjaCj0xCTT
WhIS4bmpK+04Kg1jyNb8RFkAYYiQ6olTlb5P5d5xmRKRuwFboodqJR/sOHuquRZk
XWZXvPRHnswaQz0DqKG4zKe1CL6WFjWx0wREv7e9rBZ1hAByciAnWJYKGewfzLUZ
AHAXOvE+7+WSXKzAPKeYtVj2tqqPMuWaFnN4tnv4NWQ83r+YDLI5nGjmUWdfL8a0
59SK6270b4Yk4U0ENMpFH6LVS08rEVBNBPftK5lK65hLG999T+GA2+fZnvzT1M3p
yHPdj77HJ03sTYpHUTnlLAH2Lni3mOGiQJAhoVRhKP7wAZpzrD2Zc3+i9v8+iHIs
kH2R4ZNnmz7ZhMSsDgWqgRQUtiD51kfo8QXUCGjb4evh6s2QiaYM0xs5v0ZBE7HW
H/b0T4Ac2ZEgV4/Cg0MwRbWzhk94H8PLvrYYUDGxMcZ8DhhN/+PMx8IxQjFz5ZXE
1gw9ZDEGedvu/HFRBvHATJBIGGSAyAjb3EJFM2zyJ5mrt+yga7ag+dQmEr2OHR/7
P2V4ekVYE918judOBR23d2qV/R5oL5vl08DuUsQHb48+5n/B7IsHDKWHHfY91yIb
HYWi/DVB20VHFjBR+UPh/FLZvJEV868+TaH2w9PtlS4kd6Fuupo7xB1ZU0jq8Jpx
yIpOUHqcjkTvNJoSxJKXbyrMvWgEcmQeZanYBq0CIQvpvnJquEC4zrRKW4FDlXY7
18x32TNdcdYuHKVRC2pjgW9seYK9iCvTWW95w20kwmS05VOFGt3HdkTBX47qLGdH
VIgdn88g4iQG4+DbHGxV4nSueRKoURf4tHiHXaCmFWysweK/BkLwUQbgQ0p0wRuL
buOY0o+QkXDZfb5O8CtONiSicmjWiqgK7lFLi7AtwUGtryJrouqXc488beNlJdDa
WiLtUOsNB8dTzlqR/i3yn970JYidWL3iL3X+E4GuCVaFnA3cnr72a9cl5UYQnR/T
lQ+RfTIDB727jONQpuBjgVJy5jjRnRvO2HDOcHWyvxSn775Uo7LWAZacYg3fkJ9e
9FFeZtHcKJv1oO/Q5Ym5JQxYqPt5wn2zOJZ2VTmsCdsLwRIO1ncrqqiLQiKwffOk
xQdjJq+fdh55mEW/NG6fAMX4K4/ELYMb4pgNqrqvWu7b/5lKPdfr/AD+nMgHA8T1
PU1daRP2uVUdislGHYJYjMkZ7by5odYpDuKjSlttrBR99OW/xRu4pMvK4sZakiig
gfPeevSAeMOYhVzoVODgYXvndxAx3bRmt7kmdGGdUQPRf3EtiQlaYelVps+dfsKd
ID9vqodzaZ4CacyNNKnVA3wuKjqJVmNS03mtrrqS7a5XifPCGgejPQ19dVuw6n8r
m3/3dh4doKRITdyZKLDodZXFIBfVt+jZEPy2FeWtEH65+EIgEpAhFh/zxkMiZFv2
qRwkvcc89rutKhNiZr13DBVcDcdQTE6iHNHY8+mIiE+TPLH7gs9KqePde94GHzii
GQN/JF4+enoaW00T1h4RzVFU5vXbwH5Vz2VuHwcdmGQotot1a4B48HmyNWet43PU
fJaSOSizS+QlkBcftsxfdX2BovQeeZpY7hftOYhFaOPB+p/+V6Y05+rJftO6zge7
babF4JStPnQPz4z2Xpl6zG2w4k9Qo+MIIh73Augu7X5mjE9xqb4IvnGbE1HA309m
EZSL//3t0oDz1LwL5gNVr3lHOvW5i6TC/wYDy7k5sLBZaiNNLdcr/+EAwlYu86n8
Ccxp6vi7cnNzp0QYMCf9dGCdO1kVP3aAUjjviM9fQFlDE/fsLGqHOuRPWdZ+8XBX
jQImcm+Bjmc39pMtqGOlvK85zmMbMT8M5TVJWA73B11QkJ1b7+cHn9gppVvqBSxQ
3WmyU1fFfdBvt/Y1OVPC4kLaH+nGLelAqVNcbXiecBg5lRNEI67EAmFiNpfN7uVm
+cIU7eJ1mlzRDj/ZgA40jxGrZV24wjT5M11FUAL/2j8m34pLq7lLkr4xcYmUzMhL
dz6Q18GwRQ+peCrUd5vLK9z9idGkzlzsgH5KHton1xhp5gtlaDuJJYuqOT4WASjl
zo8PaHYHcN1yCMIUUILWtKo6FBE6baE0LALNwGY+53EZIwSd2hEUbcgSuTqBPPXq
TXyWCCOdsvr5nkh3vwCyx1iHRSv2BJf7/0TOJg7MwqPcZfXzwV6kQ4zKL2gokCg8
zTvtJzv5K3VxwnzN1HdvBau4Asw01G73xetkRpUjp8Pe3955A9zawKhwkkiMMWeX
vJaFHHzPYQjrGvGa1lXgQg/j2Pvta2lh1HoDVGQeXb5kxwVTJi6em8kS0gim/Hd2
1ugNxILJNAj27KVU1Aaz5Muu98HSI+tb8hrxvNC0Ifzd+pYpRnEIc/z9wUPGxJvA
wj2GdG0hpinUQpvNkHUMml6UMyq6iwZ7mnAyeUYPaNk9M7cb80z932LLfCfItdxK
Kup+QFDswPgkrX2tXWe+pBVdll9PtxZ8hz+tYH2KG1HssF0nDJSCrfZ3VWTPE4dQ
K4srHaLsn8r8rL/Mww3cj+VQZ3I0RNHSUrNGs23LKlH655dPdZviW1gKDwJuRla9
rLsK1aM1qsm9bR11PR9yWj/bMMWhse4Wxvsf3j3I8ER5shrGRcrgFBXNinB/vsRY
1t9YDIOsxPU+zd6yllrcOBmzvdOseaQ0StO6hPOhB1BnGFUUSvjZtMSmuBk6WRaa
VXdHZM59w7BJ7kgsaM9xMqZNce9xYsWXAySGoGPjZZ+/Y8KrnFOH6XdUukPT952Z
7qAiKwSEvUxGTMb97Mms84bdH9dXXabf/weOtAWWl85NXoSHEeUu/vy4VY2a8d+C
J97Ehz6Vbv2BpVt8v+uWQMCsPofQo3yynoYd1/RgLRv++BJ2JBrZrCPnCQX/n0MY
bGavadin11VpB2SHwlx4HAmnO3KUZd/Q6VzCqnD/kyw/P+kh5c7uNtcF+FJ10Kr9
MvM1CZQbjjziX62uxVOcqC9A3+QWtaPtrgcX7ZVHWz2yWL+acg4pe4loQIVEUjHH
Mwz9KhcaubaIdmfPKz55AdFQC+C6XN1MXls0qHfWaBkq7UivxZ4PUgP5VcsQ9CoE
Fp0WdVXh23ZadaE+5XbA54W34UBgOxKT5sOaDelKM4yhXKhMMYy1F4Yoro9tYwmH
7K2z8ry8axslRRglibz1VYU8bldcFGrxPD4+hoP3X07w3CjFV0TSxQN9kUL+eFfS
+x5bpb28gAUxe7Z4lO+cPl7Xu3B2/cbr8S6uSq/2AqBZcBivAWw2FEw/0YnYDJuC
/1gCsPpdbnA0EfU31cBVUYd95VEzEsat3YSW4vMJbRENDt8iy2oz6MS++ZjBWw/f
YNYlEamRVMN7DJxUp8c+08Qzg/G5Mjs4O/AuhJSAmbdvj0qmFFJ61YWPQjfFjCqR
8eQ4+1L1o2e2wz1V7S/ojVpUoNirJTXOxabDOQv5x9iIWqgG+e3+Y7WUgUojLacd
z3eDinr5hImLCPLRl+RACr4qAQb6cKNySvk37vMbj2rm8Y3uSJhsHI12pab6STrC
k6/9DhiPQOv1mzTfZZTj6YEdc7ix0JOUJH9tTZSMiu6uG/3wX01GXCRB0hDKY/db
dwpzKiSbrHDFUHbP6hoN6jTbcaeNcXhweU2klttoKtg7Z3U0ys7l0GSlTImih6hH
jZqJIGk0jL08tQevUc+b2zrZcZL4jsQF2U0MHzxvb/w3T5cXqOdeq4HHSVtjKa7G
D44cM7CfgSEeJxb5D59mxpEOR97GXwJtb4KrNpiNJNOh4E3fVr6rpdXqlaVL6VOc
pEiDMK523WN0crendx2Gffbumr4KRlUoQUR19OhaDm6arHurMDqIiLm3I2R49z2g
G1ucRa5Mj875LceVyaPfBDEyzDqJ9yIQZvku+3szLgdquWzFrpjdL1W26mCAirqw
9U/ajtaiED3aeTWQFaW7OTEz/zT5smahnEOeBYshxti/Krsi1uZcVfva00PgRsVe
rYZnRabWBUbabQ32c22C6LUvovagPgmgXNsVHAAfAIa6rhnFhE8ILbLcotVCMBo4
CDAKne6nXVU1z6nvFxbYkkU8+tNc4iW05G0bzvIRnjkyfm5Ksi9mISLN8ML88FF1
/jGE1SBxhpecI8FUnISP6fO2gwMXSnLl3sasVCENiyMySFSU/EWuzM1nu3FjKOvV
4L6lK/my/G0/MG+atI15G5/rvUT7uaZVThoJDH1nKZRuX8wxMYm9vjcb1LHceIYG
00Aol4YDzvAs7wQ0+7VcQLFqOChlPq1pnKB6KLLaUOJrv+Whotpm9C4QbqK15num
alzKTcM+PAoSPIeK6tZNamidoVZfpoVdIY+9dvAL5RDkK1oCDvPPfTH/gI+US1Ua
HHjPmaLDuLUHlYGlnQH7DvcBtKD8N42SGL/k3wRXL1AdTTr9AHEUIJ8dZ74jMsSi
dRfziCPadPsRXcBybA6yboYKAIS+qBVd/mBEhX1oFKZkET8Nc/zFupKmNjy3Exp8
8P9UnuzznE0MlGae6Uf/Kkb/57j5cQyEtWWnawjtkK81xSMT0WKLD8mLeQY+0pOD
U7xfWASoJogUacgeRF0MnR+pj0rEt9TOwaRedJ/MSveym1qHl0nTYj6M7rsIH91w
Y6nWcRSuqSG3lSEOEfrthmO0x8p0Nwhipx27BJfoNUl9KDeUbWyXxMR9INtSu0cQ
YVEXwXM99fwCKZdAhHCz07A8WD31hJ4qP8xM5BaTPZ2NiZeSCbU+t1m0OMZ+3MeN
z3gumT86zAmJ7viNKyinC+vkw+B8qztZJ4pxmYWIHcgWdSid6V2EgfxXEt1xjIYp
7EuuaU9eFHSCiY8INqUB6pk5ZCly+CpHCXyvdgcYx1jrXD8cgzoL8GhKtWZGk3Hl
Yc6HQnZOPJauntVvQRGrzx7u01s8vJ/7+re/7I5kG7i2Ky+448M7oGK1jrSPJaah
g2H6/aMGuvklaQV48wGDqSI90JpCVw7ZisiWBm+GjA+K+Dsy06d8ueFORn7ITtBW
9LKIYYnr2z6FE0fsb8NRV1iCfP6EzL9gtilkmAE4TBNgswdKnln9rhPkk+JAsRDE
EnCdd5h01ObNaRjc+mvCGZ2fa1BIIm61ssCtH+1oODjczL1nKVF+rrua7OjvB6W7
RadCKUuOPF47wlL9kHsPm5n/Ki/vJsUOv2Bs/k8ztoTn8oHH0lSSKhLFDhKChQIx
p10ulaVxRYKJknqo04O9pve6bqGlQZG7kbs8+NzDh6kiCf0FzyRRywi1RmRnbTX1
d+AaBRx2AbKYynNdidGYOLCvdIulSwo/NMli+KR8zgIH692tHPyxeZJro4KNbjbv
+SXgkbVJvNj1Qiuc5sJWYSeluW4upkwsR1vj2m2FEnfdtezEp5LHZeivrR1pDwsA
Dqczwz4dRbkJawf4lMO+UC2neYXU0qXX0WwahcRTBstLv57rPNWKmSLCJw/brl7K
Fa25o/+qlld4kF0AeJ4cuMzwUJHC2WjQ3eD0lxeguaWDx/jbwRbaQJajn/dWTloq
XyzG4e6hs+ghKrBV6uNf/hs6hdtUdBasUW9/GRjM39Wza4a5S+tWYYxXnTbkUQCP
5s8JSLsfTr8IVuF9GdXLcFa/qMi177YeRYs95+DdSpX2MT68/9cSX8KNzeDoTAx0
hpvq2JgCqLmkFy9IDsUaXsi4dyg5crr6fYCBuLOK8U7hE8MEs8dWewhNj8uGqZeH
MtkXHRt/un+OFXLuBtk2ysxClCGoF5TjaYSoccCgwQ6ZEwUFycrc9jf1gJW6ke3w
9jkYhApThbraAqmp63O8D52kZoXfEw7ns/8ohAPUFZzI4ZkIxhyO2ceikM0vc9Db
IRacEGaA0LLrkZ4VM5UfH+XTEf6jX3xkwoVEH27Thxl9sxN1vy0pJrb4qxa0JClm
JtK7ul8wnQ5tgsYvBRN2GoMI2k6DGjULZcFswtsD1RqCZDZKMM9yN5RVqEqyp8tS
yisQXPxaW6Tl7qRt50qogMlhOjQw4i0O7bHNDPam4FnbAfDesrOYtJWUelxmGdo9
2KMScR3aqE/Y8rTpzQ/f8o1PXtXaZ9kWiKp6TYOZxI6ZzDJSG98eVQxWdgeps66p
kBc+A1t+jSI1CDdZkslR5eANX2EbZl3zxI1zlf5DCaYtdiTfiShTBNyri2CYIWiB
vDBZ5tBZLbmW7Lr5VLD5JddmVxd6sBgQyLwT2qrPF0VpA58BlAhgsLgcWAH6F6/g
eAmyxLbgWTSBxWiBO2iBbP8TAmHAGP/W0Lan+PXQ/F5PHo6by23aX4jKM5+VybzF
VAVdPCMl3QlD2CFnsaU7z392G4pAKwhIletAKdlTyUUUJQNIApDwt6Mmm9pHT/Ek
DRsjtA3cEd5U/cwZZuAfs29NoWhQigMCdyKN2Cgfirc0HTyyRTiCtV+Fbu4gjqKa
wO5C+oK6ZV3L13SAMsh3E/T8Gd65xVAec1kuwZi9yDyXnwW/dWQYGoXaNJtsvi7j
mH2/WDtRSuqZrzHW326koPnai9rBTuZFIYBPqfAFR9liVyPah1o/mtwyDLpRS9tZ
XeC8nZcy8mo/Uh3m7YFU3NwPKZpzmcgCvc03HfDziHoC4+0vTWiJHuqu3qmUAez8
pb5/gDAq4v5oxtUd3TH7bc743vl6KbxyZP68ZHyhQjnHt3KeMwWIO7FIn5uVZJHv
RPW0EcO/klpmSoIHRRK6Z/m28nD7zrC0+JOrtMxih5xesgK+SQ0sjgb8c1XNW9a7
pnRmZENqXyGnpKJzZJaaqaUYaxNFB9G8lnaXqKO6tSgFINTMioEYZIYQuqY85gDW
1XInQbEUdUk96gyLgXc07NpPpJpRyZpm87M4BniMO0e51GCrwQ94gXqjkMFLx2v9
MVWh2jCj1bVTQTxUneNk3CQN6+vFZKyywCAoIinV+ZVatF7Oo/Rx11lTwL+n4IAh
a8CztaS3A3X/1bn1hJepxi1bPldWqrfb85SXwnhN6ADirFphqO2yQKFT4v8/lMo6
1of3v1yUyCD6KsZ//darrjE+XislpMivm7y8g+utH8zjshvyQkespV0gnwIdd7Nv
nUhalVHjJFxbkdMa+4Hyy3cVaYvS02G3yrsspwjMcnBwuBAItlhGDp7sakOveAky
ZT+NXaFd55p9VphrJt9liS9Vfj/0/mlc15U8+4AnqK0G/8QpSQ/CgNwLQWpuI+Bw
fIbuyJxLB5lpF6dazM8f2xJWK9/iJhAR3qXMOuv3gXe3OmzjpNmqInRBQbuZPKfn
4DY19bkYe2DJQvPeG4qdWJZ0z+nuR5byUX7VSUIXzM9LUCQNgzKxPwCRtkzf19AR
WVI/t/uPyqRuMBkV3Bc6rF7wBT9M+CSTkkNIibpntJtLM9BSiCPU5TCh+0VZaAlh
H7xPwLMXtxKlMGCBuERbF3SGTM5dIsCcSb1S5VowkRprydWtWfez54mcnKCMqrNv
K78Z74mIkO8I06jSJL5tTWTZkUsT8VaQKQdmbIvZW+1X346YSB61IOchlmiGd2V9
pjl2ZEOyqJkx2trhFCaP+6nNFKd5f0UmXt9SOXaP3RfCWvazsfP940wVO6eAE7G8
VvurhCLwRFPMJKbMfWHKjgiElDalNdo1evT8z8/5QbrbFyiualKV9U60RtZUylZH
J/+aJZP2MOkhonICPJ9cimRy5ao85wBPM+vMk0HFS6yqGMGgKsJrI/f1mTcS+Uph
hm0nWB94bbBv42n0QGgrs8GjyYrAtkiQq6+a0byqNManljIDczWiNmjzbc1NA3za
lPnegSPYB5r1u76gzc1PCPpuP9/d08exjfUmWuTuVBH2niVeyQJCHVoJm742iiCy
qiDJTHi4GI7QNX8xQ+hpy5BmSCrQJRuKWGUtjpkpsyRrR7CnBy5jps97Q1128l6B
8gXGlhIlz0AMaVfO0H+6x/uIuhLUp3So5kTluxdkaWlyXOoG3Aa7FfB5jyTir9Oy
Jck1qkBt14VtansD7/w5KnhF4qyY21JpSDW41JsMeo1DZSzst4AeO+OXssRIyE+C
6b8X8CtcCxMWbNpGWYXdvVeNlbzNyx/EqdBFvhzDVREVCW1qSb/Sh9tsSqPUcNoY
tu2n6d2FCzyiDxry2oVADVwoGZmm249MyOFqVNMlwaPN1/gamV/pkEH7sCQaurlL
L+td/olHa7oDF+Cg8WrRfzs59fkivxH6pwJYVqJvo2KXbBRU9Hm5lGvAJEL+XJLK
tl6/hqA5YOvfl2rHqaA1oDTSJWoHJw8fJpkbfqjTbD0UGpC2FJoCKWXT3CtPDO09
j7lRZvhpP0VaflOAUvPhL93D9mpmV1XGtwMTQ59//467f937W/2biWYjxyZ95Wbv
8PefH7oJoBO7RodLbZyhnmuoX5O93lAuePJBgEAmkSGr8z7u1z8VqCuI+H6Lf0YQ
zfsqPMc//wwkSXYEa4jEzSv+LFYOZg9nN37HE6vOK/QKHsLWCSLVONSd8Nz0CPIo
9a+aaZDmelCDmgjKo616x3zlxMKc70Fc2MQmjTLFjaPJ0T2Sv4ef9V5v2jQNsYIb
ULB+QA8wEUZfmV988kZkwZLiqPUONz9J4Ks1GJ9/aqs9DvbiRM/LAdrHbMb1ScB0
u+AsofW2rrKd8wcA/RaF87taWSEcfYg5dIHhJ4dhXt+hL56eoduJn/DS6O9uDRTF
Tcnau0AQLHZjL6l/86Eh6TcaTuuK1dxwuX9aBTML1DNflRKem28HBJ3HHQ+bkQC8
t8iCRVRT9C4EKy7u2Y4RY9/8YAVLeovMN3Z/a94RPUxeQxFPo5tIk2oItJFBA0tA
fSxaJelHrKGLD47zitafJ85xq75TOpEAJH8KUvjA46tBa7ULo+dtvg9fXcg9WD3O
z3LE5gnfMhAEMhhEa2koFZWAQcJmcjMjrAqUyLoSTCKrtyUOTeE391zceF4sy0zB
xrjX/PY0UfLq3VPlAHuVoewbsYvXa2sajND8CO2LZKePHieXh1O57vHl+ZJS9BQo
ZQPbdbbqifahG+yxK73rHGKH00PjIlCT9fJuA72X66HLoj5edcVo2DrOLQcxUUEb
MN6uTOD7gxOkhEZsPWw2SPyqpPsj4W2/tm+EObiZ8BPpuaxGE206nO9qLZ7/OA3X
pNpyfAK1B9NOIm/ll+DgJ7oywnk8cXsHUdV3mgWSPvNLa0hKPmNKvvMKaNqSTWtK
65T7HDpSQGSHOc1H0/1SM94wv9Fm8+iAWR9Bwz7xjU4uXT0RBOM/Pe4vayPxf+7P
WEx81yCwNfnZ44F4pNGmYIBjtHx2MdZCOhsbc7bCSzZHvXbQbHPThSuAp7qMwvAa
u+XL/DygXJZUFZAHHXJvnT2hjzIwEEPc+dSdg+Lvpd5psgd/WJAddXNUyJHnhbFC
SZGDgb5WEn6HPWrthbpse9OLbxdl1MQW9MS+jedjza4tEnkG02eZiBdzfiASoK0B
Lq3jyjskvS0s1x4bIUs2sviHBi5s2fZnV6Ezo7ZHtT7iH9N/+RwuHDn8o3JmzE55
mDP1jp3Bd4F+qndRkzb2NBewEvYVKCu/Ol7WybGoXcQH3eyZCBq0XSgm4/lDINtq
5GZcJ8tx/MFmOqdFSqnzlc+mGUaQSFbD9U7E8OGX28XiqHH+LL3vShyK5RucCL3j
JnGLzl4p8mDmMHkR1dHAWV3OvYjsQAfzZFyhx6kDHe+Je7vbw+sfkoZxMdpiX8mI
EX0LZdcOvnR74g28dN1uIhZ77ZsSLKJ8G/i0JPhx3E7hZvcaBF/Hi5xXr1i06OdB
lq6j45rQsAJHg+6UwvGpJhGJanE3z7KfgmjTgCAHJcVI+i1/t6antb7ggv3fMnyV
XhUAvzzTHDB6BCTxiOoi+bNAT0irDpIXAhs2SRO6yPWZsr6ePQmdktCKKPWJ9w0V
6qAJPrWqFBPhEzEWWuqGX89vnG4aAb98oM6/gx5bvCv0V7Ad4YRQlBPf7Q7acwMe
CuETWsUZ6QfiNRku/SzEuIAUbWqgRpyPT15j1zd6I/Khkc9OmMKZx6EfC8PYYj3p
TJSVrdzitFFnxTUee/+57Lp0jsOyqPp3Uv8v1uXpAL5Rj/TRA4IoF4KgIXrbJsA8
lh8O7mR+dPYtzzG0mItbH1xTRi1bUSVIBKWVKeFm6Bcm7HXqUYHCXVSu+g2Ldc7D
Lil6yuBVjmN3t6Ct1rtWbacBLayqF8txFUvPTa27EtokUOqgeS714HbjnNIvVfvh
Ca1nQFgO82JNYYzDHm+5g9cWn0giAmBCuTr0TVNARmym8A0erb3OwSZ0HKsmuI08
5YEPiJNDjB8gnenbOi8P89LbSwVmKANKgHg1Ba0DTwgH/0IrdUX99mSWOGBmuS/L
C62y4NqFs4yhy/7GNnPb2bm1S6QwV8GERxYD/GUCkdeDzbLvJHIhG8u3kHT3gxpY
g/gixAJwWxSBfzwIWnV6KqS3yW/jPokaVInppi8gugxs6OYf3NnwHx62F+DVV07K
Ls7hiLxVX+npjm4BHFhRXGM/ulARGVyAJ3nc8vxVUqdOX+YJABx5IHDaS65MpVeY
b1RF2bJLSQgxNpuHONyWteQzP8nhbpRO96P1sQiDpLUCx/otnSzPYVcZUjPnCu0b
blHZyYDLpYOvNFF3KnGjUF4gYtImI5B8aUTROvHy4Sl48CMFtRBylaMXlsBldxCM
Jrhn5pE0c9x5X/y6mCACc6OTt9T9BCaOdmd+XWdagu/kAhXUMPHHsLf4AAx4xcor
hop/fdZKWtR4AULLhquJJ8TpX/qz8aOggunwQB8fIcFfzFzBtvn0v/4nWVtOsIT6
/NCjYiCeAoAHHo2+oCTdx4zWwZSc0rHQKBSfw2eXAssIg8HidecDQ7o16PCvt5gZ
rT4KPt7GLpM6e9+iCZc6ymNx8o7KIgxzTExp91onMePRMJ61FM0KNbUnFsei2NMH
AXbqpyGjvippo36oy5Oll7hWguEBXVOJe+fGLagtLfuF3L8Cf0GQK3cPXkTHp4Mc
9BpFfKuoB9qQaymV0tHQlI8BGLw3Zrp0rEYvT3hmj2l8fxvycFqxfgIcUHw/iAun
kHXAteCiVcCgcxbntXGAfCUDSawe0wU7+NquTVqHFgVeW1DMm0WVEZUl1QVaCEU4
gXxJXdMeWNNQ2bO/rReAk1j5Ei13qSd8Thy05m1nUF1IBJxpoIsfWQd3LTnngqwX
bGMTowaGAzig31RDSG19PEq8c6uZg3TW+u6vztPilO/H4OBjBoCpy5bUwd0Lt/Xt
KAIJeC8Qthd2dzrrH3YROCa5ueg/SbaLn6lVuoeLcMGJOm+/A8bLdIiRsWMjQSLk
lyBNg+O7KUIOY9b/fnOHYxvftDP/Y80NC/xMycksLaA7hYyjyzSOpsJf0BPltQho
fRL7SnZUz9pEPuzjJ1Mi25bzT8qM53MtiPS9u+Da6cwLP9iXxtWp1KzmUrRvHx8d
wBT7iXSynKGi9l0YlXdIGK0fSFaW+VYAfvwTmXoC9S4eAF/+VLVwHz8pEO8dy9pI
xqNQKTq1yOVa2qYHPiHUhpsoaiyqZCrYHqcsQOrEpWouH2xSIfzoBJswMr+77WAy
FEoPot5aJTiDUWO+qFjcVzVtBxgy7TzkmP+KJkG3NlZJFU5QdPJ2hUakJD4zBgea
wqQ3RqvGhR4Ag2PpzXFcFKuqwUR9X0xIZxPBQHC8bVrE3j2t+1HSbtetkBghK4AE
mAUnYePQ+bC/vcNctbTREegOTlzCDtI5xnNp2s8IWh8kVhZiINZY0U2R1nWSQjZR
SSDz9c4HbYELV27XCmN3ZLyEyBpsr0cRQB+337Qf1ojynesab4EsWMTj4fFkjlDB
AHYBoNFrbFP6XHqcj7ARbgsRnZ78In1R8jsu8ewLjlX9ocmiD7CRD8kU6mO7bF9y
t+j4PfDvV4/w4jnthvO68NJOzNirndQKsg/WHxTlcO3hCXTe+OUg4/a4WEehITAF
ZXrY2NuAtoximReiCjXGyBYn+qWpFU8SHa+dRqJvza7m2njl1bDcQcE5+cubNV40
BQb8wbOVHMK2B+/384QIdU2QYdFtGPshMYS7AzPraqI6fxXhOfGKru+5s7LIOrDH
oHonT7TNBXSVH6EJbCd8NANcidnZVRGu++PGx2yQWvEN/6/ut86l02WWMBRyhRSE
kZ/XNAVEEBlE1k/Wv9x7RhCK+Y9N6+vu2T9/eAtSDTambriTMT3Vc9eBcY9otjqB
YGIvIpYIJxVD0FiA2risuiYw4MmlbnEwutty0vszk6m3Vg46jiCKXatUWht4OAjZ
IfoGF9Iyj98xuSd31HXx6cotDuAHBUlx8kqU7wAZ7BKacw0QrxQ2fBh/PdYtqb4A
P5reLFC5snAuxyKnLMiUiKByViGxoP65RcqIm7HTDiTIjrv6bbcmsIOdmX620D97
6UFyTvE13MxN45N74wpLmKqx14OLrr8R2o1YjIyfqfanXWyYi1DoPX5GlJ0ctfWi
B8RYbXE4zo8x5b9eYrZusqqlg4VZ0ZBR9I1lr/yQpXq1F7gsZL2nQhzKQIQ1VWPD
YtKhWcPSqU9Wr9Tg/W/XaKiWyxx6nbD6XkJbnFyBCCqFvIkU2hkzLQx9JvRnwbrW
QEhLplUw58FHlcqnqtUWPIN6b2HThoFETtTw+41NiRrq0FNVHOcRV25AR3G7Rvxq
wwlrsiW/ADJZ1EbeFGK+bdD6VS4fV9Es167nCrmj5riJDzTSzFMjOqlJd4GW6WI9
KnbhobksF5IwFs8adW1DXBVYE2tSWKtPhR0FpqtQHrZoqX+8mRZfUm8PG5VU4rXR
k/He3H1b2NoVh9C+Fw4TUlgod+PIAl+1WX7XnLm8qZJmKfulCS/T5IcoBjG9G8X1
lTEyY3e9VQ5UcNOEiabaC+NLWx5GGwRCfMeBibmFq9LkZw6nP70vXrUkTivvlM8g
xi6qN9rMmELev2uq2f6WGQ7GQ+DVmNSorvYwSTJ1IlW2AiFrvNaFDdOIeSmvF3Mo
Doj2P4aF13Qqq9nK5RmkREqDRklqojF1dafScrrEe/6NXxIys+a8lmtCnDBmWDcm
LeL2DKLPaUXVISSoPaiciAEy6/3ABuFpOeDkHt7DcxaajMhLbupB+SV5rccVvaez
qbBfayRDAVzN2vrw2+znWEiyBJLXWIgOUt/Ux7rgCFAUkSv+5K7zSb3cNfodNCWL
hlz1zC131V20WNv2Z3hhYImk1QFu0Ro4huT0C7UIpJ+lV5GSZ3UeGns/7r2DAdgv
Jau5306uBEq8ocHveIkc3FS7VsVydrJ/vGZw5IxDPctpTSquNwxrcR+eBs0Cbuw5
JU8Jh7NF4A4OpE/dOzQ+xhaoot9IriJkDwKSa3Plg2VnYRbZ/ggfwpXRMOeFzUAn
JlhranA5V2hAxoE+CSg6UyIjduC/Lipx0qPOKKJYclFy4OQZqfQrWfUEiTbKJF2F
4v3mMZa34eb/czbvoDlUl9BnUn/0KZYodDt76Q4Bv2GSA3hRKKrnL3glc6tJa1eC
N39I8VmydlrPC5Q9V+siL7ma0iL98R88CoyuJv9RhMrTEQJYxhApwhatbHcIYSF7
opwb9hlLHlaW0WjZJlzRRaSRMMm3HrWLNEFZCOw66+xXIz/xrtBb2V/3HbyX6W1t
xVRhIAzi5J1Jr0WW7FgPLNWZEEmf12DoZQkDHzsD91gO72P5leS9j4Gm66vRLpgG
rAp5n/JPBvLCu1P84nG2k479Dd7bxnPA1II5Wb+onzFYq0DIRzvdbG9xUf3pj6zu
XeqWPcOF6USfzGzLrdgLDyj+naMO/bJW22IF7KCVhxNy1LPFyKH9/oD070P1obKm
8eZvwyT1vRxZ/5ljugXUNOpq7rZegmI3LxU3B1z88mdszIbupe2guCfdrRCOPeIC
ttu4urEI1ufVt8z0ewx0c5Q0+Dqrwq57+M/ftSpIxsgLJcc0zGcEwRUJ/KGU3NZ1
RQFEubR54cNSnDSOxJ47oOcf5r0X/EQle0o54+OvO8LFNib/BU8yg/F4hd5A8YVq
LSMmEm/BCUJwE4u5TBVI1JNz2w9gqtqhP3Ee5sgKiUV0N9CAyn0pbw3lLzKk+iX1
8WRBk+WZqM9KBgZGi7286EKEJFm8FZaFiqwEAm+dS4fS3MENrfPbOm6QMhP5L1Ub
ZT0lAMpA06dUsMlGXxs3+R9tfQIE0YNLX2YSUZzkhy2LglxP011KAYtUP2vHkVkO
0CsmgyrjTvoJRKHlzWbTQl9heIah9ZGwQEZf+VwkYUwqgK5+dt/ip8bK6UhkkzPT
0iG2PGO2sI9TRVoUvsVzmCwcbj0l6D4r2xypq9rKNaDLtBXt7+ALbIAUcoPFn1PS
9U7K5AkfKV8GMEvhXyWBMcT7aAbp5Vtl6fu8WAlV0UFXnkyAn3f/hitFpErzOsOR
dIOiYjYTesgugUd31UEFg25EIblYbP+fwrJj1rAiXSb4pNK1R2N9WXLlu4e3QOMC
0OyqGIz8ozJ2ikGeJuEg/kd/M5VmEfIdigLASyrcMmDNO/pFUuScmTTawQeKxChJ
9xiy1fzM7B0pLYbxq5OEAChDFBXtgKJeUfHhRdTcLs/nddZf6Jaq9VgiC8d2Y93h
sp7557GGWj/sTGhky0kyUsI92jSKE7F7GKm6FF0n6Ix+Z7F+0nzfn+dQ8Agiz0rl
EiS6FZH5kAiFAPMQgPognzc9rRZM3JVuv0JQgrxMfD4fciI3jfqDW/BCa0cbVy9b
jI8u5lSbm44JShq5B2KEAR8zyFgERKa/YauzJN0goVPchA9lRaFIwhr+jvMVDvrt
zvLgpa1KIC6s+rBZamM3m3RDaU2svx4bRi6T6mqlsT3YpWFgpaIIxTv4ax628Kj9
E9Mo+5FTFPugwfvsjvd7bobPqDBrNOFZWteJ1uhXyn29oZg0fHpnk3g9JAjAfTKj
QpAV/vwdoHH7MPGVnYsnmT9dJjP3BAPZzabL88YgW3otA6VWe85Llxr0EC73sYob
ytmkS1GoijRCUemiuK5f48NB147fPI4I+xGxzNx/PQxVuv7CP1skaVoBLeu3/c5a
HDRNWZo0VClz+lWeHNvQlQtTpzd0awPfrA3fOXBvG7IXO1/0mvDsilFOaYngAMtX
23712tCB1C9lTDPp2LSUYdw9VBV3ctS6uv7LxtaukfNzhRX31lDY1YsqouKfCyYI
SwDp+jLCO58tAj+mOgIc5Y3DDQUnpoXZoSEuaQu1f6m/87UIwD9ZkVLXepNnHevs
jcoQ1P6JxbfpahEr/X6ESPOfJrSVZpFdyiFOY+u/8EctYEmniBdTTl4KG17WK9nQ
oJOmPnmsEZMfZX9b21hA/TghkPl6ptRW88aq1M0ucj0qQACOehAxmR6DYO4LSX/j
Vw5gSfT+XVkW4UyyXOAKCKZ9t+PBDkTTUiMCCEcG/TwniyqNhTdjZRBZ9yIHxCpK
r45t8Z4c6venBzD9q+XKd0lvSUElL0uNe2zSGO6dMkULg/ridCj0oxhQsiC1Mvp3
Q3PHq+yhc33UTJ5nq0kIfwJevDJpmmGSZDOBZr1LXylqqx3q2gUsTxB2/npOGDDq
uwg0IRiUO59Nxaz4zsdYw2lwh3m3tHfZAgpsWLRYt09WoKRcap9R7kyYml4UVRAL
xWO+tttumwQnEPbO0X6wQZDR7ukRCH3ehtVjHjV3H9NcofAg5grDS2d/HA1z5gnx
mExtWDJsCuqZAkvACpnAqj7/bLEpam2+b6uBNDjQ7OMuYIApPj/Lnn5er3YldL4s
bft1sJP1AAFJCUFwpEjDpYTVFzi+ikXztSsX0qHPPLruF/ACRKATZJasAAFi1XCp
438B07i59lYEeS4/DneydXVd6P5Jmo7uB0lrxSfFpwZKRLSCV9jSwJUpH/jObeMe
4Zibm8M0oTrCoWrvUTOc7r4uLUrfMg/uPJys7Gi5qrBvoONjnYU9AicADDlu80ki
sg+Wa8jp+hhRPHHvawkaDkJpnGC94Y0jIe1Pf0+2dvTovOkiL7FetN1XSL3TNG6+
EQcn8zEM5Le1OFsOwe+Z1WQ8QM+HRXvwVU92PvC8N6uYvvuyOORXTKPQ1rVuRyuL
WI4WgRJvJB9c6vpVIsRJNOojf/y+sFKMju9MyuYijja7xcFH97mCcpdp+IBkK6fj
t5ci961vsEk1BF9+CPx+tLH5xOQdy4zm6aXzIQyaroPR038/mlWhzVTHg0DxORmw
sYLjvn/FdVUauyUMxhbNNg1HlfZfhjVVzdQzu+Ez1o38Vfh3Q54lwgKJsug9hDP+
roGLGtae2KW/D7NySaf1TqEIFwq9iSMZIl/jbtbBSpa2CwVISCEUvDMH1LuTbleK
l5yUpiB7v/wstnCIlowI8dl/aSQiQJK1Ryq0L4DMuUiggP8QWvnWUr4MLx4v7Ja3
/MMD8l/HY+fqHkgYCyn+zB2+osn+FFJb3DhdhbWjRwgHOa5mDwccfRa7QOTUlfQ+
vABbkGZnHM2U6GK7RjpoXi7A7mCL5SvuNYApkX2dLICNIsxHEnct4E3ylwg8qM4E
ReW2LBHVgTaiaL8Cl06SImYYY73lJy0adm31ZHidbs7aPFbR/L9UDLTlnnPLowGK
QlDSVNYb7paCfZGdfu8sxiILPch3kUQmKhGEaX1oVCVeyxtheQ/hRbvMZm9calH7
WRoCfyF0X8NcYv39Dga74PA4HSqxGJL8jV3MxT59KvHiO4bDE6OIunvxHFR5TzJk
bF55qUr9Txg91BNZiy99SExRKFvBqbIqJAKDbnj/T/+kT/NwiFzTQS+gMuaqAdyY
BEVGbVtA5jPO0Ti7JdTlQoiJ7FLMpFFrGfqI8M07Awmnuak6rLjK7TpjXkujaeDc
EM1x7UoOTKDqextRmKkadXhnFocbA6I/esETPMqz/Qo50VLaAIQfc/gg+h3CBhin
UfGeWO5EmxMYYZQAaLkM+usNQPFGcU254iQfsv1sMkABW5jxvIPY8ijFl1p5fnim
61P9jEPB32ipELx+uNhcXS+oDOZ1M+VANLvmNfQozoUBT4WZSiy7AlQanc1jPoK+
kQkDWKZ9pWOi/Rdp+BQy9/fp/uxdg0jz/RjF1G6r0UdqjCpEoJC1dnFD0UVzlNf5
3GNJbWDtJM3YiZDpDsNfDYaXO6+sZZvlDOsTaMariv8z4KeDdQ+6UziGMHXq9I3R
nP1SsRJwcpWQyIX3FlZqcgTxq5urKiDtJoqHvCWoY+Td+ou9eG0djz478K6dh4ty
N2QJizCwYmSPLO6L2z1iQu1mLOytxEpzcQKnLSgKMG835FqZJSiMae9nMYzz2xAk
X+oYb566LQ/1mcOWHH+X3XEA4e6sdLt/uIvKm/25Hz/3L/iqdP1JoKbpH8IwBq8T
7zqN1CodJzoBzIRCLEwcuM7rOwsE/CZsKpGIvh7ORrrTIdqsYWJKeIeI2HKdm25I
jludqXm8KF3GE6ycQCP30RujRFw0PQOQ+lONyukpTut+zI2AF8hrIb7HTdHVqCFV
esejGAvgtDthTI5fTB/MW/xcv5bLIOe9QYCaFyJG3C4hjqTIj6f5L0qghewFWY7/
tJ5Dh21+hi6p9c4PLfTXfip1CTv1nRI5uz04a1xIeUxfWsdL8TM6kyzTLWb7hUlC
AdypUkQUbxuhnLJ2btqb6kvWrSWLUt/femWi+xKwwNM5oFi68P6EFr6EksgEBUh/
VDkaXg+1URAf+DPz97etUJ1jv47ySpAPRHxh/BHe/6VqN/I0TA0gCRC9iA3i9qT3
modx6cOtIKKZIEElr5yyC/2gito31PSxFajHRJtkep72XD5KQXI7jxxZkG6N+qdi
J9giySwT6zRh1zD9+uX0yu/jD8AlWMdT+0PO+E4B5sAhxVdHMlfrrIAAlxs3BaUv
GpEoLX2YXJoUWDw3pp7ZDc/Indju22a/aHZ2pY7WRHHhaj7tm5co2JM67TZGNH79
H7hU25WpnxmM0g01yGC0LUp3cMNBaA3XZ5KfRHHE7NmEIQjcwEyEShtzmRTBKkxP
KKfIGLiZEHaD+lFJiNRYxp6a1J9tyNfduwiNUYXonmjPqhh2WdNFdnCQkDQKeCnU
miVErphUwj+a2H9ysabT9aX5gwvTTaa1OwEl7GqFrrvPs+A8hzHTBeOfPjWFMxJV
7NYUcyQTfOMrjr5Xl6p4681m4NfPZLFBLasRHjqEVdAbgjwwoV4k2pqhiSATuwGZ
yjPk93M2mKVsMebEnziibKBY8WhfxucoZOK1R+if606dWEVkm+BHfP+WsVrCC/5Q
ON6ZY2Sm0U2/iFS4ZqnReWMfLWKzelzcPEsJ2513721J1gHS+IYpw+pro2iXb3iT
XLIJ7Xg7bVNyWzchL2ZI0e6v7D7YWCUjXPvjRiC2ZlO0I0q3D4wGJoLrmoYkSAvF
ebwWIn9euR6sWzpj418a6CPHfh/3QNuRlrYHrPVk6OnN5RTZHC3qr/WEANHUDba/
IF0V2wDUlG4eFqFuRVQ/Rcg6amKZqZp7m05B1HcMNQUCkc9ePLsN807F8Kq2Z+MV
leREKA4nBMiwU18uyPxi3NXriVbPrKJhm0r3JtpcxUY5YtauDiRj7Q6DeKif82vy
cjmXpfblq+QknNh/43L8iperz42LyzOm43v1j7hQATyp9ZDLShf7Tayqg+k60FV+
x4ksSrsc/YP47SpZlf/BZ/XUG+7LXMtmIYn8pYLKstl89zLdYada2vtkwlGsjf/J
7wuO2l+cXmWYJOZ+ESrDcjttZNbUdvKIi2/UpWWkfq4elnxxemcsqIEDqqEzQPd8
0LmQSSUt7htNqymlRDw6NY4T3sIiVtHCT+7H/XJhFiik7RLobWViJQf45ByHZbBP
ahpzrWewjiMbE/DB42SEwyRFWtmOAdJHdhNaAqTdnVxrCD/BMmci/3igNaM+p2US
UnecOYqO8GlhrtXF7BKDa++Vd0I90uKPXWkciXuxs0LU5jb4x3HFL2ECwcCL0TKB
gnXeIh9yT0pmlDcM59JmPO/ykJ+siiwsqLr1FI4Co602/HSdNUyUIlNDGfRRMw17
WaxRg66RUefVPvji4kfVIHUUkhtFhjlF+nLTEVMBdI0hixRl0vlIhWoF43RIwZtK
vySg3U38OpTv/9gzdLhz8VYctPuJyv74DETH7zRSxxwHaa6ZdZOTpn/DpMyO4PeF
QP0kcLAmiM9islvXM+hbfUEIUbSOgpQfpm4pW12DcnNOlMwMJCeZOcKK6VBSPjmg
tpm5giNN6EqFVCtsS6+Z4uX7R5KtUSAAjl+/l1QJXhb85mjbOQx9d39elKFJRI/V
hVyQntfcEzR/ioHBlBoQs6xXfwUP1jjn2gvyo5+iwoqnL9TL4TzzmRH138zPmss6
VDBPD6KJ3wrwX/ggdGgWhOKagpcKXiXOo2ul9LIm1hV6ay45lNh6RwKc5NhEDsMX
rDk5fJiMRlmuQ45Oap6j2gJ2mQ/BoaW0FBbH8hyM56Kk7aWbHtw+lRSg4sGPcWkA
SVZw4BEKXHvPeZFG5+JatAc/yIfoFASF4QepqXJs5jSffbUsIKEui35JXpKPusdb
Ypug+URqqesAQREH4TnFLoK6jF2IRD5+d2OqvVKCtbrWuhd1yA48A94uP9+ShGfe
l1mhq4GNRKMZPb65zjV9/9FjLl8KAN5SYQH+Ex8m/hyfrLBJ/2t5J4tXQehNib6D
d7f75eQccjW01t0oir7/Hrd07bj4z3YjzXTytPouaX9UrKxNllVmHIPgpmM1b5XQ
YeCf3BLxDlKiWjRKTb3R2q0ShYsYJqmgumU39N0WH51jI+GNi/7W6VC4c3ChW3VJ
7Y33mQDKjOVGXrYGXE8WFJDWpiPtN2N3GxRVcfRQNTncRASGoqXmAC3m27/TUsl0
ZoLf8SdAUEpKCJNtKuWwKc+fwFF0d1Re9HsKsFbawYHY3tEH0X0GaHYJNU5U/z1X
UmBSZolWttRZAjHuFopPRUgASJKvJbn0B2st2s3JTNbLMBTxTPo9t+2zqDxiPjAo
ZLnMWxu7p9S1QyQQC65BrNTL7BayvnIeKASNcBG/QEqmPGG90qJHrB3sR/9XYKl5
iu0UxSYsBQoM8AcK4vGhvs/vGj/2QIxutxFW/VTH/JgA4OfyQFucfgDl72TRBhLR
5zcQib2ilCyzvp1c+HyGvGLwu33BqPNzuF7fgPlP7dNk/bYQU9k37BshxUrJPfe7
sCiM+Db4/tfR+SJ1o5cxpGt0sFD5bbECEc+yKTYW7JVumb9sK5nYWbRLlwsycnR9
HFfvnLgHktW8m9fC/pzSnXObdsYM7kTWw+4SiTIkywvkchBU1L4WprpCBxEPIAuw
rA3twNZAaop5PSL58mIeNsrYcZTeoB3V/kwFObzYJzQYAcGorWuYfasjZsDxsle5
4tTZvR3ya8OSUIy2jFrmHiT+n7DjF4VQXsrhJeRlviDLhn+MhMQN4ViGe6z7uYts
u9ZabbvfM+1l4N+8WssLTyq5USq2AdDeWEJpP4+d+6ISul9QmhglITMy64U+hUCc
5Qzs7avC5RzIHoIqNRkqqU5dUYkgAKuR3jGz8x/1liknt5ijhEURWO7Ol4MT0t/g
dtuUz9cfyRJQsM9+Rnm6+gJ0Zp4Q109F426ZCD7+57U+rzP4TKS7+ioTjSIagESW
6KZe6Oqrx02LEi1r3MDMf31lu3ZNqNszK7Qje9vaocm8aaiuqA6sxvL4zkDcvxKd
MxsJWNsm84SDnYi5a0FCMmAXeKojBDr/2/JepnLlFcJ6GpTYOopWYlMzbLp17U+W
OOHp3CDtzeNMjPBTmiwcDSWsjx1JckfH4ScwrIE79kqRpr1mlwufUV3vhSkVlhij
/4FsQLN0eNwdyeme7Z7n6bub6NmHHkljjALv55gHqMOxVYJHkqifP8xW7oVbJv2a
o5Mw69KOQwDMhVIL9jFllvbC1dgiOzWBL7Qwqk+zFgv96fZs3lOrFSupp3OCpdJk
DnM5M4Jk4k8ro6vn4QrZx0l72y3nz82hNE+ZJGC3oKqvz1ndA9jxjAFSlQkoAlwJ
oE2vqhaSok/bVgP4VT8A5Wn1hbXqpfXQf1jX1DEa1cCbqjW+LkKuNGspCjRcGxy3
ecRmdegN8t7pUSH2KzR18uLopr3mTCtz8ZeTjmEfnoS79IL18EChLbpf2duKkcHV
2OQlKQchm8bRIydT3992E7iB05ZDM+RJ8M9ocLVP7KG96geOQWPot99+nxr5oCvV
IgTf6sKCAvQbioHoBoqnTxbK7lu3hW1TeO+2zfJ89F1dbmqPmLv57XejBsqDetzN
VwqOiKIZMCv3xxUXwCrWH+07rrN61rX2iq3Pb/2I4AyaCdeN2ED9K5Bq/aMHkKIn
78Gvgr0XgtHsvBN4fl2YvYG20V1Fji/5EteNAtPedgoBgRTjsOnZG1U+xxWNC1Cn
9pQN6Wda5GFoy1ZC1r4Re0a90Y1vuC8cBlCqzVfL+vCJ6kUbscCyXm8PBFGlKgOa
V+7Ciha0Y1e/vQRqlnMtk6nIyXevUs3u9bYutwnxTcvXoFxiPZj3G65HScbhsWpO
vfLMTMW6PXKWBe2rZ482xLDq1mvXjBaU7uXH2y+f1ChQ0BOhsy7TAnBoXWLmvftJ
xlGvwnzFTmG6NDvjzOnvz/7gI9rvbsqeBnt1T7bH/5h6Y0UdA2uuAXcjuULOxjMs
jPmtUlfCFZ0TrBVxkxpOR5w5l03+sy/Z+/AIQ0US1S8LLV/2AIiDggGYFi2M5/h8
flRS07rTESfYjlooxf17lmcZyVu0dmHr1DWCHQpoYyT+GGko9EkODJN93ILcR8JM
kgh/33AY/TWaUNsFbbz4MQuyyn/P1yk+IONabYoqOnpebI7USQ7K7otK4PgV9cHc
xYJeATMLdKCAD6eUq2Ttg9j9zryLHPvbTpjV9wfji//bIQ/bD3Sj+LZQsuw+5cKr
ANgmNKe7Yhxqwa1lMNpbS/nksN4OQmEUM9d7VwIlKume9yo7ZuESlPli2dDgxQy+
cH0HH5NZG3M6w10hYMNID87oWralweFy7AMzV6NgUJgEZXkJJNETg+d89/26cV4N
KucmysKDCC40Yzoau2Tyty9uX99stpZaMJVJQAaf7AkRJpTxl+bUrI4XENro5u8l
allLq5sq0pUzM/NdRwaOlH7SfMxyZBf2NWNhaOj5laNEsBbat3on6sh9Uma7OsFo
5mCTiSdlTJwAFP0zKelOJmmlePw4ge0DXqWUfD3ARlqD4rA144EbQnv010Q7QKHy
0/mOxoSZXce/3FpS4Qu46lbFqUHTRlsjY/YC4vZMqIc7xhI0w+DKF3xCRh9bM6CR
2J14Rzx5abM1xKGqMESPQflmnV+tvzoqhoO/rT+E3ZLyTYHQh2VxdG9oy4oXXMfY
8GkPXymxeDR5vhNhBZoTyB4kGOJAAc5hKMWepFsDGQp7PPJiS61buj+f/2sOH2aH
wigsNYuDwwdVyYCsIlBPXwqOzX34V6pqSYPt2ggZvnNI+Whj6CvWbS/FHMMGl7/v
fkkKhd/FMVXWA5grlaw+sCn0bzvJugodFnA2XX4I5tgxoaE+pciwKSoIo3AkHymz
Bzpw4D++6gKc9lsgZ5IZ8Q48J3WiI3dfJrOe65h85nHFyD8E2R02hhp9+UxRQadk
7avyNi4y/0Mk1gR3WqzHtgJfu4+pG5qpxtK3NKE3OowpZqUblPJDUSuTRQBmIJnB
+Dw/CUqxOAEFfQX8upPF683tbtzZsVxQfLupG44NojkzbwqEqLnEGx+4wbftOdi8
PAF7fn8EUEdRNv/QWyrce+7S+UjWqB1WywJQ9Q6WztHVqxNVDv4EzDjCMGXDBhDE
+SNw7zykB4sw1UjvHt7qKxOS2REjw7J0cxd52lVUWf4IYqRJwfUDvBa9oGulIili
1sluF/Rs9eHea38c3koFe0KUlMwd+ByYT0n4+iQQYRx8oW3mV+lvlZaGqN/oY08d
3gg90ufiKotDmEfjATq9vcpN8Xswdm10FUgMCkGw3XnIg04hFle8suHlBFkBqPxG
bFodzBh1+0BHj3Bme2F0X+MbxBMAmUG27VVw97mGSF9rUvch5UeSDZZZ6mLL+VSg
zv7nZIgOX2ZMW5W2BGVK/yTQLWqTA57ZH/e0RDdNxVpi8e2A0gBeE/JUTSKjGdYQ
emioCQh4gacykWYwi6qjiF4WnboHQQIFL4YPz0IpsVe4AkFOTHrz5+0fSbFsBzEr
mW+ghxwIieFcGiPtVeH7nyDghCtqHNg1L+xgnqtAVkXSwGEOx1EBJ9DTl4ghomvO
gUnBGa4DeM+dvvih1csHLVwDYuwCdKXfNG+CmqXaTZy1UOzEbPEMl0rFAHkqM6/e
kNm1Bvm2lwKStz8Ylof+XH3PjJJRCG3SqWGhwYjcXaKtyZS1yBI+60tX8yg6Nr/0
yh4VG9H3YBZynza0rEkPLL167ieBHEUFPrhbqkoUKnIi3DC6GQ2yojgzTW909eQv
cKRKhiM0rRbxBgA38JmdiZ1mLcaROxFra5ubuMWPmCretUGsntP9XY5b+2qTv0vC
0IoGFn3mZZu9XU3Eu0UTezZ9h/i0Qlvp1q1q95lG6ijLN8Cy2PxaRrD72CkrcU0w
+DD1lsWnRKBcWIfEslG0XhhVA+iHuzE26E9c/c86cMAjpvzs2Xt2PGNTwODCnnit
VzGHbHt4TCe1B7O3auzJdJKSZk/BuqCr8ux/7V3Rb1axu8cC1fKcrNjzw6esu8rC
RlqgegSMfAT3iO4XH77xu1Ma0+c36DOTB4mOUn+gXcZucL4bNJMfK/+W5iMYiqzP
DJMMD3Qcx3mP0ULutl3WWmE+IP67EYaoBWTGLC57VXC5DPFdrqKkp57fJmhht2u4
GbMEUg89ifgiSQbkbmQgruB7m6J3GZsiRptc6tA9NuarqyQdzpE9j5JxFVKHzeKn
9pryjI09BwMYzM6B8XNA14rH/l3k5egDnaTpTWK3s1dmrDe7i+JhoNl1T9wKoav3
KqBXqstoZQYtBrFMu3LKjwMnZWTjjNatJPix2Sp+5DPG2PLZnso0+0+l2nMzbDCF
6R5d0qtP6bLLJNW3XdXwKu/IL4Qp0bawJXp3AUTaIUshuRdUOIyHSi2ZT6PjoDFu
O42hMFjInRg/rc23/7zBSSFxX9Sj0Ew4lq5vYxkzJXz8/MEb899ppzkuUmTzzsvx
dzC5RQpd7h6hUHU9RV+R81zbb77yG1FGhaaO2ixOpcuuHurnssFUBTyoC/vHclP4
PyDH2JH6OvpEZIRTDFr9ZKvG9IHcSDwg+uSsQ9x7kSxsJkoXnUBE/aOlBrqrs3rY
x3sWh62NBwZ4amhDG7NRuodBn/B5QQNZWeRGfukO7xfc0L1nOBRxZ6caewu6aBed
R3ZxouPYLwWeqC7zsGKjGt/7fplj4nDHxZ4qA137qcHZWdJW0zaSTXUybdA9HyXN
q2yhoLER7Nh0fWYbw/7J+ulzLpTFQgOFuEmfhe9pqbh3RsGV2fpzxp0H3Kyfthpx
suduyz86AhpmqVYWCL8bHUV8IfauVZ8PsX5qUeeE8Sf+mITRn+ZirNAhY1cj2gKV
OBcj7Cat/HjwhHvdS2Iu5wVya/TMTW3qg42T/DQOIU+5VvQxRVdcp1X+uLhWS0K3
ql4sXhW3R5ybX7UE71/9OkX7C0hvbNwDjZ5s6dK9MIYD7n47CNJPsvAqXQ6Xex1i
Ww24SxtVQckLYGHY6L+groHwEQJi+mZFMjeaZqpLFsYp4duD3IJex+7vWNkVaeSn
x77HDPT7D+uK3gZdYVqTnyDCL7QzO7AAnvubw4rLVEejAozY59VdbsT0fDqvvYzg
EwTt3xyI0XXdZGPhigFiuUD3+KnXIJb6OuYnRC3FTExV117Ilp9fm3VzeCI/6Mld
+8+FiJQ0FRq2LsBLaTMXS3FqdzxnQCg3Ugifpg/fPhMvsDXC6LsO7an2uFFiRefZ
kZrRHnfaxq6lzVFGTiXamwcHfz7gbdPi07AiQAAblV37cddC2WWdYZS2PSxs7f7X
+ptGIag8to5BBMvggMJqsrTR78246ThbQklZiIN6xIPIwrYgrg2cmW55lTB3eKo+
69mzM9LSalqegvN8Jkz7nj1QV11IK6CaAlRYkcDmhXWZ0bOlzuQsbt/BbZAvWQxk
Au1ZHoMxpFMOLd0sXDla9EG+jTJQi79uhqhxtJNOh10zUXJa9GOm4gd8vpm6B69w
A2pI/Uc2T0stPM7I4GvzZBNjxPBJfe4TAcUZaDBUeVFaSL7xl6YvfZdkkLrenjW2
CLcwT9FcG5OEWC62kD2RtFyyrSyiM0I2AmN/lOZx08QY+yWK30vUTIq+E6jWYAoy
hX9kCHMOP7K5+Bcna63/u2jg4OZnvehWYSziZCifkIhEt0A13b0lnAsNECfK6iZJ
EwFYil4X1hAZRS3JqQBvJdG/kyZzV0HGnJz7tyfPQ/3d+51w6+UCGTfxnkrbgxVb
QhW/qiy4JLjOLwWciiC5x7qfuEvPArsDqg9Hs5bf8ySLFFQk/jE0hck84LaRg/Ku
J3g7H/JsCaNu1nLidI8TZeESSc9KlymMkhxbnasRceIqZVk1bAzMFoG0svu33dF2
MaNRyy6sLeHJt+Isk1V65O2xLOWORRpive9OWLwL0y6yTEJPa9oX3qXcJRj6v2W8
b6tQKcublOtDbGyyuLOqSReiptwVSLEH2d8pV42PUMEuFo/J2l/TzYh2Aawd8wDp
Db8kyJ2JY5PooDoJafnliaFKKS+zjXGtwwDHBeUoZSwc/y1zBZ0D4xU5pUTwPsfm
KvUnzI+727pUYq4yLlruznUOVSrvBBbgvxdPau4BpEr5qyVGflYj110KI3Yf5PBF
vQHzVz1OfsLRcyXOd4lKNskaElISuOYIA0K2fXlyFpdEBOj7hMAox/catf52BNb6
5NxgSKgB/VZJxbGSgq7J2VfhizVhVDH67+X0084a2Dk8qir/5DfTkv87MFowJam1
Nlheqxc9sxuu/tNy91UVaU8hJSWs9ZjnR+Vdk/LRD1h0a3OfT/PoJ90UtrN61TK9
3wwuwJ/scZXT6v7mjxSEtBlMJ8H5FYpqu+Sd9mfERy7dF2tNrC+zkeuf172Jv4t6
/Th01pKOIMOPy+DdlZDfIBbTkZQfG40d9RBnKFo7ZB57XueoM+b21R3IzdIm2P+0
NScsi7mA8pqqOFmz29TpjFT4Bv2chl/mVQ4R4mbfetrRw9E25exJAutRkNLS4dev
cEDyakQQSw1ZpIM4YVJXSIw4R33qSiOgJb88e6oKjQABlDlO4LeNPf/WadxVdPKU
WVpQXLHfcF5cqHqTp8XRAuTemYVu7waRmQq3XK22XUWbi8Na+2wjS4g5LCea7acq
+PDcxUznZ8GT+6/JzobQn7Xd0BFwDR7G5hSpxrdusNigLbgnNHIK9xHyXFKlobtQ
f0wDXwDvnY9fPabwP7e+tZM7m62FSBOmNvPwWSTkSupM26tRXVFosGOH2WloDfXP
tLXfN50UxbStL6IFDSuwjuJXHFM9FC/VnLGzabJ6tCXK45hLXBGO9iE0Kh6Q8+mO
mxoDOjRHsbgUGQ17RZWhJw/wmAqQZgPsus0MQ8NChoRh5R64HKxQ+2m927EEF+m/
y88ExD5GD4N2ak2K6FThrEEYSbY9hsOh5sTIc22RjERAIPeGxdKXp0+lhU/5BK6Y
MrTbRBdQVGzGhzzN+UfEx8L4gFse43SIhFMBWxn4a+nZl/uH3dSWGzddLqRlT38o
n7y0U0raAQTicXFNqEszdrfEcVZrTmoJ2SewviK6pEbmTZR+zLwpktm0lROhb00Y
Awe1uBV66QP2rql9eb7aqHwrK4QHR5DvxP6+AqMjxxgaRAWOgpV9twBD83ZPQ9QV
l3N+teME7j7MI3iF5D/oh+WQRrrzKlW1SwDg8BsJKj3n4PeM0x/vPlpPG128YpvR
RoeplS/SlwzT9pr6WFGuNyBHXUUbYMy5n0fQsIEK23GE5ccIUQRlgd0C11sQX8CM
B4Bwahb5XhP7peAZkUDcdxNvH3JqH6T0ouy1P9GhtzI5mgaNYrqPQnal4DbRNtkX
Wx8PETGCJjNPC/Mdof4/4ehf7F5xsFL4NjzitWnVBGFCAEyqM6/LD0UNBP38cql2
fsN3TGhbsG2N9o6lM7oWV9GdbncB5oYMK6jspZL6dQZe+huL4GvhJgiMQ6K9ok9c
bvzvm7s56frXqchmGFmEHtj2Hb3rzR68pQYMLvntrYan8KM5UsID9oHm/20OxkdT
FaZVXkCmqpJ/2ZBtC3prSsAz4BJSyAdNy1HupzpBTcA0znZAwV2Z4GdEln0PGiiI
OCNNm+q5qIyUBAcxDT75pJCW+LJsT0t8oIHwQOfBserXQozpHN0JKSPFJ++4tjWF
+sHmG3ZEgJb/x+WLFLKwugHpV9jj7r9ilAmG8v3FJjc+PHIDn9yuqDdvBalnM2Ra
zMZU9C3Sd+ubRtrXeC/i9ECk2gQV55Qs1VivZkcKaFsJYACRNXobWzV/8bux6+Xr
QQ1NVvjcOnOOqCIEzwRoumEETMXiVX8wjkKa8G1LaQS77N1d0dvsj9RKVLRDG2Sb
LybKAplY6XojKX5J9TVYvMJQETFSB2zGE8pkjYnoRpcAuSgtpr1s4wyKrfRRQ61j
MvTaraTrWkXXZ6QGZFR3nD6Ml2hOkVaChGKHFI466Gb4XXq5o/gwUSQr+pt5hZV0
NbNZ4fgO8eGJy6lewIf1og85AYm1aRerUAa6iTvTVaJUsSUTFpqs6XJ7cbmlmdxD
A5zi8dWJgW9V2Eg4OBdsSC+5/kZaVMaXv8AYvxrquO4pic3hDLju7XQz2lDcmToC
U9IPhcJOOzKvCRIisfGT0tD5NESm20qrGv64EC1zvEtgSK/XcRbBBY/LeSeX7fD/
oGYX+tOyG7Mkrk+0acLNtSttbne+JDm2G+wJ/OtmICsRyeU44ZTId6tAC5yQKFcT
XJ1P8Gnadfrb18HkzDadhoUzQfJzOX2V8HJDq1ONGsvDrBN/bzNXB9eEnKAXKwEN
tgns47cpvtRq8GnSwE8o98LiQjZM+DEuMeVgO5x4hjsX5p4uXZLTa7eZjCMy/Ia5
4sj/ke+h7N726xBmE3tMwX2Uax+Ol60uWoLWmLWMj9sQuXzzo5nuiP8cWwdBtpED
5iXLkKnzisaGAcGYXwEmIsQn1zbknyfnUxYhlyZ5BVxsVL9s7Rx6sxG4WB5/P/R2
gGm1THtIXfy/YVY06j7z1iTi+yX25rot08bQFzUY7XmyeQgqQSYSuOImuFRRGUvz
/Jdojfy6RSIDYBvz7iMr7uBCN5CR5JIyJHDZPnrFnNxxC6ppgW/KzW0nYTYMiPF+
jQr+pbcw1SzH7vpGvEzzZ/8lEtHv9z0Mq1tSUUgjsHJm+wAOdRifQDThzyWn0xAE
/80riN9E9/DBATr80n6Ky8BTxV5krE3m8xhFGr7UpmmZC4GipgCsVqrtLoLLJzw5
+pSlIcclhNAboEcMK44gqE04Ytbap5LiFhxAMDrBZexq8A2Tu0gMmjz0GlOKcJgZ
BXIg+EPZ39pwXZkN8DyP4w3j8c9WC7A2SA/oxVdcjyqgXQHeGB5+rAmTXZGDASqP
UY4f+G0r//5+UNQyByr32jhTT/ocNQoMeGByykIgO3wPoSc0Ic8+uUZeYh6CZqQI
wQ5oura0ZBXyaBW8+JAoWkN3Tq/voaDNbue2nAxmvWVCdyCsFmKiRFMdXKV1hQ90
ysOX0FlUPvKE0pOBbqDBIcm5stsCQH5Oiu15EN0tYyUPqU3PV2X1B2NJ1sSIRSWj
lVN6niiYooxbSD9POj7HFpthajLetyMwGyGQs9XL2CKfrdrJGMqoOuBzJxVf/z75
cXJzGpLpjngai7pNs4EW89BgtLv988aEYibanQWfTgmehvgnypIC06hT5KI0nj3E
TjHdSQ3L6TwzWNwAGGXqKOAF1FyCFNo2+POSE1Es9Y5ev0ZzQsMVL58f0DzffcDn
nQHONQuLz544UjmLjZsTjFy+RgcGc1dq9/Bh/bpVVXEl2JKXNPbWwoeHdyJ8LXJb
yQVzu0r+aMreudWggSJoEpFGoLf//WSGEXgR5UANzELJY2tx1HYgH8Rv6rAWwpNn
ZnXWe8+yU4/2WyeZcys6is42herJrIWuD/lkvdlVz6c7f0OmvfAU3WkZn0RctuqI
tRde+Og0z6qVnlIogAVLfIwkFxASAStMoRBm9zc05L/NmX2dXTClfRO209tdbs78
QuwkWokXi2qEbHQd3MoO5WRu5h73ZfPS9NHWDZox4SmqruXD2zzlds2LQRB/a+sH
hWFCDZ/NQmMqoBBZNFgOFmzJ3yvd6Xc9LnQwcgLwzPwTUrR8WkvEpYiDPjFP7Dtx
P0nMuabu5peXtQ3yhrBYKaCPQstg8w/3ylYMx6uoCIl2EMmr8UldYDVayYV/7bXD
Xh0TlDrY/dq8DPbb286E2nJDR+fkAzOQDhyFViMdjyjSSZDv/S4n1JPMm9EuBQlz
beA/HbfDBKiZ5l4G/xZYk1mgbpZRf2ogIGZbZtehnG+VYoz3xgCifv5XINadThTQ
jogxrj1UtJQNfI+nq9W90A7fQdzqtFtN3v0micduzCsexb4/kj7lRiHpSzgyK9qk
cASJxpwQst2JkUNExTDqGRi3O/PxTRoZOjqqXXQoFo4w3r8GYXUMraAxMbfyAVpR
fi7qdoYCWFNnG5KsfD9SCj/iVHCFDsab78LScj75Lwc/gzon4wOE2BUtAiTvyxZi
eQf3iN5uiUcwemlGmHlGeSQPtw7m0i3yyW+HfBsHQwqHVnETL9JJeF7ZlQrVuWsH
wVmYfpNGVOzVcy3VEzzbeCZ+ZUvsDPzZ0MeaTtG7gqgfghp4+7/6CPlPy6Yc30tM
kJmpv7lRFiLjjt9kQG9Ej3SZEH3L51QKUkMtPuANEOyJAmFbsJK8VMm3iUqbH1eR
jngEbik05oeyRnzMSrJUKEQP9c4KgfkR14VEgz2lVl11JWQJWMkF/m8+UILv0BR4
7S7koZGY5sMOWvJ+TEoQfIrIucI81eoMUh17hIH8AWeGnzjxqBtJIm2YLYcktwX6
AN9syvIieHye8D3wjjZlRLSsdsWLgF9B3K5ulX+6ma4gdYYu3Yb0iP3Bwpzr8DYX
A8odh0frH2gqRadT6NzVXlz7BiGda4LvXaz/YDrJmFE4Kudc72d1sFVfbc409zwd
laqNmkG/fdJO6EpW/TbAL+9+/zDIj+gidqVGCk0F/617lPT1YGb0ay+BiGGOVhAx
1SBETE3R52ikfdiDTRJjMaKvKSkJKrCJO3AFNPrdWEorNN/PPzI+KrQXOlGcDabA
xVuTrvu9loCHTENTrMkXLiuwiMpc/Gy5z1Vt3K40fljcrr52bAH3oC5oUj5Kaq3t
t+Pllq0R4rGH05YIQcDfdm+o7CSWOhnmt3bBCPanIEVeHgKfBbKifTI8s3a4ePFe
QBM2C7NiSX4E5jkTe/8OwS9xqP79uCCfIGGjPYGV834s5V4Bwr+1BXWyfiCW7Jpn
ZL3a4H3ewlNoNIpLHVPA1KKkQVsGBpnaSEWYc974p5duHNMZvRCHIXxbxEfKlhzG
mnoXPAx74kSi+7xJMPhApGodtMqiVX7jjNPViOiC8fmUedkc825njUpAIsg3PPEF
r5lhnzMHs8A1bv0bZE1VzmyyYQJ0QckYzSpQZqpSKDmiTS3epl8vkUlIz9sYgY4W
Snw3htI/nkDge6Zv8sfAbdD6Xv/pmsvkjpfSgHYL4XYOUHUDGc6qhlhXcclGTF6l
Iyv5B0aRgiwvVm2r0aeL2anVSot5qdcI/6ZU6aiixdptYTJtmgdtMizBS3KDTnLv
hphSVae7yBPJoPKvKmlF5LJLTnlJiq8u9yDPbgclCDfGD8s5X6qkv6S8GTnNTS0Q
gAXty4oCltapSErdoXD3a0MLduSJbLQNJCgVFIrjDDwqwVLQeP6ZvXmjVwR/K8AT
QWsydk0mL2C6RYeyKLv14vzAuXrMwZ/XrHzAH3P7t4xotvmgAAgJxcyl3jvipuUv
exxX/hlJ+yD2oe04riIPniIq3pnVhMqjGKAy0Lnz2PLOo98oEQT7eJRlvznYwCMw
koM6DSP3sgkzI4gocMugNzDy4VNMrWfcKAU/Rc1B13oF4CM6B038SgrpH96sRivG
ZqDLUXm6pyako/usfaD4NUtg6IOUCWP1H4nY3LJxqMlH6lL5wZP92txXa/YBLMRn
XM/1Hek0DW4A8qwTM5XRLWO1nFv11FMsMps61mom3lnAjDRdQYcnKNbemeX/wKb2
oZJo1CQdQyjLqd9hfEovXGT+UdnyXErS4pKk87GKb1OqcjDZoEiVgIs+Smuq085/
FEuItG3aeN5sigGjJYkoKccLNwAVBMAqcJH9otZVluI6DxGJl2mmy5VArWVk1TN+
ggSwGGex7G04j/MESIsGsS5OAQkjLY8MOgq7aTkuvUs312Zla45+roK1aPZO5v1l
oXx83jgvou+kGSWksfzY2EoakYGMp5C7tHVEEWNNas9ba/rKKvGeoALqCmBM1HMg
vxFoULKZrOD9Kv3tAtvcjmw1IeaIW3480SLnkgEGE14CyhH2dzirikCkEjCZ56OH
I04nmiWxI6rnwOISSjEky8dGZZiTwjYadhw1loXl1BGjusdvg0G0evYNCcYAQjsT
6q/wuO1/LXJ7IBQZyWzJ395P0eG0yi95gJg2JawevGIPjh5Khu/MhlN2809E53tv
g29Fm461PIrN23ry2LJiloP04fSw/PPZhefRy0mz2G3w9LyIvr6BpVGg14Pv57J6
axNNrQKTWKBIcP97pRFg34slDN5FQCP8cK/Pu1R/W0Lw/VWa/5bF8pCU7tGWZ3RZ
IryH5E6hIICxaB0X+NPh7Ip5XGOFCDFL7MTAddRAqg7W7Vxb4YxigyMZLeUdUMMU
Xz+35wcU6KX0RyfbpZ9NuQtIORXMgUPGvFujIMUZXpyEwcmFyHNVfhkUAqlxSCfc
UhatdX/S7684QjXmtdqe6TurvtpC3yZOihm7PWOL0Sqaj63SJngdaG3W7mY47OjT
5Lc4W2Uf8PdlA0TvQ8hTok4v9pFPxgdIQXiYa/uGxfAqKLGVJTTOIoP3DktnEe/Q
IRBjFtbJBZgrNjKifnlw6h8w93nhhOIGqZsl8kdgdgJ8sL7RdDwg80qCv868twuY
LMA3dRKD1VeavKXNaY1EFrNAgocxEPlsaludHbu1I558I9ewGZSvmL08amgdrNxj
c6BZRg7H8c4Dodo84XI6mKR9AuXlga954koPtVpd7RyEJiJD5bcIv0evqAEAmKFu
gF06TpgExb007myGayfg7W8ADwmVICciLvA1xmz1OKcueyfaHtD9/LpBLM2TeZSH
JRo8ipYhRO8npfiS9txbcmPG6KsmnKh+9IP6EH8c5LNIcQSOTtcUm699EebXK+1A
zsucRm+hXDD2n3t6gTRivEsflKpI0wVXSEpRPoojo7UrVnuIpjO9S6MwXBKKxqyF
RcpM2Cud9B2wtLCSTVIqp35Ej/jnywE7PEZCIqxgBtM33inWfLpVUflT9l94Qn5k
v/JfvQjH0n5/KG6lpe6yWMZlhRGu6g0+fhmkwqxaADHhoMb1Lv+uPhGrFVxBnXOX
TTMnDeKnUX/mWYYkjsLEzmZsdBgi0SJaicK5XPTDYhZDpndLCN/RTIJdpsedspup
hYVzZgf0cgn8cGCJO9uPKNN0l9xQHi12UBHvIswjKct4k6UHTe+Z5T18iqBu3rde
E8NKTgn7IgoBBMjwvI/aoWnIaiu6CEg94Fs0M1gGr5dA8u8eVxw4I0RwfvKs2zVn
tYqBfcDtfWm4X12ea7OoPcwQ7SrqrKOYAwgM/X1Pwq5NpDZIUogD8+KRHhXHk+jo
Tu2bhsStYJmMdlZ1UNKk4sFsbmSmrrqy6pKooJlxqtQ=
`pragma protect end_protected
