`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GcNdhtdB4sa3JXuI8kjbF4NFpmTyqz4V0RW15+hAT0H7s73zfwJ1DcFaSxVGHfZc
YbX9HSSd/QjltWKDKE07VcAhSdKArheQg6nFmt9peTMSOfCbkkdNapq/wkfnSd+5
ygzzJOal9GHkx8hOddtdR4I6ypBiho6WObWJGUi7Lls=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35376)
jAbPIcHAllzW4UtQtmoCKgOVY6sx3rjy4RwOXtkoTuzQ5gEhh2s8/k5XV2+6iLJJ
92AkUTfi4px5R6TxIJUB7oIEkhRA3Myn0emvE6yOtlBVAPJlvw73r/lDWs2gXe0V
3NpFK7m3CfHAJe951nRO0u2X6MgP1dX5sATJlVCd/jhMiDcxZXYOQx5Mve3cexwq
fdir8RjR491M9pBrejXesptzS5jq5t/TzLnHCDl+kp29z/tcgVK5Io4eCOJ0y3OQ
HkF4/LynoGkhHqvAx7Ewhzx1m/8XUldfl/UyRxQ0JDS6nGSthQUElTFDkdp0Bnkk
ZYwcU7Gsl0TxDOFcgIWlZyEgKczuVhWlEvLEGvuFNYTyWbWEXs1EUsWWvMyKq0W7
+IoGlVy/ovBFwdi3wsWFJ8LtS4AR2c1X7nc/Utoy/YdyPMyMXD8RtMW6fwS26+Zt
nRYd2zI3ZsFGxZt+pQrjjSceLEbQqJWZUBYX+holxn2xnpzOvbKJg+WousxmyCdE
U0PRYsdQqSq/rz0sVsEBinvJt+H/QUIWUF4MZ7KjPN0Xahv4ANkwGW+sG+p6EgoU
eOVW+Od3DqON+3tiAJTowktRYwFi1i1zYpCB9SnWxCGLc8OA6Z0HDTD6+2kUvFZ4
x9I+nRLOp3V5JvZbnZC8YsJ0orO3RSeVrVZbs+nDkA9cWYl+CZX3Lnx7HRL6FJiD
Z9k8HgDCB/+1wbrcN4WzKRktkXF/xEdC3jtKIy3fyIdd/iW0E5hPk+KpAuJgL+y2
WDJIzkFEZrd9TeMjkSUvxCMiaf/zLLs7XcFqwRVwbiXd3KzkkMKhcnzqCmfgSbA5
MLcQ05y6W7LqdFLERe2cKjUPZ+A11LNro8SCr+KbjlfaU+DJ3Q6aKsv400qK1IkL
1dd0DTzTfZpP/AiPdE7f9sCC1o2mel+yqkfJH5Dx6oDGPo4y3leL1WMnYxgV4no3
D6FlLX3aQ/ZaROkI8PIIWnwUaNnbcNe4opGB+5jkodaPTI28AqADLaPiKX39408r
InINhH9vqXp9iQ0pRf3bZpTVGILodDmirzq5gAzVGE8ZdkblcJyeEZ8ZHd3Sv7xv
neGkQ/wHrKZb4AQ5cz4HbSMirTm5yCup7RXD8eiyllhegCRgVfXnhgV9ChwCSy1b
m4bAjBGmtH6zDLstXpMewdq24zbSwYSOwpDPCbPogHIqhBF9pdxB+5JAUKdHIHbE
2rHb14WhI5blOsbGBl2eF5UXBJJ47qj8vD4NaBOomLJQot0YEQB1ku6uaIslBTmV
ks8ELGT3m0/1R2JT+fPOUkYZ1WKEHq3N4KMkgt4UL/I3hNEKW0bmqszh9R5rPS3x
KniwU2biL+icBsJXRc7PsWbYVEl5jN/oCg0pmobv1TtF8Pem5j3cBwW3lpSSxmKl
JT20tDjuENi9a4CgJn7fF1r+NY2KwbJej6Z5jBStPGBF6PCib9j91SEftJziNhxy
gOctOAkU0WDm0tVnVtcFBawAcFKA6dAmHn2JRmFTf9HtVD2FvZ+y0L8jgAdAAhoW
Wgtm2z8psyZTyyM5tVJML4um6hCOmDbwKvNlaIREHcFbS4KA/5d0GVRLJrO+ShtQ
TubQvAwo81Ashl4T8Drtk3tCIYG+6KX/MRYKEma0JuBLT3Tw3qRfBfYYK7KRqfnm
MWR7NxVYQw8lAJ700vrR4WhDi/8tTyePWNlyot72CRFxaRqirbdI036sc+UA5M1V
o21BEE2bM2lM43NlUhzTMwXPaSZ9KPeKJSuj17VjZB4B1M1JeoFYG8Bkh9SiF67D
MA1vXz92sq9KhksRmmw0OQnd6RCeOsNzchoBE4mfI8KxKVdX2TDkJC4fN5UTmMzM
pSceLjwxxxnIXmWC/Eul5sp+88oChddNMRcI60SaVIA7f9nNccwAAdOu2i7bdn55
m+NrIw9SEKsIDRhEXFXabndUjgYLCVyKWYYJUdxsP8d85h4S0irCFrJUOSCypnvU
KpxEOZf1Ia/es9yCCNzFL0EkfDHNfee+59UvLzmLyVJkJnWZLacXGYHVEpR9y1rb
qcJh0bT+JaBYfPWXombPk9N9Og9tjtY301OAIIJC9daShbkHYx8dYX5ewN1J/m3A
OP5c06fPnbEHlIABqjPMeNy1CWiDr0miuKSix2tWv5V2qPkZGUGkHqur/1FRbGyP
bFJbt65+WlSrxOdjykhFgZ006Atx5KYiVQ4cWLokokDeKIAAlNl6BkJryucwcHVv
yDy+uU3muYhuPJb3K2DioLG+6HcJftkflmKznKXeqO15bYMvmvBdvK03HKERcA0d
2qf5R0lPpEGH6dS6KCPU+aFTLjzw78ytpKmBBquAX90EAMpn+budE9TNbEkfAxO2
jv5kKMfMDWSp6vCd1fao7Nroo12b1dXu1iciT1gna2Md22wKfLQQHFQj4RhM7fa9
Ab1Sfehj6a4B8QBmdiiZmGvpLbBaUfqnZPr/zduYTHRVHVTIlthLWLpAUd5YsAaI
ethcD5pmbP5udJG8bq8PcOC5svjU8NCeJ8Xcn5E+iC2L3sRlasp0J9OudNjwleZG
Y1/vvVEiKGQOpAqfDIBsT4X1epnj+VSzXWkZjlBL638N39vVTLkgaBDm8QhZyVQx
+gLSWd8oTYkxqtF0qQaNTw/u8FZJMU4QIuYQz3IlzPS3jgD8V/9PATJa4SQ6VAO2
zGGVigU69G+rhgo2FSEZnMT1AagRLRZWLwxcagn/q/jU3J5/M7PajQ/r9g9157Jj
Kj0N3Z41cmtlqDjGWXcFQg+RAxJ/a+dLvxFAgA9qZXxJQinOa85X0WMH8hfuY13D
BRoR9jck9T88CX6ndzvbHFrp87XY/S5dJxbZceOWsO5M88tF1+d+XJr3HT4ETokC
04kmIMAigtc2L3VnQjMPeBMgE7c5xtRoceLXyu4ogdx1FHMLSWgFVYbNt7YCnuXW
qlXqw8rqLxnrI+V0sMjFCBbOduzIBaf42ddZdHt623Yhz7Fz4TSODk+o/p3KQ84/
4PBb0ASWMGqtIUex54VwK5rkaxq2+bGqi6brkRdFGmHZIMshxdWAnbepGImoAWMG
JAkP8z1z9+ZKoJsZZ1gO7Uh4YcO3Dnj4z0qGQYCFwvLTyDzQD2GNUP1q+aijI6dG
pG4niGPIeWM4rY2ySdT3l0fwTO+bT86HBZGkMxnRY6m01EnWp/yrQfuhY+NTJyce
gF22Q0N5yyz1kY+ID42k+mCu31Fh+vUmikfYbftR1Xf9ansKy3NqkjPdRCxokCoi
/M3057eiQNHl3scJm5CRo7HFpX+smbtQWB+8sivHlRTiIoxqPDD6Ezpr9JX9dTxx
XYENcLQ/jAif5Y+SudXcKP7o981KCOVuy6xPdP6TKY8HKeQ84IPGEKMBXrXfQ+3/
9jdgfkW2FhjM+hOxTqEherRL7maKxioQKf1ueHbsynvFm1NwG+9cRdySsUqNdaE2
jDTH7DbhZ/RcKdQCgbPff0ATPLw4Lnag1u3FcediIgU7J7atvW8tP5kP116OmZFJ
T9Im/KBsAwhgfZkSEEU1LDVTv+tCSZpVeKnZk/FJgCH8nevyB7TtnxgGvR9XWATy
ZfYulqVxrCG+HURtF0emHU+hzGJP2nErTX8yJxsqRcu6kgQ7Y2ADMT81RSWFvAi4
fjkuLSlFPEnkNsWR17SGalrYdxkkv1Ed045jYxUSC3gGOivYYAV8uO13ZtIOt7Np
IotF/RSAUcxrFNduRwmPgvQQ1RQc3RccQ0uTjDOR+RoHSqo/RZRZODF+5dLfPGkE
xkig01k8J2n9/iVZW+TbinCr/Xa6pBqLpuShZyKIsSDP2kmCdUXzbTpmE39Vzp9Q
ydwGNcvRTM4FbArcdFdpGhQ0uT0hOowbnyZ4pDoS2lQ1nm856MJYc23IRdJGFv1c
U+3UjG4R+0laLOGqzeWiJ9/I83lYec+bAO8uDFzDPv7ynZnJ9GXV0dNQo/jywG1q
lXnoDwqUobPbLSI44Mhv+4wJ945hMCMdI2FFng0sI6nf7wj0SUfHJE6JuYOPYkF1
uXrEAz197mYJowcMxeWT2nFC8gZ4Q0T6mVi84FbfwqCLhXQpeOKMnfno3mhdw6SY
Pn035dVLNyTcos3hdpS5mDlYakYAc+3PghA3qsKxEnVk2mQGx6XVo+oPWrLEHvJo
FDN1HsMtnDj3kuaf3cW0odkNZyt3O+VHhj1ip+Vx+ndJ379YJ4Gw1H1Vwg/KPTgx
D9xYCREv+7F+YUoIY1bdSwQnLugmDE5Nr1F0I4gTF+hs3mNhB99JZ/kzsftSESJq
E3niwsZFCOIc2yYKbvWroa8e6DHHE05UAo+wzPZgkkDVfGucH6TQdz/nyNoZ7v5I
LEcSKRs9OFUmiWAHnj0qvPrsF8zWGCGGuK63dYTTgcxO0/Au0xVHbLk+h/Emtgif
9Hf2QRI54+fOnbcMgwI7eXDj0InHtiqwfeIg3rjnuiDb4dE/a2s+TqCoBQ9HoFZo
qfrJPMkr/3B/9ZIBZlYp9UuVak537CF2JH5pTrXX5066tpugGjKbmF6qzj7c/GSc
+gAume5Im+6qIl42EFCxRDsB05b73wHL6EUs8rdCWWnFJ49YV67RqcTuS8v8hANp
CEJdWUgvluQPY4M5xXA9U3srYaJoatVcHVoNuJ72rn1AqhncVTFYEB9Oi/HoxIYz
mmwCqhW5eCzgfTyRudlADsZGx7H5jYQ/J9FYW186Koasn1xpDzT0P7tajVuEca7L
pNmatGoF78mVaKecxZxIItEXPlL+QgTTiLPUPQ8JHkYZq1A+wgYobS/f0ob9PlOf
dNtYb/GsDCjWoYwJMOoFbRclOkUdcP8VyFwPW3v1UgkP5KEqUAWvcVc9yX79Fi6D
r+RCWbtqdSZ4++rJAaE52dDiq9Da55YAGZSLjqWwEu1uPO9M9Ijus/hKvP933Of3
7V2Es7UdQe0cm4gYLjeFsxme9JSphlQO0SBpjgXH2JXZDaniBg/bVcFCn7oiLT/v
pp+7+7YwcOTOee8sDtF9WG7UOq4YS+JAlOi+vS3m++zISTA4swKt+ehafQaqiz2j
7kFrEIF1rfC1x/fwuM41tAiVMHyakQroEjvfUKPDgXQUC6mMIUsHzLndJwqHc29h
SDdySc26ZoOv0gZJontS7ZcAokodPImftI8IBs6hjowrdlds2jtUn6DyYXprHYQX
E4Z4f7bh+TWAgiqeQILxBBdIjj+q6tlRePq/0faHkoL/hwITHacy5hoaNqRQJFzg
LUDi6NmcGf6QFfEo/YlZ50dwkbfF7d+j60Vfno9rNFowVx/5VzmoL114t4qrlqbh
YC4zrMstFr+rpUoqoo0d1l3mB56nVQ4Iy9CZ1CUZH3ZzuHsWn7jZpMzTvPaNJrUQ
YUmMDSJvS28AT7VGH610C2kJx+I2hdY2svjlBdQ1YBAfdPGHvWO63dx6kUNEzv/Q
HF56JoXc5bZqXa/IQd1bFJoz4swuK1cxSfAsVf69eghJUnDloVyi9oQbDILETllf
pyAkAU6HQis5ME3VgN/aQRc2IuZZmuZhpY+W6DBGOp9VEKairZ88DaPWAYWJsaKt
uHKE2GAltGSD6//JmnnxzorA6t+1Cs8lMk1YpqIptRmXIywONjtphnyBVK7G1+Fp
5lqcUp2kFhzhBc0NSaYIzHqy86nv6HMDMpXK/jTddhtmNBEhcAZxRMZsONNs991n
olDkp7gTaa0VYktC7IBFShVa8K3+syLYgQdj4pjcNduPuVl2EUuDh+RxF3uKzl/1
6OdhS30dEWcsNtDpLRF4pgCN37gdYq76mMuuOc3E/9ncPmcxaufb1AWY0TYut+m7
WvF6AZvyVITrONDDdy9mQfKcg2VQHw1+hrdbhzWLthZKH9M4a91n0EPoX8/meAuC
xagcFQkD/5Gjce5okRH0V11LbtsDRDz50SFyIUE6wtLRSj9m6TlAyej620CLEEvH
itSiiwH09vr4pmq2b79K0c4w5afR/kdHoL35PaJPlYhAZCvBAWy1mlYWsk4VteJN
scGWUNHggKtJ1xxRY67np0fglUiLSxv3tyaqY3TVeyPFG0Fyk0+2WtRISp1y2Cd+
BMbndaXgK8haDZzed2bKAvQIw6XC1ht1x6XLyhZ26xLwhIlbCS/P43aZcdNLcSak
39e04LCOysmnWxZFjbnytIk3O5IPYwwHGc3ZHI3QDaDGe5JF4aXnhGvA/dSipXg3
vOUs85zQ6kyJO4lMW7dK6fqJY/djqDkzwoNd2tYjy8l8Wpvpcx8CIrFN1EEPsyfv
EryFcHI4iPPLPpC2SUbY+F/iURptlpuYlWAL8UnqfHSZMBJsOIkjvBELx0ectgvY
r88UWIINu3uNVOlMBG6dccf8k/Acew6LoMp99Moq/ls5qMzWAgcmnQPiskE35N5B
tDvwjSh3OooIGhLr/BDiydKTjrycUYr3gW5tPpjFUISMYjFdiiodNv0fJxoT6atG
CX41fHDR8ixG7P8BAMGI8nZf+wG5MP6OfyO9Y9b9kHN1ccjenru3F7aUgJ4CSciq
cr5BOTnvZQ8XvehflTlVZFlEeDETkPgL994JmEdksciDA4xD/p1CUKlr7oBhXJIi
5PApx6MhJnnFSeVGNMDFKJJ+Ib2wHD15v1ZB//NkuqMDOz1dk2nM2PsovFxZlRG3
gjRnfmMfenkHOcn8D/1vz9x7ouDH0jgmLFMOWADUZVM1V5XfYBuky/zyPjheVJwk
poVQbDs2hKPPLr6E3XFQd2epZqguc+vKYC1RSVAhUIwlgi2ASR8UAZGI/bxqMp/x
ytaIccmUuPIkhYYAdGvMdmKsuzGqvY9fF8oadEYcUJyxpH6jyz9t49DkwsLKl/01
EKBG/UFfm/uUvRG044GJlugN/BuXLEx1xssBjkkcU5xcP5D5RFAvtvWtHDy12zB6
kYAfweCTnXcU1PRZmqpW0wWKP7aI7cZcLEzQJcBeG49mMszsN3gI7tFCWNfEbZnW
aPqiy4qxm/XNLt3nHrS7PBIu8EM2oh4t+puJdIkFJE5Q49jLNCeobwFZ9nkIw3oz
eqBBiDmdwa/zMcGsq3B5DLoK3pSAvasswHE8mS7eqSWYJKIX4Az6N0WBmAbjUDDO
UKcf/oQ5nBG0H/8tDssDDl6fTx17+RVEDsLy0cA/0HrUoyXYzWasjmB5OFQnduZt
lqcBGVpyY1qiRksckifkktAq0nO7ATiCp6aXLTOvVaOjrI1g+xiaL0ke1vUhm+Ai
tdenz30SULks078lQiX2yGkKIX+MJ7iI2nq7Txkv7kra9t5C1XF8Ub8nQDeCdmmo
za+4DBWJiLRCdXcKOWrdF1H4SAMLaRr1mTYJxGPwhTBjGdf3aS2Si0tGUyenk30/
MeJ1fy3akaTf8IA6qtR4kYes7S6kOVe5g2Dukw+bGe7BDPvVPZRCmxyv88vMKeIg
dt6uyuiRQfKfrYkMPY7rD2T7ZTsiW4FssZofUX0CWtf0D+PyN+Ny+ByOPjnAe0Gs
ANMu2jvvwLIT2B3i6BvCsGmFuZ4qdLGac+s2YxebmX8q+f2sbE9E8MbdIRQUEoAY
lo9EUSNlDcczoWk+9U6Gse/qsAI/h63m6VA9rTv8QDOmqMp4eurpuICTmwfGtAM3
L9GR92YqOfOn0fzp94UOqpwCr8/aIJEAuvCdHypFr5zv1h8TenSMoUaG3ae3WeOM
FmyGdqooKNei1wGc7nsqJHwYvNTHj6tvWSPwR09QYKmjLyKF9xh3jvHeIGFrKaUQ
wJOju/WEGZuxhcD4mlCb8g2xNEo+FhW6lEUfSWaxNFXGJoyV/5qXdXOrqsPW7OtR
siinfr3I2Un8d/4HsUC76bfO6CJ2jXox9iRtV/uKfBqJf4VqspxjL26P/ukOjlMz
RJgNjt1TS2DEJNDnuHWFyw64PBcP34O0zv9ipF9Jb5iPNgckTEyRlv6q9KPAjqvz
m3sltPUEq00ZWjrxNmPpaqVrMRoUtEKX/vq6a0em8ByDbCgAT0rrTN2NyiRYsgX4
pm6TIXgyKZcn5pDincc5QHVAxw8+VGe4hbnXee4l7hxHABtVA2ME3GqJuVPCiNWP
Ct22OjJjqg5gjIeK/UEsbbQ9tgTNwNrrayD4ekbmNT6ubKvsy6l7b53aQWM6vB3W
IYMXQa0sCUOpYSeyotMXsQO0kBts2bfITF0R+xT8fcx1dxyNx5gzoc4NqBlSjQHu
SvAz7HR5Y2sW9oDWOclM5DudCFQUxNjajv/kFso0cr0DDtXHPaueU4RVlK+whRTG
cATF535z15nWD7vQSnlh2lAGdRiX4wOZbO557e6qZaOlr8yalGD+g/Yx8xTO0G3V
CHXQmSLa7x2/HNcUtLbybXNcERbbDn0/ynwEyCQ0bnPbxmhfs5+Us91C2E1jq5YP
+HmHEEcIbsnswpFaJl+17a8BxvJmp0y9e8sh3GlAi+14I4oq29oF60VdbONNaFql
3H/9jrgQ2iBXHvlw+oUogec5nx14qx6iOAiN3+5E8PQX4LUNWBU860Pl4u9cdZfT
5Fy+9iCiPUB9bqSFfdFfYHPP7bFcVubjxlxb0Z+tCMjsgLzakVZcEkVatiTFPOMi
k97VmaBHclVw1iQ/l9K47gZfoXcy1NPFCCIxaVTZ95PdhDFO6a7n6jO5YbjGaIoW
Fkvu0R5A20Lc+ys4e00KJytXCW8sZPdurl6FMgtWWk6mNTfd2ivGnkqEu2ThCc8Q
z6qXxpvbn/S2sg/dhwLvbg9ol7k7QRvIgVy7Kv36+fJ0UzC9y/q1RkUF27YpFXWq
q0b27cQ13k8QgMek+8H+RXP/jEEVwjEsI2I3YlR9y9uZKVNpsg4u0WCWV8En01S5
2CM0w2zVdQf72Op1ZYhpBXtzzgfTzcHvpJi06nOE6C3owxtuvmqYBWTVxX0vmKaX
iRJmXt5SbSI8yeLN8CZ3Yva9Hlcjh8JF8ScmOOLJqU+OUJZ3Rvb3o1J2tiH86eq0
FpI8At3c9hq5aIFagmFbglvkHooFnwBOnluRH1gPHP9Ygwf/kkZYXi6fMrOB6NEz
D9HtNrRp3K2RXN5s4gcJkBq6+I9bmQEBHmfeLdXsqg4KSUl0n8N/Ph88fK4mjZqh
Pqed9RpJEvt7P3JHCc0ci+a9jh2G5EVe3HdADLhxQbCixjswjp5J1QKpjP+pLZvk
IbMTH7TnT5b2ZSyQoeyT4ruueHg3nwbqJ5Z7OfxaZWXHUtx9EJUyf8FBFOSCcHSd
zQxc3UxDmcw1rsDuXjr3NM5gTBkH7+sub4BDGm5SvIdY4/uSPFWRiuIthruZr/Tm
w//KWxUOWL/FwKcbYSUwWqp1ZroDm0nCmNpb5v5nTQsVm3us0SM1cYqX1IBNrTX+
UUJ9Qx1gZZq8L1Hv9AiLwPfbeHfQDhjytOmzkZOMWB6hU5HJ7O9rIjRvFUWNXOYT
PcwNZEf2T4vo0G51wt0LKvX4y91SsImGJPBtNajA1/yQ9mvrztzgMjZxQHbu0mof
+I7Jna3r3e5xMm5az3DwWh3/0C8gS71aT56PqbJUwBDlkCZaCaam8iU5ZDLdondA
bhX+wJFqapzmu8lTHWfv7FoWyXtEUGGRj6rbRLy0PecLIYwjbhTvjgGmyg1AUuuX
i2JkFewAvzsG8pawK3KN6WIUqNNFmvFHX21vhkAzoXwOCxPGiT0RJKGa789gLjSW
21XPlejO0KP+p2i6P8kfdEo38BeJCUg/HdCwopYcTGtFOsT7c+wHSXSq8p9AhIHb
0l3at6zsKzbSLylouNPwEhZ/zWuI/P/UWDctdARFHAXtc9aAgNlHR3uCuN+xz0uG
Vz8JPw99fGm+OrjgkIwwBWUAqkz3aAmFcLuEb4K9qPXrF3NUb8Biq+Xbb6fh+aw/
ydIM/NiOExP3PUiYhbwjWtCiMUVHpTnLy+1N9KLBJqQKFb6OlsAA6r3PB0V5cUJx
2zBxfAMR3Iqrl43gPsVsK6hP9EWrBbiJsl/8/xrBr4pGbECBMNDB5FcE/HGIHm+c
1iaVn4r9RjRkss3/0vXYjJnLvWLcseuundmA81n4lRBXuzYpelQmjNF5Bf5HD5E6
/FeZGOcqhVj8jk5AfY/lQgOeFPqlJ15hNRrg95iSrT5I4juPuvSwHPjwZQ4CczoP
9BezjhfK072oZKEuYor3pTc1dOHZx3+0BBn6CAObZXPdZR5aYQCZ9xlAs5XkhCqy
eSJEuI4pLQotLd+c6Gc68Hgc0xoW+R4DePlzp70Cforj3MD97GU9TEDFNK9Aj7OY
zqf6vabP+mwfgM8hcTMQp9ugA46k4bvXST84yWlWbQcXCHY1e5x5qqGO4NOH5jHI
nlbEmLXs3HcIkyOouqIUFouLWoGJZZLR1jYgW2ykFPhCH5PTvIB3Kv8TTYbEm6sw
Ov/0RHtm0LXQR9Oj0THivmyAiRDoHjUP5vazsOYJcrUFKD8aslHWr+WxkOjcEL5g
r9lhSlNIrU7HeR3rBZ/h9WgE99to0fCCGFwhDVFIoQlKaMwcRZ1fWFXOozxJTct/
aCkMERWKy9nxNXqDR4GoPQIJjtTvyyd4f6HjdPXLAPTAU4csybaOftWoghv+Kejs
zOTm3FzJL7/5f/tnwyr/wYlM6p8XaxQuT2aXJQ1ZpqKiXrTs5oC29zgj/2Op5hvp
ORhAZxFcVd9YnukTSub7+UnsfoGLVUCp8AE1tvOqNsHeVBIuLgM4Qeb8JGXUBf7H
zUZKH8oL7rJBHd/5r1NJMX2WBB1HUk46Tg5XO4BqYvo9ZKRoDZ8OUnIGYikHJAzS
N/2tizrIyzamAr40rbMjqz3M8kuDzj3XILlDUP+UVqmm9hj0Ot4+xMYBhGmQc2KF
JVA3UG567DZxP05fDOr4dLuQMctyhn5s0NoO+aTjXmG1rS+i0rGDdV0QqqNc+ua9
SgDNID5uOy/J6NiAh9s/vCUq4n4KRhW5k4gSj5JG6iolhjfieKdsvJ5YPmT9O3ML
2hlKMNOseW0IfRPVH4zoDyOrsOGiM5kX9QhdkwxY4FbE/PXWpjz/Ul0/XsVKdImk
jG5YSSfrwCsqSBdeD5SoLG/6AMmSIin5tHb0BFuCurILE+wdjrZbjDqtOUisyB5H
MYJ49doucI439WEkRGVnEoCyS35pUsn26m0ZXuERRqjZ5086FrsgiQ6TSHAPTxNm
92fd9H06fqtoQEc9a7QPgQAKb8L87JqIqnNgz9oJYlFNM+hhKCGovGFah1Nr6Dsq
UaupMuYsZazoYfX8SRlQWJdCqFZZuYbTnj6z63DUtz2ZoG3vZ4GE8TdwSGmsVyvm
rT5OP6ieQECFec3EcYz0qMPSITc+mdv7t/iK9Epi8DeyoZxUuMGx5OSoOVqCAuaf
kX8pEoYwi0aYUdwaeMf4rURcKI9yMQO+EJ3LGNcw+rSlknyyv1E2EhGlj18w7K5B
+M0D/pTbcxwuuzqs5vuAgz6IQqGKY5Vh/pJeq10QtmNwK60UDx4JD4s69uv1reVC
ungw4OoYLeEKPResd8zonLzXqsH6fDtRtDOaTaqQWcODExQ3Q6T0E7JMzTGYonUY
vJUayH7SwgqOp9+yp8KBlDrSogU0lRlebm4Zv3dBm2oYL6uYjAaW2tvOadZ9AJ+W
lgKVyFwlAFUmEwviMv9cQApHceozekkkBIRW/pQKwsUnVFGFZVRbFbb8F/gSDB1U
OD7GmG0UjFm09Al6TaoF7u28uwuqv65/PqigMdlNJeyz1wqK868JQFnVn1gIw2Z/
4FG/rKvC1fBKu74p25abuIu6VUecMX0xByOOaxLupkvhntd3wxuE9vZlz4KVENQ0
6c66Cg6WzrnQQi1pbtf/o08XXk4oOodPa5gPNnHFmnNaNAbNj61QnutlMROJY0jf
iQup+oCM8aUpL3JhedFykvKiqHMF6bnMXgmSM1MdtZkunS3oUertYfXmBx+E+BAc
GpGRZmYHhjWPNmepN+A059XzFCsyJG+dLicnbyb9HWZNWPrZQT+TxlJQUKWsCptC
yI3lXZ3h65Fm++89+Yf0qAVyxx1N1FPfV8QGbrtqe/LL6KWQ3WkCJc3sr6p33DVm
twIwOLslBbJxChsa7MQkEkiLDsi6odiYw4jBI/X+er7jsQGnhm8WAP45R8EGGyhO
j2D0DoZf5Mu+KmvKTYvdYDk2INyUBwX3DGve0g8Df33wdJUT1GIeorjk8HZxcL1c
dYQLY7xr5kpAsNl7jNoa3x6YmHba0nTnEF8p911NkHpySDegAvJ2UlyDByIIiHeG
sEDuCh4fxWcGVL3q+gRZPxqybc8CW1v3aE9/68UJWSmExMJew9JiqE22s4zcZi9n
jkYL+LTvJ4PhpaUkMkXDNIt/Xd/DeBWfkUeJJzuyFmKfT8hi6okR0JXYXLgz30YJ
SIWOX3W6/XQ8Ao2G0dltnwf7p8otEyzginiAVgQHemul9S9HsQWUXzzUHc42IZzt
XYXQCWj+eocSx7U6+DbDs8mniuv7Vxk1e/3VuBlkQiJ8IWj27I0n1nJxDpCzFecD
NFFonZFzEU+MLsCvo0YrGncsNR0vzeh+e8cR8ROTvm2G7t2LdKUgRE/1vt9WLCeA
rLUVZxJxgBEp7d8PbM/xbA4x+j9IwIoVFUAQMGBvNPiI1lsLHH8MkgoJhroRBJw0
H8+VXVLnRnHxY6stjkyeDFcZu/c4tj+dzdsUeo5wTJpD0LsfmrUUWoWz4IS6Ptnz
HgfTTz3MOTkU9hCh7EhF5zs4z35RRlYxIDkE+KM6j/7p816o4f3Rj1gxtMcioTTN
to/YH7CMT7itsrOI+DuSR9bp2CZG29yPte3b+JNMmTkcIY8tPEqX+v7l85teBDGn
7EYKGkl8LDHFqi5WMNy6MeesNCJQNtivrdLqFmGudF1pzzCESjMgTVC2NYr3mqz7
npRqB0d65T97UVbVZFqrpAtslsIZc+HXWxsE/qxR5IClssiUZseG/uXnCqxjlu1j
XW6tJYWjNzNmYlQfnuXJhqu5ZOFQEzY0OPVlhkjk5Pv7VeYZzHg0ziHzB8q0wojB
VlDoqJ2NcnV2nrd33DWM7JQoAuPNS10wPzFuNWB5V4Yl+Vilj6gNXbsK3/VVGBQ2
VDMrT6YN/xdgls8/nyzDeMrLToOch8cMUqKETI6WLbkLj+HCIsPNPFvuBkbGfeAF
hciC08J1vjhTn92/UcHA9rhGXEYJBA8BsFtoIVO/rX67T3ncvCUio8senAp2GlH/
4Rl9wtTZk/ayJAu8rvwKOUTC55Sw59B7tN+mrYgfR09Z3d/McMw0v02ADB1zy4K8
04Q3ukWEjo9S6Xo011QikVA40zjqZdFhHxTXCHgr18/ArJJSEx7gct9thiskhs+A
0hNbK2qNaQtlHnRGx2DzXJ7hUcNGSekG89/xk+ImzJldgM2CzDxAoktKJTZmlG4e
rn/dFEuTvktaa1xOBuoHBkPEWhjZ1ODNATkttz0e5p9jwKAzejko1eVDrqPkiiYZ
Yh0RMxV4ZCMVF3pGrzrylvU/WoK/Y/LSM6TezwRXXg2znZniwFvh5PeU92tOLoWp
p0TGQzXgejWtUsaTM0sTthWoy2X8USTPca2g0ivqcD57ZErpfQJcR9+g0pTo55c7
p3KoT/f3/O6jg1EnJbfGuuXrjHtcEW5d/dKc97wXRwI37nenhOTl7mtOhckZYen0
tZBnH2xV2zJKk3/WjKwgpdsLTttnqRnNsGhYcNzdz4fcG1ac5fFythC6ErjWsHLX
JDvTbvwkkTK7wvT08GR51lf68GlVUMAQqzjPZ3SjiZ9tyHpXkT4YBZuZ1OQCxVkL
DJ4M5lr5VUBXe5WwI8RtMLdab6EjHqrC367oldGOEBnAXG/96+2JTSX+34mj9jaC
c2PvTM7oSGrB8mKgyp7ZfAM/EKokWZwGdkHk8RaOungzdqizhPaQWvTJAj+qlSQe
iwzEx6wk/Wj9Zdd0PaZk9+au2wSCI0g/52yabIS6uPZ7DwGAQREbh4S1Nq7Dl2KQ
kJKD0gq+XORa4o0uW9rLfiK7ejghzHbPVoMXOPU+x0NEUiO7KZVpzycyfR8B9uOo
C3h1ezTaaXLUhtXmnRhm835Io3UApJoD8arwfoq1xyjEHeyyOUTlkl5W4YpHuJ0u
AeiF0cqMOXZVZzCaonixyE9g/9TApTu+U4lqM9rPoFySviWxvMXIoNo0HqjAqJ1Y
WY0diUUZpH7F98EQKNvTovgDowSwqYz2N7V51QJ+up/v9gMhHbwGLOhKcnaU85iL
nFu05URkj3Ul7KgOcnMjFGiHWTZuwfGlX88MhIXcqTid4TyZdw/B0c269tD4y3cE
BbQen9r8oXG36PwXWgXP/xkL8oEJXjUN+oirYdu6HReVd2M+QUPujbv/+kJG5SnX
vlA75M3BKb7dWxgko/xIP4x7KbmPJdFqLmyqR1JSMnL2Vs+UskZcsJTeGlP5kh4d
9Hh2BHApb3J9kwyr0f5RZ94wK11FchEh7VWuiZqGYt5ayzIWisnxYMt/v7wPMSM1
FwnVvnUOaP9gDXE0ZHr9hCZ8EuFzs0i1jiIy6WjSnz6KecxFqdbGdbrady7P0eNB
9SvxljdAP9Doo/74ESSRPoRINm1TO3EjpQkxJxlngRZh6n6gkirAWGgczbXZVfOS
Az9HU698Y4EEG4nL0VOmgKaYZyzk5/X3CjShYWBBb7Ek5vqkGtIDl4KYlj5EAgy4
h0ojHne2gPGYTRKNULi5qmWErngESfqpd4pOnS7MIWwC9F3Wpr1l0D/OAMrtm06k
b292m+ofA3RnHMzy8M5Hordi6RorDQfIfnscsyjm5x/Q00MeMORw8vY401wD7Pea
o6F5hfsMplOnFuvIW2nCoScEtWq5DTyseTHV3mjY9D7H6k9/XGIELISk/wUAMiOk
nbtReVTQbJpKm0Kk/BXx2DtML8e5j4egF4Rg62kReP7/SgKpWdAFD2Xo/HaKKXp5
Vlosmgwst2UrhEK7o6eoAdgm6A4wncfVGAhnBqFwyrs0I6kuaf8GD4h2fM4O/dR5
Kh4kH7QDJdqf/rzH3AovBBnUcwcrFFP/McDjBfOrn11hpIXfcLUNgZ0wd39JjJM0
q/WoWMmy21Kq0AC+d2wmLj/1C0PjsdqhK6Aszd8tkHgkNCClm5jPOISHdKOVGX0E
Lm3KpE91DwADlpBnuFu57621StE3aS3gwdqr5r1jLbrwX8r4UtFJS0PkzojENExI
w3QHAnQbtqZbRZPiysa1N5803ZhfVRa2JQo+VifbjiMTGstbnVnA0Tyn73chc1px
+bD59G4jDEpplMdoAGv9D4vzVlyeaJWTXtgZTfubdSPFVx2FpTYorFnLdKd2U+yL
AqPtXorsD+JAgw0W3mKytu+rdX6DOGl0i0eDZpqeDdjAEgW9vQrL1LFMlAjObzEh
xE/XQxMHodAbqO17pmIgHlD2G2uRTfJpi8PTimEC88c7URzTUQMM0fCMv90xBFOJ
+MSvR0JBBMopkTfhlrvyUHuFcdnMYtEAMiMIsi00ypIHTQQF2u4TeBbxP3J71nPM
i+0gY+DvJH9p1NJJYimQH0vMFg3va+bj+nz4OobzdVqppXGJGwBvmboDYvJKhSuM
7Xe8Y4bLXTU/NTdPey9B4M9FDSCJi8hp32b83K+Vi8R94N8f1cmaGv50xsyYK1ac
YCS7084CXHey0wUZ62PZy1hfA6JovggaUAqtPCLtgFgWV3uklA3Qo99xmiyPL/Gf
gej4okrs0l3FmT3OlM9gBa81SzIrSFpb4Jxvk5A+g0y5fjxghXZ7Z4Y4w8P5/QPE
qH1HHI+VgIhJrr9+nRFVBFSeA91KLhA+rs12/Mtg94/PnltMXfTT892Hw6RrJZW5
IDgeCxkj65hNIyoMGq9JXZgNEpjDUBuCECGF0lzRaTJxFh55y4hNW4IB+CDYJzuj
XKAOZOfvsQXy19mAmvrPDE9mkGZ42REePkgfDb9V/ZK3wAfXxqEIKq5YYQH0Tue5
WlAT6YBEM2s5rGAvHbJEuE5DniIH3+Ie/qpbXXbqcSkRBPn0rz3bbEpwwUWgtqMl
DhMnRDVB6D0BhZd3doO0IAgnpbqdOrYpYVGzwgjtnqWQvPaM2sNhWOeGFBodptZr
RThtpdzk8H+NEKCT8pUvRyyfm4dNSrXteWucYJTgPT11GabXAWsCYtmoptRrGo+0
htbGNJJ4J08iKlQezURoaPaaGV3PgllZ5HKS0CdF8f2mlsLTUj5AQhPYzyJhE7ey
zPPrwbFk5B8Bs3dzrog6rhTYZOdtFIgthx+UpHYun5MHv3T700j9kPmwyuNf93Li
VkRN8hXA47VXV6VIxYGOXgKgJaZXsCVqLWpWYX9I7aqFEJkCxLwvO+1WO+qTorwk
MQugTj+QKW08jAW4hcBkeAvoaWYQtv5UP/85cyXWcuYOusKxmMNBVlBBh0Hm+/LW
WNB7sIbab6BlX8MemT6OSvUN13enC49z225qVZJs4RhyQGOFkokXYYEkBRPGmHhL
0E505aozu568jVaXev4YeVBmRVECfQPUqAKLO3shX+COn7mGyAllwIq2RAhKnJEP
fHfiaQI7KDr/lhKksdjVqtdPC3ODQKhp6ELdt5lT4zly6NxbQ8hU7OvTcF8it7ab
NGkXmI+Hm1U1CrDLa6th35W/gujPcD0joRmgR6Sjdz2uHlt0iDvKiwgg1LGlnZjc
x7X2TySQkfpqHVM0SqbKBMIEed4wvT9xEyLQVUr+tWjo/qc6Jx+BmQsYEEgUvIZQ
BTOoJOBP/N2bmFrj8HVUzJEa/ugw5GkzmYdskmgcYNFW79iXWb8CXin1S/tew71W
uGSE7CUoSvw5DkHyn9b+f++fz9BwCtFVhr+F+jwNa5kLonsK5LI0hL7rg0AUq3jG
VTEH/WjNHhMQBLkDoQkQf1FKX92fJEIL4RkCBhG1QqKJ+kSluxsZebFBXUbrBOYA
E/66SYawBzNGxA0n24hKqP/wQgwHwbQvkuVcZ2/6zq1wyByhKf9p4JfU3qzu0vjL
18Tm29+hLaoIYByRjture7wLiAZgoDowNogRBjuIzcRaxax3Unjt3VQ2blzOrmqt
RTZrrhvlqKG7Ch9svBJmVgtghGfK6EFKIwb0NeD6pf67UkUFL9r3R3yPyGEB4Mhl
uNrni1oi3f1C9hcq/YtpD+v+B5Fjln5TKMchf7HORurxnUjaT6icfpasTiR3sxLU
68nGVtxiq6XQo1BrmoIylLqjmlrMPVpDtBrGpeMc94WT3AGEkahS1ZnL+uC4ymS8
PYJiWbIohxAWXzV+eaZBD3VwTCvjWOhx9f1HLF6eNJkM8q9dm6+kK2eFeMA+VpjD
zDR8qEVcCEneguhgVIstv/nTzJtsQHJVeMSmtQeoqMen/jo+RivQIy+uH7k/iDO3
9cHDQhXtAgsoEG/HPlgXKH28+odpsqe1aGDGWJ4kb7JvEbQy8j45gWaTHJin6KiJ
iMsOLfeDTsO3KpJCKrXlxVFPGe2JNtc/nD3RwN2/Ylab+0j1DzVX83WQI/UFRyl+
V56iqXvjq3Gh59UgHkKKTTB3cpFCMqmshNy+0/xze06ieGEDdcgbJjbYWz9sXg2I
/K5emMOCgRmHhkK3CXvyF1LtXubi6k+mlqVdPXCRuBZWq0GKMbFOUGbd/1F5id1Y
vV18jyr7mk7hFQ+hpgHHz8/zy37eGNuyWqZ8lh5gBl5kKgtv9VvNawShExL5cirN
Sc3JUE6s5hGPKFhhcrDmpGOhzsZ44JvVo1WossJmxlBEFuJXN8DVVb4Qelx6leH8
j2vSQegeutkvSkS7xBBMFhqZtW5smMyfyFgSL78KNLFYoRJJUKCesVX1ug+O4mJI
pjGB8LUIh0L5LGkWnIiu9qdx1rjq3Wtb62ajvbd7tteSt71YzlLu7R7ZNn9GLxM/
9e1tkRRSpFsMOs/Nj2Zy23dzwxJyod7WiOlEASQgH7Kqz+ZnHGWvpBDFaq427uau
HqTrL0cQbR51ap6D3rUfH0S/wfosBfHJ70mBIhq+ReOlj7R4YD+X2DgrF2SzT5jf
xGJlXHMJlPG4RzYCCWTPzDfAJTZpOOudHeC79/RwZ7XWSrFXxrmWecHcxg0BmT9z
A5Ldtp43CwFwr98U07ikFCz34nGcXDawca12kBHwyLhuVnwYJdyO4UElgKR5laKq
q1O1JErRGLW17n6WuMksnDD6yNa52YqXoorAwi+wLL76Q3+2jFWc0o8mdHMQh6xF
Vj/iK3Fg2u26Snno4uj4O7AFs6qh+7nfdW1JMvVy41vQpf9amATFsLeyEV5KyNWs
B1DuQ12YSQNIwCUZFoHpOcAXlgVxOnU0zlShU+MsZPKaTB+H4mUcOTnNmvz0f56v
zSD6f14SE0F4owUnk72CewTFGvCgV3HRcbG8/R4pEE3ODVVqriQ68Y7HuJOp5qBj
WKw+ltk6C8aZxYYhHwMbKxF2MGsEcvjzzDUMAerVNXO5joNGXz5pOK818ID1p+D0
Ql8it46hv2xhKtHT1awlTYBBqTWCeQAh2ZYQoVuDrVsz5cxYF/9LmvktXn3ILTC5
sWhLNvZZxUSft6yYGn/oHdAyGtbqq+iR/MiGjQuWuRgVTjcp57cAjSzk7LvppCxY
GfskjudKz99/kavTbbmuV+FbISNclRdFMho/28el0XEcTQU2UaZd4MOnUqaOF8jo
c3EwCP9Vjaxvzjo25I3tCVz4hoJYpO543CSbKEonWxiH0EBaGIxjxkxU1J7kKctd
wBvwYlznMybXpQ+PLeiJ4dwdqKAIM4c5p1LsONNF85JBHWCHvXkIHlwrd59AeHug
uCeLRS5Rx+fE2pVviNOcbw8nTEGxPm44WlniAgg0oresiL1N3B+/sejrTH+SNYTC
5BWlXEqnwKJooHEE2F3qpsqcCCvn/A24zGlghntBSITpIrIJJx2rfJ5XemmnhHU1
bCynnF/zXo/hank9+YyX8f6NgQsr2Epx7+/9N1k086D2XgOejLbHczE2kNOjTYHi
4IsIgV/SIS9KIDU0hjHK2t8psQbfzihVLJuKAO+79F8sXyVrHqzFIJAgNfbwb6RD
S42hPVUr3TyWOyZyYPbLGSNUTPiZCzYqgIpr7qBwAXvcHdX+OJHQLi16/LWud7dN
Nc6ym9wAE05SREvtRdW+v24vRC8On2RsX4zyINGjIJI74JAPytz1SpCuqOfW4hSu
jvuaCw/ivxaUrEzg9DNdiKyMkwcNAKYeCFy6CK/Cdw45hfPGbmtOA8tMKcBS5YqZ
zRRcflTud1uiL2xDPDhYoLCkKAk2ga6EEZmFXm9BdBhLg+ruglGORPqACEj3R17s
dwD8sWltljvGrIUdvotakXERu9dm93evGoqEOfya1q83al/W9g04ecI9GdcC14kD
n6oSmQyEmtdwt07l06ldJCLR+1Ge7RfIdoglLlSJQSc7bxhiYrnHvGP5pbcDs7WP
E62pxAJJIcCfz0BpN0vpVenRQ1sAw2iMX2Tj++mRYV+wSPgyjd8rQJKSdAzTBmEn
eNVqrkSyQyiqfvRbcYgcYyluAhdUxGNxErNS/bXkxearZCGSYiJAdh7a4jcbbRgP
N3pl2BYjSu2NEi9yczpJYUugu7h05CM2kIXff1gtUe6V5JBPz7kPfWq/ciB4T8YQ
EoMdDoEl7XGiit4Cn0tt4YIpjfsuGMGOJwxgbTDzBKaKrGSz6RWwd/kqfrumgVYu
zkPZQ2t2xDz+VBkvNjuOUQ73lUvfBF0E8Y8pf0WeMhlHoaLLvsGMs+J+wyqNEl1Q
Ch1irAAyKgRB3yZVFkIDPdof++DnmdQQ/vj0g3s6dw1AgIqxgoRH/wS6+eQ4QJ9+
BJyWi6Wq7AdAmdZW6AHs5/GakyrV/EnBLfFImhvUiTJ54qwiv/XVuRg0f4byIboP
d0B7aTueODIhfo9Dnf8+AcrIZiKJe8HR+PgoEJ61QsXOCX5LyqfYzEoyf1KLFGAB
0n7CBxPoA5gWOo8Av68nlgn6pQUXCWA+OF1Uk6WuLoOPSZtBFPP6lLEet4e/U3fU
SuAwVtLW0VnRLo0u69xcwUWCDuOPYPQPGJGOzcgdspovvPyhVPbPIOiGfipEC9C+
E0X7KWLhfi1LXVuwEsDFi9+DMNuo5KrLj8lchrkfovbLWwkr9/q7I3m62pv1cPfO
URZVabIUGaznLOAwu0rfNdqqg0+Kxpa6VN6ixBjJGQFgnlxPI+lWb2y5N/5ZlwVl
l9xcEnTLWOpbqlc8Q9bwd7hRVYcJ9ymE02KCcDoFt0uFw275jvQZo2tL1AI3FDo+
GZell4QYMF04wi+/lW/vx5GnBEPNUitzgZyZPC7pf4eTXN1maBcluJfLVZj1L/Lo
e2sxoN9BDbGBwC7a5h3isFikYRveKtbSRRn+duVpVGcHWTFDSuTqhGnvOyy/Qo0f
zF3rPRP+T9MT1l61CAipgOZWpj8RK6DLHhsRcubEc6Ca6d8gxAcKujkFs+DeB7Ho
9rzYdi+pne8Fp296FG4f8+fm0cgnNSS0UMnVlsZkpsnDMYy5E9+/plEvY7Ro75b4
NkOwzdTaV/NXKiLnPEBysMy0X0wTajNhlVdowyi6ekLi2cVAwEJOSWMJ6q+KqJV/
ho3rh6NZVN6OlCGzMZoFwkkjRg6H8pQYDtP57klz/b6itZZc9qJdmfqP+3F2N9fO
tjvnGJ3F+7gmfsn9dV3QY5C0QuRf6dBzxjrrK84NSZdO47eQ/2w8a+CTtEJrI5Wp
B/gUpNex9Mdgh5ciP58DwmRoqfdjS6hSANPgtp/1Tu8g3SoNPaj8XaTgqJw1ucVn
EWfj5HrV7OicQ/IBM11DZjBsykIhDpK9pLMTP3aLIMQmuUSwS/o8PZhCfr233BUM
qIoW9cpfFQh8DFm7u0JFarAcfkQhmTIjzNX+wVXpfc9mZet3ASElCXK5URqZIrTR
ZC2I5dLQoEhQmVaZ34Q2heOrQugcmTCyKssEldllrizDQfSuzYM2ptJJeJpyBWop
C4YGLGBAx43SRuaeyTLlgvs9XGjllFe5Myolnd5Oq+GDj66kgv4h7DLXIMuSIQvw
N7PdM/JLaft8tRwKN1cYy9CIBZXzyGD3vWEb0DMtbINjpBIY1C82++OIopGAOQh4
qJNTahgqm6Ob6KHLCdm3opq/gwV8Q4PG1D9U6CZfqL1cXfyU9iDpqidTzyohSQPk
AMt0RH2HJeFpekJ8q1pOD3sHILzAHjM4K4pt9EofqOjUAb5LjqhcWh0xZDpe4AOa
TkXHjcoa5DCBYOP8l2r3rDYTzMyykPGnFOi3D57CE1kvzu1YdgCV4VYHlSd5hf5Z
3bRQ5rxMrz4uv9elGjHe96FJcbYwxDJq/+/U4ciFsey0T47TcdJWAysVWRWULigk
4fsaeVgJEAwwY4gnqY7a2CCFXAOtrZ5Hj1qD07DIgf4M1+hinXKN99I5defK8cmu
8QCyod9tG7TqDpSbmwf2vFONIvoWGEnmkEhk+ilC028Mbicadq+QnXLis2/sa2Jj
n1ptHu4zQSm5gJD553fQVrPOKQAQQHD31Qcxw6Z2RfCVMOGipXN5XCdBrP8OMBwW
JBN379jxtRmVCtiy23X20UcdMdq0oJva90KQWl1dYsdAP5R8Nst+Ri3kZ8W8Rkbs
SnqM/w8YZ+o2g1xLtonv1bzU/OuWK5BKXNbzg8ibXGBaaDH4VRGCm47u9gHzw1fe
RILPA3Gyi/V2CE62cl3+bOqUw5i+TPtjEkNEI0OYBOikfPeaI1nhbUQZDsGxfijX
KMWoIC/L5M7mR+poqnsw5ZrxWCd10KsFKmWiBwiW8vaI9qWHzhJwpWPBR3Hi+UTO
oI5AoqmhQmkgjiL2GQ/fP7iVS4SCFEV7AZK9Zu0ImI52KeHSBqQR6mwi9Lp22M3l
03yXCi8zxDSA72OlZmC4gsmE1KaRDTatXOwU0eKYxIWsC/AsUISqZdwXCepSelCE
cR9D9NJB3JuiZ+2Ku5RzEFZamAoWKIZnO7uEA7P4mhDF4DYT5gtqh9xtwsL1qV90
1d4pnckm6qjy8ez+rtZe6I/tseC7inoCJHMv9xI47yUEgdtVN4p3uNTN99hU5MA9
ps/j9RagpH98GKrgzmHyq1cKD9AtCQMiMYOT41tFOvMSh65cZKpYWYgKdY+5h+Yn
ItHKp5/nawPFCjXzzIy3ZmkyBDqZI/mo8EkZzYaDCi3p8nfUEzTAm0ahkD/1rb97
ob45L/gRwYP7GO6dSYMdBaNZfH2hHx6rTqRfi3hDTL+MAknXPyCG7pJjOqcSs0im
xikBJeLC3oE0VnQqT5XMv15cDsSKigVXMuBl1mglWc+pHfiyZE2PtRWFBGoD4ya4
ObemF89jxqxX3WpRCXyb0bFae2ARrmzTW9qpUIYaauPbTA0HRx2mQ1aPBeWblKjP
Pq5zCwTZdklko8RRppOPthLh7FI2BCp/iSYIM+QGLObbZXD6sbbz8Wk4g3rb9/6Q
HiFob2DejXzZ7ACxk0lNM77rSuet1VwQAWksILI1qX979y7xezPyetc/AB6ypuYi
jyq2hxp++2zMIRIvSiEOf4ZUKPIjujMpQtVVu+lhJXFbmycAnvVQUBjvQVjwkpXd
tSFcGhq7WV5rZkKGV/cKkUrvdyBnm02OA4UihNetIVgipTHjuvodgS/r2Yxz6knf
1OR/t51g0FXyysvsyB37RrZyxTnQB5Wy/ow9EDzDcLgoLfgVDEwVyRL0Hb1VHL/a
FJFgvzLAnRJWQpe33N2M9y7cuQ9E6o4644FVCFilkCHnmR/lBMvsLjF7h7B6CYLn
8XZLW9HGJRwmrVOb2GZnWs2aKLp89JM3q8uunTYwk+wUFqSydE1intCCZxEKLJZ+
oq1Lw14poAC2yGFF6XvAGZtB24xQL/89TobT1b0VgbRgc9fd9EPGpCkIaXJrRtMY
gERxXLmB+iYqqbLqX8ZxuNf6EQb9IzhSikAQhIF9lWojjeYzuCZ3KNfZ2yaEvwC7
LLq9jbWa2sJGr/6TSjmSlao3j4vjkVXpHr9GzBD1QVty8y3P4Qca2zCeeCEHpGrS
OmxPs07LtMxtSZkNaiLI6aKj5bx7MEh1c0JZbGxmdcotja5EdVBUgvKnL0kb4XYF
Ykjp9j5N6LZlNWmp2+QNljcrOqxPCd5cDPEUPg0LE5I9B0z9b8AciK5mMOccl1Zu
bh64s5EaC152yUgxdlEmQ1AwyLMoqoENHOhkzjeRHjAV9s6w3cF4N0CXWiz+seJd
t71ye9sFpmaHJz+Gks3NlXvPpJAI5xYuWW7cNUqAKmXs8aESrD8PM8YZ8Wd9LbpE
fmbdPi0KQO5OhP4JzB9rZqu6NP8Erj2BlRTsBajDWxYYj7RaDp6ocO8JsVBGxFRq
gmuPMOieQx7ezMyv+tLwA3QTNbioWkqdIBhejxdRvOIvKc9umCdLJ5NMAqkivhnp
yILQLWDN3VclOeswl41eo7g86ub9jcSFekQtR5Zr3x8gs5xCrjEVccKFOJ1fOpzy
+7ZyS0EhIM7P2PSX9Phc2GSPsFnqOU7qXcv+usNXvIXg7BfR5k7L5FRcA0uoYWHv
tcia7Z+yUZbeIymUlBLKHpmcxGDLgqpRhbysTHS+/f+G7sbBKK1gWZSy7hAeuvG7
WJZHgiyiqAo9vbejnF2Tnu53YSIhad4HP4l+bKgqJuOVeOi92iuQui0RVwYJym/X
5l3wmyWB7LFez8GvNaN0+qb02un79ybFVWzY7DFVp3hIKsdgHEh59i1dUMSoIm1Z
jvlpqliQMcyInmS9qB98tXjRmXxGq3vAOpBkU2CY/FhVflSG4ImxeyRNqQy0eYEa
dKpCB7+e6/uzfGXhN6EloJO4x7Mlu5yHZEhaeiU9yrEC8NIZdrNTCJmbx6ka6Cvm
PWzD8JKwTPBNutBFq/KvwD1DYCtaGeS3JQZ0h27bM/i8Hnu3GLWucrP7+AvkTpzz
0PbsGkaOOMzjYmXONSSdFqHeJq34EINP3gBZjJMVYT/f25Eg79PcQgig1+xVga6S
TROo4TdfXZe+PzeUycfA6yajhGa4mke98kOZo3SPEBPFPGONf2i/vLq20gdrNR0r
Gd0VdpdFx/tc/V2GfA1jXVa1O5k5LAWjUcliLEtSrVh2kg85yHPsvUs8oPyiXlpl
4TrRD5CSTqemBKicHgFzqAKEMJH+8aaHLgFK2Lgk5M3AqssmUvm3VaX6W5qOnTtR
tqkwbNDeXgKNjzHXpbKaT6KaCHMe0TQwMJxrmsCQ0T5kwxkRacMwd7ojajIXEKWi
8wY/pOk4ZexblAMePBOYdM3UeANwPZPO+5g86ZHkUUKHkOZ5VRrLrQXB+nfsItzx
XQZE+aTqfO6+3Vc3medBOXkRMPVyYc8TsxMpLpsf4V0qFbYlLNDK502Sx8Mvd40S
mJKFOOuOusUeVqY3e2i88mjL7qjNKxVEd+gpxSgIb0tBKZ1PwYKe+pHQ089wTSkx
+zJEm8naSRUcjeP4I3nu8C/8+bOlRTMSvfCtGX+RQsbXpgvgQrpC+D590YjehJQz
fiIorNyzdkJ3EGeRVqEqK41zNf2eV0Pwd1p3QH8PJ03lI7hPNJzdFUMs0JL/FRrG
G+nI8Nwnye13e+0vFUzy7FRFlTPuVuIQzc6JspuB4NuxdxYZ2BgGWHiwF9jrmEE8
td67U0616p1EPJ3oC0tz9STEzP7KTkt6wOAigf2N8gF06zo6xp8QvdRNfsGCB3LE
iAHoVFM1/PS/Tm+ypTH0zvbNgop8D0WhncIyu2/V6ty3SYSUvh9vTEecJErd1O1r
RNir9GbbIDG+2mi8ZRoKdk0ETPzE7QLVv0BC/beX2xX30ER/R4ktzpP4nDGdcEks
yFjGGRI2NWFNZeIwDRB6fLZhX26+XXHSpUYHQeTg4SCOKA9GNZQ4T3CfWN16wsr8
T44jnLQMNpFwqWFhQu2emWs2v2HqaQB3JxNdVQ6DfDYX3gd9f0KdyfI1lAgoFLQ1
ENPlMZBSHnRQN7XI68EpuT6vgfMdlGiqgLp+yjL004aO7nDwVNQAdOdbjsE9YwYc
ZDxFtjQrOmvMpR1AoKjHJaT6wlFzMkyUaaROEG6C5nEK0RYoIWCCPjimSrkEA/0v
NjYoYSI1/Pv+9uuu2XJ8LxjbYjTxMrYh5PddyECZpoHcsLGnrS4XIzjlmD+Zm9Zm
1rDJ5RdwlsHl9nRFYC7Kuq+QALy81cj3DArwvRvaV3BrMoQCayIakS7nGdHqSeOF
nsG+1rgPM6p/4IkEL2KjHpQODg1rTn4uZfTO22YYmqG7f8lvtwa5u0dUcnR9b7XA
PY/M0RoW1lFbNvci606FYnCgkfQ/m2+ADEQT+EEiv+QNR7hGMO1LmmbyWCplcjuH
KnIPUCwEFm0h5adr3u0KJLyAy9Ww1oEXSbZbo295nAzuJE8fFf5q6CvOQkVdkNtO
6DsV5BoBIiuemc69TjaDZikcTIAjUmZ9GpHPmu84EkuwQasm+7/laY3pQzlaSlZ3
0nbbfm90YE91pvMwcplk2cJSEVTjOjSbQLMH1McxCTML4NlT3RWlJiSoRCAZWXh+
dEkS7wpHCfufbCiuqJ38u3kWJWI2kocmU9G4Q/UZ5gB2kd1qK0K3FiQpXMmie8Wg
rCabFYi9uxLs8ks9j4/pVC44XDNncghXgKeBA9UdlLFkWIwfdzPyZk001efMgUzx
HfDpFGqYwB1bSetEtkQrQqWwDnHaJlTmwj3Nlj1x/DCS4LR7TpQe4yt8dvMAK62b
sb0LfOYnx1djDHi0VUV7g7umPJc7McOS9qqX0QaS6hM8f5/MxIz4ElN4AXTbIgqn
EnmXTneRvOOCIXYGMbAyccVB17ERcqpeCQoyORZeEABbUhNq23ZtlrXprY2gj61O
2hQ6BcDvthYpjMr3eCRfjE4JlZkAngqWZdjQnL2wR4hMhYlaWkTuTfF5G/z4zHpz
HKPRwIsBebbZStyi/7WfhEHUEg3BC2yILvSAdRMW7gdjgdUySx9+xJCm/YY9TIYg
HRn9u37MsLRXZJsv4wzaJav+7vZN3xhV6YGXWAZXT7xMekfVhVkUDJ24+ja4YBCO
TSSQB9jor52Uw18+MDcwq71WwdnSCRtSmUKwpCsPorRyfLGTwkHHiYzbgQjZMTwd
aQPXBjvN01bNKCrQZF7AFHqu3gUC8lFLDG4lWWcSl3wGpFSeRwWzRRiF0Pt/SbsJ
JRcwOIvZzfzx4ETWDZZlzxndB5eV+NX68vez1Y7ENl+SekVx+cXLQLyq6DwKtF0f
OF924gi0fy1V9Ey9tMUgHxsG1wV001XF3B9lTn3ZKGr3766PTlPTNdkWKc2gel2f
0ylv2NcqmF4T3/IzQOkERPEL9AGLLFigC9ZW0UJbVG+AE9jPxlh8vE4h869DmgJQ
JEH/of2RwbyTr9y25SQmfrT3iSOp3mzYvKzetcx+aIJsWbtXXQh/s0fx+S85ZRVI
3oyKf4zyiWg2GBHsRC/wU07JWKdLNTYd3R2Z3t5OixNmOHaA9ztqnvauttWu2cBa
dkb+OoccyTaQB06CWpTz4ENeYMGBH6Q7Wpiko3WZAhv0cDWTYZa2xYCtVb4SkXK9
1QMChviXshm2FRCw3nnNvSTxuXqAqWie46TaVqrBYXhkEN+SwyVb7KfxhFgbICgc
uc+BQRmgB9ExaUWa+nscP34z01MOfCrkymSNmeQPZU7ddHcnI7AQb+afQTUnnEBV
j5bo3CKiti4SYJjwOikJV6n00NU1Kq3dUWClYJMiVJYerKrjvM6b2x2K0RQHph3Q
U189Sk+ouEdMAXNF8LmwdSynl4iZRex9MpKRlj+WSNRdtduSpfn9TX3iHY5C5mTd
7hdF8SBatPWOk6PXXiZCGBUQSFjKTZ4sMfljxmBpADGs5bdyvfFfASrEhjshqbtn
Q0DwtqzIzg8fSTUM8AzkXqrVBkDdMtMlEUJ9FsDtrWxwxKiuVeXlf2yduxxy1dU+
eGBhmGi0ZA12KvVRoWW/XdhT87l1MNQdBwkwDDJbXm8aDi0PcefgV9UFH+WTHMG2
+p5Ry/t8JNELdF6fBHpAHPPXejDBmHhv25NatQKCR/TZigXA5oWOmyWovBcCHrhd
+emU7tDF3g1JHk6SztnOj16wiTAXn9lhiaBsaxUmcz6F4pB7ci3Y/bwB29SN9Zgw
ROe4P/x1vUppnsewoluapcfMPPr1KVj5G1fpHVuc92KJ8pakA0ABomjnhTNMaYap
4pbws/eR6HG+qdSaeLwtQQrRmaWzzDxf6HNrJLvurLvhvBDKWCEJZkpCBDCNDhNp
jOm56Fq06RXCKX9Ss8KdIMDV0bA3GsOpwjN5vYlff1m2SBBdNTSzyL/mNakV5c6W
1FFZOESAQwwtS2wC8AwULY4psYH4gR+h+Ksy1tRIElBWg+1kHWOdWj/JeF1Wg/B/
vvzHXiYd39894d7bSbAPlhxFm79ohlv2hdYPnJtVLpBgyhIwEzN0n4qgsFcNkUYH
i28abOUBYMRRlonDUZgdhFkcw2A1sVDBozwVet3P8K+SrXZaK+To6ySwY0A1x1cO
WT9YhKGcOJ6BiFaUyby/iXa0piTNHSCPnhVVSLiofmXbq944y1Rvakeq+tutDA0Z
+IQgp2MGnMvBDHsYzGBEKm5oJ0NbLIA+pMMrDp8Ew7d6l3xcx3T+wZa+audF4SkV
LaYAuTNrDaXyFCA3ELoVEGIJ4mSgomOQbEOoDv6wX8n4Wm0ofgPkIKbzb/vX0byj
tfYo175gDN45qR87XJk516NrFJeBN79x09mbPkrLmFqKze1h06Z9Kh2jfV8kgCoi
DX+yvpzJvWHl0IPaOXS1kuvmNE7NG/YzosgGTQHi4QFxbPvZxXUOaeVVuYOylfXN
9Jh1cqm5PTAu73OhQhtteAKxgRVcLayxl5ybpmY0L1GaNlzNOZvH3RFzUldIDK1O
p8GfzCOG1A65Z2/I/QVrga1muQJMavylo7h+Jn5gJ9uAfVnJgr5BPZkx304s/+ke
sC/BXmBH5ryStP4o/bg9PSVJ+IWsm80ePyn0ukRODPn2b6xmRob0KmC4T/xfPkFV
G8p0Qgc1/rWVjjnmp3bKuMifhU30oe8XfH2IKCYaDNu/2EDJWbUTbCR9sCREv2Pv
qX24CERMFe8YaKIVyGULtItRJJC7gUatHH1isN2SAYErU0xpRnsCv+ODuyRoCedh
458/Rys8BImfvKCAU/SB8zdYT0Vw73GIuXNEHctFDZtClzPQEapseOwBIgkG32va
fOAk0OH4CtcS5sPdbA52C7Imki45WfqkqonMF3vBwITTY0NPdEsIQXSzh9ze/mdM
5ihatg7MWiYqfHl54kl6ESFTpQSwEGa3hD1MHAtj2VCkm2x0pmooyzhQ6QeUnhV7
BYYN3bxW3EM29cM3pCgkGlRAEyGXd5gowexPLBe6jOyxr5UV9Me/8UvCjSpU7lXu
Lwj50687nmZvGByqtzgMCr0cc9qHVNAIpUZz8GteYtC4n35C3AjVTgn6GnQN1O5a
rWQRg9yH7P/kjrAojgCfy2YAIyWiX7gzFAYffU3Sq6Lb9hcU+pg/4WOR6Gae9vNg
DoEi8QHdZ9jyLbcOXl5wYSpBUKgbBnQUtfRSQ8ouadPcIUIDv3gxVZ054lOJsEqs
GnYUQg0pdBrp68KxKzvNiTugdqrAxLv5vRyyud6djFRS9qEWACrQ+2P20eRpNTDC
wgu3SGvnh3QgIWlK8F4f9foc3f9EdK4zpVDiVvefiFaXbBfyh+Ef+5n5hf3IofCA
0/3Xb1qfIG3dO+VnwpamdCGQh/vVrQq0XsR+2j3vooy7iJzAasb17GI6EXZGBpUB
jqREDh/aaWdYrbwO+kw9PiG61kEO8ed6h23rkWvim8NmfO67U5Y15dcKXrq3ReXZ
A3+hwFZg4C1mv8gmW8R3A/fQaTyYzC4SxEOA/+7xlm6MYbg/7Wvr5c4aHAEdizIn
fJh2wtiaRFbo36zsYIHvRIAtT81cNwSPbJGwfZxOM2jldYxzf90r4g5cVbxpGCwV
oyFvb3uGHM4D4iIE33DWRYL8s1cUGeXO9EQej7ifUMIrSTmPBSnEZUO1aJfDwb8k
1Qj0IU3EtJZa3G+Cknbzb9e49MNsLsiVMM9g4526EuoiM1KNDUxZUipDCqikgfu9
vjqiaSW7UspP71gpW7XptBlHO5P6LZ4DkVYaeD+6JtNyi6YeaprYDKFhkS05st+h
5nQg5PcsAhHaVGbu6AOs8B8SQQureKf+xLRlQ5Pm2fonnGBdSp0mnDiGlKQrslFp
rXEIEjQGW7mdGcBtMbglCuJHRs5txnyMkIscaDd19wCKk+/PiOCPEMm1V4Kt0zYC
qTwibxdKiThtJgbAzc3q1b6BRRb3wjGDQv8jkZY7UppTcKYdg2Ev7RGbtPP8glTo
MlhdkpDCF3pR/CDDjVYyhu+gNU67wZDb2klxTawJHB5orMX8lMVNSRcOzGWhtE9s
7w4xCFh7wBGP5eBJuJYBg6py5FogOairE5Gyd0sZPWYBA/qp7Gvk9yS9f/vu5Uv1
P23iFqhkvTXCzRpGs78Sy28hctEbR06jf5MAsEjaWOjN+DdlaPBFyWXHE4aGr37g
bzMO64/TUt4KoRRaMpTjqccJSTOv8wwjIzHZXQkGKUE2pqD/FSj/0BpQII1krezX
s88nwD0kPblnWVY2BX0fyVDLHShaV4f446dLyjtQXjQ0X5s51sTxWMVj/cwINwdI
WlIIYqiCIfUUxAQdEf1YBGEedgEj8xezO19oiWADy8UWXDZMnOuoaF621XNgjVm5
EAAkWhf4WLhgxvRYDx1S7ELTGGVj6w+KnrSDp0mFtSaTPKP1GPi9UYtcmUyDXPQh
+ed5ktlnKNrhTMF09zJ1ESYYUhUhWjJglv69qsvacgzyXKCwyRvhIZJZNytueiGk
3weI4l+V3/SlF+vojmLqeJBfp2n3InNsYwRZt4GKN/IFpQqYDcA4LQwBbgQsbquQ
SbCqKOq/lFv+ij0b7Z3ZGHGeFOhCSZTXuXZ0IFUOtEA904nXYierFcyibFpMSxQ6
1zV6WNX3O0dU6g/1EtUSAz/T8nSOoDsWv921gppt7BcoSmtyzviqGdgi75Cc7ztv
D3lWBF7SgiygoLVJCl1XPf0nnhmOxffSPLpbK8GGX6KHnp8xhWezTpIDPG+qnAkX
W/QQJZwBVBSDBXNHE2cC6mvBOTLjFFpe2gGpBbI13n0+ekAZA85K88esIrU0qSDr
GuC9THBq85wBAGTS/e1XX6nFRiZ3+Vw4kxcWlqeLIRak3RD6DloxdJNgbyiZRrSG
gX/5/P/9yMBCD0VtX+OIdQb+whlmrUWjFlSkNIjKHHOQ43rlsdrbV0HT7nWsBxGa
C+ny3mafT7LtbHv8R6yH4I6SRB9ejduTvGFx4u8iDORgfu+fqbbAfpopaxyRrBQL
ftB4pueNosPbUJEQDZj/j3TEH8+jBAbQb9cnUdHIcSp41RIM3Tv7j1GK66qpKolm
DMV72uAUQmxRvt+d6CZPfkSaNzMuA55fvs5l7kVRK9z/VbR1bMn6NoTp0+wCvwRT
trRmrwpYCjLWUr20CpJhAwY7tGx/Gk0vYORcgG1H3NL7idIZIZAXWDa6hBn8dGUu
Nze56SPAdoKy2AR1z8NAmHveDZM5/t8JC8e3o0DaBskKB8j0+9CGwCMNiedveMzW
2PSJKdt06mlQngws28nVOZBx37MDyUVpseynNFJIBYzXaEV1jG1zSRlQunTYxuix
5H5V4f3RzouPHlXm5gfhY2BRd5ExbOBxLKuhxdXTDd4HvMCgJVf8jdppLoQSGSw3
Qh1lpKBqtl0O26gyChmbYNrlNmcxnQcvPlSp7guXI3XEN33RholT9c8vEx6mr6Iv
G4woPrbAq+yPP+s/piBlmtz+rllwBDzpLN6RvfIY/etpcYd5OWL85x85aQ+sXyP7
A8nIB2Upi9BfirAwwsgsH9g5IwoDmnzOiM3sC9GgxDVCvmwILos2jCwRH2PIkoK1
23kSfwFJGe+PeVCX6RaG+DasErXvHifK+cu/CxsJXGKUcqXNfK8cpR9/+zXlT4lW
vQWHi14bKTsuojgF2r65kJ5Eoo04E2Qe4rMSkUJg66fN2lOiarKBN/Fs+w9J3V3N
ycXhvXf0ZAcE6prdNOVBcG7yLKMdiqdtUtaJz4+dcvbmhWE8AiSiOU6gg7QfOKiH
BIlUMsINoxd+copMPtB0WbZW+k/PG12Jg/V7ldjIuq9xj1wABwWMNKY8nhpPLELe
J8m0iRsJyOuu1wLteZpMuaMZzu1XQkjyOj7RQG1uIOmyov8uPsaxZN1ReerkVopi
PCcFMmTlgCeAvGJcOeR8lj9O4z9QM3FTy8ChAiiax5zBxb2OEFbxY8UWjwWUQ5em
Lmx7qNIjCwK++4uk8vaNMR6H83F+1+R0s0aldSiHDBx8j2rFt7Aefl4b80FU0VQ+
9Lo7R6EY34qE830YQ7Hii7a+ZVmZ6up9T1OpYmOrQboefErx3fbCxg60TvNY97Kr
EHHHKAXgY0PFnG+kNDz3YxcO80BAuaV+JedwljJy6luv9lQccoO+CYlRgaunAZqG
l1vH9Q9+LTIWdudaFNpED0JpPuTIv4aE4Xu5DCyhkppeJN/QfP/VvLDXtG18HH4t
BXXwjFSoA4bvlF5rQ0on9qfJUKNRSipgRtn8IqyYjnNjlhfE/M7bowp8Q4woVRsJ
y3HUNivDKAPohCUNMDAGSDGZ8DTKnumoS/PzlfvKGShvnBTgQ0hQk1kyBNyAYNnb
fKC1ii3uc7Xxv1cnctbX311IHcfYogSMjTYkS2m4BXqJAjaZwufLpHXArpaUDKIO
wftVy5pz0kallq35SdJlP8ug4UD0WbyMD7ypil7Ua2UjEYT7mLK2OSZML9U9c/aa
wN+o6dANnWCq4+J9Tms0yKpQXpG7+zrYByClhGOOuOhDApwHRUg2qfEF35jtGRCA
GNj6CHepXaXhBseNAfGqRzZ/mZuG996rRxMVWRS27385wUluSWttd4VdVgajnu0N
R4pUxRiirMRy9Gq3JeSmolVIgxNsyevLuwvBr5L2a6OAbQcGdDyPN/X0v5jQLljL
ZbdFjYvxEnaGJe1XEWzbpUTIHdo2ozIjZU+ao1FIXvZ/Yo6d0Ui2k7wbnnfYuCTz
YY0qtKmvQV2mTTiowlhHnaTF03t2LrLjU45NIljEB3LcE1MQoHdTZpcEZwEoGEQG
UowYgYC7bpLNdiwZqXhHH2R/jh17J+VVpNBfT7YsJZMaqysSYTzUIklVZdwjAaZw
7gySc1URr7+0qnkU2UfOylSM7TFAZNNTkJMgKeuyh1zWMdNr4Gn46VVRWgtvJIv3
fKJ3K6dgQPfeylQmRnzHU3SgbMYb0Mhceu8xQi/gj8riHK3hojhoxzFEb7m+VS8V
8NDT3PgZu9GBf1vYxao22IwPtCWPsOmJpR72Cencezwlbsi37PYa1AOEyII1Gtwo
bXFxCzLdJ1zLNmCtp0eSvDxUhAkwtWWYLOtdblUcr5HzdUNo0Y+7bDWGUpCpuyC2
BqphTegHetOYbaNOavFoz/aazDAa9r9Cj8wJaEQeKtOVBaTpbPcdYNiX2Lqso8Ad
k77FEydsrDJI6VgNPxGvVkiFHMRxEyIKLSBvF4hgYbxM4Mfo1QNB6X8ZSFcX6Pmx
SoP4faQ0SiYBndCdEvuC3IOSOJeNrSuzBqs0JkbEM77SEeiAsz34S9IQoBLNoY33
K5H48hxGqIuilxnT5IVY82YmMDwj6xg9Qzk7QFAMER6W3AoOeFHSmK3GmVn+46G7
phrB+vCCqEeupgMdIGMI4CxHyw4Z2t64CoLHLJaGXeKXEQDxwKSYmTd7bNxaKuC/
/vhc3U+8XyFR0omWLZbk/vThQDur3fBpOBEE8u1Netn7TNgzJZI3jec0gdN1+j5P
qeqWVCRwp8f4gmjO9bkGADUEXCYWMy5erk7phWcqTWHpUS/c2ftpWqaVME1SrmEC
cwnSRKSH+BT6lvx/X7wcnvOhB7rBwTi034pyWyvbkrVtoFcSwBmBqwyU2TkZLVl7
JV9vjhzfUSOu+HywpB6m7Ut008M9XXgOf/qYOh3+qhM6psiFqOGk1119FQQuWOf9
3SHAP4wR8szCHaaOsEadY4PvOiXyntRMw83kIhvN4ZmXDLo1r1b0s3U/G78c+UH1
5a9wKzN9jkVnVnDLSF3l6plRCzmF77CsQdnFQFjgg44U01OeiIbg62wxE9oA/TRL
EEwSIHs2mui2lRONwmjuReV47p3npXXaCb/FoNb3JptI3dpHbDzylZRnOjLWfsaJ
ZPktXBaBcLe4oY4/Pw0Dr36Qyn8Ih2IrS0Oh7B2EObSqIcpSzThBzcw7hdKv3MGB
VYW+DFX2yi6OPC8Ays0QnluiaCKxCjmN4IAGYL/y7tNNzw4O+Kfi2OLLYWeD0LTx
47OQmoJktHGjiDn3vKLvzRvEWb5M+TEtP4XshsOT4Rn30U4qBhcS6geOKDJCL3IP
svJpVF0kQtJfLwAIW6R7yCZHIsPYPeJ828hMMeje6J5VXGzkMWhZ3VognRxql3Es
peUUaeGnfiJcMTWSX1+eTymw9grKIrjKKIevVp795icqosOS590Z8KVbFATtrqt8
1oyqNPU5M21CXwtENXh93KRITjbQ/8xBMOJxV6xKfPLfuzx6A3/9gLzxht1j+/JF
NI0zxQIymxfSOPsTKa966/+bbe9V0HMjGeiEL624yFndlzUSH62wCldmzJrjjA/z
Q+TNPD8n4qPtYoOWpEvLMLzDwFKN75+j1wmSV6jiLpE0ryPrIaeOWjYtg+6zdSyP
Vwn8zOXwrnchLkRyHtXnFfH8z4ERUgMb9JC0TjFt9Wjczd6xi/GrZvtDXnqtKCGP
7OdqDFxWRxViOdShKdwUQ4nTYzaFEXypSIzMsxo2EBIxq5eXAKDlAmZ6b6ue+qSu
kGB3JtIfhORHnvGUPYDUpsARtJ9QA61wduNgcUzAVTpbnAzbF3r18PzsCOwMlQhJ
M05kIJDtXRbBiv/QagIXe+c9ml3o6G6GxxTDIJ8gk1pJjM2lvCSwvF1/3BzTAMYa
YSYEgaG7JIkiGY5yKhGdKPJ57KCv36mUXRYM3iC+YjGN1yxYdEZBGggYY9/o+PBS
VmDoNayn3AT5otMuFa1VjmS1i1C/2DqFLQw8iH1ZmLssBkkehJKtv9GOFo9hFA4c
QjnMbgEOg9W9P2Jciov6fNmm2o8Q/DXkLaP0WcThj7q0mtdGqVKFqKXj4e7g9Irj
Tu79r4A/f9eogzDlL1jwUJCmmJ/Qe3pPEPba74CHYVicvyU+xDAqbWZ5tYBpWoFQ
7qeJpm/fyNWveu9n6R4EG3wqsCwEAnQr3DpnPA5GBI9wOtXBAVikygf16DiDWY2j
9gmBN9KiQqtfOEaTcgnTtbfFU87QMjyykaGzPEBihcH7CgJW/WL3gi71Xk4mEUh1
Ifqw0c4JCsVxY3OwcUhJENXH2F79xdXF8cAUzB8bqRiy5dMLSN+0pt0mYMAaOlzF
lv7fRvSr5RpJGOGDb9NwWBI7hyj2NMcTNOwrUAgkJgJq9HeeSkCpuUBcQui6xkV+
WxPF/aJUa5ioCPTRJ3zY4WvjCaucbneNNZFb4v2zgg5sJ7MBkO1kQlj3J0p+4GlL
ZlQrbHbH7Y2GEltm5nUrzXDEtEiGqRfWAt5TTY8Jt6OxsP9JG+1Cd2FHSzAIRobi
msoCX4LO4ZEjyQ0vXa9e4xLFjTcUMQztePnfAoPJXVPzO0YgskcWA/gYE1/GTcd8
EXJteAQ2M13fD/nnhE+kuw6mx2eM26bI08XekDriLzjkt1aGoLapLCFjTdZMGu82
aQ2AhhXdzCahMiKVNbmDcN1om+U4K8r/4zb/CYospJdlFWwzJXtJqYfumNhQTa2n
lrTUIzVMHLEAD9rx6IoHt0So6W7wrjpcu+rRaUR9PKc4jxJ/CXmBPTt9r1IScEWD
19z2/lOVheE9Ulx2qW+Q83SznsN2fPml+2dD2ZG2og+mum313eqbdoErrFzJ9X+4
XtW0NaxsuxrytiGABfd4Ph0rZgAIXgCAz67QVTDbp7Bsyp6xTMVd5CFBuA7sNt8q
8PfyGPnphkAZjhu5KuXgfUtwI9BIi7A09kUzCRLAMv5YOEiUouM6iWkxiVCtCNW4
qfAwFq0NfM3WGqHWFUfVAOJ73lXXXw2S+PZ1JTxVDpElXo5bzWQfrA/n8bdRaiYP
vHHIhk2NYQ9ev06Q8Ah0sq3MaSaAQkW1GxM+yNzPXFzhh+Aoci9erb75EK1MvJOV
02g6WN7pXdm7ZC9D2EoDTQtJ+xBMc83Gg0afU8r2FJVm316SKEfDGDm8d10sdnpF
GLp3QDb51xhbSGjmn+VQFCrceIzcCNY4ZGya6pXhl+doy1A/w4y33BF9ZzCoSFms
dRjTmWG3IFpFNlNoYZmqwMBEOE9mFu1Cz9GuR/fQnQtwZRbmiKuuBaZSbXDXT6qx
CU2N+S2Y00eaLOqIA1M4Usd3APtB6mxvFobU2ovDpXQnVjSfZoq456zAzy7fq+xQ
YtuoVH9Wdya4YUrdOtxv5RE+BxknDgaktboxroi2aEccfJZairyejk22UNp0vUuF
2xvg5FPAwTsTc2Hh6T1FaG46/r1IzFVPcUZuwO4GvP2JNXp9g8+o+w8HRqh54xhB
RlVgvN+Hkb6RXvFURdJxOtOiqy1SYr5BvOmSEClRnjENfrKsa9L/3G99gyKORbrA
96qoNtJz3SEulG+RxAs+XaCal7CwK43Jf71oR2VSJ5Ek7le1kNyZlaCqaHVI1bcG
Yq78ge2axQEFpigUFbDqWj7y3hgCJa+T7ShYJsDJXiS3AsSvoQ/0x0WLVpCgTV1m
2o0w8gTaA3SmaF3A3GXH06n050gC2N4hfDoGSzEJZyoAj6wFVSQUq3kiO1j7atRM
ETGqfMk67Q95iYP73HKP412J3C8i2HLGnmdzKZMWm+qoR3b07Py0OiTlzZt4ILZH
Xy5ClofAwtVgxweTTQ03ogkcCE9NWqVfOUYywCVxeii5JeITcRBZKe8sKGI0cb/5
JqMsiGxQBvbwn56flglr/JgZwjXff1MU5SdocIgzTefihO7OAMTlPaeWV6RF0CK1
8lBAUKj8gEw2nA69ia7F1EFkX/YAcpT/dRWHZRLUn1vJLK41rpQPwImDspYjN4MB
dNF3VRcOXzhqUxtf5HOkqk05XLD5SdjIX+Y1QDOrgujs/rt7cSQOYVlscNq2OsCd
2QVpMoAm/C46re26DC9+BXfWhPC9eBiPPB1ttOcRbUxB5YR9ipJsn9WeyCUsaeE7
0c/FqnSlkAAFDSdDQZNTrw2WqrzWTJD5CNxICkAOU8a8t5u8n4Bo5l2/EEDOq0NA
T3i3FAwBORKHz8BzAF17PCZAvRGvzNW5chmoOHmja5fu7RSoirgj19V23bU352P4
R0ik/XsXDxWWzYI3uvec+7b9BcetR7jhJ89tVUrjBTuWd1NKoJLisFVoQz3rkEjy
k3alxYpWZdkKDKt7/sj1SszcjBwFSSPrF1jrMKNpI0GGFT/vZaZBLTRkY9C0JgFE
mdOnUCV7tpN9hvWeuA/Fd8e6DBqSeL3OsthKfeygMIuoi88zgo4CCGJGA1HNwLlx
A1Pmu6k4Jo2H3zUiEErC1Y1sIK5DnUstnbKBhpVFCNIcGPK+OG3VGHeOWDoLneLn
eXuKq8AdW/s8SXqw6+EQY61xcGbYedAUVOH1mITpsOtJXEb9Fdl+O6Id0wk2bxXX
0w4K9hT5PL7szB8ZlgP7xOe/qW3+xnG4LLGRbuObINv1Xjb06b3GXqsh1cjX7ECE
asOIWKWwDbzNSctBSPg6Nzfha1TsA9m7XplLNEXFq0B59Y+x2Fen8PuOHleUkf7C
WxvV9xqx/bSUS7BVtFNx2l77O8OyQfJ4OuW7IHO0kFmJi/862h52QTU2I1egfv7O
7MDx6/edYjl1x33Z5oX/P8phl0Z99OGI9iKI8UyCJAND3uH8d0TKFlBZF5QP1BLF
FUhrjyIEdC3VMaKz24br84FqbbjJyFqTZ5bIPgyiwYa72sBeNjRF9ahwXte1uMsm
bxJqG8b8BtNCcZ5qvctv0upUmiHhYAIUjtIrc2+LCNaPZd7IEtSdQzKYGKUwohw8
rgY6W/p4qlJi2XHWb7wQ1CB5chs+dz4cZ2t//814kOeA3/Xv4NVH9WtDbN/yDAqJ
RfCBrRKH/+V6/f3I4x7KoHVuYtIDBqRjpI95lUK+KqDhujAOiCNebXr6enAFI8C3
Was8k2ThBA/6xup+WBiB+irYCozZTqrNyFpfK16G2nhocTFI6zg0vqEUA8Gncpwi
5xZAgAzuCvV8Z+MEm3VsVO6+MyHzp7M4L/LLC3a5gdWyWzABchjiCPYx812xEIqg
O57rAYeIg52u58Y7tGa1FrzZWCUcuAsXBS/HcCmCvRc/gL1RrVgRQmbU5rdfCYJE
frwvO4XCs1uGpR/TTbNyRv0XN0E8Sss6xd+2AvD+B3Vk9FVyFXwHK9m+qnsFxip0
F0j7uxFTT/Fwq4GfGVT74lxcV26oaP1uJp/WdYUZqfmrJnHUOEwMoAtehk1ClJ50
TQCCUXWEuIHgrdDpDbwIGurmuX8uWnFTPpRVpaUTGaeEvEevb0o7Nw/E8HeYVSx3
l3WfeILTQcz5IfdcBlkDzTdJ7LPIa6ux9p6yij6tPU2UGC9e6l3gfAXRwIj8Lb2b
Xj4FteWUDLsA56w1GcdyDTzTOnzstA3JLbXwCTkeO1WlM6TPlPzkARhiFt8Sz1LT
YJW/6P4CV6BP0w5QolpdPV0TR6POSZrJeivMJpW/LSH5RYY7NnKVGfUo5amwQHOp
qhLYIOq3bgaQttn4R74ylFqeBDEXEEBNt8SocW9/P6xe98iCwsjyFTH3Dd1wSr+f
EQ1cstYLqeLaTgjmH5Ffza5wQQYBljbCZGSdsb+Ngl4U41+0ivlw9ZdZiEwe39Pn
qgbYxPc921oTuecnJxbvygYG26O3HJq7pOWojWuTogXQAZZXHLPxpBi2KUnvBFML
XBclbD30d6skm19x8XTLUu/eKHe7P5q8kHhasucyP5C5zWbkFLu7/h6vJF6+tu/z
3euYLysk/HSuXNOM2wa3qUfq2Fokmwjzc0dbTx0rG8u86Hka/Idq/b3mw1q85G3G
OcxoLuNF2IVqsLG8nwpJOEdX5GGjFYZ9OBgoe/j2rP2dXKtdowe6MS+v/TAuWW7x
h9J+4bc4qOxhxhfG7DvYhpA/G/ikfQrCThdFdtx6OaSMBY9n+35UafXDwGnUE0Ol
UVMB89yK9JU54q2YBbXl7XQUs7zktsIEG6ENkCg2/2xHRxQE4nFzaKxTo++HwZbv
uw14peeqMBl50zNRa7zwxjNx0Nn2AjiQzAAW/kRvsGMFePMFJvTO+gJ/CSatAgBw
qsSKJnAlTCHJ6Z2IAS3NHngWLPbv8dZw+oI0yD5XjdQKZofQLiTiNMKtZd6hNSS1
XEKpB+63EGWYueIgc2I5LVDcuz4aaqg2G9KmQgUMo7gH8lg+ikj/J3cEJER9T2Qv
RcfszZkXDpr71cX3nfOMZI+yI9xu1rsM6JE2qyEnxuPPahOWt428/B9yFB3ibn4m
u0eNwphvVZcaYUjjrWU3R3uDetYz8sCvKyvPLgZrQVXU6Vh4R7aA/TTAT8KZVJE4
3vxvcKOotPtNQ1bRecLtUIPZw6ZSXI/7kzVq30UQ5yYD6jwP/9bPxytzNXSpadDI
rwjQ+fTBQtr0WIGps7wDqGqW43JZChNXf29hrqgUJPRWYVflmEYEOufg+U0CLtco
SR2GNJPCkxAN+DiZ37u2MDUR7y+EPZqKp3t8zeWgNV4IXnl2i5jJg/guPlS8waLh
1nQb7/RsAB4j6DB2NEcfsQq2lYU+D8JW5H0CX7fLN4Q59Yz1Et5h/aL6jd576PBs
5n+WY7IaBSiD+ls2z5q9OyM0TR7YVolf1KlFKEM8G6ZmueCtseVhjeqwrCWpfgRt
eMDot8vdiG2b54JdUVxpQnA8CcluGtqrRnceJI3vSXrTX5YGSAvmPm1RvuPh/eXX
TXkolPMNx2F6Ptu3e32JwkqKdlpyO9uBq8R7hFva3NvgI4EjEyJnBxbIPehr6C2D
m9YrgaMWA9BEVB4uDOhpAvyCZV8HZcgqfBVIQKB+i7NPLpk+cjlFrin1VWLzGwwr
EUui4/xOwmgtBEk5q1+EmstQQwv9hCZ9qeupwJ8lAAQ7mcmzu4mWyS7Yca80+6I7
TysVSbMzYilFkEC3A1z1I9RYRqstqasd30MlsTRjCQx4JXIqryQdjWgzyn9dVwOt
prJPLXW2ekoKYorAZmwirtOe294PF8hh239OBYsHS1JFRDb3xQf+x4Vele65H4l9
+3woOKHzGIcTSKupJcaTn7t/5Uy+pG7q7F7tP6F3xInhqGuoW4eIxAfy3nqlCpA5
dr83MJkw6fdyNAKPKifEjyE39ATXbzi7GaK/99V4yuWhGX0oo+ywqIahhyaTJhdy
Inv44N8Fqa2CTsJHPi4dKlYTNf4/lOpxEDNVbpsz/8Cs2r8IBWqJpfWcVNrM1wuC
62iQ+fJexz8zyN4Sdjt1xwoP09ld/I/YhS/kOpGuPdXeVWKJBgsdqdj/w+WFGlDn
juQ7R9bYLyUVPGNmY9BXsbK+nUmA/jQeMhr8jFB5AG3Kt1i3XqdgpjJxOKlSWchO
a5jiAeSH33Zk6KOPQtcwLQm2lPThLxzYcEfrO++Of7+Y2kM3XiktI2DeW1trLzD6
hCV5XWBgmRL8QBLaPxvCWbSuaz6vXnwq8nbkCgynMee27wmoblWe2qlIwND56F7r
WDnrgHohUviWGZTIQEK7V03F2797mGjM9wSG63HL4gnNIdwXdrW3AeYGDdQ6d8Wq
9XWwiL+z7mOM0Ah3VIVLw6ZDUyLYvvinfMkUjYi0cOfVJRuKoy5mzoMqxoV1UQni
rz9celxzJ41Lqmzg4aQ+PmzBqPbyHk4N0UxFcmdDs5YS8XkVkCdUnIiKydi0zofn
Zer6mqvHPfJn6nrvIjZtD1KDiGZk7Kj9xMGPOCCy57lV+tsYTqi2l/XcET4mEabB
aTyzpaVpc52peZ4kC5G9gMr0i+E5OvUetxKCUVpqaHvADlWnaUSpMfoeyCU2DLJ/
Hr1F8owkEpgLiKaXKRzELJu4ysAz3dqg9q8Tnsgw9eWwjV5QmNfrXKYz6WESKWLp
VJv9e/3vZGDaPaoPStoTzhTOzIOMgolw5+aKcIztVjNgq4B7oeH0KhLkerO4VASc
Mz9fnn+31ovDZOypKNM+u20cCxymYrZoWG0XvvA9jBIs4Uj9mIEQWWanBvFNjbYv
FD69uUVJaDvk+tr2XBp/APWKMAkV/1MHE29zcKdlmrDado9peIVzZid733wA166r
WVsd+kXkCMLk1baO+Tg/h43qeWSixbiXokaIpJL/90Rd4MslnL0yXpL9tl+ykOk9
W7x1p6lWon6v4JLVwFqtLP8fKuYnHUTjHVE0Q525+dxM6Kcfy3YHOaue7V0eXV96
4XeJuSvUfdBZr0/+EZVlhREUgWqjptnZfHrOKBzqncZLPqOaAXi+jkYqPeCtXjdM
4++mt8V7BxQQxIoDR77rlz/+Z5VpHB+XkMgApcHXhxaNzSqE6mZNafK+KGBy7to1
InsXNm06B9jQbFNcwQq/kh8ULUKLOE742H2EL9B60Lp/QczSCtnec1va5h2R01td
D6m2mgo3ntBSMDddTb3zf/LyjwNVJX3zyhyoPKl30VacpnLdcAYL5ve5EZEe+LrN
d8wt0OVpLxyn125uFWyMnhbjXdAkSDJRP4QRc815SFI+K8urNqfyTL3LH1R1238M
zMWjd7uDiyBgOnHquS6S73qHbcbn8WSyjsVUJWK2g18ONYV4qys8x1zocmRSc7Yc
rX6Ud+BIlWcgee0KfwJcEcP1eMgQdRDp1V9SM9OzyixYLSjtVfACAth3byt6Ul+W
rTIrexrew4t2kSV3IiQmjZvA+a8epFQTo/gAEboXkfwr78K1g+84ZXcdrBSt+IEZ
pvUb6jruN+JqyPe+cLQqNnqIN1oy156VpjbX/mWV69/KoSMfBzwCpi0eNGmujPdg
mr9KkHbE2JKEGOQ9uAMLKbB7ciS9h8HeXb7ybk4/AZss+nVL1Fu3z3GFJAG4Rihj
Yenh3CriXIRh2wJ3D8i5imnMx/t2eGqSIoBQ5lGh/b76elNktTthTuYGkiKOK/mD
r7u7Csfif5Bz/IZPej9hFb07h9o+590wOrcOgi/kESPKxQ5E3Bu9uVs/Dahq+sh5
uqpXQ9yX/VkbfqqUZy3NnIX4y7VsyBmb55aOXB8Zfsgwl83Gj7VREHnup0X787wJ
TrG7ENFV5p/jQwZD4hRMAKU1A2YotU1elDCp7d02T0kArTfRCc85YOfRmzhCZ5zY
cJxcmXaFpczZtWNH4LnUWjP+jWVf/qtWuZt+JnQRejpRX5zJ8wAjW174JFsr4iVI
b9vc6QnO7e7lrKeXWTJWYPs9T+ZJDuoLiBnIObqgmrUi3bXZw4AsJ8klmwVjRMZN
LWmwcEs3nWJ1kmKuRgrJ0lh9GhwkLbO92QScLHo2YWlzJezuMfzey0QKLxtbqvje
nQ80I8yJLAKGsjgl79cvVpL4h/f93b0rLnDo3FCu/y4PatFVPVCS1tTf+XYRGdKM
nq1DUb6xn3hRAo4PDNnBTlHyWsCoO1n1IrJqxnONToPsD5RpViEUW9TEPMNP8mwh
AMMpG90haGTVDiIvCNzZ1wLHz8MK/oN3k2OwmjKebrV0lIFHo3fx4TU3la0EzE3H
hBHBB+ogduPtVNMfRSPyjqSJa0lrGcOHIN1RzdSJC290aQ92gTLhjF/mYnggNC6m
Tc2eOz81QRylPU2I6nxqgqjFMVO4ARe9Sw/PONuzolYTZ+JZ4/BVjqTMPism/yx1
PYT30g0WPwM1m375C1JfF1DeU/XlgECFlOiIkCoGDyflv/GUe3A1HtB79g50A5I2
3aDPmI11Aru1aYza++r+nyyEfeDm7gEvz8yC6nRwmbXDvNykJwYiPunwMYqsraYQ
K5dwdjp93YHTCmeZDT/1XHe/m6m3ScSCVr9/5gcWUAvzBTGUR6mWLO0ImJdBeFKA
ZY+UrV38L0Wxg+c4bIwNiA9KOXcX6Hvr5mXd1YLUnEdKQUW/iyqgMH/ED+VVGj64
xpyVCzPdkL31+87u30UcPc4T6LoMA1UXxhAvMOO9adBN8ojXhezv77Rbp3ZKHKa1
BIN2JUaPeU2uxyKw3JBiSplAAXXhvTYjumiFn5CnjF7dJMPEWbzcsR4qh5Ou3efX
ka00gdADAThzvjkxC+9bK5Z7JcTp/QLc68VwROTx6EgjJYWcNN2zg2YbAbfum/ec
F+KQjMnkEupdQ1XiCXhLOWFwYQa4y29ZrNznNRQpXznF0Cr4GMuhFjlQob8mouaK
dTK6Nb0ItcXEDmbdeRTT9tF0P83WbEPaOFUUyASOb6ugHFtBy7bWI3f4hrnL5EBs
TLWs8t+X/neNcYkY6vaAMzDSQb4W22RFj9//jSPly9oelMf9xELEUM3oFxSiaxet
1Ye6IVCROKbKT6c1//T+3fgaDdM0R3FW1VgQrgu1dr8bklGLDjprSRcHjmS0bsOL
UG+gyiK/gQZpOHuzsadbbJgQtNpjrdfftetKwRalEkp0hEBy2kNRVRv4cHEoK34/
7TovMsPPzSTZHWGKLA6VFUZ5dY22L5kq0WKkiFq7qpp5tTD9ZCe/K2rF9oKP+N2q
0/X0un3SWmEKioY1FD9+ZPO/xzk+qA1FP3t8X4044Hc47+e/qo+ZaFsGiDrcPDDZ
w/ir/ksL7PAoyqVRtB0SuCdMQEPHUcYAZ4XsylL/OHATu8+1WcmmPnuSJqBT78Gt
OlafljO1PM92QfMwP6f1YuRj0zQSJv/6oLwqEZxdRDPwDngyFVV1ffun4b2X3OVr
7cicG6hw4lKN0Ue191Ou/HBx/pb4YyITMFPvpJV0mEjbcvSm0xVl1LIEX5IeNREX
gcq0wDMn/v6dR9xld1udYuwTNaGxJXSfNjtM9Kaxd8lzkTrG4WN72allcujEWQAB
vv5Zpd2dw2fEsKzec1wezTsSior0/5rs3yrt6EIUmxMzAvyRcsSHHpyCqJQkw3kb
VaFfbfcqYCZkh2lDBzRRTq2hVkJZtmLEaTILhP1PIF9NC5zyp1futUY0jZRL6+8Z
IcTtIdOkJLJnQR1h5r8/bjLpFh8+aTBLBRQs6mieBD5L7IA7OTtUu3TDrFEHj/uD
LHaAXQmc6com6SdFRsTq+bbk/3fnG0zyMCgPSfjoUhiFqM8Jxx+HmlRTYwsJcHgy
7KbdVrGSMFM2lVlnxYe6T2O30ZGX6lKGzRSCpZlfjMv9hCrG3eVrG/9fNSZ1VzIe
F5tFyvo+5MfqPlo/QKQ5UT4V8kLJHiW3rGFlXdIo4bl3OsDc5IE4/kBZJisuucvE
fm9c3vIe3wFYkK0Eoi1MZbkGmIczJt7fePHzO14qRoQUl2cMwCSaRinBhpMKwH2S
prtF2+G30ZSdtlpD8PWQBKhGVkesBWDD5uSurtwUIjMbYEyTmG6/zOWkZmLBCVJ4
+0PfTac9mxKzUcnoIGfWkQPcsO5NYIk8Qntt7cR5gVF8iBTD/QsbLBbiyPnx3Sdv
cwdNyTSeUu1oLfz+7T4ww6tyAubA1w8/n0ZQFlj6gQXYPfzOewcWZrexOezWorgj
T3KHlJBhyYXGWfonXCjDhgqU0RAr/IivN13/JKarB3qNoCQDqcaT80JF2IkwsBVf
SRZgrpXHAgk+nCAog6z1TUccAN98nZQgRtv2sfQu9rqd/52ZHPPyWzF5IBoA5sKr
9An4yG1Eze5cUcd0ycTcoAJ122ZEAWMV8McpO63QikBYVrWS2BdYgSyPOwpo0CbT
FaxGnz7Zv7Dlc7PQcVet4vfh/+ykJVwtoAI37ko9GRNhVFGxJp5/uhWs3llwXl9B
9bZlwcSLF7kZ/SlbQEneqyo274cILY79069aJr7QeKrM1eCj3bwBql1OHcGGAmp7
3qJ5RJG0j1SPNbF/+RzTwCULRcWPAYsmUyWCoYSPoQ7WGdFRPYVsl5i+1OOoyo3c
CGeT/cf5gbQT0I0YK4bmKjeFu8yCAc+QIivOP3upYgcPn/FCK6TvxngTqD06xR7N
YoCrhVv4xmw7eo/0OUmJFBBmOmna51neGgckxp+U+0d5t4e1QkTCWeGrw19ObOky
AZiDDsNBgIjfj72wWlNuFvzPL1caztrt+kjnyupocnjohab/32wsdPqimMNSnWbe
FvXE324gfnGt/P2GFNy+sKOrYsuuLcP3coOWwqqvfnsLJcA4zCQQT2EepP+8o/q+
64+1LLOYd+zrR2GPd+iQFOKc8p3CweQXgzZDdoSQNnghEM1O0f2ylTlUgxeCm+7v
YAeQPdn4Vu9xGA8ITsTZgXpedMgCq2JZJBQCp7JzkLkc8aoa+J7wErAJaGx3oUlR
tMuwxx5VFMwxGV+zoJbEGiA+kBQhKFlRTtu+aePwk8KPMNSlFTPZaaQrRw6HCyEj
e5P9MxzcIDBkNyY2jsitGa4BYlxbYpYedcC2BAOvFVZkXz92AHLc+xfI764uU6nW
k1wGWGl/RiwEYzEIh9fAqH+0r1Sb5k5RB7v70zBy/Sxm5AlQfxsJaV9HQTAG3MFj
ITrh88bjVsgL1mBK63ox7tH1qNI6IZo9dzJk007xLjjhMVswv3dVyt1G/kQvD+l1
KFxyWA5EDDxzrMMZFtcCRnwse4+NeZ2FqQ7qGgT5xrnG52Bsyi1v9WrxesAEYMGp
RHh5FugTx3O9dpHqeqhJRLv6LASzd3QUN7r9NEZ7Ezj3VNyw8UjDwJ/jj3Yt6RrS
hu1TX77n1RkfAXwMOWT0EAiqK8SZCEat9Ix5bMj12JvuTzT5ZdLE8fhLdjmJCRXv
3zud4CyVTMX/2SN/siQx6fRaxCi64x+B4/Bll1PUaqio78MLTq2OPUE2awWz9HaX
T1xhYFEhcdsTfA6KJVxSf5mYB8xZeTv75pZXT7M8NO7jO+RQLUypHSqkZp+osCjA
10dek35oQJ11bF3x8g7iFzL8Jq91zbV9lRZ9QGxZOVh7mj5DH4sgNR5zL3WTrQj+
WPWt/rqndc4FYw9S/uLIF+YTrt2nEXN7gVGvHM+LTcCnC12vLkecjow7oVKIAsHO
OBnZWKleHwUUdIkqp/rZ9piDqURqib4tOVzJyUhWridY3c0yBpy7tXupiMlL4U43
8vwWeDStbF/wMVltSf2fZeSQN0bjuR6zbq87m6206oWY6HDivbtWQ/dsht8FWmlx
70N7BAfem13OPSVZuTlfKBJBhWJMgss2hy0IDkkdRtkuFrXNX5JcYyu/6puzTxRg
Ddf//xX4oUNR9erpO4olvQHNERyd6CdzLTiNG1huK8vr8s6ItuLLa1yETia9mP49
yGrjn/JTugXjiPYsq6MlNqnCE8a67dkYLgH8BauNLHott7wE1JEFBERfi7WMihMY
twFOuuS1yA/uNJ1TZro0C9iDaZZe77NIT5I/MHOJGRz+O4cU563s5sAY0wXBswhz
WkpCDaprS2awOv5aeCAZ9S751pkHyFoAsAWUkzFJmWH/nb2EY3rXDVGX/V0RIrqm
6W3qkVmxMGakJ1tjR3VnKY+qBaBNVkEoBdcmFchttgri07a7hh2jX14aZOhNogST
sxZlEYjB3LlWrjPaE9XAintN1wW6racIuRPSPGLrdE0ItKJ/1qMRclh81Dn9gePV
cuWFKuzSOWu1ggEdyO7R55kU1o3OnbPeXahm8AQVUkUUaaF+jGU2V6WVXpAWApUO
9rFdcwaW489THtRr+ozkFrWA/32ROJ4g5a3FgS4XFeq8zVJ5zA77CtAOfXQPCyEG
JGY+d6IBsrHoP4L1SAioFYTebpwlqbQPEHMFksfTAPgqWIMWf4eZ8ZTVTqEIZCOG
GNBsDe839ErTJ9wiqZ6mjMOLsGF6gi8oF172mOoJ8qnAB83mQErxZ0TwB6BGRQNu
3+yvnJRxiLkxQOrjbtPT1XIFHdwLofS/jFs0Sm8AVVn2UmJDCsB6hTAWLZgRvEBA
B4rH60peboeWt6xaO/gos2QoLpk/yL8r0kqjcGlF46dDtne2NNlmEeLcRaLMv6ek
OaK/7q0teQrI63q2KM6ajfNUGXSE0RGUCfIub7XVIvOqDzrIwN1JzbI3KjIN3e9K
khZd2S98BwhoGUN2yM1UexNjg6yjsG6NDG8InuNJJ5NGWnsUzh8QAvhw58cB/4QY
/weG518EsjdjzxqYuQONeE0zh8RX6JPYkhPZCRUU92VEWWWsdobgzGyzTQkuB8ig
1yTC6mx9G79Ui6Lhoqt8mTd4bKqaguyO7U2XwtvY69Wv26PwvbSlGrCuPGrSEj8O
EZQDo7bEpzFOncvEAFxsI8BkPvb6FJgd+S4wcSZIe6EniTkmxQ4aqBMAJNPJDUdF
MLW9pYTeupOdtaPMSQdRnNXGMpWIpqc1F06qNTIdtyLWyUTpP/GaEjTsDcdtsGQe
/ZOTuychjBMRUEb3k7QLIi5861e8/wG/MeJy3xZVY30YBl7JK5USggqDOejhrxsr
iB05lv0g/kGmjJDoO+hzXJXXXbyGiHDrpWrDyflYYCtF/hsmDWla8xcXTJjsgBA4
KVZviUDR/UrEcOmC8GQCGcbsXoPM5a9QASKUdw6bB7rHnEee58b0bU0VyVvtfZcB
/U/HjymomA7dQH7YpdkFC9wr9dptWD0yj9C9ilWvytcyf6nvtkHYqgxPDOLAi/tU
7XrejkyAFAOLvwIyB19Zc8z47xH0augKAbT5/q+8D+9fB2xmSHzznw9uS49RuoT/
y50I3dhqzEfY8bW4aRsCuWnc8fv5SMyhU7rgTppEMQyuvVUopD4FDVTjmwGC5H0l
ZX4FAMsT4yIjK8+cSjDkqu7rdjm4jOYI7g9gJNcH79WJ5lszR+2vKuXHqCg71+vC
4T6zJpyLXwsgRuINP6d9163Fg2h9JDvUGI/7ipXqEjwqra/Qc3Qyw0iQMMN5ib61
4MPbzyaoLuEveFNl8ScwNfPuX+cF7kHqu82sMxookWNYoZgaArCxetlNs1AjTaEq
7eyNBmqEvEtb4OB5ahqHXxR4JJZQ0YEXrHeBwJsUawCzyYjdO/Ou+z1/cVdpgMib
a9wSheBL34cOdhrxcIsRddFgilBEOg+sk8FLNg42U3Al+f4v/dGsx64sM4tGVKWk
`pragma protect end_protected
