`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h93LiVEBuwAQQf+tbb1wra+kUd+o0x6j8Q++ysKpJ0XZp/iBmyNjOelmlWvr57Xk
w+taqjYeaMQPcFI3uT0WQprsbqQoRxgC4BEoZtxtmZ+ZteGb5PdhULBL6jM5DulI
O0ULSaFzDmrC6cdG5JuPH1q9XsH7zr9MI/aSfj1Pegc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22480)
Z1qBqjWxQ7rih/jUzgQFhH3Y+lW+K1JE0l21NTeKubVGxEpGfEs7wN+3aYSf0Npl
0MxGTPAaREsDAihtUEu9Gc2jM7Pkfd0Gt50xE62ikyZXytqz0XfXbu+11bHh8lYt
BFceag5qHmgO5MNnwx/HPWQVyK8/D9xD7HAuWPhXvC7mAiy6bZ3swGFMoR6X14wa
QdAq/35BmSw6tmip0GA+YcvXz5i0+UsBw3niCLlKuG07mBw5CSqsOBmXdD8dktXr
QtZf0HRHmHkvAWVvXKyQnGSj40Vd/3vMnyVNjipwcPMeYjKzz/kufhIjPv4jzfW7
wJbGwQsNb8yuBP1PmdWVyK1UCYgfh3jyiUTAn8o+pLIbhP6gcZu6xuh+j8osFRRs
IsfrpCfArwRds+Rz6MtdeZ5DZ+obsWzMEueIp7ceCBoUkQgMpwe6eSxr6lc4nsSO
AwHMTzXYIb0/NKingIFucQ1I9Y1ZSAzq6wvcROGMP9NhasMGMZ/SAEhORON9iwIP
YbOOwCkWygroaTHwDXiK68ZHkzEJ7jiK82h79NcsFwwyVAEwDxWdsJW3lB7AW3tN
KFuh+I3U/NLineJpS2q4YjN8w5qX0PO4AdjfQlB8IxoilA8mTZfRhA/4cBRNtunQ
M4auun2C5kSX09AStRKSxn4KofZ7xWkA2hnB354Akj9u2EfG7C5VJw8kF0DJHXwZ
SmrOtlm9THQ6vFPquVfJXSpWZQd8HoZtg74jXoB/m7oUASkn03lFosu4E1TYI9iQ
JICVUvgb1I+NDYY/+onwNXN3+TztaxGoZw2J+0UnoYafG/6tqk9nvmLNIvCe9ooN
AO8EnxZEv+AwDNzWSpRUIwy45QwdIYxmgovLWxMaL01aQg1f107rahF782GIkDUl
hECk11TfyzktqCkkTs8Z+lx6qWU/6FH8CePkkUT07hupfioJb1/FACi2GUNLrWC/
oVIpgaPj8TeFjUcre7SsmWM5SDiA1R1grGrt79VzKKdH4VSTTw/T/i1jUfTqHAyy
NuV+EsTIjWAoiGhFLb4V1Hln20PPOUXz4FUrpV1goLWQOYVtabp0TCx1QbeB2kpP
M8r6bdED5LfiYRWV/z7II3rh/lZak5XFDhUCYzh8h9TKykEhzG8bj6/ZMYB+UooT
zT13wmDgn03eK9BBFqLik83K85zZy9U4nulaYRMVPjkS+2tKi30QxCA+VjIHsKne
kwJZOIFaFNazemrEI9mh7fVvrlKVa2grPQTVXU1sf6+Fj86+/yS3K1lfsarPf8Bv
VlDC+mlNcxwxzJTRvBQL1kxfxBUz8qA972CzTvZlVzCZaKpXZxj5CaKPwkttjl8D
I5msx8p+NdPMt5Yqf4/bV3g8Y+0/d4KBpd1km9s3VxgoLzFSxK7u0RPh9VaSMetK
jT1fRIcgucDWUDL5KJJC35ot+iSLESNYsklgo85ltzT5rCg0tuBUsJklNBwlGFEu
wJ9df6399gkSJpthw1ziu3yy77CrrM+DURGXecImhbkbsmSH+lmDScTowP1zHGGt
fFpFAnNVwrwGRwmhJcRjDPbsoJLx9C0Y3TUrMUGpsLsVgQbSKZjcVXKVTsumi3N/
2VPaJOxcOO0t3/IZeRG/LugAHSSGm/hbyU10avpvu4DdsHWtjlujFtS4crAiWpbc
8Wup1pxqci20zDUlgxqPJ4KAX94q0ycECo1JkRhXiqvx/7dPTJ+YtrfQhnNZIP5Q
iejPgORyX73zK1Wsl0dguCPEm0H8GIscIhXrDVsgyo6Wrwsljj4riana1rMO3Wjh
kcItdCbhyKV5y2Q8BfNl7qxK9Q7PECH8/+LVquixSOx1A6r9JoJ8d8H2rKBWnNCS
0INzzQCm6sk+Y0WCjBmMiJlAm+TyroVWjTAjP4tOf/lkHtFvKO8gY0A72ShH0ncN
QL+pN2jjaZa2yRQkr3TxlaeW40wosk7K2c3UhboZtyNfJxywGZG0kf4KGM0QHCcX
baQVK/DEeChDEwJNeMtwm8sUHzp5+EU2LCiCHAJPERtb6VqZunBC3mOFZLRsOPov
7pawV3qcqhPd8nTUKqcCbhPYf7Iz5xGm7zeoBWi2xzjROH0UuWa172SazA/lEaEP
3Jv1G3OeHDg7/t2vRAbgVCiiVY2l7lLycLOJKSfyJC2F5P+F5HvRFtQKSDT5+8ac
f7W58EKaWCmCocEbA3Q4MfApU1hnN98AE/H73+1Yk4K4+t38LeZeQndk5dKeIHp0
LC3Jtxp1W2D1dTp3iFQb01APPTJC6BnySPN51+Xk+9my8vaTMFXDi3U/IjaEKXIF
oJWfCjsZ6cUI2vde/4jZjcpqTifp0Yfx38r84PhwpkcmMxoMS2G3d9CNpwd3xHC/
G2xH7KQcKjBCyb5PPi0bmwD9RIAIsvl0n+K/9uIMoMB0sZ6940/IH54l/Gco+zOs
CxL5+mKPuidF4SsnFFNHB11jMhXRRh3Ie2z7YF/hBrpFlEBOqNsbPIEOdoPDuy5s
QMj4FrL1tzRc6LANnPDNrV/FDfvjFcIxKC33xPZpb+0qH3NzML8unZsLNoybCXk+
f+mEPfx8fgHjmKoSUvmKEFU+UrUCae33JcymbjJ+cz8NVzyfMq6G1BN66OWLNeoA
/KJ4qKOM0sBPWskMv0QNTNb/ZO+r4K1T+tKYXNAteZDIb8Pw0PRKactUMwmsf+av
vZqBPBy2VntJrCT6NameBKTcet+/K0yVzU9t0sx6Mffp3UT+n9wF1mAJmcjnU8gU
m7c1jdVR/5qkKKL6VoyluDmOm6BfgEqbAQi69tmiMG7V8Z+r3hgwW4m+ZPLR7drT
15iooJM1oFKS3WYYjNnG42ZLkepwLzovz2ORi/Bxx8qQo9HLxKUeZ1RO37VMh/5B
YFPaaRxUrnf8arIhpTuZexFEb4J4neF2Ge92KWY0dbSW+2FmaEUvEiJNme7v7jdy
K2Vg5Gh4bGapggsbdnPiKISs9hD3E8fyOfA1mwQZzIuV4LU+ycObSv+MUjNDcMhz
vDXkIVl0w7nDSDN8NGquitH8J2284jhZXqbSQ9MJea2ZOmzfirCVVe6muVsZaUuG
mm3B3lKCRWEmX3CvgpMsRTp6XRLwu1Q9A+IGqSK4z0AjaLeJLyn36jKsSc1wnC1C
JD/TnejPjKMdE7F4xRtvlolUVvXcromLIhQAM0q+9eJfnFFFeFErlvnocaI63zYe
ZKGGoOYgFtI7qwoO9dkgAPoGN1nA0yeVOHkHGfOpIlXc0eOK50Q63k6xHUM9NI7Z
Xvuyn3mrZo7On88g+FV2WYDcsyO+UnIYI0tqyNy9YK0p2wQcfr/rlCeDY8OO2Ib9
aN6XJrm4lqbADm5EzIuwI88098HtfLcSBSTt4ykVA1BEhS4E+VD4m836pkfWHwLs
d7e8Bb8OqHTdmR2WKLjpKNiSDDlIdh5EY2/bjtKIv9bgs2/CS40CjIZF2bV8oRX/
Z2VQwaVxCE8pCx2WzMj1/H8K7KkX7H9sqavHuyNk1OB4wOZsOcLLsyDBlY2YKwiN
iR4Av2b1tvAYDg0dftuUe4txuDfzxTiNmEaOuELChVbVjRAyn3ccl5HzHis2Igyo
aJmox3tplc7jTFd825Pt1tm7nrErxPMI7BY4paT9p41Mlnd1Ms/IRuZRCMpdUh2Z
SDJpXhOQOM6rJpa+H1czJk6nA9mHtdFDQpz8fMo4z/nPMRqEU3Y9nZCU0i/Wt1vy
ichqBGhu8VXy53A0tXhAZ/JpqfvN+dX0geyR/XB7uhho5lzeZ4GcpA17fQ+2uSDd
/KKm+j+vJQwKrYm88CvMP+ExiZvaH/uPy7s8EFLgbHgDWy6S1ezj0O2XW1sssU8b
xkG2GP0/C9P3a7yHDke99JKQt1SdO/WQg9L7YD8XoTgzvyZWHeTSHZVIfkguGouK
84pa1Zv9GO7yxnF+Z+/ghpIPogcCa4ykmcPkkwK1JShWveNeuBoi9t63TpI6Vhzo
96IeTfBGABfORapqC4t7/hFNB4PJ7jSQnpjRajowEKkGdXBFCq5wy/rzGVKif8bk
XsqzoNoiDGGSnRG53zbH7XbbKtQil/8MGhEbSxFiWZfJfIhH8Lqi8ztzXJKMVOBA
4d8Uijxgc25Gzj0Kyxha/FJOxfx6RUHRlunT+dJ3YxUqMXsTvGOo0/pfIl1x7Ytf
rccmGqbSMozBh761fmc9NBekj/oHzmsW38imH5l7nMUXjs+KmxBIY/c55oJKCzRn
I8Yw0YngL9XByOKM5rRIvwmZroqB2iixOVFpldnRut6D1Dmn+piSHCmfBE59jS2t
G1LHvL2U9i5nmY+khsyj7wi/ydm8Mi7dCoQktw6yLAsGjiGqycaFYU7u2Tu4Ntwe
i7rF1JpAF5vWHKk30CrBC8DB5cPt5QzLAHRw0iWWfllUKACWWNEBHxvPeP2xYS+P
T+9gp3rdA/Xc2HVi9x6Vgp6iyY9dS+UrKyI16+UuVsVpqswqcxuXayIZbF0RZ2HU
5SJ8iA+BQmk1JrhQ9txjK/oknYsqdbC/DUWnepMk60kcTYJL0u6jg7XLsi4SAMLc
yY12ZyoIaO+3OuyvhDNdBRrVGBbvOAK9V/KhEpil6ANRDe9uttndni0q9rzp/Bxn
hKuGJlBiW668+FU2CCNMuiyNLjYZepnNdTzb6jiJ4nXZs37sp2sIiVLGGJ+TPH7+
A++QPZi5JThKOx9upMIbj1EPHbHS9YeyFcG2yX8OggTwgWPGbCTPazBcfUKQBjs0
LYTIhzFrOsdz/aE3mHSlNjac28RDTmV/iwhPsCiMaGmkxqUnj2hnYHz6o0EA/HPr
2c7HJYX2Y6x6uyW8ca3WrBnVkWQq19+NOo7jdiYAXPZA3LUMjIveEulNWo5calwL
AU6qesPlPRvRu9rnAG89gaUSHixmcl+tWgp9/YO8aY4h4OysLJbofs+I3870hi+L
Ufkhk8GzUBmWMVjX9kle5WiMpWIv/WOsA885jrzO7K0n+DTie0okzzsba+IwKozK
NgyWyBsPEKC4/MTN+kS27IdImm0CauoGrbcinusaMBAM6v1q6mgCVFW1FAiGKxQ+
kKWC3m+xa0OaU9WJHFI1JF7w+ag4YezZtCYxODBhDPK0eWAlWEwn8RjMh1Y0c4q9
vWR/PlG3ztC/j4I2eCYTFFqBuounUQhqUECy3WMzK9eABi5OfBh3BpIGqX5da0OE
fklzoSGSg7mEFmzkTDhv0GL2aYfSS+cQ4EcMwZC6auF68IXBQjMp7ihnv1SnbpAl
HVjSEhZrSkA03A8Dtj8I9auN2OJdJgZBF6KoVel7gqKszVM/nRknKS2qzT1Pyh9B
J2yxA5N1IdU978Jnh2V4ZdokYH/N7/YF9Ik5sKzRuCTHsm9V+TEV17JUK9gtkRnr
kXYpCQdzS+1mH5qSB+ZTWynV4ffnTXQ7biOLjIIw/eRzQ8tPYri3P7CgdPwCBaeX
KXHdjSBzYZ6ZF1e4uY5aP1T2m2zvX4+9vVJ/syh3Kosc+mccxwWFccq1MXw4Fl7M
EDBeUPtdX2OA4g666YoCuzH/qBCdr1NOKn+3quD4RRJAQFsaKzJYp2dvuI5cIxTU
XlvuVtDre7e5sAKg6b0KBLTC8IZay0JC6NxN4p8kLRoR9L6jIBCFRAYWU5cxoy2I
mARLO7cIYWO2FRhG26X+Z7m3c1FKRwFJjc+UnyH4v92z/9DMlOEofa+yfCCmjyFr
eg+whBhZvtMBjKnx7rbusaQj97IcIQVqBhl5n8etbrhNWh/vGEvqwdFnN5bDsA66
YbyhuMNZr9aSkNBtRq+JmYkzZLuKjN5P9FLPUonPsKwN4L/Ab8J3NfJ4fbuGbTI/
hY4dPj+p6CMsNa57rV+5VsWM6KUwziWdYyL5lnM7aL7HeACGJCxm+rK+6PljLXAm
kbKVNgGxp1s9uvK1xpll+TKtObks0G/5eT0afVIGTVsEeiTfy6p42a+quGeqZ1Jk
gEOn1x8g7Sz2kkSxMI+iGYCxGE9XzFu5t0lWDlSJzOAx9SjTd69WCUO35MSVtKPE
rtjhFvpgvtU4hqSaNMBEZ1SvWQi3QKDHx6JvXP0SmVuL5gwISZJRSu7bZeyFdN/k
4HPrUkuCmWRDc1Jpco5utvqDXxmCGH6D3//XEum0M8YzNas2q8yyqVhlcgj5dvl0
PeOkvJf0Sur/xjlz/jil2o+Sw+g1oF1IGPDHrk6Q4fa99AOvkRuGnO5Q5OuGw67J
x7yJjapi67AXjxm+bSHKwPiCRz0kmD7VSjOOCbOc0EIXgV7yGuzB6OGlf7aOGx9W
CZTodlp+c8bRYjzIg2upBtiMGY62trAM6VDLAlV5QsW3FCYWxHuJ1T0yxt0rcIQB
4xEXVi1iId9ayhTX9+ZQ75A8TeyFFW3YKFmCGsBA6MNDcKQGtsbJKDyzCgAKyzkP
q6gjtP2PZVZrYsD1f49nmj1V2AajLDDyvyUfTs4NOyYrsMpLcoQ0xkgXZUPLDpX+
SaL/dFGILzOCq6DnWkzyUdssK10pTwlk4z1Cox0nvT/kdJB2to/7MTEITlMZB2sC
bKxCVVImEitrBQjy/lYUGng4QqsPC1zIsIvK/03nWIr96JmUlwvwd9do0mtBFKE3
XMA5CQdP09ffasACTfBnoBOnMCsmt5NOtgKooOQU//2kwmFSNQTX3GWdaqvGewMR
YpysvA16TZCcEzVocvWi9D4b8wR+k7/mNDO+tei3HHN6yKgeCBDVNXMLp1wt9ea2
alCVJSFz9izKNNpE93PP3QLKHk/eLf3voaVNRJCdri7CeqcF0BsxUGHTnwmJ31pI
n+chAYoQyriNLjzoJaXeAvSrAiIvywVnCGCmkTZi17hVQ71Xt7lYxZdhtOPd75gc
eELFz9Of+uZLHx4c04OnhSmMAClrVczyrmLRzoI/2kLje3rTI3ABe516kXOIcJTh
sCpB+pNCSvjpE7L9lrVSZwmoPfo8bbl1Io5OPvSIuBfJLk6qM8x5KDXlWO72nUUr
gj8rRrWdLGXOqnPmsiK1CNX3YMXYixhGt+r6hPOG56m8IeR7G5+rfZ/KhU8uQHnj
RAJSzfraXW2FPs2pNso0jrxkaGYAOFRddzhltuV1olG9aPOUuZRzLiXa1kKB/h9G
OczzaCNnwVzX24MZZVqfJJe3yQieqjrcozU9AQx28KB47bK8KyF8Lu1kP/OtH+xK
QSABeWs9hOBOx4jHOXvPauVI5qnmZCrjvoIu1zKLW+723GhKHLPU2fWEb6FYMxpo
DZ8Gan8Y4sHZ2FFA4tDzMPiF/1cPnsTGwQiwxmJHoCK6K9W/qtplPiJiwxBerclQ
+AB5fjIgx7R9MZJSOwIrO6I5sFhQCXngAVkFtTA5uUmsyFJuabNrFOr0xQqg6NoP
jn0KmtHkj0nKn7drXLhLDzwp8h8Ue6u4Dc4RLKi5cyhz+Bgjh703CsicB2SrmPK7
PZfE3KGlYUYRYqi1oVjNuAOYctuA4McdKYTOsaCTrFalNy3Vqm4sN8xgsFTorpgk
8iCGfcejBh1QZy19SKSa9AWTIo29NR0JqHnl0hGQuimOZrsnmIM17adrfRRwrk8x
RBnnHU90QRwKWP5Iu5S8fluqgTJScHK18ofMvRE+1AwQ1tlXZQD5g2WA1ZZTPRCd
+juP0bcvcuvpoYrlageHxyN5vs4imnDm21g15IZny/YGvFLQ33lYtc6AT1Fp8FWQ
FktMYQXOzim8zQa6CCzCQfFmDfntdVZODw0ABjGGBahqxwBb6l+GUodNEVgjCfYv
9yL++DmbjXGbJuR2yS8whR0j5VCYZDaCWoFC0trCL7/wxM6A+i82aNUtMvHNeQXz
mHtrOOH4xCS7LVUenIWAQmCqAuigTihPIlR8FbJ67aw8cA0c3b3pEag4zA0Ox2rZ
tXO6jKYudkgMhijfo9IJXOf+Drn11njd3QwD4frGGpwkNCIaa/xmrZ4pXl7urTo4
1x/NTnzJCAB0G8Pz1GZqAdkvq13WMRH6JCF3L80VFXgR6SBr+Fb/r1tTNdVxjCk6
D+g0n0F8RisVfOKcCz4cqLyawiHDmRZT7/6NwlqhaAmEJu93NHy+ypMSkikxjB0M
wPYfLmWhSwXasi1mIErwMqZDR2kWrXGSYaJ8WG/kqnCJt51ACJd8wp0kWAQsGTEM
VETWwn1HWAKAGbhmRfyzpBFufS7ZAEdd9WUHbD1mYqYWAyuGsBPmrFgyIVTGXeY5
SALwGKsYvWfpf9qWxIC2gB+4ovfrBWQR85HYeKdD/72vkE01PlrTiPI5vrqvJeqX
SeFPe587jk4r3RX/misetC3tBezvBVDAF6Bt6rAaWeLaO5mzKEgdckvXD4TrBhkN
yu35Vihqsw29OZLF9X5go+2fSH1SN3VKfwc9wXX4s3tcABJMumW33JxcoErkhpP2
+AL2rocpFCCx+mfBfvjhe7NtTjI1MS/e/DcSY6UKG0lEbUqrFQ982X+Qlzo06+wJ
gkk9V/9NiwEt+gvoNXM6KKh4k/p1P2PTdSl/CtThyBavNKegeQF7qBDz2/h1X9Z+
om5EdzxbOJGfw97JvkFlKa8YT8odpXUcj1xp1Fr0wKDPdinJ4IH5SdNMuSQMPomv
Otkzf/1rF4vbE2Jq5dBth6t8lmSUW2Uk0rZcLoxwGTAMpdgArxJukQ5CQggmVDta
UGSuFQae0Ua0YeiOCSHjULPztwhdJ4R1S9gGOb14W2HfNJ1WQikq3/qjVWxQVpvj
D0pm6FhFQP+WAyWG4OAOZ1eGMjSsTN82koxHskb03JwNSYAnnAr4OsATG4FfayUH
GJeoRNrV0EULv/cQyZch+Zc22Ebt3iuma8PYS7pnFeJoSzjaKm2iW6oiwyt4DHur
b6wTie2bO+G+CksFXweaNi2ecrnZXBHVh7x2RvqIBD7wMK7SkceAgiykqP1AnUEG
dt2yfH1gN231zPD4zh4UlKoTrm2cmp3OgfDpcOlzkXEN931KQWQnf2+jom0rKXhe
SNELkvbRiz8sXNVooS6kKjOJu2ge4ykM37HjadaR0XJksg8C9MDJJhEAS0ELJd0S
rucc9hOAxtRMY1O9QSEa2r8GQxUd0O9UUN5CTGwDF0qMxPs5DFCG/8LguDEI1c4f
2iwJz7DSsWtXn/pJ5cRWgVtsSVc5tOVCH3jctN4GRJwST2MTSm3Gc/J/g9luF/Oc
Uwv04oz/dPjiwRslMWQaRyHHDsSRqEV2NzdZKxAEH5QR4TczFO4J2o60VkpECvUe
HbW7U1eRUw0vMI0oi49t+AKuJE+gPb79PmIe7hzFRrjCdFFx3RvrjIlJ3x6FpcWz
LR1JZpLJRSS1ErS+htrUOvnDmGFdKMWTlEuhaTeHxjwZPDeSPo+X++YY9DYOi9gD
ENYiz3vyk7z2o50gOTXjpWvOSC6VeMpI1KEVBn8Sg/rB3QUyFCVw4czEzD+DqU6S
vX8CMqV0f8tfiOGhfyS4vuA8RIeEhXuUCZHlcwlMJeXUph5KHGhg+1npnSVmhT9O
yWWZPrI50lB95b1tOPs4/YXfeJCxYer6NcmrPb/u3gBEvVfB4BzONnb5KWlQTgtf
4EwuVQUay1irDimabmRc0w07oFDbC/+GLpMTeWTTRSSJt6sXCH5v/WKWnF5tLE/V
zCXI8245rs77vcJkfDimJgI+OMjiZYO71s4/HsyTxnQupFz7pFt/eFDYb72H3xRF
qT5H9TiujqKfxMVDa2CMTs1fc3ypiUvTRnt1hyIYuR3lllTAobPw9lTgP21ZfIkL
eCMj60RKfXgzCJK0Tc1w+KtYLwijjeunAWz8Pfn8j3n/9jfBVxjkeLAkEjFFLjN3
KUADKO5V7Mm1G+LNphVBwXqLaxdz5pbxQbJbnt2hab1+wIN0Memdr3wha59rCdQN
g74+p/RapVxBX4zxY8iChg0zAfPYuamUCQU6qEVnXe7+2R+juGLWtOrLpoVPoQ4J
K4gYkOTjJo62BJa4LYiup3i+GKeMUZcNjMBlzFvBM9PpZHYzhBlLSOaqzIU4T0v2
6H2wM3QjGMJYSXemXdHRSZaC4Dmbh71S9hX+u+vPtqDx1zo5jVZibP7Smc49auAA
JOdiRnG2QzUN/4d6c7szRLG8JZ6tK9G/14Jj+HaUdVBzEWvoY1akOhntEgxyBINH
uVjT7mlFpqwU2Bo0rHl2eOSbjfns/725DbqBro5bhNnfB8cnurAzLeTnu0tf/3rK
qNjHenxDcN4IY8TFOOQxM8L7VTFEiBCqhhcU79O11wlVLFG5qedSalWacYpVngJJ
KiqvkHRTctSFmNva7lXJ6U3Xv22SXnwur2M4PM6RZwsNrmzp8Mr2iSg7VjHhFBkE
feNtjfRCrzl6sccgkrGHIX8Ba80jnb0+JU2POd8IK+Et1j7Hu2tH8vPPKosQwCpM
/mV+793rbWLx1T4uiiUAray4Rrd1+k3UlkN3Ck4v0Sql4a1L5lXphFsL3aYQRrfr
tdzP12wqIGl0XORDMleH53IiEdmyRHIp/oc+CtfjCPLrvuSthfsJkLIwoI3t1eAo
p0VGFHTuL+kXmONW+/3ccKOIUsl7kny6et7hZ/VUVHU8t88q91HpOzQ0bKE+KzVd
uXkVaBedkskZaBOJsp67N8VIIVo5qUTCsHrnE8jAPHyxTk3j4fguHBdsN7/ja3D1
4+877RyRs9lihxNoyQmA/kTU43CmFGjE/o0KMYmjRTpgkmuR4npnl85l4gA0DHIn
BOV6wHkmywf8nmGXbCV/Za6jSZe9kCguXLDjqQ8429gLQe/MN1FHcKx1zuCOx5OW
0fpfyFrsW9UWfFMRGxmzTnNraEAZ9BkwgB9MvO/kvT4scbNSNyVxoukAUFzs9CV5
5ffof34QWYN+OcwcElt1QTwstFtxwP+mIq5S9QHZW22KhRt7ffKnwUJVA712KgIX
ShPPZCnYvqenkQDkCYt7iUhM8XEctcaQAPPsgAiQnTMEZ5UQbMOfis1/PZBS8qXd
DMWXvzDKEIeN4VftWdtoWsTLHc3foXkijSpVESnROOih4+LBPB/S3Bv1Vmdvjww9
CFs6OaQ5Z6Ydrppp+ifSJ09etMuyZuhHmjesCVKpWNrFEDmF5fwaoM3w/LkFNde1
uT2r74mX8R1i9Gq++XWVGKp6W+Dn4Dnm3RpGqKwSxR6r3G0zLX6IYOvQ7mSvtScd
311gWFwAC1wUQAGRlOfZf4oHc1Gs0j0yEqTTUGJqh9E7SP3AgxlbrUQDx7/20d+P
kwC39/RvNukilmAlowtp8sBjZql7jrQRHsEcXBYQk+SCzdTdJPyefsC0lXhez83s
dcqzuoXykpCVk0z2ivlGZQvFgH1m+/MTybxYA8eAcIe25Ums1zF8HaM1xnzT2Ry9
CoWonYADOAAPopJLIq6Xtm4t/YGZqExBF+Tlvuzu22sLuDGTI9sjw0+NGXg6yXha
Ao1hHwbP9jdVfGsw6p0DCs2z2CHrHtr6igovY2w3tTg1A/VNwhW5QJ6okNPoRXHr
Dr0sml+NK/IBu+ALejcMk6u7tM/BSwS3UXsrQMHzD49wsdyahPtefZj3oPgr6PuP
Guj1LH/WdNXuBgIAjbUyqfAUhjs30Jcg0N//DJ+GGx9G+H32afGN1Jbj3n32XZLG
biebYq/3CbkXbuz95LxOXioYcjTRJWndy53+GLWpDl8XVohYtjrHvOzCT8SNuHDU
wvx3tsLSB5bTGCGXgWzLhULFNpHQVSs1nZNMSVwfM8unsHTb5TJvcaPuUdA5k8fp
54jZTKNf1VTfrQRs5LtMd9z+dGedmdRqDLmYEmklltKkQgySLXmeAHCFCBjav2oq
bt/MB5PQKQIrCYbhxYinJuiEK3gT+OHADuweSvZMGONoXxwjoq2RdkI7qdD1uJds
C3NoWaSwEL4kVo5gJQedR14H4TPCYPoDPuIcMemgyB+k1AtXk2Q0nnTTRwT6RAGB
6DDWcZ1xbsKLuDkfXbNmNtJeTDYNJbGIejOU9HeYpf1nScgTvApAxXgBKec6LWcc
vXiCGBnk+DMVMom59wb4OBkQsiVs2hNmKejlDCFl8zJvXvKaavxMjeC+R6DF5qVk
Mq8+O6IKQWdjkxip6l76hyhoEsRvYVQoqwYZPwUzpc/80niXbTEv4IVG/sOsurj2
id1wI8ATXbcgT26YHWHrPooOcEhGZnSLb3VTnEZi+rca5suylL243MqwVip5Jqhd
okcfLxlvH5BRM5oeeaucAXlX866FH+CFBvOr7Ck/+CMedxZRPEuuavsKigkwSSMa
OZ3z68zMgxfOktBOnghkRpDK7pQd1dGTlnsD3biRYks+YGiVzuQ6zOtzDwByDHzb
zcGez9WVoFcRndrZUQGQIRe5VXxAHS7Dbga5hnYDYOUjoSP+3nZNtqAh9c241wBR
vTYU1DDspUT2/0C7QZps71E8Y6huZn+2YyaQj0UNQGGYdh1DZg2ESKeb5lgBcMl5
u18inNpBKNcUwbFueC04WfTiKwUHTNa4FUjKPmfkDbGAqR/PEfOOPe8EQz2tt3po
O5DF1nGbVsnH35Fj3UHCdWLhga208MTK1/DvScBp3+dKLVvxYnHSW0n28JIkS2QW
KQYu35wIXDrpPozWx1CKsydWnfO8hkzZWSqUI5hRpnBHTQTY1EEctosKfMnpG2in
m/CSPAr3qL+nL/ffU+SAvCeNTBcvZ6xKpXNvbhHj9QVZOnR0x7wQFpVmvBc7mhMV
yWjtJ0PjOxR1kodDcOavTXZcjHUFwv1FD9xhEpmAO3CP61/BnjJ0Zmlmq3S6Klz7
UaNUZg3FCO/BfmrwZZPF6XyjIIZCGZvZOOKu4tvzF15IFyi3ZYfvozVMcowg0x4/
nNOU9KFsgnZs93kYM0VO8K2mYv0pEL9wYl4iBZ7Yif+v6P1cQgoDuVEBg8GA7oWJ
gUbXGhl68cSXG1ybMuLlgEeGbEmqdwNslCulasS7UBZcMMQ2sf0RWewAU4RajWQX
cL3sTrlizO8OUFpan14jRjcTwt3m3O69RskRecFu87vq1qKF1+mKmTGTHkJ6euWV
mfZpzlsNEm2bXyJgOIvYSmFcHhXjj/sy/kEsGzpIFCXFi6gT7WfDBJ7YxSjBAYjO
rdhtoUNs5OvsXzDyMJVICw8EFbT7nWXA3Fhzh8k1oFTmXrN5G+niWoUNBxkz3fp9
GZnwGNVwT0Ovxxt3JdkfhzHDp70ovTuhoGPRHOVUzecsly7pggZ/EX/dF9W4ATQp
EQy/hUA8VwZr/eUczz3hXPLcOFeGl5shTDpijmKeb4en1m2n8IKd8b5knuYiA7jL
XH3Zmet/Uq86HbGB7+YRF55XkBnpnoOC6Swi2s21ZggR3IhD7xd+p1i+kNcW99Bf
VFPhoi7ZtaahIv+jgXqqvjuzUCINjse26XoDyeMaX6nSyXn+6m1Gq3hifwYPR5nZ
xYymOIxb/5bRPuYzAawWHQJphd2ROP0ix3RGIiYZnBeWUCzG3VOB/a1/xZP9+bYZ
7bYutnEwOnd5tf41GfcTotYzIebUd3l3AoB8D22ThfWcS+4b8r+/lxlqMEvMg/fD
djz06EYCrsxcrsmw4FzDSJ7D3ADhqAwIh8bU8h3cDG8/lLPBlyhvOLoNor9hPx8y
HM5kNkBHj/Bc3EjnXnMg2bMeRintxgyHydVTQ9qIdqs6cwDs/KpwxPWHgawi1F7n
Ke9Cj9aQGXv7rj2y+9Lvc+X9lp7MB9UT869W2e1qRQcDN1jGHNO1H5vbuTUWu6fc
Z9h+9N+ab7/0RYeLYby0WFrcMgBtkcxH92Uy/6tesJEWupgDSJ4jRsHVdNJifoo9
i946zMcSu16XAtyfAghU12/t16n4tMH35JKbgWqWP61aRM6WjTR0dZhi2QgOlUpS
UjfHzpe7SfKePmU/LOprxFLX1mEuaqxugl70BzFUAYpB/dSUAtwHmofsxfkBUbbi
E3CcR4RBMcMSQpPqSXvGktSjPXk5iNGwkEYXKt1Aruweq6midSY5dWAIBYtU4uBE
5wDPSPWnoK1oyEqSLETKhPR8zjbEl1d5ed41/SXkCkXKBDsUqAGVloDZyMtvRYf/
kuwFWUsbcD7ylyg99OFMau9mVI060u/mu3d2sdQIfJhBwGbLmRRa3LuJA8tmRULK
7KH8B+BV429GUCXqDnTMLtgelE6vtJTHMt1fdrWUwpz6QpQxN5fLIZIvBQ/chXBS
dFM1CmJ+u0oBJCApz3A5EZqFsAGo+R5B1AgUoXPfBQu0L+8c1DMt5XfrD4lGPR41
c+6u4xfhvZPKPJPJZXhdfewa9CjcoHWYhZecMFOctXsHZSYy7YYs2irmm6ycjV1Z
H/faE0tfWKucWLwolUAndPUdwvxrmSQgnbyVJLA2KRsxy0yK/Uqe13yQBYE5Jj8e
5IhCwKSL4TdvdM2wO/ABppF0TilZB6RtGupx0y2eYU4/XA4DjRIaY1nMy7XLhGXR
cm3KW5ahXsf4buRmzmo8cWjCkbSxMmOFc7J0T3cfoWWnP8zM546DvK4c/00Y3r4Q
8Q/Tqa3FbPKYDRV3rHQFrXWy59aHwQdpwuKhPnyYgw9zHYUlzT5WoQwP0VPmhPzr
jTc6QItZzrbokYB7tyg5gnJCQnsNUzc9shwSIeLXDHsotNoo0ti5kBJYoPkvQ+/o
qqgjI7mJ2KjAKy9wwX8xq+S7WBcyXBtQ00iozDUj0okGAXktYwDhQ18RvGebAuJN
QgEuQhC/S3VFqPeM3nui6ylLHQsPgqbVKsl4EPPVWS1X8cJ9fOFGR0CfVUHLBfGM
hBn/rx21eDuAHFdh3dLXxxYJDv9E0m8gROI4ZfNny/djXoX7Oz7heQRpoyoPr5zB
ceALyMtAaUkhawlD8z5hsOK+ZuHNUobumZYtcEUUMGIE31cpOyHDSfVC3O1BE0ss
jjIJpMYhH3bOsbXswJ3kHbEORLIhLt0Ba88A7aovJHE4BNtkHM1/qZIB9dpK/XFv
fVMXv8dcX1Za1VnEAx5Bqy6Ncvy63S83nGtc+mZw+NqOhWdZVqKbSGM/1gsI095z
6J0s8QZfY9frsSI69CVcN5YhXDWMI70i34FWYWc2gB5eU1mFpHMJXLsOqQtTA9iW
QmG3cLRplbo/g+DgrI0v0TUVYL4PKP66E7UeRvlyyCpqtqrJ7cudMDdNT/jpVcm2
imshn5utr5sJtmp61egXO6yfiRsd0ahRg4Wgazznmswpz89RldbCJ0odld7IXVMP
xdOmS6Ek3R9QG0UyYNdzQVy9EWtAiI5uT3k2cQPexbx92DGWGuiOUhHMvfHe3+01
/ga1XIysyYOQbRplz7CxeHMMS9xI6YT+qk1Z0fXi0Sw/vabMeqLlCMwz40bTqGpE
nGfdWF//7M/337f47NaunI6xXEwn2/QK8tb5WlBtjW4svYa7lY91N+ffl1FeudLr
goI0W2IU+BPbc3xvmv83YtLoT+BFeUXpIaTlzmeSF46Fw0OSAC7U78MURQ0rnlVA
tuFxHLoZ+uNvmjLXhJeQ9Jxg8dlCBQbmI4ccE1fHIPL0/xRDfv/lu24WS5hhQ3mx
7lC3T5RgaKWqQKp+NE1+kuBr21Z+LrgYz6BwciTBjsQCy6K0SuxMggRGIVs1b4ZT
zRylNfgo04qOvxpeTAmrjnIZjXL8Vrf08skv1/e76thHI/b7gQ6y4Q7JfJBqar5T
mAcvVy4r/W0v0JtE0IWzUBKKVdy+V+zAx44eFkqZS4NOtZ/xCtNgfgCnw1ycJiom
hiOICUwHbJFKVD6ANvkJP+rC0GX1fNzG2VgiDJ8dB5RVRyHy8JRvxPBJXSdAXWUR
e8B0HFAfFMcAWnVrYnVdUhuvzq+w3Q9HEFXc4rQjnMn7+/kdl1w8MUwo3bA5Xbpj
5KxxFOGj2kPAm6YSGCOabU8udS6Brx9M2TE852MKyXyBRCf4/f47Cu8Km91EbwKG
F/SkZB1FOvcjdmVnNvfdMMYiWn0wyjZVlhdehNnB3eIA4tjL0uz/AEEcA+0NXlUf
P3W90jKgiBvuYeQR2TOsTGwhRqjFa3ygBhsi2NBpROelsOjUibNFM6c9LkINaxfD
2dETFJnD9rbMKfwYW2RYzUhsiQA3DMcZA0S1hY9GgV9tBvEar25oTa/Y643VLLoO
thV2zxdtf25MtqcQUWFJQC6R9VKhVT9axNgio7rPy2K3eyqPAw6vPuFxFXumQDOj
g4Eb/ym/C0Wu+f3JLldkqmZVQxIgCpareP9iJKnJBwEOfjPJOmPbKhChrC5rYSn7
/TW1I4m4zFUEnLb0B0ktQNwATWM4gMgcVA266fdDlCAikm/wHa3QeAjTq6+d3ETy
k8QE676RMi+9Yk8QnrTuVmpSr69uGkEn5gLFIT48hTG043vFJejgJONILCYievTj
chC24ABdDk6zAg47wzNPCBKLH/Yys9K3CQws00EcKup3gZPNht3DErLZ5a4eslPT
qDve268zzWVFAQ4S7UNW66id8TlbZzfW7O14bH7s496J40dDM+4NaLXWjUQhF0WC
QVBwmr7T+HSaqe1Zb9oOx7dRtpG7fDKF7HPpgtNjDWDEeeJ+ZC2a7N9H6uyNCkS6
znYHGsihnZ5gcjzwauhmcDsjlZ/oQJyEuzIWwOutK5Z+U2Cr5yYOnnq5akfv2e6E
uqdvC2grG5Oog4fuxMISRbcr9421sFNUTtLnPRuu//cRAT8zLJ25Q9Y3OBpJIVfG
zODFKDt20AeUY1n18OYwlzPUogvE7j6dXyVBN8COBTjHF3FUoX9S/4ukwo0nbIqd
mvn+mwTR5GY43408KMXcFhaDk7hxoX3MfuPXRbKJvdaj/imPMiaVavgAzmVq524n
uRIDHT9gpHBKF68qUYGgksCTDJTIONeqMwMCcXOs46Az7bUbfAw1iUyH1Q9Qs9np
HgL8eH9HxHNcVZE37HQLOFo2xwAE56DPhcr+jPPm4fcKdMMYFb9/eu5xpF3tXs4K
qbD5IVdZ62BOGJ3VrRKJgakkzFwSBn3lChj3LcjSE0u+/hYU+YlCwZ4562TmJLFk
urx5ZIcVhvO6YO97L0fTJi9eOPb571KcP0+RW9p5/+wcnltEjB+oP+mbSVKtLye5
JNTqTHYGJgM9DIMmnn+RdoSi2dPu/PzrFzqWlu/XmTDYU3Bd7lylhpwfBdKLj+KF
/YxQapngNckC4MlpLCqQIS9SRoNfF0YGUJ3YlPyi/2mYQAURcXZYCzcAG7K/SGix
8IRgaqvDspym6v8tozuVYeAaUjSF+fB+KcxNc39c5sNwitl8OhOdUGjFRhjlyFcQ
gzcqAuXAwe0zSEAM2veZx9xSANmPMv8j9O0FfxGf7CfZ3XvbUO6PAZvJf/3OJG9T
EpViTS6Wgc+9o5Pa7wCWbWej2gIbZBuOQEYMz/r1WxxABpNAhYfjO+l7Ncdm88H7
U555DRUo4dU6kl0icgmlqDED7XAGuql3+6yujkOlCc8Yb+cYZO9lcyl7h8uZp/v1
yj4w1JuerTwkIl3YwyW8KGbXoIpATlHNnvZnXRT1AF+w6hG+HQJiCpSDinVOGfi9
z8HIRMtsoQ3zrgW7G3GvltqOPPqfgH+1oYWjlBP1gFqyWa36lsHy5T+8sw0IKK3y
b/W0kHWyVJ7DZACnaN/0mmdpHZW0YemnklddGSXalPQOE6qKGBMcqp/S/1u1TiS6
Qjh+SrBrOuAbqht+fzBV/kRBRRldaPzcfNDEeEl15pLktT19MCRheoLAxiAD1oe1
ygPC7nS+8/TIHVqmx4LnmkoKFp2c6xxC1EU8GjAnkyzlt52rr9iQ6dD0KN6ijNcT
Pqu3NMKxrGZL1oVlBILtMqXSfzpNHETfrFE2wNEY9KijbPP+1Hx4f5aUKZoE4wq3
QtiPxcOA6fJGPbOyNtTx8CyMJ+dBY1ChORJlHC6P8R3ENEmvU2RYFk+9ba706gR1
uggEID9g1RVxuP8lA65B/OzOXchklhdOdsTg7qBa5K1v0vkem3O9YWeIORqiwYwG
BXV/2K+L6/RC5PDltVvStN29KlAPPU1i3snpBQMmGIaS8+Rs11IgQADXtaeQ7rh6
dl1EPQ0wa1xOrOFF3M0qjV2Nj3rZLzbHDyagOb5gfPvCSY3Vt8lr0nXNoo7APQ1x
rZv5z0iLzVLcZeMT39NWqnnGgxjta1lQkAiN/FCLZFlPSwASh24JfqrIlYb2IRxS
ZzSZqEGMXYF+Cr23VgWlE68X+i87V98rrXy0lQLna3C3I08L2LEtzn+OL39NUQk6
aDG0grzl+nZDlHeE5xqSx+ZRN14ohgtmVX/TjP3sfpkU4mhjrATLsVEtD4wop4A8
skp0pCaaJpD41UtrIoopJbOdgulhETOs4i5gJ6edfMocDV6MNGiUthtiubQFB2Ib
mVEWIXDissWmKr1zx/HFOBOgxV4ziqNcyNS/kOl5OodztQjE1XTxb9dy7qH2KRgM
o91K80P9WI6EfdOyxkgg4U9xfqfK+Rqmzz9EPqWrocvfiBOgA755C42iERoI39aG
NBsktg8rAtqkqWx8qvbCGEPDec1BYjy1nm3dO6+r7fvmKh0Z9qG9Rl7a9vrM9s7R
/Lkoh8OdcRgy3VdwKa7M7GPHjyC7+i7C8Z8D8ef6Emb1Akgvc4sXJfSof92fYLlO
iU/1KTBfu+0UTt+HBs7p445bjsrnQy5e598KZN2Ozjoph7OIgNqxO2JsuHdzSKc1
ukupEQzO+1MIhhh/vLohjFPE/a3pQteiBJkBrYZZdq6aL5I+4VWTzcGz3BNem0r6
w6mXvqovVQSjuUYu0uUpMo6m+QdnM+KJ60H4sMRzPqc0LakbMWSj955YE5HVld27
gPNP4jTbKMhKr+70ayk1DU/XWhlJUtDhunlxVDRhthdFtWp4hACJ/GTwt2Gi1XYc
n8+oD2SuB88GAwqkro+6/N9Wv1wDYhRgwuVpuBcWIAPtVPixD+OipBfNnSnHDcSv
PltOG3haa1s62xm5xMwueEbB9mzbMciaeF4lqFt3ea8oeee17rdgv6pOYNwxO2JB
Feq8nN1FWxmcIp/Cmv4WpLFWkiT0z7mBNMDPofkJ2uRvde/Ojyz6ZEGVanEtJg3b
47A9+UfbnEcdfstZYigxvkYRUYQX3cgTVJq0F/eft8mxzR0Eiy7by2w6f43M9/jo
3Kck/6wIYH0wYZNPhYTn5yjlI8Q1lBog9y6MeJt7nVrr3urg+AgCWHay+acD8VLj
ozUMdTJWMLlLA+RdTaonTdHAJDuRG6AueoBWXVVa3DbsKrSHyZf4RglNIfoyx+wW
PxhWcvQEtqslJMjWcO2TGML8g88cLHs8w3ZlygjN5ptx59nTaCSPtfBCdIuLkVhX
6EdIliP5fSI43KemUp5PwO90dMHZQ3DKQr/Ng577czdfaLGXicCNf/KyvIisf2nz
15hFag1v62MEKxJHuz3Aa4fGyysnkk8HcbeEhboJKpo7jiaF1pX2zjRR3nsGIKSO
1SbsEr7azCsl1sG5lCwVNymdJfKx9qtiC+GBkEPTYQPJ9zo7vr4lMeYzeL3i9sb4
dw5UAbzXNX6vvto5voaP0BwKbo/x8YW3tTeqKKlZrEJ/W5dzEjFRGjHuQmp1tqAl
Hqd0R7UIbeG6seM8iuWDey8j9RJMnAEnrzcBow8iVtnMDSCDRNqItPnaf0Cmh2Fe
98uSNdf/SIrwgvpyM6z+S98ZyKYV15AeogmyO7nGBRy5Xs7WalJRo/JeDjkwGr0r
DM0YxMH3eiD6EcqOifUy4WIRUJXldrGXgpJR35hJDQovd7oEe7bIUl+dwmzTdJqH
lDXnp4zukM7wCybP85l58gvFFYJ3f4epaamwjxifvnyE4c69L43PlJxmsGnqodvS
rqp8uTSNHEyChsIAtmyEzc6QqstgipneKkRRCsXlVjGXAt5ITVA8BhyYtJlXaZXn
31CFz1iV+XBebVMixb7UIw2bRzMnYTnpa6+UDb13XOsxdvKl+5MzKSzWhnQXFjp2
3bitXhe3KNYKZwPDuBBP2WV7/WfC8mUz9FyMz+DP89wTOmun3nCgDYk5X74/QLKm
lxM4+olbP+u3lVlnTcVUvGrot56/wvVuhGhqR7l7m9jdPqsVbQChHduQnxB4raAB
11FG+sVOu0w/7Hy6wDqlrg9jCrRHxmmSKF+VRXFTkboOLWKNvFIPA8HAPXp1ZOqU
hKiAZzb3YAECVvwAgKgA8pZiU20465JisaoJOTrEPOP0DzB01B7o5Phy4vKnlyCE
QFDjagHgLti6Nf6pa3BmgxJnRL7C3j0FXRq3OBriX4eTRUiPr2pr7pUAOi8NRa0f
6VTCgdz+AJw/G8Fo2GKaRmd0XnZihGXt5gX8ue40XhxY/BaI0OCq/lniui4+W3Tm
/iUoCNSdRGOZnWxnvj56VdS9NxnrT8SS7Nixx1VuvNWp+ToCO+/ZWuRozNzD6rmk
EJT7HADC1/8KEB5ZHLcWG0s1qoghgXalLv2R2ujf1RiFkUVTmRAv3800PWL9NCZJ
wiQyoYtA6/7Z4dEyOaCsKDVs3cHE2LMcuCNPBcnWKcYiTHELIBGznmC/1SaKLe5A
u3xKFUZNrrMgS2K9xk3h9UtJMBaj7zU59cuSjctGh798mLuWzvgeMYzx+5Qx6xW4
hEwyRW7xL8sRh9UM8p6i2HeoxUg2M4XNvaqSdkdBhG7iPJMpzeCmlM+dH0lfiYLL
Y647VmMe8jkwcVLopNKXKmbgxli+zcUJLvEq5kxvQJ8Sey3Yz8JE4xSrUM1OTVBX
WgjxjzP3nh60TiALOcAMP3t+qN1xJsXS908WLOH0Ginax8Qm6l2Uqw5ul7Hzg2rc
AZROH7ZnXXyCYjB3yDp22Pi/EDCFoiQa+BJx0oYJ/i9JA71klKmaGQnJssgU2jDT
fFh0nAIk/9Bmqrsqnoz5JT4OnO6JJNY2KLObLI6RCthoid6Fb1EDNnY58mCzBrK+
oEEKMndZO49vjfqrehnOuqYH2KMRZHvG0o9UVTm0NMd7HLzN2a1XKEeF28hCoqa6
kz0aP5+ZTOO44jNQ6jRNAy6vsZU9dbHEiakTGe734nG0+ZDtZ/2JepApw0FvMljz
mgo1q972e6foEoTOU9k/MNnDhqdZRiAkmpjLL+QpC6MW27a8MRi/mFi8LdFlu4cu
gmvil1NZfGo0ejqkts+HoLLhjBLzz0d80hw8iwCbaVcEpQWgd3YKgjX4U9IFTum8
3vpUIx0wJSdQ/WrZB3SnWvsg4RvRwLrduTgsCWpHP5tek3n8oaLNlM/Ox2TpstNa
W3PAvwVtLOURzHz/Gaj/Y+A10z+RkaPih0g0Q4Z5FVyuBAF7aZUKYnaxa1kVHcx5
hpB5N9+noIaEZi/O86duaj1uf3sUUbZzHS8uGrLDZ3+iq8lkbJ3Mc/HD8IMznJKq
9WnpOuyC8P5HgpqaaTj8NxpTU4hVqn2oRHmDHb7a6gVOX/ghkO1Cglg3MkY4f1K2
HLFxo74iX6G5vIqq2qRApgMH7FgSyB5J1/DBu7wgFM6sU68bw/O91zX/q16DMAs9
fJShhS9b6h0GXtQ/4woQULYhmkfEkt5dMV3wp3wqa5CBELHIbtA39utErnnVtddU
wZBLTJerchyB9aVfHfbUERgeFiVz8dMFUSxZV4Oha07WaNYz2I2LBrZh3x9kALCq
G06xBAvgitr4NqkSZo/P/tvRtiXQ298WCKtCZ+XXT6nRhw8SvGSebAIjANiu9qa/
QB8DvW0y/9oTF+XqAhFm0IhXk07AXtVin0TzuJuJe4kVfmaJmwcFdO8J1twtsK6l
IH4m+VPAjFzipqzbCqD6TD2gMzd+gBg7zxmeqzWa2RTr7LGgz/Y27T02xJtk0piD
9MSHYy5DKyeSrGAT/Cuhyrl1/rY2+tMn8ui77nDWzmSJL7U579qeImwHH4Ti4ZtP
Ky2BHj8IuU4pP6KsG3aMRPcIybP4TCkpnL0D7H9t9bQmdCkLmoTQoi+l02/T7BCa
w1Sxv0icRIGUJ8qGzmruj08FDe/H+yIH0J6oQC1mxaQFksngXOsxTzjpRchqlm9J
FAJ+r41782qHcwzy1mGOOBCAl7dkY+pkKceiVybdC9TfNIQSQUyMJloBv2qZuc25
B8S0+00wnz/2BNjRj43OH6SajTrFOtB5hTdR7KOWfI4JOQIH5JBylUifAW8EUGTG
SfArpmRVI2Vqjnyjd0cBoZQW0hlpadk46eUskVmumlLX/utfwWY4bOdAMQC77NEZ
1ZNt22HqA1/SllF2vOGPZo226wfB1t5/xulAy6iUh1LiHcmcyDtPUrZ9CpOPDJFH
Gts2bWvKpQJlidakjrU7WUmGGEZ0asw3YkhtFi2ukQd5A6zU0siqRwjNHheIxMS0
pzUMIxo9kFWZ0PdTOT7aCOk8ENqTGAJHAwTzXZIfvg7E9Amrkt4+WqW/tJ9OgJdX
rS+dG1ykxkMUYT5vsDcwfQhts2GFSaPmlZwmBbehVWyz8nMhhiqFIIBHShARivL8
SPf7qt1yzD7S+CkDdqZ8s3ClgjxINA33Iq3JK8+WQgylenp7lOHmOiLvg6EtyqcL
5X2rcOrhAZf4jAMVwBjuNygkp19karUyOzmHT/at/kuG1AzwF1zPtRH2KrAYXRyS
17XRMZBCNCFh4fnWHV4VKBXriVxqN01GVEBzTXgzF+IPOyr96ydxViV3zhSMX/ZS
RloJ0pzPdGJ2btVROnMPJ4hN+6sEUPWAHF0KVZEgZ/V08c1hUFz+1Ny0ZmVRqFpa
kJGxou0dpRQstO7mwtUvQglDtU49dUmGRvqBDiA7wDCuhF0+0nawE46iT8D0vuF1
84eQkI/9DBnp2rc1jXisRCKws+fC3l69zbZ9iClXF2KKY2s9Q+VAyRL1T5Ztq0Ni
eyU4EtLd0/9EhoYZ6pmndsT0mWRn2fMoFbxwRS6Gq4BiaIoM9z7lN34XyKoZpJ6E
nyce3hL3fbP774l81GdT+WT/9hApoeUbMYO1VYTa26rzvoIqMZnY1wRU3V14iO5U
/DJA+3SdJjs52Ro4XcxYP6FdzKf9dP8i//93f9PQltuTOOFsXw/r7jEf2AJ6K0SA
BZBRQny7TMcWgzuo2xQrts9gwPIQCsn+E1FQiE5w4TQ1x7AjYCC90K+kNa38NJXL
C4s90lGvfx5sh/lcxO/5uoAVOzAVbtlqPqZL7uqsZchUY51XKxc/kBncO24p5cx5
0kucj9tQjKTXRv04SBC6B4DyGmsFSyhBKIMiX4rUEyIj5Z/yHVd0aXtT3aK7/JHe
ckcLWq495E7/KHUTn/Se31PnM/9mT/mYMA0/MVI1PF5wERV7KN2mHS/zt6s9z1Ow
PE8ErOOhgybEk787R7tRXHyTANy+EJikriV0WDhlcznfHtz+al+DSZ8uYuA4A5sW
OlQ/BWQIdlhNOulohOeq+jFZMlnSmdpnWy0Ytr5GHcUVsD4zMF/b3e8j8kNM/p35
9wbeipRE61hHrzEmqWH+1EAoafjM/k8dXvfeGFlOqiZO88TLJzqaU4RK86vdskSL
OojkcIy1BMuwvmhaK0v/qlKzBoCyCbEhk/Mb+kTwrCKx6BmXMIvcuSIhm+agFS2O
sQI4WxCD41NWXnpEEykSJc9zL3HFdP/9b3Vma+bhe6EI7Dttgbc5yGJ+669w29kX
ZOiXKMZDKNbZn8Y/29O6KhNDK/gh4IBtym39BkxkBY/ssQOFyf9mKzX5QwVA2suM
D9Zh5iDS6Uo0ZemV5w2Xwlw3Nb/q3w1/S18Kh9irkVQEPFoNNhyGdg6+0H3MtMKX
xZq5MKYq+WvUKwp2hwm3r/0AM/hYIYOgifruuWn4qw653ixM8T2hGys/vzf8Oiij
3+LARbjesz4nAm9Kj9EpgZZ//7iuPKboxkeWu9jBHu4iGGx3s+CYYNdYza430kFf
FtotBJoVJ6K2Eedlv0X3rzBfp3RspUKYOpiiEWcmvlfA6uX8p8Geg/GjMemaJ2eB
X6likyGhGZVzrSi051bY/+oD93DylhSxoeyiUm1SCMeuQx2f6pERClVKF3NCs7V+
vArwc6vFVzd8b1Y6UHbm5MjmAHbwE0L/jeNV/vj4zLw7UWb2DaKcSoOyQTHJuKwY
wVn5B+F4IolV7aUIFU5sHij8/JvNH3M7jxR/3OiSbTD7Rnrwwmz/cbu0O+4PRSCM
F5mDzX7XNevL1NaBBfhrPXqfV/Me1T13ahhNC3emyLp1kW9urjQycDzbDm3a9nF3
10X/svIBs49F3bOzicEZ/wjyyUAX1kCxrf56AVITo5GVySW19RnwTV6V6lzprsai
qZstdRQhD4fkEFcJ7+0y/8CObCxlvobD+de6gftLP+LXmv+3WQlCESlDTNCXw/LN
tZzRR82SwTyygVxPqZmuUVtV1JxKLXOoVIdh3eA5CQ8Jna2bcwy13cLLalBmcpMH
hYWZp4fj3tAatOTu1fwEOF5X8WGlQ3hYC6V0ucVeI8gOz+IT2r9r5CAEuHJXcf3L
1S1HYNzpAsGRX73pgzVbUnAEcInXiPvzXRwzvcrJaVrJRKJk+8TchwFUuaxH0CjL
1WEIx+hac2Rj4F7hvkR59DyKZxH413jbAU0DKhkOXfUj0DJZPfNgV8zaBxYYwGce
VqbeAT5gQvaftTYWX9UcD1grBfgAn3uYDlEm3nNTdUVgp+TVQ4+G71+fchyGXvMo
o0XEPS18mE4dFojY2gPmHnFEPmL+XafS+9nUW/RzbTXieTUD2FdKgJS+9fZzwyVg
8DBNDC2UEW2p7nfEflWQUMxGbKDZw6OrQtIqJC93oHHFzk2T8AdR04ONsbUu7TP3
y99YlRdpJTpr0PoeppJOa3dVvF+sB0Tw7s7bc3PXE8IlJZgP5/aPpOMl4lSWPI9F
3U3WE3OyBvL/X4Elh7K7qm2OIZ6uyWdF2gSe8v64dTUIjN4/fL2N+64LBvyeWZmh
NsvL41kXRrFj4N0bx3aGRlIS+ypHRyzyq8jXA0PJH3xC2wUb6CBzzFf/nyfkRz4D
06eRojdWN9BrawxrSQBgMldvyBpTDfwUp/a1jd+qcdrlcgI2PYKfFIE2E5VpMOda
e/TpcvUkybvuYQdnK0EqFrK/zkJh9436vZ03suqRCX97XCtMuCCQ+sv1FtM2CJ5h
P/SFkWSb53yNUGAjACXBJz/Y36p9QW8fWjBZQOUr5mup6OMh6urwuZGveZpQBLtl
lw+iF+GeRfVt67rr6+h1PyGSoPB7F5HjRtzbHvd8PTOLhHU02L2FH6N4eEQ9OvbI
ZI07JNpw7GkoLjdg6vEoTO596ojIuwubYufRysMgWYh0e/y9yveDjLo0NDnJtFoF
q8W6SQZb5QDCqV9wiAYDown2f7FXWOQSy2wZmeJcyNBEGulzWVsjbXNQ9SPuSmC0
nVOlVKGlOJ0b3ZDKYWUgNG3WA65BsYx8/WONxS95iNGTtG9RwIUJM6HA+Xc3oth6
boSOsrnWEVstNkLauurm0cd7FWl9sDMFxO2fY6P07K504SaNesA+YXtySuyX/Y+5
PqbWXVbsG5QLRPkC4qBJtv64frnNwwC4az1DdFtQidmkNg81wfDbMpF8by/bYv0q
MVvMnfbvm8tDTxoeFlx/Ta/SVA5Cn/6houZRrj9hOsf6U+Fr+uGFail4PDgrqQVj
eypcqlBa3WNeuDN/TaUkXq11VTnA5zjsxQQYYGvLjyq+qQ7H56gljUtezwrB9Lch
p1sNeds22bS2ulsB3hQuZtuyucMoaHIl+aPxaWmR54DZoWO2itAoDUYxvwR8o/ZF
wVgc6P878nOWwhJeV5OX7Z33rzfUVDAbwnZrflWtNISut7I8eeu6hrCtWhvOIJNE
ZQAYUaJsMCzfzkB2Tnzg4tEsDkHpYmoGPYraiRa2Y94QV6AzOePUnQVgQpU73kFU
dUiz3MsJOSv3lrLyvASxQB1hQk8PKdjGZyywBudV/qFB+5M6vZojkafOrBhyIiT1
eodSJF21+ysa93XyITJXLBymG91fFVn2/DE9pXg9jTypA29AROlWboUHukfYXULe
0m6gtbEodPUNIYbuBL5xOCI7tL0EInw7AqjoSFdG1Pij0A1FkYwUfZRXYqOH5VGl
Q4T9RjGfOxZhBggrO9z/hiPkwotBBYCGcDClBaaQ22k6wlGo4MgOEmggw1BWj+9Z
kWQhkd8mBqcRxb3D8BEtz2QP8V0WY6euxrvgLyJUju2YraFElZlkEiaQz17CTz6g
IZQBgoiXSXchW49WiXpMpbfEdWC3+VS3ipePcE09FeyqF5XPQlDEi8XE6enG1FhK
G9K+7IW24aALA7+gpMawaGY4K+Za9Y3mZdhNPFwZRHwoTjYZdDgkgEa/cWSafALO
mFFpmjrkKNunQmYfXAL+jDnVj59Ufr2/g5oGLxHKAgcIiAwVuKnwVDYX+pwdQZ7r
6I5WYhdpZFFQwDBK9Oji16DQUAgLMvagLckIjbjAekwqd6hi594a5pT4Ty3ySXSe
zZExH8aC2xF9emrM9jQUW0DRYcdAB2CdYvZssJbRqvBvWzbghdj0I48bToyMWaHD
mH/c/7c/ShtpwVHet0fKctN5KqRo0OSx4VpuSCvkmViPutIhX9ZJYRjvKLF1/hRX
W/1SRVW5IvSN6CPotp1CpHazv1nvfIu/ikHHCR0yTAJ/eBgSpr1fEnUQdQnv8rgY
MjbNw5v1LCHJrwudZExJOR7rmZZIzwtPNXmKsdQYCPbwdjZofajmI9zyfGhcLGQB
isiGS+H6eL596KLjb2IH48K1cc4sSj6eaukCYoUUC15JOvOgMxfSCSe8reA/k5Hz
1Eb1QPrc7s3gHxW30IW9xp6PkHJu2FxoJ8QkMrYwbbPNf2AnUCbRU/yGZ6eyVscH
iMBaqeXvwEruFBzBZuDoq4+IZHmwk5tZwHL5mEesyC3+bV0GJXhsNDQmg3pqJAW2
Silq1AZsfd0BEcHcBB9Dn7vhAEut6ypTk4B8R6aHUJgDxQ24BeAaJ1WEiQ8kn52n
XNf54ERGDiXg7XM1hhCA0Mv800A3qtpDBJPPCOZWuX5XIXf6V/mS0RTvZA+GAMkX
BB3YBo5e+VoaZMjvsqknZQh3j9BiDXzAx82Q79X6GTUl21AVwS5xTZtF1zqiuLwM
R5iXsdwqBzrytTu7qO6gS9kydZw3nIoYHio3znGjuk6R988CLnrMic29ER8oYSH+
R2/ezhTbbgyBaP0niHZUtLMD6173flVBxw110Q+NTEfD6JN7wH36e6lmFVOOmqkP
GiZmBTR2UveKva6KB2U9pR5G1qt6ugDbaMCmkBkXWOn+/HhXUmsnCCS6xOp8Xysy
CoCn91hV2qCjpijOfwqNRQCK6FNy67u085gdPWz82UhtDXeIHvGwi1lwds9Yrdwf
rBA6gMYCm4lFwY3KIBalLY2uUcUUAjbyAGip1w/t23D6K7FC64EVLj7jI+LpSIpd
xfc3pHzrXyNbOR3V56UOrHKm6HOc37tOq1dX7W8ce39GJCnMlJfYRUAAXvp4beMx
tLXJLT4msWxpZbxjLwnJ9zmIU5S167CTx8/9nLLFMbHJtbFP8QtM5aOErUENHGNx
yEazomzs+Pzz5wjdS2wVXGLb39ISN/wREBn4pU3Y3b5LAhzLIamuaHFzPoI+NcPJ
Hqz8z5d05JugLWh3sjZ2tZ0JnCEaIk14raOdRdeqAFBOeGfRKkURK4p45HekyycT
EH63mocLRujnf089rlmuGTJkMACwGB4XlKc0xgt0+DBGFDMrxanWNalSSjGyRBgG
jZLfSlum/9EOpxWoAXg9yYzN6OBYmHCUyGFD1nDvkEAqH/i0KYGWDMrND8DqvE8+
j4GsEGIcHSeEkZSIUo8Fgf6h9AqNn1SGscqT47i88j9q0priRnDasnc7endsJtnn
eyhJHNDmaUhBYT+KzC7CDLqZgUFOWIxYPs04A5j55/vl7RWOtDGYTqOl90CZGqdI
mq9otMvJihmi2QE48XZ6Zd8cPrWxoNN8UpoY4lsBz2V/bWmAUP7vwJF9vspPzywi
76119ltgoyj2EqR6QgD48Joe7oD6UMirXNnWMOa7V9ecmooFRKujYAuUxwKVk4t0
gwpvhkUgkUy+k2WigWAW8ft5CEc2UkUyg/3tMa4Bh8r8BObydY08xKURvZsLVQ3E
g3qOXbN9LrQhFuV0mhzWUA6otkSiZ369lfsS37vWK/bXA00vOG6/vpBNvMdf8NS9
hCY0NIunUP5+mqyyyIfxZktX6FIOCWwuQ4GeOaEjq65tlnO13/VTVhdp12hyrUMw
4jWqN+vv3xtXvON0P1C41Y0f29f9p43t/21OGoNTsLiDspK5QnN/SXxeT+EdK3fm
4stcvM8uZp8dfIUb0mv/RmboYECduzbAnKp52K+8C0nGxfGKbC1KAD//AfrYlbkk
veqBtEI//lIa6iQXnssWSRHUpKJgZuzQ/9YD5WKphMg2nzUr4lJVpPWMSr7jNw13
sPDePTqz/KqzAa3c6eht+WR7PL3cn9wftN5XxFpLuoyWmVtSRQUs/tCvWDzLm9j7
5KBv8i/dWmLrw0xR6wymrevySo1Ocs46gu7p7VaUUzDtSn/cWnWfoUQsWqMkhxdg
ZwhAAcii1uOFew+tjudkqobPTz/pasoyF+aOSclzX2XZMKAuvTOL2ljwbxoJgj/H
EhSUCb13u0PeRFp3Ox+1SpOgQJL5KWrZTmb51dl4mxDzpIfYw7eCoF/Ui3IK+god
OlPFEfoiK9ZaspGdo22SFCpOaeIXmVxHIkvZv4AZ+qm+KEBnBc2xpcDVzchS6qKD
xVxfnsMNjRx+tog14QE47PuXPHbuwIgMDnnOQMf6rzJTBjYziPZuRBPK9j52zVmO
aA0zkEvnT2hAPWBWOLT7YSTJejsmk6MY79Cna7sxRvtYHFiILf+m4VpFSt/VsP4h
ZXru/SwZWvCmcmWIrUg/VLnkj/5q/xDYjqBzkr+yiQkoRRu+smq/8mGIYscQyRCf
86YI16Yor66SeFwNkg8KQCOSvdpcisPEFCtwafGmC6myNceT4fXDBuwlv3A9NEuz
pG0z/y0xfADhIYQNJ2N39Dj5c5J5jOO7OX5mM1SYL/KZ9AnFVXfODY2FHmXfb7QH
fLvJeLpr9Wlr3/iYrx9ry/p1pXpl1DRKLpXgBTyHbZgilSDfTSRk95c7lITpAuuL
+K+j4YhxZeiyJPRrtwk078qIXQteev+soRk3DnTgayWC4gdfbsU/TMLlXxRu74U4
ZkmDZOynN+X4WXTOVfdmLz5S69z41ITyWxCbnBB7RnHr5OBewqEIkike5M+VNqyW
eZ1z6SmO/ZfjWyE40n+9mS2vPCJO84JduRE2Qa7BdHq2++VyN9UlG0NkdtQbMP+A
1jJK4OLzrzF/ry4DC6Z/olsckWgEQjaK2WfjKCczK9N7UKu8GAcjC0cmQbrlHeOH
ZZqPHrHSNcyvRrvELw3qg6NC2WXQj88j3JggGzq85fAflk8/pdEdtmaha4o+ccvk
3iPQ59uwW8FAxKiVhZOfPX0qdjtyDN7ROVvKzdzg5GZv2zAvn5Nqb5MLkjVuwzV9
CM3+a/ALtFY6gYU1sAtauX9TD624+9r6ugELL4MueG/R1J14kte6Ffz4N/6dpHqZ
NPGZUQs/hhoackws29Tbn1zsNuo7sfGWTsVZGRTNGhcQE3BnagxOvyQumad/wmOG
4G5bAl7MzEjRLs7iieNoZOrLbGFmoDarEfLlUngDjU1CyPOVnQrlwvufVRgFiTJW
m+jAphb5mxpXIHdtABf0CESNI04o22BJPVAJkv/HzokHLB/0wRjmOpwpsZbbdtGK
LLxNCDW7xVMqmPGFXeX2dDSd469nQoNQaWyz0M9dJs5DE5NkSjYVxZMpdWOWxW7H
IapEOAvAH5IYGJV8enMyu5H8iKP3tMyht9soUUor/pUM/PqBvwcxBeWXq8knyLIy
Pgl7ds0MOOT4X4+X8OztPdjVfH1k/fZEMAjbfmQu3vtE0Et2AktJEcuFAe4vunAm
jHAX6SalPcAd9qUh+zozVmAadVx37zrssrOseXc/C1iJ6a8/yJQQWFmqNmYVS4oF
FBBcXLW32Md/wz2hq7edXw==
`pragma protect end_protected
