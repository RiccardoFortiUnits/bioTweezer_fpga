`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZhFkVjVT24iBiFZkhl2IHBMmJzPPUiS/wb0Yna9Rti1BuMJNcMEIMfh7I1nE4qox
Sl+5llOWMy/F1NmHNzY0syKHmfnHmcoRM8B58Iv0JSh/Ox2OW+NST2mDLiK2NXmW
NArYip/OGKoQGIXu1GY2h+vN00c7NVBarG/D/m3+aq4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3792)
X4dWSPVSVmIPrsuRuVXGuvMoZHpMA38CqSEvg0/9PVlaQJwkJq8ufCzIl2/rXCsE
HXwuTy0CgpWf0Fkloj02oAXWo3Gk50lLVmlMb3HydWw3xq05zkjVVVnMEFcVU9oZ
RLAk8+XT8fL9fRGMbz4sh075YrzBjhX+ajqUCWzlPiPzEzfuQHeh5cHq0lqEJH19
g6gaGEaRck7ZnZpFRiSPCwduq7rWejbF1otlRYDp1MDWuWdfdiNkywZE7eqDmu3t
ZmBJSK7pBwdb/KYe56hkkbdfGqIWq2lQjwB7otpbZyC8ZodcQ11wr/6Kxb9nBynZ
E3mfjPgDVgsZk/MLbywnf4xsIW/kYc/8nsXMFZKXcCKpT6cvEHCUvzzdYX6yNgF6
m8kUAR9gLvidbSQk6kU4aYDhslUNheoC7Gs5nMmVmwrr21WOjnEIzB+d/H0pMl7K
UwXl82HFIcVqy7eY2bYO8xAVtRSe5CStjFKLfyDZfENFBoFnIKeONrP8ARNYyZqK
xuZAzGpSz1ZUMNoBNZ2GRmMKJS/y52ID26SFKhFjojURUxaoqj+GX97OjRlhPZyK
kFho7dZl5J6GMtw88TUf0UAVk0+t3D7bAw1kLPeHht7K3SotL3CmM4Y32X0dDxX3
dfJi9oE9pDxkBYNzxhwgnQz38Uc7S++1+RMrpWwxq8F18BFbzLTaZaYPR6jNoFY2
MyyeXU6C21Y/LYszZ2IQaO/azTge1n5Aw0gjhPd5E7zuTLU8dVIKtqwQEEzVtBiQ
jWwPqPWYwRVtwzQcgTTlyv9T8bvTsfd6qYAhd36ltq+Q61hhvLFQlOaWcaBJLJCT
0APn+1zzl8aKC4Ww7K28BklbsWktBLHDVxceXST42T73pmrhH3LCkPK3DQMhYZTv
g5uadr+FeveJb7VLy0IBEDInRFhvIHHHl8W58VuMoVTDD0wJAreCSUamop4c1n3G
hCRMNfAmpOyPWaum7jURSQKl1Zitjry/ypz6Wm24MKm3t+0GpLuBJ55Rx8hCYkuK
BqG9oiyPo74j6P/9/CpC1rmcvanPGRnPEtteI2WFgLiDsIHdKhxdVYp6cZ5RgKjT
gzsnvCay7zTv9em6Qz+HAVGo5dlzH7S5rcx6JMIAwr2HSBmPuTewwjZ6P+V5HmLS
fdd060Yhg2vfYtSkgO2ykQyfZVq4Qgpr7sv1lvOwNd/2l0kPc1XdysWOktZeF3yd
XmvWq8wzUwGKAFExgn0wly3x6mDlGLnaI2/j398Og0692wJpyKqQSQxZzVH7Ydrt
vigOhzvGFWNZMpgsDQQK4wgxbm8JlD3aKcr/HhumjAAdpHJ1T7SfgFXpSVBwiEbQ
ENZ8duUUukb+1zfWsJBcburmeGOihLt3MID+n9X4S50YKsMvz0AjatU9qOCK55G8
XTKvIu1hszgVzKmDT9kb5zwLTRfvtv0oRbeNmRPiY4cX7brShhCYJEHslv/QbZXB
aDpGyufxGxtgMNOt4Voxk1XnbzIGQZgZBO0YDwi9upc2oSJIG2Mx30FcWtP9uCjZ
WrIMwVK7V0b9fUifOiOcqpW+x+y/W68HDV0UZ5KJEgCb8W6BSREBTglERa2MtPA8
Wsugb0MnBidO4gIdbKIj9cSraDy00hFAkVSvTK21y31KXUcJ1smL4RNzs5fUu9Ss
VXSXoxfM/ney002BHCIywtd7lPkjT9knOfm65bqnhf2bPjvkdGEBsg2KBqNAied0
6OcjpDiocSU1sZIaUDd5N2St9PvIo7xlkPicSVfL+ubUnuNpsvcaWShlMjk4tF9u
KYep0hokZzgOY9l1ZakyOFiXdyTsyY6iR6V1OWejzlYreDdYrJheNwyxRM8kboVB
MZg/pO3S2FWxw0hfISjllRe4Nyx2eP73p4Ya98gHa92yZXCb2nwXTJrwD/muxq1n
1yGgsJtcckTpXyyYLCEODxWG9FlXlxCj2M2b5G6pjjwtdVznJ3HEAH6iudOG8gok
2WkHwfw4pczakMP9ngg9++TFpm9f0zmsS/heRHzmEt/HlW9SlBQHFLqGVEVUf77j
JW/uoBVH9YRWWdNiRnlkWG+zKpU24Jv2XZp/zIWEYdE3+0YU3QD39e+HBldK3GOl
Iz7f/IOPr2puLSvL7vtkZ9np1WnpqT5MCNev/E+m1/fLJy3qXBjqNTgzIVL7yD98
BVRSXxp67Z255ZutBDxYX/6qmUxoC3VlwakxZRU17VWdg8eu8Sn2LL6dUe+BRQzi
mJKCYC5RtwD5jw7deA5lmkCOKOFMCXL3EttFXry/0J/S4VGN+MOUhBfLdkjIaAcu
83m/zRccCaMv75Wnk6qTytng1n0PncT+w3kfeOOU/V8L9ldd/mHoF05BC0MjM7/r
1Qy4feFmE0eVY64lg75KzHfOPQdpa5p3lvUNR9tY0r2YcQFz4is60IWCYSI7LGWP
xQSJ/3lW0b0RGY/hc8OXXmwmWHqlykK3LcpwV+y8Ehixsdv0cPLmcwsW8vKhs+3H
X45rihl/kRSlMV6JGRyQ3ttRuGrM+YgUvRCVuIOz7OX5MyCTb1SEXtacajdAt0d3
FloA1KRaNixlTf4vdiflZPyLtfL3PKbaOOdJwsyGoL/5B+ibR4apY4Aa/Zykh/02
ps2Zhb4g1WTjzfCBhGfeyBF4OW84JPJhCcFcAEEYY/BbvcngaTa5h4JRrJeddFJZ
tOKAHPINhJh4IOnmVA0zZ1rJ7jX05sIogUluZDgu8z5SaJPU/9x2phJPWVmOSoH1
WNxX2g0mXNF0ZBJuyku4QJFhxjC3uqNf1Uqx0vulz9zTtL7yxihp8wFeUCQbopy0
/j53gO+ynXPjVPEZbBQWJV6Y6l6/bzqV91FT3yKh4ngzugGKGRWFLYFunqaroSI5
lqT9QgfQDAlfjEMBmKLz/a2aYeh8bPH+V8ZQhupaEHPR6++cU7UBJO3sQoxxW0rz
EWYlEY/xZQNtqCK1H9+761gCmuLzWyfF1iaOQhYLg2VEP/uFMsnQIle9ObMp1w1Y
jVcAm4/DBmJ8YkjSu0nJO9P2DSy2Amy+Y46GfAVj15kppVjfjqfnkOZR6kX/2Hpx
o6qbqcYMrdkLehpeOpV9agFFxGqFopVJdFlOFE31iZL5AB3vKFD+BIEzIIJFfe6g
O5ZzhwG6OdwNNCDZoatEUo3ynhHSkY2EeKFeO7bf14X9wUw2DcCjaq5IJ9oCxCsU
oYhtiLKBGoXAHfsVZxcG4wBpRasQ7P6s81zrVVlNK3/2xmoPLJVfRdB8zONPV1tQ
JmmAv8WHUaDMI3DXGgpE0S+WQhtEbgDKwByiBEtxBp+y2I1CuZw+KkpremSg07Rf
PmDtvv6DUx8kS1bGvM1x5he2psEUhcuai/0qJxAoSxuAvFjBxUG16MSddvMbRjsc
ATGlSw3PtvOFAhWAQjeVmaqcbNDvF5KeHSWdkrEtElkX0rpSEtE5CN94HHULlDux
Y4sZ/w5DD5j2vcRXHux4v2ZxANRhqTsbVPMbz02WPLOXdB2oYlacNxNoM98i3ZQz
AFlBsoFBTfm8ByY51We6hMh35Imi7OY06lRyMp7FJMz2BbnfX/puVPh9aN9D42co
NnFvEgSQMTfMvHa8ywiFZ55ZoRqlp9wwRebDvwxwadY3R8GFRnDNqMJ7+4aEVvO3
ekFrQOT+1oFcYH3KhgUiqwoxTrnrNS6V3qWhjGx7CBf9nUWSCRLSf+ThnVstrbD4
q3Fmr4WF/zG0EePYDy1BhOJP9+LVhCML+QpMNwCUG3gmuNKrcofhi88/XY0HN4JK
V0ddULwOit6OrOEHuJ3F4KMmGaF4VPddCgkHoJo6JmSoG+v43WbdfVHKVKnn8uhF
vKbyIUmf+TWrIt0Bb9nazZ6TGJODJY83yT/nzzel3C3BVFyEbza1qZSLfFDPzlkO
P9ITRc2P+iqymhpjdj8hLpB69is6lp9wMZOV011jOQ8AzJW7yf1zM+D3ENLOwe6V
1CMIv6cvicYPXjeolFbxuBZ8bLifyUxz1sH1GhEqLxg0RfSg8EOPjI9+Ap37iaSO
JwL9VtGkHSNjHs5mBdfe37uiWskWk6wodyo5d/MIFPFeUBE/KnqXh2hEytH8Yxur
sZF8rRmllydt97LrD/jqlRi75RKnnPcGnPj0+7mau6AJNZaskNGXAg3gKvJc9BiY
yj1xw/nLFoNQcDmUg4JiSKUSGqtgINbrJ6ZsCybS2274IC+a69CF1wgl+Lg7uyrz
fP1ukg87R7yl0VCcaF12v9dBPWc2+Zbbam6cSwOoIDEM58KKjtM6Kd0x36Hdqc7m
7fM6Tr1uMA1gPprRmENrH/Fj39YT3LCpP5IAOZ6wrmNsdAUQ19iajBTsiokmaGkE
YriljeToVBuzNXZiTgSdvhHOkKCCmEnx6aHe3nA4lgmhsO8MzF1Im6yYFBpO8YT0
ABEXgh7YsvFiORQzozp07+XvCMOoh7uqVXlUnzbBiWnXBnGSAsx9zKE4TiJi6896
UNzmmHRxzI6oUiZ7O7yJueeZhPvpmqCyQg9k5fuCL0CFc6MAAfSA8tX0zJrRg5QV
OzoMwSAjyH3pna82lEhAruAzwWmaScXw/hSCfKK5CjxTD7PyP8flnBWI8qc+AlgQ
9/ycvg93Xj57Dkmq8smuB4ISmMnrMXMHjV2jcvTO8kaC56VSOu+OavUFDGt+LBqh
ne0mEFPuwPrVzsXY6EaRmnZutVFVcPBBipE1okR6CJ6UfmxYW3jT+DrTBv0AGKBD
9daLzD3qYHWIfwJXC+Qgu1ZRqkLE9P2E9KkbZrUmnRIPpEt8zkqIEto9abVq7zYn
wwQhaYaAcdRw7Two31bicYuYi8ZPQkVvxNuWvfGRYy2AcfDNfSfXhFsqatlqiDqy
4E+XwuSQf/AoG+T7bYIKaGvFKhJKbloAqx+Qzj8xbFlRy2e9R4rtUjUYMZSOhO6e
mJj1/oLA09aQXp9deqxbzmsCBz1zyOPYyIH5kMKOPwKfVSpQ+vSBl1602rtRZdEO
/PDNI+0jXLgKvzTkp0Gd+Cbvg5/aoUnz36R5UHdvds2uQN6e/yOIQwxCFqLbsClf
`pragma protect end_protected
