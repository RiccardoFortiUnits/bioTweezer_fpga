-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
H6wLR9eXKtgXYjmvXVfGnxIn7j5QlNYf2Wh30fyBIOttdOm28N0AdC1zpvMIwgmbPvk5todbjy1Z
FSDUnmi9PHmNo4OQ+Pbh5NTNJh2wXRp+/DezWQUAqs1ttFFVjx/46Q9XTGUVZe6pPaDXIQQlASAV
XbAPzJKXZOeRp4lojoZv8E1FXzmspud+8IcshUs9D8mWS08Pf7+5fyqP2gK+Djr89e0DTQaBZ8io
PC7ghFv2/c+Ofnf83+I3wcM2s/J1LfAciQwyTVx2/ChQfPbgHBJDw6ijvebJcuJpQdDyelmU6aBe
PEcFT0EqxMhoHV493AIPh5QrnF5sPPaPwgdgOA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3792)
`protect data_block
xexYL4HBQoY7gETwvVORl8CyeDtZ6XgyZSOyHmzKsXQq3xuk6MH3s3v2HhFfuPcQPoort2kjx57U
0O5M/gOYTbACYOKhCLRnuTRFDBY9MfBRnP6CaQ7rEc2gPHxaEZrZZ6skcjRYw8rlQ0o3sUQUJ2Hk
93Yr2D5oWM/i0XHDW4gIxrdGfkacLmBtTHfXpLhpk2SVrBu4mtePQulW2qXlvakWaEcz6AzEUyZz
KZmUanmxmGV6GWqjtzlfVfJUjNdpNtjCkJ9UeNO9AkehfYGl3akDxN0I4sGXBPrFvaDUz7kfpwWY
s9xakk3j68+mdXRrWlawpgNR6NxIxWtp/JMRGVeRXIhUZNM3cQUpyNIGYnVz0IYY607OewFlcShB
16csOgbFhV8oL/YIGqQE4nfwjiqxPTSn7elqH9XHVnj3tzw8cn3hL1VK0jUt2ebhGKUWHoen6Izh
D8+38qQc92LmsAonZ5cDyBrfnSn+xl3KHTmP0bdjGnlam3HegTdfbA++KJ2zNO8mUHzxdiWV4lg1
GHZWmDXYoEgJUbzT6ZvauhzmjNZmvLXZFK0mqSXzc2X91WHulaU0L5aV5svquuZvJ58ivAnowWYu
y/ZD2eigDOCfACQR9yRk2clwXLAGuJrWjFRC3Zg4xpweyZhSsnUE6Nn+xa7B5T9VMi2zUO4XLSqG
wbOZXs1bcz8bkOWS38ie0XnXDO+/C2Is0YKLWMILhLgzhPHp3v49utf1Okwa6ifUgxV/6e63ic37
xtbDfDlnvfztmTPTcaG3H0zJ5z5Jbft9Yw/cZxpo5rbZUlrsfG9sWHt5N0gDkfxF/CLHT5AK0OvA
hFIuMKMI5OpeFKv1XS1KfTZBbTcIMwQ2dlGhVUB2+/pJpJp3AxJK3CeD4BUbQ5YKBbi+5cN04W9p
SPrg5BRyGiaw+IvBSteH+wO7R5TsPk9HE5ay1fanCZDEYr2Ffdfav3/Q2g5Lw5JaJ0+vLlIYEKdx
uxTk1jfGiA32EtQZMmKVsRu+Zt9MxwHBZo0L1eAuVR8vW15rTJuARq/ZCd+FpJL/rrIsjYhoPzew
O1roDB18qEoMyGlChpU5SwTVNTUfvPr7tAHWhmGK+MTApMpU3SCeF16JRYtpisrGTm49clBj6Eh4
XwxUyfZvDBYIOmVcn8hplXJO9xjU1hEuchFzzR+HaRH140Pv6HZavwGb1QvwR/t/EkdlafKcFPvM
JsPihjbwU/CW9LiB5zd/CTqZaI16xzzmxXdqYHA2gCcV1CszObQ1YNVEaVeBgY2PxyeJQbnTZlFH
xvpic+uKuzdtKjLa0jz0OAY4cLPNDD66HVGVi8ayGrx1EoU8OmhMhXOmyBoL+PGSkWa7Di8IQAer
I/bYQBUcyK0QNYWqvb6/05QtpqDOurleDaFI6WNY9VNqKqkktzxaEpttjUWdroFFAFNHr1haZf7z
a/hHZPwHd9stnFu0VOxZykqnvHTgxJ5d/we7AHLTvccz4fmGWixcOP3vnt+CAumiDuteFfUDAXFr
RufAJl6jK0ligj0fMLC0ojhLZHZ5njbZlRa3GzxAT0ovXhK5lDF/7ADhXn+eSOX3UF3A8t2YZcWN
uROUMJQfgwJMoES8jFTm7TkuUdsz++TLg6d3L1X2jAp1/A3awAhXxYO75n9CXzG/RXKq6ZsRLcHX
jemYf9d9vyZGZ22d9MvjUGH5yo/rCpgAFV+zvjHfRF5lsNPAq3rRhAGNex7mrdoF96zyUGGB2cAC
6YliFGVwc2gWZ9251MUNSfcNcMFCeJrnQTSwZavwTnxn6WbeA6kRdDI6+T+h5d9tIUe5OVeGppIO
f7Wf6mfrHpqpCij9VpGzh8B+nABPNZ8GPCA1A6d67yHR7dL9iJGEpV0ms+5X1/UZTZANUy7oMppI
XBLNbEGKAXsBlIQvkdL72UI71Q7ldSSLogdLFOR2OjxVquwStijJ2oP97byviOR7iyhlwhM0sLNt
AMxGjfeawbiGz8Z+Vyc/SUReckler2vpgrjBJ4VYV1RUaytm4N4YEtwI60DSWqwDGWBOyUm9PF2/
AygW4+fLj3+971Ghfagut5yJyEfN977Ce3xykjCwyMRqh78FZp/4wAGokY1VUaWu8JZjWzMzKG+o
lrVoJNomEvoOiqSeqg2rIm7+ZU0CP0BYASxqy3raRoR+8buksLAVIItlwigd78fTWIO0STOCOTL0
UlRsH/wASUyDtE1PhUuoilTBMph8Ve6zX4DPSvnm8QULLjk0i1NhkgkI3jjbsR32aQWAOr7RMDIh
sh4G7QL3oa17/C3QkZEEGOYZDq9U+0l+BN43ZRZgrwk7IKEvIeAgbz5QSx+jn44+y8V/dg6uGxj8
PyLnKb6E3n0WpUHlQRrJR2YcYJ09ezZLynnPP12uex/x0FE159jSfh0Ny4cuLLHO9Thj2vZjTbw9
H2YnPVLRbXAJwRbm4840HH8atLh+eX49MJ2UG4XDR+abbpsozTFcwKME0q1QHq/AmP4HNAu9wFam
0xnr34ssvAmPeEbmOzPgf60/1+tg3NjwEHH+pSLcL3k7lBfzaEigL2vZyBT3p4fdfpm+dGcHaoYI
a3yd0VMfPY7JS3UcjQQ5RShfTL9cLFr5GI7I8+mFuyShceDGbQgd6Wg9hztSZvf39Edl8uhEgb4r
Z5lMck7cvK7rJBQ7tRs7+Gdw7gGp1KnZhWLdXdyAkMBrQ0m6ZWWn3/FmexHgu2K5DoF1GdnWGeZd
o1FT96BxWaDbD+HQ0c8F7gIF0kXMQA9VcAxsDR5LPQsapuyIQIVyx/PtKvgf8db9dSquYyzgvCP/
pC9RqRzLeHSmjEnBzfTzP1gvjWz5VQVdZsFOTXNGTsjp/Om+GS7gcCPKhF/TIXAEvjJ/WJv78o8a
pGLvgHXz9ZgMTjCzy50AnmK8cxIGU3JfduoaDf5ELcs1iRQrQDWjuxbP5BSAZadYN++Ezvb9S1sd
MADTb1Bn/7tFSCjc4oaU0jiaV0d0Kqhm+v2iH4mbBzGM9Hxz8K6q48ZRCqt7Bbl+p68MNRLE9Lz8
ZsTn6i4VP0av1LYXkzBZrn3zU0KYicaU4wNMHq1wGFMXGsu9NLtP8NPZzT9h7Sjj13g2ItJx3/Mz
QVv3btp3JBPHR0wLFo2HAhULDDQKUw1Tj7btwuavKqblj+jiPVsAYq1PN8G48VM6CbrnPG0RVLbt
yv0xpkRfbUu4Qh9eC2dprpczoyBGY2zgYqsiUhdakqqN147AyFuRCukoBnq/n6tBIMNpUEIZJ7LP
z518HPJ6lJQRdiljHV8x963O3VnlgRLiKu5BwV5wOBV07vu2ZQ4w1NP4I6gFCwZfmPOClFaV5Bgl
K2AArmD/LsQ1/8zC9/aKomza3Y026pD7uE0VzoG9y9N59BKgGzQ+QIK72RRVY5HrGgHaFefy4N2S
GDrYjwaUdNmaRT7ENt918D22dutYfoakb0rAHlwNAEeGGu8LV27GxCKAZFpKdje9sTxANuFYE+VA
88lcm9cTHL0G6qGboFVNsegGbB/XoPgGQFtbi6KFBFjlxRoGOCaYEMQIb5VyZIC4TyQMazZJPTJJ
PuDKFoJ330wC4lJxKceIpdwvDJtoFwM8DRxwmJMI/ROH9XwMuwasUnSpN06i9TCNUu6SSGrXqblj
MYEm86Pf7Bsy8V3iUkTfehsXoIh2CtrITkIscC9xBrzvzBJO0KbqERVSOf70M7k7KiSO6MVuAGc5
tAMFjrxEqZOREKCd6YyJ8qaJsZEklb/OjWVA17omyC/vnSAoGiw0c749HLbEEov88a70E42V1e2c
nHILAUD4XvZXeXzPGdpjEMhbGRHxgakPHde7mbkxPMaeqXj2BOfCYMF2WmEKy+j4kfzE/sRv7Jsl
ym6bOrBnfmycb0zIYNPRDtYv7JDKohalIlw26UZikLhyGTMRhbzbiQKZB6qtcQpRCzemxy1y8qwe
dYu7BjqlIGciFcxfWA2QHS9bu8bsCUsot5VY/ATkVHCL4YjrmN/qnItsWbRB+Znyy/1aSo6FejNc
o8puMjiujM8sQ85NBCyYrP8e7zK3rqiEAkqjTf0Qge0fg+cI0BURXgLIkZXugQI9aEAmZoj6U06r
+NCuNnnUZpg6dIQZBHt/niszdMnHne+pLlHaA0NlkiKzF8DuxPUe6ujMC2FY/3ExitSL5DbAM70+
4re62j/5TvWG8iF+ac1pfkiaROYAiQIwzpCZrLAdOSDmwhwMspSE6Xuj8nlpqDTokqbkaPdI5VYA
c7mRLi9kS2DRgdHZBq3EaYgEwhhQqb+xfgMAMvM2RixP67efBX0Y3auANynuvMqk70iNRHj8Z5p3
aORRtAS4dJVHupXRfSt58ZpCa1iRMAaCy56ocB/X4Z090/CKzW40VBH4qXjPVv4ud1mkcGtIlsdr
1T6uqzQ7oX+JzL2+neVIwXwb2u/L7DOMk3HXBmKcwe0YvkBgzMfvGl0r7VUVCa4akdsVZ8MQtKzY
Tg23iJDWaXgrVv69mzvjS0f87oftpRSbkwZF1e7hDYVccQGrtSFnh7OtwYjeZjLBjJyrGgJld9Cx
ptIp/ubP0ZjeuOYgGfbLBcGv1BEClFDpuD6MpkLfZ4EgpVTj5/jy5uy7ySaYYhVgl7fpVYGNxngP
SRaPWDDIW3sgkYCGKYh8U0IUwBqRysEX4OlDEPEjKCx47L1aKxO5m2LuQGkqf1nGxR3QShokT20b
MF2beJ10TF4IhzVED8xohjHob9PCOnncYKh45/gjSEANsV2lltRF82uqDjZc4HdIQ0nDGHrABZ1Z
h+z0Pd3UhHa1v3r32EFzF7vUMsFwVSYc6cVw7kgOrMdAiupmncm3kPochqpDoIB5b9Zx6yYMvwRC
OYVwKoFA6uqRBHrFCL665kIvrnbYyzYchVi3uJoXE+GXdRm1rgThK+XS0BWK9WHw0gIhdc2Oeavg
Fa7LzjJ8TLThzPl1bFOPuaeAoAXaVYwKH5fHzyLUNmf9KBVPbFu7fUWx9S4m2z2TEq4e3+Y2br3z
CcDqfnt+uW9Ws8DiMFtxCwNwTqmNlHmF3Ij2cOsD
`protect end_protected
