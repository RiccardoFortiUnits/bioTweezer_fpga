// megafunction wizard: %Triple-Speed Ethernet Intel FPGA IP v22.1%
// GENERATION: XML
// tse_core.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module tse_core (
		input  wire         clk,                //        control_port_clock_connection.clk
		input  wire         reset,              //                     reset_connection.reset
		output wire [31:0]  reg_data_out,       //                         control_port.readdata
		input  wire         reg_rd,             //                                     .read
		input  wire [31:0]  reg_data_in,        //                                     .writedata
		input  wire         reg_wr,             //                                     .write
		output wire         reg_busy,           //                                     .waitrequest
		input  wire [7:0]   reg_addr,           //                                     .address
		input  wire         rx_afull_clk,       // receive_fifo_status_clock_connection.clk
		input  wire [1:0]   rx_afull_data,      //                  receive_fifo_status.data
		input  wire         rx_afull_valid,     //                                     .valid
		input  wire [0:0]   rx_afull_channel,   //                                     .channel
		output wire         mac_rx_clk_0,       //            mac_rx_clock_connection_0.clk
		output wire         mac_tx_clk_0,       //            mac_tx_clock_connection_0.clk
		output wire [7:0]   data_rx_data_0,     //                            receive_0.data
		output wire         data_rx_eop_0,      //                                     .endofpacket
		output wire [4:0]   data_rx_error_0,    //                                     .error
		input  wire         data_rx_ready_0,    //                                     .ready
		output wire         data_rx_sop_0,      //                                     .startofpacket
		output wire         data_rx_valid_0,    //                                     .valid
		input  wire [7:0]   data_tx_data_0,     //                           transmit_0.data
		input  wire         data_tx_eop_0,      //                                     .endofpacket
		input  wire         data_tx_error_0,    //                                     .error
		output wire         data_tx_ready_0,    //                                     .ready
		input  wire         data_tx_sop_0,      //                                     .startofpacket
		input  wire         data_tx_valid_0,    //                                     .valid
		output wire [4:0]   pkt_class_data_0,   //                receive_packet_type_0.data
		output wire         pkt_class_valid_0,  //                                     .valid
		input  wire         tx_crc_fwd_0,       //                mac_misc_connection_0.export
		input  wire         ref_clk,            //         pcs_ref_clk_clock_connection.clk
		output wire         led_crs_0,          //              status_led_connection_0.crs
		output wire         led_link_0,         //                                     .link
		output wire         led_panel_link_0,   //                                     .panel_link
		output wire         led_col_0,          //                                     .col
		output wire         led_an_0,           //                                     .an
		output wire         led_char_err_0,     //                                     .char_err
		output wire         led_disp_err_0,     //                                     .disp_err
		output wire         rx_recovclkout_0,   //          serdes_control_connection_0.rx_recovclkout
		input  wire [139:0] reconfig_togxb_0,   //                                     .reconfig_togxb
		output wire [91:0]  reconfig_fromgxb_0, //                                     .reconfig_fromgxb
		input  wire         rxp_0,              //                  serial_connection_0.rxp
		output wire         txp_0               //                                     .txp
	);

	tse_core_0002 tse_core_inst (
		.clk                (clk),                //        control_port_clock_connection.clk
		.reset              (reset),              //                     reset_connection.reset
		.reg_data_out       (reg_data_out),       //                         control_port.readdata
		.reg_rd             (reg_rd),             //                                     .read
		.reg_data_in        (reg_data_in),        //                                     .writedata
		.reg_wr             (reg_wr),             //                                     .write
		.reg_busy           (reg_busy),           //                                     .waitrequest
		.reg_addr           (reg_addr),           //                                     .address
		.rx_afull_clk       (rx_afull_clk),       // receive_fifo_status_clock_connection.clk
		.rx_afull_data      (rx_afull_data),      //                  receive_fifo_status.data
		.rx_afull_valid     (rx_afull_valid),     //                                     .valid
		.rx_afull_channel   (rx_afull_channel),   //                                     .channel
		.mac_rx_clk_0       (mac_rx_clk_0),       //            mac_rx_clock_connection_0.clk
		.mac_tx_clk_0       (mac_tx_clk_0),       //            mac_tx_clock_connection_0.clk
		.data_rx_data_0     (data_rx_data_0),     //                            receive_0.data
		.data_rx_eop_0      (data_rx_eop_0),      //                                     .endofpacket
		.data_rx_error_0    (data_rx_error_0),    //                                     .error
		.data_rx_ready_0    (data_rx_ready_0),    //                                     .ready
		.data_rx_sop_0      (data_rx_sop_0),      //                                     .startofpacket
		.data_rx_valid_0    (data_rx_valid_0),    //                                     .valid
		.data_tx_data_0     (data_tx_data_0),     //                           transmit_0.data
		.data_tx_eop_0      (data_tx_eop_0),      //                                     .endofpacket
		.data_tx_error_0    (data_tx_error_0),    //                                     .error
		.data_tx_ready_0    (data_tx_ready_0),    //                                     .ready
		.data_tx_sop_0      (data_tx_sop_0),      //                                     .startofpacket
		.data_tx_valid_0    (data_tx_valid_0),    //                                     .valid
		.pkt_class_data_0   (pkt_class_data_0),   //                receive_packet_type_0.data
		.pkt_class_valid_0  (pkt_class_valid_0),  //                                     .valid
		.tx_crc_fwd_0       (tx_crc_fwd_0),       //                mac_misc_connection_0.export
		.ref_clk            (ref_clk),            //         pcs_ref_clk_clock_connection.clk
		.led_crs_0          (led_crs_0),          //              status_led_connection_0.crs
		.led_link_0         (led_link_0),         //                                     .link
		.led_panel_link_0   (led_panel_link_0),   //                                     .panel_link
		.led_col_0          (led_col_0),          //                                     .col
		.led_an_0           (led_an_0),           //                                     .an
		.led_char_err_0     (led_char_err_0),     //                                     .char_err
		.led_disp_err_0     (led_disp_err_0),     //                                     .disp_err
		.rx_recovclkout_0   (rx_recovclkout_0),   //          serdes_control_connection_0.rx_recovclkout
		.reconfig_togxb_0   (reconfig_togxb_0),   //                                     .reconfig_togxb
		.reconfig_fromgxb_0 (reconfig_fromgxb_0), //                                     .reconfig_fromgxb
		.rxp_0              (rxp_0),              //                  serial_connection_0.rxp
		.txp_0              (txp_0)               //                                     .txp
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2024 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_eth_tse" version="22.1" >
// Retrieval info: 	<generic name="deviceFamilyName" value="Cyclone V" />
// Retrieval info: 	<generic name="core_variation" value="MAC_PCS" />
// Retrieval info: 	<generic name="ifGMII" value="MII_GMII" />
// Retrieval info: 	<generic name="use_mac_clken" value="false" />
// Retrieval info: 	<generic name="enable_use_internal_fifo" value="false" />
// Retrieval info: 	<generic name="enable_ecc" value="false" />
// Retrieval info: 	<generic name="max_channels" value="1" />
// Retrieval info: 	<generic name="use_misc_ports" value="true" />
// Retrieval info: 	<generic name="transceiver_type" value="GXB" />
// Retrieval info: 	<generic name="enable_hd_logic" value="false" />
// Retrieval info: 	<generic name="enable_gmii_loopback" value="false" />
// Retrieval info: 	<generic name="enable_sup_addr" value="false" />
// Retrieval info: 	<generic name="stat_cnt_ena" value="false" />
// Retrieval info: 	<generic name="ext_stat_cnt_ena" value="false" />
// Retrieval info: 	<generic name="ena_hash" value="false" />
// Retrieval info: 	<generic name="enable_shift16" value="false" />
// Retrieval info: 	<generic name="enable_mac_flow_ctrl" value="false" />
// Retrieval info: 	<generic name="enable_mac_vlan" value="false" />
// Retrieval info: 	<generic name="enable_magic_detect" value="false" />
// Retrieval info: 	<generic name="useMDIO" value="false" />
// Retrieval info: 	<generic name="mdio_clk_div" value="40" />
// Retrieval info: 	<generic name="enable_ena" value="32" />
// Retrieval info: 	<generic name="eg_addr" value="11" />
// Retrieval info: 	<generic name="ing_addr" value="11" />
// Retrieval info: 	<generic name="phy_identifier" value="0" />
// Retrieval info: 	<generic name="enable_sgmii" value="false" />
// Retrieval info: 	<generic name="export_pwrdn" value="false" />
// Retrieval info: 	<generic name="enable_alt_reconfig" value="false" />
// Retrieval info: 	<generic name="starting_channel_number" value="0" />
// Retrieval info: 	<generic name="phyip_pll_type" value="CMU" />
// Retrieval info: 	<generic name="phyip_pll_base_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="phyip_en_synce_support" value="false" />
// Retrieval info: 	<generic name="phyip_pma_bonding_mode" value="x1" />
// Retrieval info: 	<generic name="nf_phyip_rcfg_enable" value="false" />
// Retrieval info: 	<generic name="XCVR_RCFG_JTAG_ENABLE" value="0" />
// Retrieval info: 	<generic name="XCVR_SET_CAPABILITY_REG_ENABLE" value="0" />
// Retrieval info: 	<generic name="XCVR_SET_USER_IDENTIFIER" value="0" />
// Retrieval info: 	<generic name="XCVR_SET_CSR_SOFT_LOGIC_ENABLE" value="0" />
// Retrieval info: 	<generic name="XCVR_SET_PRBS_SOFT_LOGIC_ENABLE" value="0" />
// Retrieval info: 	<generic name="enable_timestamping" value="false" />
// Retrieval info: 	<generic name="enable_ptp_1step" value="false" />
// Retrieval info: 	<generic name="tstamp_fp_width" value="4" />
// Retrieval info: 	<generic name="AUTO_DEVICE" value="Unknown" />
// Retrieval info: 	<generic name="AUTO_DEVICE_SPEEDGRADE" value="Unknown" />
// Retrieval info: </instance>
// IPFS_FILES : tse_core.vo
// RELATED_FILES: tse_core.v, tse_core_0002.v, altera_eth_tse_avalon_arbiter.v, altera_eth_tse_channel_adapter.v, altera_eth_tse_fifoless_mac.v, altera_tse_clk_cntl.v, altera_tse_crc328checker.v, altera_tse_crc328generator.v, altera_tse_crc32ctl8.v, altera_tse_crc32galois8.v, altera_tse_gmii_io.v, altera_tse_lb_read_cntl.v, altera_tse_lb_wrt_cntl.v, altera_tse_hashing.v, altera_tse_host_control.v, altera_tse_host_control_small.v, altera_tse_mac_control.v, altera_tse_register_map.v, altera_tse_register_map_small.v, altera_tse_rx_counter_cntl.v, altera_tse_shared_mac_control.v, altera_tse_shared_register_map.v, altera_tse_tx_counter_cntl.v, altera_tse_lfsr_10.v, altera_tse_loopback_ff.v, altera_tse_altshifttaps.v, altera_tse_fifoless_mac_rx.v, altera_tse_mac_rx.v, altera_tse_fifoless_mac_tx.v, altera_tse_mac_tx.v, altera_tse_magic_detection.v, altera_tse_mdio.v, altera_tse_mdio_clk_gen.v, altera_tse_mdio_cntl.v, altera_tse_top_mdio.v, altera_tse_mii_rx_if.v, altera_tse_mii_tx_if.v, altera_tse_pipeline_base.v, altera_tse_pipeline_stage.sv, altera_tse_dpram_16x32.v, altera_tse_dpram_8x32.v, altera_tse_dpram_ecc_16x32.v, altera_tse_fifoless_retransmit_cntl.v, altera_tse_retransmit_cntl.v, altera_tse_rgmii_in1.v, altera_tse_rgmii_in4.v, altera_tse_nf_rgmii_module.v, altera_tse_rgmii_module.v, altera_tse_rgmii_out1.v, altera_tse_rgmii_out4.v, altera_tse_rx_ff.v, altera_tse_rx_min_ff.v, altera_tse_rx_ff_cntrl.v, altera_tse_rx_ff_cntrl_32.v, altera_tse_rx_ff_cntrl_32_shift16.v, altera_tse_rx_ff_length.v, altera_tse_rx_stat_extract.v, altera_tse_timing_adapter32.v, altera_tse_timing_adapter8.v, altera_tse_timing_adapter_fifo32.v, altera_tse_timing_adapter_fifo8.v, altera_tse_top_1geth.v, altera_tse_top_fifoless_1geth.v, altera_tse_top_w_fifo.v, altera_tse_top_w_fifo_10_100_1000.v, altera_tse_top_wo_fifo.v, altera_tse_top_wo_fifo_10_100_1000.v, altera_tse_top_gen_host.v, altera_tse_tx_ff.v, altera_tse_tx_min_ff.v, altera_tse_tx_ff_cntrl.v, altera_tse_tx_ff_cntrl_32.v, altera_tse_tx_ff_cntrl_32_shift16.v, altera_tse_tx_ff_length.v, altera_tse_tx_ff_read_cntl.v, altera_tse_tx_stat_extract.v, altera_eth_tse_std_synchronizer.v, altera_eth_tse_std_synchronizer_bundle.v, altera_eth_tse_ptp_std_synchronizer.v, altera_tse_false_path_marker.v, altera_tse_reset_synchronizer.v, altera_tse_clock_crosser.v, altera_tse_a_fifo_13.v, altera_tse_a_fifo_24.v, altera_tse_a_fifo_34.v, altera_tse_a_fifo_opt_1246.v, altera_tse_a_fifo_opt_14_44.v, altera_tse_a_fifo_opt_36_10.v, altera_tse_gray_cnt.v, altera_tse_sdpm_altsyncram.v, altera_tse_altsyncram_dpm_fifo.v, altera_tse_bin_cnt.v, altera_tse_ph_calculator.sv, altera_tse_sdpm_gen.v, altera_tse_ecc_dec_x10.v, altera_tse_ecc_enc_x10.v, altera_tse_ecc_enc_x10_wrapper.v, altera_tse_ecc_dec_x14.v, altera_tse_ecc_enc_x14.v, altera_tse_ecc_enc_x14_wrapper.v, altera_tse_ecc_dec_x2.v, altera_tse_ecc_enc_x2.v, altera_tse_ecc_enc_x2_wrapper.v, altera_tse_ecc_dec_x23.v, altera_tse_ecc_enc_x23.v, altera_tse_ecc_enc_x23_wrapper.v, altera_tse_ecc_dec_x36.v, altera_tse_ecc_enc_x36.v, altera_tse_ecc_enc_x36_wrapper.v, altera_tse_ecc_dec_x40.v, altera_tse_ecc_enc_x40.v, altera_tse_ecc_enc_x40_wrapper.v, altera_tse_ecc_dec_x30.v, altera_tse_ecc_enc_x30.v, altera_tse_ecc_enc_x30_wrapper.v, altera_tse_ecc_status_crosser.v, altera_std_synchronizer_nocut.v, altera_eth_tse_pcs_pma_phyip.v, altera_tse_align_sync.v, altera_tse_dec10b8b.v, altera_tse_dec_func.v, altera_tse_enc8b10b.v, altera_tse_top_autoneg.v, altera_tse_carrier_sense.v, altera_tse_clk_gen.v, altera_tse_sgmii_clk_div.v, altera_tse_sgmii_clk_enable.v, altera_tse_rx_encapsulation.v, altera_tse_tx_encapsulation.v, altera_tse_rx_encapsulation_strx_gx.v, altera_tse_pcs_control.v, altera_tse_pcs_host_control.v, altera_tse_mdio_reg.v, altera_tse_mii_rx_if_pcs.v, altera_tse_mii_tx_if_pcs.v, altera_tse_rx_sync.v, altera_tse_sgmii_clk_cntl.v, altera_tse_colision_detect.v, altera_tse_rx_converter.v, altera_tse_rx_fifo_rd.v, altera_tse_top_rx_converter.v, altera_tse_top_sgmii.v, altera_tse_top_sgmii_strx_gx.v, altera_tse_top_tx_converter.v, altera_tse_tx_converter.v, altera_tse_top_1000_base_x.v, altera_tse_top_1000_base_x_strx_gx.v, altera_tse_top_pcs.v, altera_tse_top_pcs_strx_gx.v, altera_tse_top_rx.v, altera_tse_top_tx.v, altera_tse_reset_sequencer.sv, altera_tse_reset_ctrl_lego.sv, altera_tse_xcvr_resync.v, altera_tse_gxb_aligned_rxsync.v, altera_xcvr_functions.sv, altera_xcvr_custom.sv, av_xcvr_custom_nr.sv, av_xcvr_custom_native.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, altera_xcvr_reset_control.sv, alt_xcvr_reset_counter.sv, alt_xcvr_arbiter.sv, alt_xcvr_m2s.sv, altera_eth_tse_phyip_terminator.v, altera_tse_fake_master.v, altera_reset_controller.v, altera_reset_synchronizer.v
