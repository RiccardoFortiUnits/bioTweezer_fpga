`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FIpkWyuatbYxdq27kcP60dNRSknLxXn+X89/0oi8ioHE4JcCxvj4tVu3wCbRrvfz
nfoP+Ir30Z/hAOo5T9X1saBN+yyBdtqGGcfHwRDYYhu49piBnV9Y9f4JjnJmeGNt
ecemKdc0F9WrX7Ms/R4eGrPdRMBznMCGPBBOf/T5rgw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9536)
ubnABvmwhRdSqhnJIpbjG8eZELBhu5p1umdmBZ9hxnVHnKov+8U1IQVlYAMXQsv+
T5AIGAK0ytr16BRBZs6OxK99R/GyTuUayT4p0hwiSWF+FGgqXXLKFWUp8lO+bbQU
sXDojtbL7kZFSQpxgVRgmy6USvIz0XgQUj5axG+YGdt5o6ClwnAvuMqKtxEsnDK4
FzUCXWuUXiHCxaJYM3iX7L/gulYPsT7ESMqxcz0KSMdxm0JpzwYJDQYkhMuZsaat
M+ebJs/jVsUQTcYSa6TryqIksv+wcNOMMLEzr2W/8TRKQS4zX799NxxqBSU5yh6a
H2iebZeJu2UpS1+o3gRfnrFyqv0SMR28+Dy0MRwB8QeEljpck01sBqmkYgb32PBz
2VK61b5r5k59lOS7DyK7WOlxzsRuRVLTeEZnEjYdCxFxQv8BHUWWz5NwgtWJASnv
nX4STbZULdQMiD5EoSKkpEstuzPtG8AAMqGF1E5LvT4bIggwUWQKmDYQQvMQARgf
3ApmsI9kS5ceqGgrEEccEPzlZEli0jfxkl7VtESrxWVn9Lxqfm9Vko+60yHSyAHM
MCPd35Gzh55UbkPqSmjJn4P04R8jJY3t31+2x4miVhfyfdjTtcivTK84PABG/Hhy
ZX0AU82bVl+vsGatJtVjlUMCxQUQU9SjznUxWmCdER817GRTwuZjekeSwM1+AGW4
7tusdY3HK1C7cgRVFOxOg9+dDiqwNtITqwq2zTDVtf/52w/LVnGIOioPOyps2LGQ
zefnHHn+zornJj/fjJt/rl2TjFJFDhAZHVDxeBQldE2IM8TXuqq2P7g2IMPPkzCG
e7f64ksdu97fjFbgVDg4TJqYj5naw/C4XUvWFPr2XXrDfmdHbpG7s0AI8jle+/RE
8eOUGkpiVcigx+SW3kZhfU+PKRrQRxV5E1Qkr7OcCYbJxivHq8UCS1MzpfpU1Jrf
Y3cqNr4MwGFtkLPTvumtSQePe5sa7wwKue12Okx5x06ukogfx+gUWAWztijv4gIy
lAFXcjfHXnWw3GrSyylKFIT7GJv6kduCIUc0WAVJGqKm4oyQc2t4V4Y5YzL3K2Oc
3g/aNSWa/v3GSnarLOFmo7oqXTZ+bNl5uC6hyhKXYNMIyVt+CIHGMpCT2N/7T7S9
ou+VYyV/0BKrnIHZXKA0d5ssHf/hGV2VV6cpckrEcX+eipO35UfIVsEDDhQzLns0
3PlI8NxNW9+9D9L9W1gUn8r8zVQOLMinChwUir8T66Rzsatg7buTwRjsyvTOUjuL
4N9M8FrHNwQOGK8NpbRg0qe2tyPhwobAvsG7vmwnyGnvsDHRe9z7wQ2th074m/jD
BnZBXkEUGt5VfE8fD4cYd9ngneWFxC4L//fVzHZsxZPkMlKWTwDE3lycYumCfI/e
lDB1mEl/hOLj7CsIlxAkQLCDOsY7lWQopqqwRJYnP+qvrNJ+fQSBdJ+UnKqQdVI5
8s92NTT3XZnVcgP5DdCG68HhkYEJ8PBoOzrvIk4gC4v/nzCzf2sAKHYnP3c7UhP+
6ZaOXMzZpcjrNbNeXHJ+zGkWR+RdZyk7JK81hiQcVvf8a2DlZouiOe5dDrF2ORcK
mil5vzNwRlkPbjejEp2oVOseYe64bMjEQkKkSbDKoMbPV4GM7FAX1NvTyyv6KY6H
bRkRgBm6AnK03RC5UU+5br1Aw8xJw0QmSUNBlTIc02JRhN5GuIZfmC3mLAn8f2l1
f82XaMHTZXp29hb9FW+hmrvyjZfjBwFtchu6rtGGYAeFDhiPHwWzEm6n6FwBKvzK
s0O1y70KGV3kSQJizuwhN1yBDPQ+GSpVyDARoP4SRCyiu2ZVmZEI3WWBFHMKrnHu
ietEPOxNn25TiPWQ8FktAHSqKM0QHX70l9ooTF7+Rf9brhUN7HLpu/Q/qI4Mpei3
kJzvKW64Yyin/NK+49XHey29GXzMMYVthTnUVSOtUlxENRgffHNVoYkj+jj3na6n
y4cFZnLW6liHrJ9OGM9xn+mE8zmWn08X5W5l6qrWhbVaWSEfk0V2QQq2b0WUNaDm
mTl9jyC7xtFAl7c1nZMdRZgsFkmXIzRJgV2H0nlkILIUQZxnoUW2H9G+b6ERKV9y
agGlJL7mtbkY85MSVYWNzYXJUTdKqXI5Nd3LL14wWQGHcd6ZpA5VVNYww3gjHPgj
3dleRhuWtT9+NiMCSPj8qORaaqSAWnEsdkMsKa3KQLqFY+MxuKWbxrP27FXGw2NI
IBawRGDHrv/8kixVPnsH728ea5kfKYLVSg45bOm/q8lCZ/xznLvtKNJlgx7BC2X6
GEybsA3kgExGY6mzs+jrnvVvT4YBOrhXPWoNM39At8DvsXtvMt1R9hJrIRC97Oq1
Q9nMGyWSHQ091V802TqyS+cDZPWGqVhBWNni56OitN+MUocNIJGtrnDiQF/AOR8M
xH+dmg+WSZ3V2zrzopQ+/OTFfNIwqNh85d7MRYOe6ZZg0frspmaV4pzIqOsayzVT
qfns+jqzVH8JYCMsiG6zIx6UGlTkqvLhV7i/SGWy8/KBVNNO8jP7kCuVTaOK0wRH
XdFV4323YnSOx0jkivubbNd6oW31xO6CtQ7FAG8s4xd5x3dmYccXLToZRNbFTHz7
5HVjKA67vd0nlubjtoV6cp3RbPr8rVakwzfUnz7BJ33U/lH/tDHTkNhQQzcvqbbl
0OS+D3NGGFIa1IMhDzT37EPgyaWd1hUN3xl26JaAfMSjoo0/85yEmBTI3tDJ61Mj
abo5KXhKFobreOLhg1RGjTiY1WhF7QMvrAnP6XwPGKi5duBsfwuI2EcueHRA2Mp7
sbt5UJuv/Chx4yly/R8oxXYzxaLXOYzodtmVA6+L6ewZxquFGUFf83/pSGQUW0if
C0vet96zK0hD0n+eoUwLdsONN0/eVp4M67cj7qPKyQUDG9t7iya5nBH0Meq0AVpO
6uG6ARApXOAf9r9J2YBva9GL20o3N+RerNXAbNvvXCS5V+I9UE8pNTC6JTvTG7ID
yXbUtKaiGvhD77EIyqcRQ/rZ6DgdTAdOm+7feqRnvAs7GQmtZxemXWrWn+YYoqZt
NdVuN6rB4WRf3yyeD5JrYz3ORmGhEYYo9bK0/cRHBrmEDkg40t7lI3XLP2bVWtHJ
pTDDCkygo2nrMxrIh9H8Dp4ImC9RlQ0/JkrqvKcqtldqs4jKFrHqlYSUYdBhOcbd
ZgVIHOHqRBUCvTN9W0hoagD6mMB0uyxdIW+DwHerCN2lBVTFmBPfNALntQnXidXr
s/CuSqdSD3++Zq+lRgzFMvDQXoltMLNPC8RPOz9trGsem8kM3L4kV8Uk5IS8uiTE
AS/C0REOdXTn7l9GnhE8sbXERuMLwqgYbemszK1XCN2L/uyf8/n7AEkyz82SBeC/
43VYfvo1E0tlFbpY/kiE2yLyVLEmgWgs27FK/NW0wgcitcqQATYMc2pxCFb4C4l1
eOFRnnMxhbdIqe1cmigOJluevFFH7g5FGBwEzcz8Y3eADiUDYwEmI+qnIdJZn+rt
+KQc17/O82fhpDYTyUHl+ty1uWfo82uy5XMDdKvZDxRzmh97x9kRM5HEzY5PgQlO
ISiKpjx7e6ADBvVZ1bBYqc6taIEx4EF5pcYzy8jZ8S4l8/wvw5tBXPpS2348XPr7
x9C0ptx8G2C1RTm9tocllh5bSvP6JySs6z74a4t+/O1HfFOleKIjKtO65rizoCtw
tdb3EAQWVMjwHVSUnFp43FzKReog8W3RxncIdU5SySOjmeeAti830WBOqJCsd48k
emQ3b18z89zgvxSg3VVha3wTq8XGaKdT7AkQ4ZKk5kDK6HtDq2byvAy1HbaN8rax
eR4DVKwQjXwn2zeu/Cp6iA6Q1B+bYZOgDrLH4oT1alFc3IZD5bwlwbr9/Tnf+MxY
kN3nOp6od1YuNCHHGtI5opmnz+E0d0OKd4Q1B3RnsIsASmRwArMcc10XsNZRxj6Y
kHmTQYhqP6CfQ+3LlJVOoG5Wd0zYZvHrSIIgVGwtMLJFGYUZnQRYEq5JON9jiY/R
Gqjo3b0jTSX4fwNw8v8TW96WGxJrR/YHw9MAK4b7xyv0An3cr3+xKOdZmIvQud6h
JfrrS9npX1UFT12Y2PPzlO9FJQgJIAy+sAtWmhNr5Vqn9LRi9ZoRxHg3ukjAdPEX
B2g8LwrCEl5HHNcpCSZqQidwhIQCoYxnoUWvUHyslrkrWkT6S1jiXXzh3Akh1UB2
sXDrhJXBvGIInajkujCxY5KSzxNYigyK9m+mqtR77iWR0PO+yY811LvWHOmVXpeX
6EuLz/4Ao7Nrz5SMT/bR1cVc50KthzPFfjLhjphLjwjaGvTD/YaEN1Zn4WH4G/xb
mmHOu8zBhgIGHjsF+oJqcgUvPRozibv1T10zcx/ZjW9xu/TshR/6Si+mp63+C+Os
jRvwtVbojwGI9sp8atUGB/ZrR5qXOG51wMKs5yEN7nf6xVabZTmmpz4wugp9pUwq
kmMthRyUt5hiHpXt9CVBoiyZOJlwZtj9L7gjg70dDEnSwHMrL7yaiyhPtFTrbo4o
I21C6pcmcBYx731ZaFpiNoPpY7WQq52/BTFCa7e86t4c8PkEeLHuUL4OhMstKcYt
P+AJ6kR00QosdutfEsyy1syet5iOUDCF37NM5sNQwpHa6W6lp0bSiXhWUJJNIk6c
z/LjoaZ5Cqp9hJ4lcdICLrxlNwpYKxAsArToQ83ce8E4CPDWheu+XIP2qeu6W3l+
zs51ehUG7gclLksr0nmAB7QggqN5Hq/G2bWkvlGYTVfkN/+zRIcvNhrAnpbXDsUB
Zr7XFvsdxkSdpZBOjgPqYNaBAMqfeaylp5I9pJPwsQNIpJ00AilTYEdOz3yFwKB3
+ZL7f31kH/FTRuJMeeq8qFtRRYubgNRC9lM/TRnAA80fe+ODR+PQ6FlFKMQ3GDe7
rW67tk2G6LalPFx3es3wj9iVI4QHoH3sEMbPXnoMbR+RW+JKsqRWycpIchmj+fl9
prakw24oxe0SaO99EWtI+f+NyVBVv0brdgvHV9wVVTtR2+i1MCwXkkH5WyvM+SgY
NXWXgh2wZKHwm58zxCVLn1sAZQgFT5NIlTdLKQpFOGa9PHMnIA1dJOwF1kTTGBcU
gsetyc4bd1xHl8/X/eT7m4dIqUPp5+I/uLF9+Z0i71e/Ink1LENxGBchkrwhFlZI
0/WAzGXE6+GVrYcFT+PjEBegY92XWw7cJlY73mq43i/mQMV+drYiTHeAMgJx1jws
fFN1MmRmzuhbaagHCjkxzV9DyXOzYDkHdB5U5m9fxhmNr8O+hnT4knel88cy2AVE
gOPmjNDeNjjlalREnxWGNOyVCwHZrXvxCYfHNzv1an5u0bb3F7TD4bntjAioqk2A
A6zwS727ADVR8yY5LFt9mpgLYtQxke5SmoCOPwcR6AYv58D6cVP1fOnLSdNrOxBw
F3j2L4L2A9ZbL/8Vgx8VzlEm3SLH2Q3JOlo8QDNeRH5cl4TRqMOzMAlnrL6tBrsG
23KcoYU7OtgbPz9tfR6feUiX4azvCybIhPLQZFnyKM31OAOJKhmXfZYtrJFep1u0
9Qd7JREyJSW5A/1+ZTtXSs/tapdDJ+uxpQIw4B6mmObxl7N7+4Tip8yLdpofbB30
UpUNMrI52Xl6qNW1Zwyv0H5nDlQDRfYkoTeJTA5qJO2myAQzwoJJTVZhliW+JUVZ
3Bt4aczRGB4WLOgBfYuIjcjvIeExu5kTWLnSyL+1IRNEalOIwNdWgHic8TkCXQHk
6WVm5cMYka+3yLCY0BD2VtyxDdPkULYBfqW37Bim/9ELAwqJeC6vpYRf0SfzRHC0
g+sIgFmPPHnPRUpICbcxw0HRE3l9KWSWvwEuwudFgWIpURPP8P+cJriP6gwRK4cE
K6Q0vOq49V0OHqeFubwJ2/ydbIIAItpSNFNoB3T11HsHivuP8xF8x6/a5Q5Uew3x
vl5IvS+PFq0eQ4lSKH1r5DJeb/ge1775+ycvLs+wuo8pi8hzTG+ve6zZrIK2gSIp
Kmgoc9G/dDWQhVXGjnScyuQRXOHfb78+rGJydOYQsNp3Pu28GyuMmSuExBXB1I2b
tYzCcDY5Its4s5PIjr2K1kiiTc7XPCzjSPFkjnWvvibRB90mBkSXuGk7sESJ2MUx
+X1H/ZSnmITdg3/uJGpc1ZrsWKc+iD09Dpw83BerDVYxjXTD9Q27fZL9Z+OaUr1G
/Her1HE0+EhnoMjoW2ndoBuOnrOzcrkeM9Yvf+ELwZuSK6TIQK34s79yXyoqjBj9
d/OTsJxOkHWtt0nMraHRc3JuEuHs5jm4IsgOVMC0Cl3yIaC7vjGKtFD5E38Sw+yW
CEXgb++s6OxxG64fxnYtreZ9gWtJACycEj8Wm1W4LtLuoElPLTz5+cNhYLQtD+9Z
Z6Rn6uPBXfPZsffWe4Y6uXVObyyqa+ni/MAzXk6iHj+QSiZfT8lV/gy9UDejyVIS
fnLtIaMrrg/FIeNFMM7g1EnJ8xC5CSFTGRv+QSDBTmEu/qwbU0rJ5odYdokJaNUb
EzpPfNPVOEEnLxpzkww+P712eELaSwvTso7cvlM/PA1Gp5Aw+vCN8y//t+5E1ieG
f/9mmvg6BmYQ2CMliwnDr3WHbqQlfk4zs3eyJlgf5tLst108z9AgJeny/+NVnmae
4c5ufLnJsJm/qIUmCQg3DGu4jMkhcJzCXa/8nTsc9axxOQnBiUHiZMtzH1hj/J7k
SPPshd3do32ecqoG6QG1RQDZvNsYquY156KwuEIofLDQuZDJzbAhImdUS2qGiH7Y
MWlR7JMhP5V+rFrGwi4AXcLKVCYlZKiW+gEHyMel1mw2Q6I8Zz7fWucGpxyDUXOM
l37hj93kYDz35mO2y38gkeP7KWGJMFOTvffQyLNj83pBdD+QMpCL4KjuFUFvmwsD
ztXDzWve6XX15laB9nesG1xlBzkxtmS8bohj6Z9MAW/taOHmrQ60HlLrcvtUANwe
AjN5hskHWLQ8j9BFQWDB1C8fiykPDrbE9m0+eWOgiwK0EHXAzDmmu5i24WzqnhLL
jD/b+83LA/wYC/Blx0DQDtS5i6+BcY1RCxKLu8pY7WbKwln1Nq62Lq/3QaDqsiRD
dzq5guKqmTpKiOSfvjeZhIbYyFFgP1k6ivtky2mGXrHd2zIF3IMOJ2NBxNOOBSN9
5iSoa+GhvC7cg98sCPrdeDx8qMXJYW+b7nePb1MjE0oPKIFg/ph2nHsDhe1Xkfkx
3kynlCWIUG/94yaFXpIlZy1Npn2BA09wogYBB13GYUpBz86oN4Ry4lqvHTM124hH
qJjG+SZj+5uWz05al4JvDrEssV3+XubrfofjVwwUD31WGx7KgdwK1oa97dj/8iew
s8hh7CEbM0j8oB7cQ36PotI9eAicAgvTxLSsdp8xep/zIpiJXVFzuKlSCZEYDZja
Ed0rec6uRLOR4LnEVHhGIldYIpUeIhxHJV4ddxZOwI9oXWCzplldcBk+QOHXLvmd
iuBTTlBFYShhiZ/BLbnDf2IcBeZne+d6RRWALSL49Jauu6F09OoBu2CoCu8jYBYS
hUjLY3IFHiKVYO70kmyF1nrn4ph+lkOaNexB4l7ZPYBzW7f8qK4wR60ucQWh5zaV
KUWxiqMUBlqUif57IHbj9NS5Gt3YzTQM3fT0Eb/AyICqOPtrqbSwfTSCuw3iZa+w
f4Z26iYU7+hUurJ1dL0XN1Vp6LpdKdBI6zRNwu7pnClXWAU50weKxYCP8YgL+fYf
p0zq+3/VDnzfymQ8GIDtblVBMC6zOhGA3KiNC1sM8C+1mlgvc0crMEc4PI0h+Qt7
M9PTRC/fst+MONXY/oaKpu2+aQVoYVA/apPnSyN31W7A+J/0vfeD3wI+vFh/sJdM
VRDC+O6d7vDBC+rqP0j/PB328z5gM2vllrGgIroKoK5X/eEXgzrg8NLTZyqWjFQu
/GbTMthhGk5fQeaDwEhqOMaIQ7B9QD6wr2wjTRLPShuBZiWzse0kwzoph8XVpSv0
wKoe3Tmfn8AS9qGORkyPSe3txln1T5rSWrrEdKCqTW/wRgDVOQHh6mA9gZmYXqWC
vssmy20EJeDM+l4jm7+Nm0tZ58ztMR1v+8vjC1vMuSSUlqoaJ+xw1xUCEWykhBaZ
/E3g7vOzxdNpQn81ZDd1lhNOYpUGdezuKqx9kUtQXgI35kyrrgJ33vLjDGXhiIPY
bbEL3CdEvlRPV8ql6rvSjo989cr9+Ae49x0MgH2FzSP6j9mA9ien8r5Nk+GTfh24
Xa5LHJhxae/U1TbCjfglWVGviZK/tgXV+acJRd4DnEqulPKldQXLgVeFPq/hh0kR
OcugqHBzCWVhR9qnFlEtLiX+JJIIUtVZeLAw6vYyu6QJphNeseRiA8tMkc/SdXUc
KGy6meJaAEr5EF8IWQd9LXy7yCT0yOPrCU7ELzIO3RScu/AiyK8hxa9ICWlX5/l1
iEmeyuBMm2mYLmpDTyK2O0knw6hCCvg5Rw4rx4xdjBSmV/mkp1GnTEvzq0goPiCw
Wu20Ah+ZkRo7kvXjoyOISM9pp1s15+VN1uNGIbrqmN+BrTULl5aVhmm2M71kkheV
ozoLr2DfmoxQdtPQAXG6UG9P5Nmd/bUAIG1B51UbfcV7KnpQ7EpRInm4cayn3NyP
m41ni4FruhWbN4021M09GaJg0piGRLlCDAujra/hFzlZMDgX5ZKfqueZwXTNRHP8
rdgm8NlRcJoApWQypTtu546O3xDIliwKvnstb/tPoQ92SQGlStEkkvRRQvojdhjc
zy+4sFXwLzTp4sIFM8gHSIO6qm3D+uyHhdHPj4tOEgg+ksr+ycKaV+kzL+sgYWxk
qafdsxGig4WQxvdo/xWAaPtTy7NNpBzVFpl5LN/QwlcPpWsw0Y6vF/UTJYM6jEA1
5YN4ZFseR3gVtMGesSEYap3vYd0CYBIu/luMZR7yPhFZDLCU4MC9Xy9pdPwgEUzA
5wHScIQZZ5qxhHumrj+ThYPSm0mBuKzQYKi2DyDXQ+rUpKEQKLtQW9HcUkK+mbko
RP1FH88lfmatPy9aXg7/NQUzmTrzX8RHBo1alf3eCPg5d2gQJy3pHIcJ1+f5GJPb
JqNZpKNcmYfCz+LH9Jo8Z30A9MQG8clffe9+eEdL8D7BKv/gTpu2aNxgf5orPfJJ
0xdBc5PgPF7D/4A0VTXxfX2ruN6FJNpQ1rwCsXs9SxUCu2K0HQIrJ5ySfCykwnhS
9fZwyAtM+8WREo8+rDYGm6tljOO6V1LAQnsnGCR6AZL55jjVZAgOYWJ/EvtMwBtx
3/eKfv6kxnZ006xK2J00OMor/Hsa4uZc3iRZm9maeiFPJ+MKZTENAFOQLqj2Pb7Z
bZi8hzFkxBthDi+EjQiDMx8Qcly4olp2hwur7XmT6y2G4BuKyE6AoZ1y++Aahpza
UWfezNmZrjpHLNStS7nmpoaCYmW8xeOX0FFg68Ds2UPjOmg6mXyJPdY1kwfNuIPl
goFMyip/rM9qbGH0+v+NussbPsOqoHaFuB81jtUQ+F6yFoyIEYIFLUoUhUYXOO4n
SlomHs2PMIuM7Wj2GBoOpnidV6fx43aQDV25YHH6FOmdpT8idKh/+NhCj4fuS3nh
DxrTKL3QRKXquX98SVKKOu+tk0cXvuzMl/kh6eDzhw1Ya8gPILb6xCylUWtzHeKA
RDzXHh3odM7mpdK8dWfaJl3xCezI4Lxq2JAMNOzswLVXUs85UzyReDb1KckAeipe
fLG8ttrp12i4yCdMP//m5qlKkn1ANFV+/PogP2fB1J64orUEzj5HbOMkyXGL03ye
j68gCu9wGKElszBajr4shq0uavMjGYeeCeBL0QaTejmRt+eAv/ZdOzHgnif8cDky
dKYMPNH/lWyOa6UYzi/BIPLq94OIf+pYnQIdrUgs+a/jlqK9pf9a6UBh4r+cNuPv
Xgr8LV2zZn1QXvKS/m2T6u6Gk6X35WvOCHTdnLryBAwq5B8A3CI9m5qP63rmAd4s
6mcdaWwRxT4dg7h20BBnlpfzfR50MQTFgCI67qOFwNLttOUJJgFshlodTsn4YT4j
y7Oj/ETejcRL3ljCkwqNWvEqpivifFHpJdxsdMy1YB9CGHDayt2pkNYDQV9aEU9b
tcY3xxlTWyTjXb0rq/7ieSyovHzFakjrIwXG4u8es/Ncn4wcRkwwfE1NJDHnBvqi
dFBIacf+jB0K1bDJcDIVJ34L4YwiZradu5tjogy7VSJO+UCRJsc1tHiWjIbKVSw3
M+dK/t+mGsbIwi9M8nELjfPDZwx8mjsu8Z8IQsTWR+Hi/l7oESuyf+qz0XCGOqcL
Oc6CYwzPqt0NfNCqPATrqS4q9WlTJQfVSdzc8gPC/IMGXMKLGg29rPMwsCNO3GYc
TSduAOkyxWF8E7xp17Qfkouyu8JB+y7WaPcwjq3FMHGHcO39/lR88nUvKy4x0cUK
MSYnxACuWMVouMWZWESVi0kCf7uxXXEayPTFFOtGzdYueQpZEnxy/IwML+eRoisC
x+E8K6CyL3r8/MXYuuF2t9M6rlqe6nLvwKRUHT2MX+TBNwRz0fZsWe6rokHLE/aD
UepaoqdCwKFUNptv+o6S/mBbVjrgueXUP0ikt8m1yCUkCGtjuxHMLwnKkQvFqVS7
yWHFLltj5POYwYxqvH7GxkwsnFhakqCr4qesKxJ7rmjvy6a/WANiQyvVP+UU5qE3
vF8IZbpuNYJuthi2B81EW/7iIRYKkKoaE7NLASc/MrSHsE1io0AmEWc2AenR/8rl
WGLR9xHqGBow1VzY/IPGYfIvKlwUxBc1kgpR+Ii839qtKff/ktqF8veVfTv+lWoD
ZTZkGg4ssrYKKj31ib0g81BFaDw+UyqUHHe5VUl3/ZdqEsXTZyupFNbIWlK9t9o8
7gO31KpFRfULcBhNhabmawprZcsVF/oSIEeZYF0MhMFkEvS6EVCntxTQmqpO1Fw2
9Nks4zkcfWQ1INKEX6vFEu4ES8GO3XXv+prAAvuw0VmZE5VzqEH4Fp1YMcz3P+DU
EgaB2SxtzY+DOm9wA5NVzXIY7bb0cvSvWx/IVftCNzfFHAIgAdFcyxG9gru787am
6atRoOWwezDiX65VaKg8bkQr44Ufec/dhb95qFpJLPhmxQihjQgSwXQVesO/7lRj
WIGnta08QW77PgAWIflrDJ3KcqrkU7FA/GlUBAKm775YjPlP5hTAGjWA2VE1yYTM
/vmG1TRMFoxC60yBk7pSAbK8hoM0aaRXPZYb3T4kRzrbyQnMLEBjS3lO0OqkRUdn
uRNrPS9wM1SavHvfLjD5uHC2eEpzIoAp1Ex/6rHqWe7mjCAz08nFkxP+XKDuCeWY
fFYrpBPtu+4GXlg7rob62EKVtQ8e8eeY0ro17ZCEdo/9mi9HYGsCn8sVnOdnkggy
C3YNIS37QgFzv6vhjDhVLyIOa2X10H4/USVbq+uwEMpUGRBlETnLb0dftqBx2dud
MtlbNX8VPwvHlVyUZDn7Rua6ps0ubpoIjRIWJDtZGdS5+mzD3m1Rdq9QFU9vBMqH
Ckdg7VZE0g/W74w7uahHRfg8MwXOW1XmYGSMw4H9kq1aTGXxhKCPEJUZx3XuFVyX
K+VfAfkThZA6Dea1CUqJaS0xYdsHWhED3HXhjSjwekNVI2PrE91i8Y1nzWeRtlLO
2clZkna1tFpQ0hXeSaeBfxcoviG0ySHYh/I+H0YH095RzHFZM4PHBYogU3MHRna1
Vsqwp0+jd5P9uoFHuBDJQjL/1k6u3z2kCmUfjsTAsyqw/vkUHmkW22tuEfCICqLk
npIUld+CB3HkGgTQQH+IzC/civDicI1e8VooYqNIz/d3Ktc6O6XipvUTOMij1cwb
1W/wjTwIMUDBOGWLXjVhyuDTsofWK/3BxWlrDKURDPbwbnDiFR9JLbC0c2vSwiBB
x0w+rGFTs8ff7HL/H05gVdfOb2OOhmEp5eYp6W8E8hKxhYOTCC0NQijnVudFElOo
tUBHNcli4M4/paETxn0/1KWoyjCVNEP2jb+TKFxOI5G3aroosutW88kgWV9tIsr3
rwUmFA1/Pv3PDkB04hPbfFmh4HOeyylhnELC7+AnKGeM5j/TOxhRSw+kCuNviJrG
SvD9EbpUiqIT7MfgxceZDQVVvz523tbBD6UmEyJI6S8Y/Uz4Vfxw+ixCosMRXmlJ
lpFcJHVuzoJ5LVTaere0FPyQXAbiBYKMPc1S4ZCrtXfUuA3w5h3a7OyrIy1jaz0e
fIYvVZxszIcmgzAB5d+VT+TEEEQYzdacSu3ArfH5lWPVQpD/XZLDEZ1kFTv/ipEc
ksurnyGI8L56NhZajOAmSqvwexlh7ZTdKOW2epn2jLWMKpY4i6bhTzJJJAc7M0W2
RmvnB001v9PxHVANN8c0oDfaI9WFfFSZ5JT/m0L3FvIvbhOlkQKrkGixhbxluuqN
0P/fobql9Us92zk8Le+ZPKxhKiBsJKYWQWRGTz8tdqyF4UuraT1uL8SQQRH47t0h
qf0SeW7Z8udnmpf//XJmQfCMjtYupbqHAwQAv72J6d/sMKv0ByYftSWPCwefSJqE
Lg00FC6SHk20MkKuHSo5TILs/PX+ia0aPTTAebDt9PAM8zEgJQAC6lyWEVa1GYM+
OcmbOwgq3ddg301S6CjfxnxReLFghk4X0capX/bxBIOLPdlhWp8w621YUQOOr1Hs
r57DAxx69JTBrqtW/HvAJehefJGV2tjCqBL5TY86foE=
`pragma protect end_protected
