`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GA7X0aTNrEHPsQUsWWk9hzWgw+qzefVXhY//Nr6GpRRur4bQGpXf1rs1Vo0FkXDQ
5J49Dj+YDLVkmf7fScXm2bgeWXVq31OrqgfUPRkHKZ3QUtgVYi9ip3GgJ1N6mHkO
fWhVfptsjI+xRGZFC9xnCTyGVa32SItG43zdPNorN68=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9184)
jIE0eJP07RB7rOfNLSdKxUPpKzi8aoNG5RCTdGNgLo+0LZ2S+wU/n5KuSkm8MgUL
t7Hq5rsxJP+LCK0r4nF/2sljw2Knq8cewAY1k2I46bSih9F0KNB457fgWvg/x5+U
YTDQEkKqNS0Djbr0Hi6C9dvYwKqgL9zFI8HTHS48g/85+bdPD3VpEVq6YtEd5fjP
e+pdtJNXxiTXIsoYYVMsFtn2jVP1pJ6pGcqyUVw5eVAHy8ljexS0XK4sJjoPUrZe
xqcUigYASBgzryGeN4VvuRfDCjs2WkYt0049qXfPQ3OKxSCKpXhWg6A2pH9kU7E0
OkbJJ0Wq0d3Neo1tsra/bGHQIc+FZ8N/8w+tN7Tes7n0YJhhJerVemJnum+2ylCw
araMtUZh/j+2RBNHzf63z9JVEuWbxCmHfSUO4ItOGJHkseEv5TvUZVm9zY/Jb3ib
+fLI4WuwJB49/tUZj8cJG1/E7MyVfK7cF8FSv8zYF4SWr8/VIpzoaZ9eMh7+Rq0q
VX6if5LBomiyuPPO+9PFBnAOakZJy5LiAKdH5yxn6sVN3RK0zAwGLtKNdrXF9gjG
43QlYs0Hfxze9nB0kJCY2aPwOQd7NavvomcrhGBZRVX1wVMzDdLGJvjCOYQ5w541
9g0M30yI1e7hasLo/4NcXb0XemVUr+fIedYzAFqEx6ZiyIz2BTGLo7MxW7R3nvin
Xy5Vh2qaD8kWBX0i0qfqAFNL2HcUmkxiauai4bDTUj9FWfflhZwmofWQtpZrJETO
wJT7kDnmGi6svZ4HfFoWiFsQ4GfsQxctMsUHmhZXETjFw4DmB0r3CqYG1Li92lec
UCZREvXtTDoEx1CnQnsGls5JRYznAYxQyRfm7D/MCLRhKAC7+LAWN+5YuXDP3Uu7
BYXC9moMO7ttHe0daAH5E3MDDN392tFZmANXHxSzaVKf3ScBD8LxzJXC/XecVehG
kZIiae1gGgAn19YGGNj7/ub3bP+rDijcm2KZs2szFDhcM+HiP/odkC6+QzVq6RJN
0xdv97U8f5GMdcRcsDdUm5msHciF2AGG4tjnUoF5YuD8P3XFDYFhqk6z0W2yIDXQ
1ckMuyoyMPA88ikaWqVdDEc0/6gvriYZ7w3PxzyOLNa1cyfcS1gKrypsqoyvzLET
99r1oyTxEbruzRltHbTg/dt7fP/RpxjcS5KeCxacIPx2gc80fOdyQSOmh6583lB0
3TlapsfAxD+qQHLul+1hi/xIsiG+Az0ASYIQP83+c6PSOLjdgXaelglTKeEcFi0z
MQCZmg/cSM+BFa1Soefy5DX4D3zadinhFRRs0wdTHJNEl2KR2CdAsobGS5I/9FEG
MCFuJ2D2Q9132hGmLoL1nJX2jJVmfQJNDrQ1cD7J8g2kmduSKjiKZ3ZIPcMUlPIh
ow586tssrCZ3zmBVbf9Wx/zbHMQ8/zG8nMlp8qBcOwOpe1yROaOddwO1xbpk8Tgw
X3DRt9ZFYZ8ymtyysRty6j1/dQd/AevQlTLj5AsJT+KVgZEEi5OtRDZwvzQwJEz2
isaxWSam9FXn8CEwXXeMLM6EH0I8Bw58sOFlVYw6SiC/ZkgbSRsTlQf3TYcR4hWH
vmVkGIPiE/dqGH/clAq3NquQQTkD/06n7gmLRWHAqaSRk3TRPGegrS9uLCEhxxiR
cwOyQjr0NgEawUkMOCcwO9LFvshf6VqpIETxnYYK3GvZPOMJYbRusjQVXfoCfYkP
U0XkO831ZZYkcZVyi5OqB5+b/0dx9mEDHvnaB1UgDfkeoAr/HedWChc5B7Tc7ls6
1LOiMT5prrY8btBJnXwkO0Ve0xFGgjwocY8JBfFTXzCUjJZXjyllPJIZuUg/rGbW
yb1awFa7/o7PwRz5FlC0j17i5z5eEFUsuR1UNPSCqC27FbMvTpu4kssvOj/vs+Gv
a3jk19DB6wz3P0hBL5A0MT6CYDKsqaInw/+NniP3ykaboyZ0aa02axp7jfKSZHTp
QrNTKLg3bBFbjhgkqwOfHLusBsBsz4GgDMQIZIdHgETgLJPH1M9ZfBKUBmD8mTdA
8e4vejPXRWDSGqaun/+qSODDacgXBgcLoSUIUmDyENHNfm5Elxx/A4MJiX0DmICL
GfSYIZq9/FDU4PUdeOkQI5hVaABhLuesbSqeNpRAHqFIBfReusBtoDDm9qeib5cX
iWXaAQJfgq6NzWJ7A5MZW+2XyX6LI91Uejb/co1LYZSps1ZyhG80tcG+J1VWGEHO
o8Ixw7diLFuRTymfZR6HjXB4Ez8DrcaC3SKPT3SjXCCvJRF6lRFU4g8Ysug2c0KM
wlwysyWXxj/v5jy8PxQrwCUWzZOdIHglUSgPLuUdPwz2vym60jE6FMA+l+Ab9Jtr
1stoDs0lKBXMcpvhFEcCJBpBc+RVREUeKHtcEzItYP5n0wp02WWC/TQDR6aemzT2
KvU7bRugZ2K+AncoU+nsJ/SwTYyS28XcdnoW0Tau9MyBDvl98sr3I9q8dYwoFkYw
PMd2vVTYVKsitnoFPGsaKF4HXKEmOuj/NozztNN+KaxOYWUMv0IXT5PXR2Bn4DbB
c2cAi3GHzcCVt930T5IBJQorlWi//d9m3rqEewIvqqGOQmDerZZ5/s+4aD1E1M2m
uwi/V9cOW6yI6dMXOw2rzrLLosfpzQDu9VU5DbI1dBpdO0iVPfsTqiT2pnN0hdrF
5bJCJIbKCBwBLNw3k6k50T7eLeivadavytq37aAw7RjAaeFxYp0js0XzMN88WfoI
N3z2irJNS6ojihoIAfyWDU6jq58g4S7EwmORblE3brp9FARdnWz2uaKUjJXH9pG6
qOJopLHtq9cZBEq9EU/0S6UsFUvq1dDd6KfgIHMcCeJWY6ixZXdnqX/l4CZj4Jrb
iRGwny4N1wMtvUt3yDaVrJ1GrsgqZ8OP9ctc4durW9Fvv2V4+Szb0xilcT40MEej
tBDdvKB15tOORyylQ1zWAE+BqQ++Q/nVS6IyEN8tO5laH1214Cuy7fSpwbnLEVMW
xdWUzwVjjl4E8mszWYz578IU43aZBSxwaKiF3UzgnEzQmwoq4NfUYUm3WQ4yJnOD
bbfrFXGUUvaDf5PzpJeMX6ACm/8bbIGbgL0pA11eqoQXfKQ/ASousfJJXc0p8RM0
psKcDNLM8TbWwKZts2Snbm7PfDQxh+HqKDNhpBRoD+FSG0X/u1o7EoxHsZfoD8S5
OlOknWOvEws/ffPwhOug/7T6+wljBjC6pIrKhhQ/eLl8DjMJrUPcZ/sRsIlnVN6v
Z+AoYP31mjVskfWPdTFWLVUulwjNOp0LARqHGFnh6vldyvrtBFY2EDLjZ30M9hE8
lI/uPLWheFS+XHcyOLjOrpvikc9uiu7zTihYfNSpFB2OOvfgm4kNcawbINrNfEJP
g07ff/Cn8DYx2IHqoCa1/X7RzjFSVeVYmkGuSHv0hdB3LEZyhD11lLrINq7Ds6jz
3pZVf+/J3hJq0J0aK7W1uE9+Nr6CYUeVfRu+veB3ra6kOsyf942uZQzu8etoK47Y
cFsYuFJvLeK5EduXt1fxHRLBou5yg3+44XBIKWTx8l29+ND3oLfQHZ0vEMItBLbF
4Sad+rgkIDbYPW0I/sYD9IyHLxWuvTk0tTqA4Jyuy6moWzwKaExbBBtW9MGP+N/m
u88BP2FGkWb2mah0HKy0jLOOdby003AI451mfXIpYFzus7cBouaBuN1uuFzRVkQg
1INXWoIzFqWX4v5oLwVTvt2pIerA9LTFoKoihB7UrHftY7ciLyUVb2ONB+biyK5h
4e7IMh7NIdCLc9BcEuacoVoulCmUPSO3k//fG9ziywEyxxujQOrV3pjOsen/pHV5
NvDxcy+w1YmnbEIHU3GbxDXB5ieMD5dd5VC+6uCKiayBlRFzOUb1OxsynVqf/k3F
g7D4FNJIIhYVollDmJCna4NEYbRYg2zHg+GDpCcoDgsfoc2nVRvX9alxI0xzKStI
LixeUi7qTXsG3SmK12d4yybEK+v+GUyCwd3enCzu4fYhtzatBcBYdaR0LwxrLx9z
BLrAGHHy8KnjyDAVxIaSefZArcbHxaTNRNgwcwAdw9t0iPT6owCjQAgtFFVAhHUy
6X20SACDWGWTVBuGXKX3rYPC1W0WHUacE+/FGbnl+9Iwpa3t8Vw8RR9MnlwT0Djc
tA4FDKY0T7/qAYWLc2lsYpaepqMcInljO19w2A4QeiBcFn9CnqX+7edqIWE21NQK
7vbPY2mTwIz35bm/+xegcNI2ubLLYmrNfiktRMwh1NyiLKl/jaRv9FpCl9xlOU0R
N1fxUxLC1cdqOxoRu51oV9F7NOhR6/Vw7uRVwu31AqJAQPnnurBOiQ0NnQOiN9H1
uCCUcvvA+5lHSTp3rss7fTjpaZwI/d7rApqstAf6/Ylt7hmg0NjmmmU139lDS+5k
8DTykw1Uvz+8MWLXcTfGWrCEw5NwZODWRBGQyuONlpWhwSy/jTI7JHqCg+I/r4BP
jOE5xYCtpU55c6B5nrvcdN8Xzg4nm5dpE/ITXbaP/GtfnKwaeq4qiCnnDCx7y2U5
QCoVW/Vb2bYtxTy+DSNaDLRKHCS/fkCL8ARHc1s/YtdVc9Hh5GLB4WY2a2Z4n8Xp
2+buIzD1Zzyi3mvapgIxkFbhnJE/Z5qi13T68GBDfL+fWnyt2ynyWSHPV6Sho/gc
+axfawX6CF9fsXMt+kCc+NWaXM7NQZjRxh25XmwBANpwKVV/4s6o89UiHZbPoREn
VbbFCwtOSao6h0QQUBFXeNkL4s6r8JFXcvOwsnVYY54gBzbcEQ4PE0lJ9Fxcksno
VCpGkF9m+yjz2rncHrlbBQ73+Ax/pIxrONiWSqCiNhyhIDW4jIJeqULm5bZYQns3
FBiK7DSVZgGw2OQ2UBOPr6G/nWs94UpdLBt51huihA5+oETzjy1SVH0tYpcrrb4c
V52brwErTHDE64OGsnChBqTHEZBz3iOXxHzLMNpaomSlSrHNEgLVBjl8LT2N2vsX
4PgKKOszsM/Rk2cNgnFaLv/BbEuMt+VTOsIQPCcXeb1J9aY4Sa4pmWBUkwxkeviJ
UQPwv/GdJAC/XxDR4jirsHqhhBfjhoOv/LBs1ruqGH++6VDSoOKYrK9b7tSCQFDt
M9mG+f/mBHHa1Yje8hdzgQ5ejqri9YOPD1KPdXK7bS3lVfOQ4T41DNi5w8LQ5Z7+
3+lI21+WmYLqFndkpXguZAUX9XWugxGhvupYAVHpgvrb95dKJidIlR/2NXbqs/18
uHiHV7Bull8lyrfXDj1UmRPCAwi2RoIFCZqhgpjEoqTe+quKVf8LMrGfauJXbjAA
yjHg8hC4TKl8BTSicfBxbBNxeeCzcrJoxWuG3K84uoqT4z+Be3FhuusLYLliTJ5O
B08Yxj6BkW0VND3xkb2LO8MHnijIc3M25VCkANK6lDS5CSHg/h4p2Wg510Bi2RRu
QyRAGqXlKZDotgW8x1gISXoh8/kMWAckbi5DHtN1P9Xf1DIs5h4bF+djseLlpYBK
H2GAKOC3cUqGFoNXQcLlLul8IG1oUFuDdZtk2ToxH3k2Wh9CfU7nZ/l6VM9hGCCK
Gppy9LpReOQV9tDoSmYj68HUW7+tYHPCvBCCdweb+XkzxkOk3fa5mELkgvotf3rG
2ZbHmR5cZMDiXf5bMH6RUA7k6MX1B8S4HUmQc6mu6FhOJjZ6zOpIfm1hTJstI1JY
3GbnjUhkQsWLh+v5bouhjfeoZjUJays4jjNjXU4o4SxoJ6gGhyB4jwnI6EnbWbXG
zUmpHjmchY5jUdp4U2bUwZm6W2TTFZ/POlkK3GPtq/c2SqdiAvOzPMk32rdwZN4r
iZnzAYsMD1W1JBEAUTVCTYoiQDia9YqXY92+MOZx9nStlJzGmGsRuU9VP7hicuhL
gVL7u43cEXsZtPqIvu9HgfOu6jEz6MN2ogBvO3pB6zRBnfdLJKRRhSPIl6fsxO9Z
iVyA0z+WmGYXvbhiOUpoKH5mVDOROd9dS6rx//pLwPpz3w3/d/RWdTZUIp2aZtjl
xg13R7/cDwebghENZ9gWYAc8QB7vLY/4WS0KFYT96Wv0LVdLoWDfsmOrWAWtqaDV
FSwvfcuiu7TR+Q3Dle7bTvKRXyD5vYpCENBxcC1UiYUGOvG8bt/TxPeMWo2Y/InJ
VuboCIDgZrTPMs78m3XQZtw2Xx1ToPK1zDlx84CVHabHJ6zdYbWhqbTGP57QB6Nf
tNddK5hPYWox5208LIlIFPiwfPmFPVvQ1uNOPCcxc2C1cOdqykg+WxtPJXkFzvHB
cJzmjrWkAYSgqd2HSIRm3VgMZ3LjoyhGHBQUbLupP/0o4/Asc9jJMsxuplMpbHTj
8Tm2118wSLV0wAOHIIw4j/wT+Xsc6PHxIvpyFoZSW9r7B8ic9sjWl1pUO7eXjtF/
8cU6CW0QQEWLdHE/illrkiQnu6YH1UCTa4inHnAPlZanGEuy0MRZ6UVPJS0I4U1F
hfPW1ai4qe4reP8dZu/GD7s3SLZFkrU+8fSTl7Xvu1vQeT6tv1esPjMpseKzpO8M
GYVgIt5UrQh/ybu/cxLavQ7g4bXLaTrhbJE1mCdCiZRZ3qDfbTLKWKYeoB0SAix2
oDNUNC65qzYOT6ci1NgRMs3pmSIOfaGNT20NIrdADEgiFQ8aEfMVN3KI197CgMbs
z2kXJEwqqXaktgoZ1o/sr2BJjxZo7h9mSJAi4QPaZrLCMHBqBbGMOpUUCD32Q0Dn
/flAfiNpkgmYuwfuyuxnkubWkKV9U2Btv3fe+C/GOsbMdppITUTlUxskDDR67HYj
iT5LuOnJg/og4nPE1G2z1jseo9huk8up0M/+QigZTqtUzrw/benTn3o/yWdsLikm
Qu5mG/gkU8CYtV9KFP4qgq2JhG2HzdmosCfhTWOs/iGT98Yic3vuCE/OPTw7wLWs
CLqbU8+VTcYHwARp7EoTegQ0d6iBUXK8XvW37D/iFRHBJjCEKNT0tGc2aBNLVZPX
YuA1Shx4p8+dAP2D5dI3pq9EYWExf8J5pJ0N1URxr0gxqpLPs/rtD5V7/u1iAK7/
+Pj09t1wTbw+4A/oL68NR5n8ptQlxJF/SkQNeSgqTdNxZsTT8D3cAkDmwjw2kLTy
CsSsCMZ4DuS9aQlf8vPdgcDlt44iRjFDBfFpRiLzjeER8Vcwqeb3FCy2rMIHP5wW
1GmRWlFRTFRSAxgm6gbxhL58FA2PCmpTQyzjooDn7g28v2RxsRH3vh9dU32igeJF
UYsGoUvaYV2WC5PpoOJytUZnFWXVgLHzHXPo8kRZ/mrGQs9mRl1laLWDdJaBTaDr
Tr0fF011oaa/hEixLsbvkwWzGI9OwMCef+P+kGKDBEkg7nsqvTWioOaxQDbcewqD
KvjiDcw74AhlpnUviMpCdtYZmQ4SNlXQFqVB305yYCoowLaJPxSbs9vh/MWEoU/r
eD1Hiw/K8iUt7rPPK+lTSwTnod57wRVgkyMT6R0MqrglVoYkozn2AA47Wtth6MqZ
ivzq8OANJwh8MfB19L7MOjGpip6qBEvD0chZxsWr4yL2AAAcD741TL99ZZM2EsTS
j9Mf2tBcYeLdywTvoBufUKyMcag2FUfOgDZHPEUEfEYTvkMPnaCtoYX1OTyV0pof
X0W/zXPCx1gOwwRme3hEQRLMQEP/5BrdDh6mE8W2SXVxfb0NojmAkuPhdLT5Zj+k
M3VqKUCSu9wXuhoRo9JhNnFczbJzfJmzspY4fq+RWDbVIorlBx7W2W0cvxnFFIja
yxZ15ibPp/OYOrQhCA4+CtRpV5P4M+0JojX+QbM7qpBg91+QHcpZiisHlKLXlfU1
8c0zZmcvbqmeX0aitlV7bWWfWW2/GvZPMZf4LAxcCurF8ptwBZfv5+fjgdqx5aRc
CRPjOVhoqApcRKphoZ1Jqg2AvEv7eODQ4fKviO0AfZLQwItusmAJt1ZV7USWXxRM
ClMEAvwxpasq2wM8cu0rus+JFrsR02u+m5ziSlzyJXPBnr3+16FPMTdXM8NnQ+kn
0pIj+IiOeav/j3/YIdXJCgMFN3L4w8UDmRQSXgn6TSTbYceBEHSmm9QPaM8Z3h7r
Z4c7/E5NF5SrGpB5bKjrCkAI3aG32Ft70+JZL/C9/8a5XKJ2X7/6Hltk3xsayVEl
PuEbTsNI9J4NF7MkB6TVXSUG1yK5LAMTWdGRQmwClpCZ/NoCt0Kc4NP8ZTXC9j1k
tl1RILgZLv1pFmRK3j56qh2ZfqyitdOV5xrrRQculfdIFSIL/VxA2N519YYfGPdB
Z/KO2mcpkvzsL1Hdzw31olpX5cOywpkHoJxjSkeWOw7xfORLWYZKjUiWTk4KXmIw
0NwQusiqXNAP7qS4mppP+c1VJaKHaFHMEFsSjTKl7XVsNotKnNLJ/5El9AcWi8uO
vsatHLSO6lIZbjmDM3ykNzmJP3mMZc8w44qih9LJA3ZwBjyc/dE5RB4y8+KgIz2n
LjnwsY/FPL5X9hF2WPUUBjeqaKx4jyFaa+TCnGTHR+p8rGV5fc61MIPRU7qPME7Z
1w4DuLqDi44E/EPqo1hpdLrHZmAA3bRauosTgMgGfjBscoVCUQMDNLOIjITUB71/
oYeKEIszZtO2x22hoxcoRF/MhQE0rZNbzXLZekBtQB7ArqSJM/696mqm372DffZc
h1//EKqumha1O2SAAm+rNhmBYZjGO5dvoIryHv64zTpy9NNX89l5eyKEnAX1eNs9
LU4XjiejUs3uQm3b+arDxbgEK6HsDMI8sz1KRXGrw/V8Q1UosvVxYyHvfN3Gf2bU
LppPj92OlXGuTWPzPInMumh2/WwGZHpAa76a7sm/9H6438593xAbqlpi/kX8qQU0
5H2ki/1SaWlODTqoDoGE3cltzXZcRkY6PSzAkfB/Ta5ZyAcgSur8YAKDY9ch0qqF
h1XZovTEJjAfQ6f3PfS4cs+UqvSrkxhbuvNRLu/RO/aQQycNJrkGdaCRf6PNCtOc
mG+GyLZvr8B3Rs1KsNGvOiwZ45XuD3izkcC6ytM0RQvCDCTmwqlSRu319EESV+NN
ikeGaK2LTV8B5JFXE2EKrPeN644zEBk6Pn88qT8aLlHWwBSDezmPMvQS2qSN1SCA
oF+khjHNhRZoh+hR+q3YG92iRtS3OFXsnLaPPsXua1bKuA6nZgU0hbGoRTTbx+35
CFZX6Z+b6hXdmG/WWbPXX0IxcMvqQ+PTiyylnIEv2coQZKFg4+HY5BMEnMP6HGr5
6muXr9sPvVCSXPUfpJx+mp+VRFLkGOcbWCXgXuiCMbvNvze64kIsu5Y4GCxxwrKa
se9RvqHZn5BzqOttggCKyVTRh6iUUjwTcdJrUKaaXWazFZiVQYTgqXGNTrgzzM3h
h+de87kxZqG5tSUmcGRT6j46beSKjYkY6VNfvZHaEpTAbHA3tSwl1p9MgDtvYSRJ
3TOnq719q6vmhrR2ZEI5KslwiaYtwlpvCRdaC6qjLo8ph3HeUA+jPrmXHD/oYi8a
p+zi4Go5j/vfSaKsfTfHcyenpYugEpNgFzVliUjF4W6lI1VwLrJHDJyOIcloQtYg
3GiGNUvRRZNgf+bEv8M1BBFtMCH0MJcMzzTctxMvJk+AjFCkBx01d/e0QE6B09gH
KvkNw4YUVyxPLAzFv72ubfkhKLfBmQ/wGnCwZS5T/UKw63lJOp3Plc36aXQSDcVD
b574KCTJSpqYaHT+s/Z8rXvnqrSn4feZ46r8yH3tC1/4HXAsWxPsrHUw2m7k6Tcw
nhYQ6rI8UHS1Iu7xSS5stIf4QJsXOA7u9FU2492FADrcRDBgd3v4W1S5Ne4wnDMD
DS+XQw1jCuhrAQElabyamW/NHeuMw6+MpNWLLSNydWhWWZaZbuP3uKWUFn+GJ5/N
nxrIrI2apSdMYcvV8NhCgjXw5ARLYs3cJI7P1VaK+bMfDLmJgbLZCNhU6zixwp8/
0fZTS+fIoY7z/h1fyi6Tdd/edAG+T9aOiu+uLF2Ebkj//PPVRTj1K033S7U+8jfz
Lo7sMjAkMqbZW2Tb0VY8xOf4JqCmPp66V34fPpzGD0vxT2Gb7UiwdQM8u0kQcn4e
WexbmW48O7YerrTvZZ8XCRKehG7s6GA7LqpXWorisUSyB/f88hiJH2nm9hiITWC6
8tRWJa852C+r/b5VWeh3brgc1M/mymDQWKczPK08bg1mrhOYYy9siOVzRpIw9VuY
liiLdLBenU2oGpkFqhK7PGIg0EOxhxy3v6MwD02dKmHdLGgC/qTSdvqkVvbmnYAh
iu0gL+xGfI8PW8AL7pL5yopsCcCI5psEznczWTlps7mhoG/3QO08XY4qDPh5ijlA
ugnFDHrUSYOvBW8dZBgglPP5bSh0+r1PE8nPoNsZLZe29ITQ1oNdYIUZWyO0Nn69
ibrEtpf4rmDXXv/iOTrPuIt1DUkea1vaF2bsvwMfo8UnQZWFVDG8KNfIZzZji346
MYACVqRqUP6MiQG+7n8S9ZUJjvazzoH6aRqjontHriqLKCBNi3X2xYv4l7ZnAN5X
epj2pEFqFCK95W6XSwF+tXidvVICQBBYxC1fwFMCCqsdKaSjXWvzoBNm3Z0tPnJf
DGR+IuFJkmDKSp95GpZasJEXcEbRLzM013aLo/o8GD6TLxD937KhcEUa9n2KDrqc
FCSZlpJO5auZUwC+6J5bRBTL6qLBMh7Ob2LRhbKuz5p4ZBnsRudv2sn9+ZGtqYLQ
9K/ojLJ7XspH+Cga0013OocXuDK8PW/Q021mM7jRDD/rWrZsW6xsloJsn6A5ODJz
/PkR5bwcDwPwPkWtsJSXWXNCnYNw/WjsIPYvOx13JNsV/Ow9kgKWNkszuGvmEdB6
r2cSeICS63tFluZNFH5dODjSJgExHRFzqUrCsBcLI6rm4R12CR/r3Pj6Ih+jAnWP
AZnabVIYh5e3bLyG7GetAZRHOQnX/rbZOhh+mbkhunNYPlN9OdacyI9H8Zc+LjQt
S/HyGckGPu8LFqAy7envbX6w4bi7iWChfcj+zUHP22JftqH0pNsjR71nG4ud2dJ3
C1MzuFlrOXlhb5/ePQcmzR2sFSz8IYJ9S2yHGJTutpEwdokwavTIGhqiIFmwiHUU
wQ/U7FW4hDOL4OeKyQvKJOHoIsjYW9ISjymIgKQPPQ6E3fZMFY+C5juczYmkVzEe
SpqazGo0eE4EgX5yGe7zBEHgiWMQ4o62nTeJqd6PMksu3EQsfycG0DsLt48UmzYF
qQV84qgnaMxTHEabFvtJcgEzHv8Jyy0Z7MMN9IzUSX/cnyO3m6LVyF9Wb97sb99U
vEXAWBPnO8KioXzQhFsrRqipGkXzpzbz7hIRIV/R+xR7X08j1o4JL27gyoJAyLFg
n/yAX0EYmaoGZgMY0Bke6XCzUrHiQhsR6Dw2hKcQxThw7X0XBA/SkU0uTWUg95U3
cjZ35WJto5u+d7S++A4K/t+nRrucou596PP64wR9Lbr9APnPGYcFLYu5fulqs8Tp
UpVeww2a9a9tO60oKlSkYNsjg6BgujasBvH5lhAGm6ZYXKLuyzXeB8UjFHZ3exFN
mzvVezf3Xh/55sp2KZnliT4H5QXj+Vo3UV4g1wmerUoJ+1dQ6l4+aOrbeoboYIP3
IZKYEKQvtcutVgmKzGX2LiTHWCEiD9l5oe7FGnVJKSpmrTFUjcRrIRu/vBnq4OUS
+/1E3KFSjoL0Jlk74HreIruOL8u3ZMj8pK9cOk1zZlrU/EC2Qb/oK99H1U2Bgov5
8cRLPg0nifBMlVzw/NKanYaPfs/nOMo7gVdNhu+tfkzYAw5g+9tiDxVICatgTtOw
yrvoycw4HHC/vIOCy2VXWsunMPOEJffdORQ1ehtcIgDteC14EOp/2GvegFIXE9mm
O8PGrIwN86/OX3K369mbqR9hO4q0rSct6RdalsEeCmCJGIrWI5KgPr2Yg/1oe7TT
DYTa+DAkBMJa1+IK/1JggcuqyUlICfmCG2Jgt/AQ3S0RvwYUgVyP0RiqvF1Mx7G+
zeTQQJ0f6XyktQ76kaGolZLcn+JBwWAmkuk36yqEY+ipH+XWZa06Z9w6btAage1a
ievfXlSCzfwRy0/itAq/slp79sLNaShGptwhRW3IrQoSlu1lizc7tg7CnV3b0ywC
a02KuqwZXyWTemMYLa+RwXfPi5ckiboK962RTa8NcYH+1fm9vIIYbHufT+LKxP1Q
ktf4owZovnEwQaHomPnfD7MU9meOficX3BuY3uNB6uuSAr0vWeY0nSxN5RWGkO25
kejZOcz5GUnoeyp1EIMuwA==
`pragma protect end_protected
