`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n4k3VWYxHeT9I1752AhqxTMOBcZywSOB/u9n3fLvmbngE6ExaWBo1IUQD3H2CHf5
y5+yJxKgsGZRuaiu/cencwx/8mX8DT4CtScFslwY0BWFeqvUQmcDfa4vFAxzDC/P
6Gkh/4M7HDpfzgR4D3no55krYjdpAXTQTZfjdug01CQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30832)
rIiSB5/Ech5uLssJGLJMdgOos65YNQBKRRdDk0rYBmPAoL/UnrnugRGdai8i3JU/
cdBwlQ+iV1y9H2/KZAipx8ul4lio8E2rcUVCc5qRu8H6xbYFbKrGI711DS1N3pLa
27eUoXUiDM9lEXAbuLzfNLWZgBJWAww39SeDyJ0uvflEB2RXDIYa+ma39+e2exx/
3IaEghoi15pcaeUa8xEcnFju2g0sK3Eb0dh9WkbaXdLVyZbHuj9G1magN2J9oWKY
YIJeoee+ivbmBgEH+enguPpEi22PvBAwJGayUs3N1ss5we1trkOZtC3vgEnZ+ZMJ
d6thrQxH3fX4Pmd+KgdsR8IboUJZWPhpjRwDtgWbGQ0DYNA+/oH73W+DBDRFaWEc
+BehYPk+KquIoqpoeMyvL9CWyrZF72sVtGOhQDDfVguDJlJwshF/NzNEiFQsoCQ6
75/tNzMONAbkVNxvzsxQPnmg3mpf6W5Eqh46TirFRZTAuI8SD5xZevgbzTulw675
1ph7S3GZO5dIH7+7ls8dOBIvIgM6EO5fXH/z9YBAWLj8SkpECPLdo3+U/pJ14fI9
b6g5FFuWt4rwdRiqWn8zc70SND6wIa7ymvqTSaGJTNaraEBxOMhzAoVVqwl/rq+O
NnD/IxfylgUXklZ4352Q0ZzkZq74xTcylxE5orOeejlceRf+ZCVQrWIfeG76hZcg
ZridkrMXl06Ys6w/eb4zU/jdnEG3jjTcDbSnQnAQnYjt7rAVLceHkN5PXKrgGsAO
xbhd0v2txBvGoa46mmiFH271h1UlbC0tHf5pU5Dg3CbsaC1nh6EtKn4A9///Jkid
irjZNoxR80LhFs/JAGhCpBTmTDMf9mXPdKjQvM5r4lAiUgOBYO1Ty0o8FQ03d2Bl
a2kTLKbbrOcqpdAaPzbx3wD0SyFlr2aRDIr2Va7LiSGMW3Cq8haEQLdgOfud2R5P
KiwedNzH0paVSW6zHI3lkBRFJtG0EHl7njyfe1THFyHnm/pFymJdSGbWy2JTlJLa
OkYAJkEuI69BQpZw5Jv5w2Mes7pmfd4DxEr3MnxMXY+27HBPDjM+jfQCBp20z57T
7sk34d3ju9s46UW4tma+SXWlk3mG16kYJW0vs/dNo7SZsIljrdhco+ed9U5w1lIL
bBaaeZ520gVKWhxtTpp7q2WryX5Ab1TAAcOAxT/UXAc9rMP6aN6fwZhY3iDG9nB0
19Lmo2g20ee1UeVdxBOT8Ozv4qzlH1WiXzmgT+ZYxBBFnJU9sZSADba0o/vgK0cT
3yybVwMf/cDfTEDoJh+pdvPNIZX7If809gGuux89Cidma4UCeZHTFf7Cs2Unig4/
sK8xxnaPFrROuqA4J7ATnM4YVyUpmA8NPNPrjDM143ldOCBt5/vvQ93MhsZHSX4E
5xOBQ12s1Pvg+HUmhj8IGvCVcKbOFque5zbsDRZa4iz2QstcxRUAvYzdt3qhufUD
EX0rQY5tdBw2eZklwnYB1Lv3RA9iRF8TrJ5Um2Eg5uXFQGYMgJ4nfavocqs1Zyp/
4Ln3hpU4+tjN/oMmbCAkrr6byFoyAnNbq94BpgoEEYK0mAO+ElW7oQlxQiwsxIDY
YocKP4jcOytiVlvhQzP2+EqD0f8FysE1+FoeQUMN/CcwYY8spIeBgm72Wj1IeGFg
R0+R4E+eJW/rzuUc5CXFmJy/W3v/8OwmYi0ScY6i+TvbTw43JCWQd17OKtigxcKt
npVbOX9qZ4gqG3QyYzUZIJAbpbduYWaboU0ddnaqMh/5LyDVSbMYbzngQhbFOngj
A/PmPA2V6AieCpNtaGmwfSo98Bmy8d5nf46+7vnvBOnrwMiTTa2TQc8qyggUP76a
eb1FMWIkllt0UPuM1xK6RA7mCKCdtqQX3FaRnT073Fp0PV7jxGh4GUODriDzv0Vh
abq7hmNuL/dcGPsGPC1OFfn2SnAPThHJr5wxz3HFck9DrYItgLBj2CDzB0PtidAi
051ptqgEj9ARz0JD0AEoLNhLhyDi6QopmLJj1t4/gOFj54Fe64iv2L9DWfMYeOoO
G/YHbb/jF3IQkTDMnjBjeI0SN+P8BkM/kVluLNJuRYesytNbbheAS+DL44hP70od
j2ThVe/5vNZ5oEVmME0T+kOZZ0DAYjJqPtNhi3fUWs0ciBm0Jnps5KOckIgGczHQ
wmjKhD7yNq7e3vYGpf8Bgof3tSDLw06mmvzO1PcmmVyOWFH0FWTuWZ2WkU9PfUEo
tg864EzocZkoTHl4F27gQz9NdXB0qmwyXI5mkfnUNyDW03VRAMWRI/9K00+pr7Py
yRvSyuWyIcvuPaXVYoP+mhm23LPUQDd/yLlpQgFyhUKMBovtnUnhdVWn/s1iDpXK
FmadsnSFHqzpgJt1MLQw0rPA1Imvg0aasOHG9hhDyrb0zKEqpi8XYOOHxzxqwQUZ
t7bz3Qpdyewehw+z0nZYzZSG4b9KkqfIuXm5263HkIe2L9+64EUweZut558vE3G+
QYsFymcoVD43N8BOjVhG5pEeyt2qj5CfapuGOwkwjIMDzjDNZsiPni37NMbbbCp0
n7M+bTDxKOSE40PTuLLxFUBtKHHm2Uh8MF51JQMMHHTHE4bgApOMvA/0j9/wx5dC
xAEVqtffaXqpUffR6qL29UuX7rdCGaHOjCm4z/XRHpKaXk7zZntvfYOWCt35R0jC
JjEO6UVNmGbXOCnHiWJI02r/tlLTJ+r8yS0CH6XWXpHs8rNrxPxIwDhm5t7AuAZh
WR8MWbtxhUH1LQiVoD4xkk7K5E9Z0YNUNDvQANwe7xXdRuwlRJYRUtdcL29NLrPm
bacy6QWbQpQ2MABlgo+rthaLEWGm+SVAXXclwhQ4ysGG6jq3A7QfmbA45mGNt8Pa
xVCyYjx3e6ybGUZtgHs3rEPgwEo4hxVefuKOIju1wrB2HvKfw09F8+/MyMx77FXy
aLTDBlZ1W3QsB/z0fJIXVfkKn/XS5bTsUyNLvrYxQfsyIh4Y4KyiHfibgVzSqYr/
X/g+AEmc1nRmBp4xtqw5e4g3Zl7AWQlEbZLsyWPVR0K1KczBC6HBPlrZiwH7Yf80
DipV1JYSsYxWUo8ZHQJrK38M+5AMOrpW/wNjESQrgf27k7+0zXK6ahp2JS5atd33
Vl+E/yBIOEZ6wwIjHad3NgYvVWPXosX3BFZPnG7BYt92noa+609bIalLagyb4E6I
zx8+xv1YtUIdbiJoEETLrAvoLBIPtFWHMAYjRWKj5EOt+0csuPCRcK7mg3cFDVhX
SCgDS/30xX0re0HkVPevDTcW4dG0AxsK/SUnRVeWZ2eFO5GxDLhA8iD4TRtvJqsS
fodSXaLssgN99FMCK1x04UyBpVJZj67WUNx/V0OtoIHL4mfsUogS8VmIjThN2b2X
BzEtCVAPdXiwc+6WV9RpcG6xMKxYiOnuVI6VDo3eyvb8WKGiRdWDp7pFYsNFsRmG
yKq1/uGBcvR5KMhVoM37np4f95g41rmaPqtHyOViTGE347ISecvHpjMra0vfUClK
l1dXy7tsLQSmx1rFqF1KcOQZaWqIs4f9hsvEVKmBdogLA6IiaZ2i4HfRFE4Lr2H+
NEHuX5v71eCTmoDl0iuuee07lXmkYKso1RMbgF8h561KaVP8j263uvJuRw9V3is0
UhmTzZqXLyip6B8fhUPICBCkFRKfSTVu9OfXpoOhzXuCUcTww3Bi5F/dLCCzVIQq
2W50M1zqSL9Dw9DdarwhLwNqAmUNYFn04B0AHOPyRDBtd8M8Uj2MklpYI+WnUuZz
S5lGopJdbvrOtph8+DXBSqHNbRHt78TSWp0034xQBPL1CgReKkai/65RI3MNWaXg
2Nr7O7kGZA51xWQsvDRUriYR9glgJcy23dvwokYgzbRBOZ8W+20lB5h6bri6KXvg
KUs2K6abi2j79BcsZoKzBNPg+nmJyd27I1VUYJIBWOS7Fa/mHc/mDs5EIlYKAXxW
3Ppb5uWN0yBoOSCinfIyJHjWqfvegIflyyj2tXzQR/3wK+rf6Oe2DDnPmy2HfKjV
7JouGpXf5kacBOZItPWKdiLRfMYVA5fFeQAy0ExXg9cbRJctJlpiCHfNHv2j4/0N
IFMcherEfCZeg3hwNmOHG4ScYaWtT+pt2aoxj0/Xml+jkC8T8SnW2d6KXclkR702
o1RivIFe7pCB1JRXmN7RurFZ0zrjZkT1Tw33lRPKDMq/oKAYQFjLtvFCaJ8c8bcG
Pk3nhrZye/NSwkTeGsIYDAZlGz1/r1XYRVQ2aVAW54KB2F1Ofp2Z2qvX4kgxF3Jg
QnG8mTRwcIA1bY9yzWUjT/kvk/IgtdZm+GRxt5amf5Mnfvnumq7KTOveWWymNvjY
jW2Vng9rOiLW+Unw45m7O+jY29hLe3Z0Mbls32rsFRDK0jCvHLA9H17mdl2sORyo
7NN0HEwSe8hAwxdkO/rVosSixpwZ86iQfLI79w/yADeDcT5oFlaRgaVvRGvkTrxh
kQ4NByKFW+CtGvXofGv7B/ENASrNAFZjIzPMY61W+36zz5l2602tN7C/MWnVO1Rj
iJLr0F+sLxRMLYmHw8KCOHNE4zAh9BUliCKpGHd7VSkWR9kGM966jEz8Du5FSP4i
4lp7fV+vKlduerGhRL/O0Mm4tZlRXQqqInKFvuTyCSID/Yj/AhoLGz34VsB0/i2G
057brrzoLEgqFijKBDNLgfjPqsWyGaLr1ljR2kOD9eahIuwTe7Bg4wNxQii+9POD
mLdwk8YnOlalsXmD0bvk2gR6eluBZ+MflIXuwbBvVIG4suwDn6qZ5a3UsuVSJLhX
nu5DOcy+LN6XWWTHZbA8V3gvz82E/0Y7L4cTKZtgGYSzapgB5hvbKHbK+xmSFwBv
j2rBC5vWu9APQn67lX0ZwqEe032dgRzEkzi4hzEizV2CXVEZJTvHRf6P68hlqk6t
BlOZMCYc0S2+tXd/GAX1fZvM4FeGzUsSEQTh1AJBan8hnCFUY/aTbZLrRcrloVqe
6XnG823S3+Y2MsnhKpjoWcMOIodK/QR4RO3SIpXtyf+TZ+0KnoTuJ3U6EjoDsBK5
VkjgsugCZRw0ehfNuVJy4YwXh9T4Sb24cEmSPlbsUIiDvcbTUGnZ+pa2GPr+lHum
D6cwIemog3JDChE6i7b4+etMbOgEHSkTZRUQPx6/UDwiXOcCAM0WU48TEGyhXD/p
Fm68wAyHKjfoc1cwKXxtbUhMBSSpX5VDupGil18fVp8hFue2tDWzMDsTg75sWIXs
mXydCGQoZsqGonyBmBBNvMJGZ8y+gchMj0IQYtvvQ4HqZq8c/Nol0EC1f4a1tbRz
OauYtdZ9Y0plzNIXRHA2eaTc/88snJwoWGJF7835mEgQoQhKgHYiczvgjAdpMhaD
yKlJbE9XmXaRR30hLkn9dr3ZxECbsbavDJQCSW29Z3HKKK3/NhezfNJRfL7dV5vg
Iq9yMPIKTXe9bZHQa5kqUnkSWh+OMI99SGeQo7M7nyWcq1PhGZ0sEw+TwqLs7Lw4
ecHuY1ZD3feam0WYu4Ub5r58s7p4/VkBfMYnJqQlCyJMLWiKvgV1Iqc5x4ZBsSQp
/VrS3rLn5+r6JzSOMLISIqdpqTNuutN1HEDzlOePD1qgqXifhyW9nyn2BW6/5LUB
g3v+uentAtJZgfb3Y38iIAYYLh8HuutYfzj2mWB9bmHin6fd7FbeuydaHYaX+M3Q
mBWGjOY74PrvqpOpnIhIwhQJkNeP2BZlR6HzIJ+TXO/6sjeEdFv5xbzo7nyeyc3V
TR/9NogFD9/2u87JBqFod5JlphKxgKfI79/Ht8Hg7Q7JL50PFatjbmk1fmY1DOZz
uebC7+AHOfP1B7APAFNTOMoV4lG5JaAH3q+9EEZlDfkBqOoLl2ODT4SS1A9Z2oKV
wZJRIP9f5Rd+hiKvO+FX65RmyI7gqigvUuNR2hBDCSFD6wtDibWRThLnbeULoS3r
6nhaFct31vKuAN+aNweK/Kuwlu1dKXah7Z0z8dRvsDoc/t6ntv6Ejx5GR6VX6s62
+dQ23OuPxV08dpYknszmDaWgzZhJ2Qbrwc/Q09OQtPm6HTwUgS0ZAA/SZnCEytJK
PavvUkPsKFG/QlhwZehhYM64AB7w+imwob8gQFHr3nRdES2W52GHcts+1zNT2liD
lMN6EIBjf8HBbNPiqHxLTV4AwK9FDGmgqf/1imSIRqvPsLo91gxY2jGKuhlZwurT
WvtWr8G1SaFJHJ0Ex1uCTDwZA4p05AV2SLp7Xtcozchs6Kh8W553+iVxQiXajwfx
GxXwusyc+f/StBYbQrZIaBivdnmDx0JZh0P36qzbTIUcE1SGbJSivleY9dLkLlEU
WpzFtIAXQD12anEigNEgVIGMAwD3CIdWnerSRGlKFkzdqE7kmoMBXCPyujb/iy0b
E9ukfx/W700GfC5POZpnBTFlxH4WPsG7Z4ERniPWp0ibwvBZqTqFiErheee1XH32
O87OSbI3CRxtOg6OOB5kGHCp1kPidq8tpcD9GVeshSNNflSoOdf56pAWxbfYSBNw
9dFiAA3IvSeoh6ZllNRHZnikCyTettPHnMTvuWsNs4iuysTZker2twizZxBtqls2
hRIckUL+QDxYDyhtPTSTsc08k8bdJNG0gNX2GFbvsBPpTKseWW9DY9JFzlVKQqdR
ufOFfR/zGSuyk9ACuSgG2fIubUB0IToehl7X2DADhFrUKsx3kd4vf4Pc4LPqhh25
W1InvaiZgZFz+gM0s5KrSXDNAXEwr4EfbJFMtF1R9Qj4Qi+bIhyQ+diVMB//jzGZ
QPPXb1ZFlXa1Z/b0x7XPCe8hCOvrdma+TcGO+FoMEFjimb12nMGHHFzNFRzA7aJt
bCCFYpuDOb3AW/9RhOir8p4SLePEY6H+CLkDxKfAVAAE+lltDx6UzBwCBd5sfjyr
Y96/W8jiuNryFm0k4kE9Eek7Paq7KNJ9R0q1o3gaynKEfuzU7ineMXn5Fj7ffMjn
QuZFP0CRxZ5C5c1I2fVxHIBjs+nnKFP70+0qyPfKlMPZDotYIWXhPp7mcfziP+4I
TOnHLAW1TKg6Ub7+adYM+aa2k1XGoK4GMRAn99HJIO6shepm1bZkOjXVTXgaAVpZ
/X94lNWH2hoDics7e8g6hsQvZDby1ZZzESNgcD9cQoRM2gDBV4wij5FOYAsJoL1x
dKL+1i1h5lT1HumURNiXBfa1Iz1Z5U0EUXl07IMpZRDGRqE7CWnSgsWXkWLJqyxn
TH1tUSKGS9I+bidiZ4lvCuRSxxe7iROpPlW8bmq9iEOevbTKwlSKL3BEGcp74c4y
ZmDr5Z1F5FpVJD5bxafh4fKqxS4C6Zh52Ivcm86SeLJUWyepjr/Jw4k3+2A4xhlj
YaDlLsfhQU+FDmeCOTiSVwm2nfOcf89jBaNU7AB6pLaXjfT413GvXRCZ6V5c5e6R
s62M2bUpR3x7HP+lEiCkXQM8DLjW/PD8h3aoMOmgTjCQAirMDr+INKUnzrWJ0to/
+cHzlQxgtaRTXDl5K5Fz1R7PpgSdeRLdNM2QZJKBF033b2VeUuZLo0kKQApEh+ho
g+i8kHTHf2xanNIrEJUSrtP58jJPZjWvaCIVZTkHEMpDr45tt1i6SQt0qUbq5O+b
2UnknYaOqLyIJq7vu//wYDbfSfvAGdftcqJyJ205ThBfb/be6VRHENj9yjdC2qKB
yPkU2mWtjRNbukXl3t9p5mmDR9G5PfcQp8Whl1imKFSGOJSs35cunt7HLSsYeRZd
nq7TSU6iuVDc7wZ1scaEeayfAzQyGP+zWR9aJknleVj+86D72k0fvLfjuhQAhtCi
hzbUbvCtbrY7R1fA8hCiwobDIEhTLKWfNcGgyGXEE8ovTopb3zHcG/qPtr8+CuVr
R8REcSKlsuDyKtTO+R9/XG+yYs/SPF4RmYNxph1ppQQFYfCrZYwlIbY8gsuPwYI0
PhcW5HNRsA4hfpnO8tE63G3IQleWS0Qx6aw6j2f8KW4XIVqxHPO5ehtexmkNRC4m
4SQtwQe3EM15ee+g1oyC230uwXKJIQegYwbJTS2BwO5wEmUVrqgV7k6kS6Xf7SXf
7iF9pwcHxAiDbm6CjTtdAmrpGu0nhMOGSqefVixt5Olfi9KSa37clny0syBisj3U
X5RgOjuXsllq+dqgVmGJPYx/aKJIGXnyLPqQlO+aUIenZ9siUOnPgmANp9X6kqw5
JkyljpEp1rvbCh5iUmLxsj2XEppISp9oG9D/Zzz7Htd0g5heZ+pQOQuJXJUtwgCg
+r0WJaQgPk2gpjdMcAzTtDhhH+82dCQgEVujPzx7p6uLsWeLVTINDQq0FffeLinF
Tu1jgSp+hYGGWLM5EDJGjEypoY41/61afuG9gF1QJi1bCVF6FK/b66rcHz/s66A9
D+n6l4g+PO4EYdDRom4cK+qXPxS1A8nzKHZ3ByBLZd2yR2SfEJY94QzFhxGoaDvX
8Ytat6p8RU0RWZlPdLmjnyvL2EssdDeWVx7h3C+qOp7Z+qui+1L1ZL/684kuZHL1
iu1Xe6bUKLVQu+AFwPhrDtIN8pfkT3AA+OXoEvER98tgDLuG8aG82AiGTp5BbJGM
rKBfyx5j1StCmlJg+lT+RnTjiEeUnfgERqnjtGV5dKYBQIThnF+GvnMebipjBs/L
3iCgrU2fi07p1B5jcuX8POgk5oF/cbw4Hdodxu8RKY/5bStX95OZIsjHPWYP4UbD
NuP/Fx7vpENzK3sZz7hDvRBt0NNNoxhNtCyhrmpWP65MAfnwgwelyRPSTY1b1vRx
/hWRMpsPfxZff5YGSZxCnnbrSC78cIhaInBg06oGzhL2DrzoUGIND0ZVCLNA4Beg
cSD3uOSzsn0l+8X/9xEPKEwu8LkGt/vE0Sa96mlcwODUIz7HSqVjG0/cilN4MVbQ
kDC2zpKDx79irO1Kzt1bMSuNf/oLVMA+Yi94pT1fItnF+E/1h3ZGvu5OzWHyCm+z
pdesLQ0FwSe+a9hxwy2Smof/OSgQrEzy93zdbSk3X7pGC2J81aJR/+mK47Ea6C6V
i1XtYOCCL3rb3nCO/Vok0mx04w8ucSwQlo42vvWzcRxGA9GCueiZm24jpdEYSarg
KBzIS8IE6yUtsRnHW3gPo3uYStFEX2cMKx9knttHZ77LqanS6+1yjqu3OwLICzeY
7tA0ZQxWioAZasa+0qowgD0mY2Izq4iHCo65vmSUrD4EGaOIT1ds0jJScuCL4ndG
I9WwkYYw/YsSyoLnEC8k8OEy2Nuc7PFm634xe4d3hY1hiwgfOKdRtN6suXL8wZyX
7aLjs+A0vrPRE/0Qn8oWbnmRPuFWcUkXiR4ESPx5RJQvJU1YTui8P23S8FIAYH3s
jDPiHGwBJYOC+c7yXGghwenUmf6JjepT4DwPMJc9RcxdQ/8nW8Si/8TZCYdMCrmc
nFhBok+lxyNAbxkvW/c1QtXzM8AvG0+/ZSqxqQZl4dTi7DJ6p8iRbDhZjxK8m0Ik
aTMIEG6UyZGa2uTmaWubv7YaEj7tPRl+n80fDDn0VHSwBVChO+NTipGh8z4Z78zH
uQXpRlsY42NFSlzFmCu9IYjTFoHSfQMmjcG2/xAwhGCFJQwWahtFwe9Rup1bxPqC
llt62KrMjakgg/sBA0SKqxJXDpAiI6mf+xtu+P+xaMvDl9S234hrpJmqSSjKTU0e
+MgETCJV1owBhyEMQDuPUtcxJCsYqNE1JGc8HJeumKLrJNmRS8StvRL927dzlXjZ
hpJwD9vYd4cS0VECB6IG6PnPdKC55Nu8zTSa0FUmX+fYD62u5sKs7ZdWlliTZgL7
jOTUljwbxq8oY2Z07WRU1pbuep3vRCnvCwU6pLxGqQS5rTIwlFE/hHbxFNLra6Vy
pjCMUal1oSgqxpgvVESKMQNOYsRaGLs5IzADpIOn/etZq3Pb72KUt9jixxEcUTJ4
IA1QHp3+sEYA0mi2ntSmRYzJwXmGOsf32q5ZUe+PtUkWS/29op+nqPVo4TpzYxXf
3zqoesWi7CDmV3TY+ESWV0HUD1yrT0A0eQVScXllNkFy+0oKx76ru5bX3h+mMXDY
1gwMoECbxvgMXvxCJjs2s2tXvEl87+NvchXU7dRnm015xfOTlYCca8dpBM4btKZm
XeZZOrtphv0kw3F0H6fWyW81Y6uGtAeBjMsLz8lqhJan4E8wXyHKAn4LOWsX36gQ
XKzqORCxMgrLZ/gvE2vsKqkQLm8nowdKv51FD+FqzfXc7M4syflBZ8k4WDqlPxQf
rPs8aJyL9U0eA6xifhwmKBLniFjyA55H4zXVHKxCYWL6lh/8CANJn1oEczIf7NoS
ZQ05W1XBHGOzxETa207pNmnd8aVvELgxZN71T3+zOebjunq88fKRkSvzERt9Wwe9
sN5Wa+kgj/xRF9Gtput3W5Dsj10Xj0SCfWh0IAvo6h5lmKmxHXJEhMT6Qxyv8k/Y
S6vg15ZCuNUF7lWiaKtLNVswkhz74KPVvYN/bxI5f4wtlt0GsmC7dmhVtw6aYwvd
TQBjImW5g0KQklJP+b450Iz4ewB96NKVSGlXHybOGXHxNwuX4Y89fVbep9FA3J51
C/8yx58+vfgfzDAgXfVBPARY/tUNd+aSS8c17PSCfwaW+kyAWLztQ0b0kwuMrL/g
Dd2VkUjn6gLNdDUjZqhCPtZYKZeg0sAYIx5jm3SBOYfE026422xVoofxQ1T39YOR
aBvxC2TPTdGKs4VZoiL6zmnxPuYT/VC2P3djKimY1xcxgSrOoqw/8geCEjZps+0+
ZQv9WHd7C9BZPN2v9Kf2AKGfRa/+R5TjupGk2qtEEjzrKvJtNWstVMc4nasYYFX0
rDsEhIYVodiuL9nd6n6to0NSKT0WhKrYqDM4q3B1h0Geik/uFi2xfPAbeiESGA+w
Z83GugysJByKa3inB00lled25NpcsD92SsQzg7ypmtWEqQC4fAbKsiUqXzroUSVm
mfE7tzu/n1jfcHGkyQnFPyRoVp1xiQu4l3B484mtUb6CIk3E/kupjio63wP9sOZJ
6Xl59b7wqf5qTmYZAI+aiQannShcOzCd+peeExPgsMPn9JfadewW1KxkmmMH9UtU
w5zo3CP7PKgMH/DhMn1PgUo/bUd6MVi3u5slrrM4B4YFsplCTDKxfkSyK9y4bOZo
RBqtOEGNxsSlfpCivc6QfSyYxsueXHaH7p0aHLT+diXLcMEastLDQZ9qLwIRm2kc
YS7IuqqwesI3FWg1zM5fTrydy9AR77/zWR46GA6fxg4Cxpe7dyOF9NOg4KGiQl5C
qO9aOSHwov66B7C6UY6GlkQq+ExUR55J7HBtuzrRtbS3ih60j/xYv4UM9WXg7Be/
bx+GU3Pz8Of8UX3Tls0ZD877kkeJvZYMKsU9QcowpIp8lYdSNRrwEOzMF3KDzIBX
GNELrzGgPblbEIozC/91jUxSeVNXtKXeS6O6GRW80k8l3dMOYrlU612RcPrMygCs
Qgp1xuaCOd9szooSZKFMEBZU1l2iFAANtb9nZQWWIF7G06ecqFJogqL+7J8518Ny
/P2/So0/a5WfF75/HHAj6uR7t9kTYwNLcB75cDL4Gdo9/M88B74RRmLj273rji0U
JowueOdOXr6ukaoEygBvOTae0iui4KR0227gugUx4qWMurwLjTe4hO6XT8s6eT5c
zxajVrWLGg6QV9Q0mH2RB6kJrSK3hlecs3E5f6GQjDnY1y5J/jn5KqKncSoGjZZl
rgLjZzYNxULinUxjTIvokGIG4cTMzTKBOUUgXgA6W7o5ThRuWb95WKrqEya+14pl
HZcEQmb8WiOX+LfMKE8woue0CfmhaHg3M7AcnFOdDXhVzj0n6tzAwNZawPAxNOZf
C9S6YYDVB3reobCKFeVvZvMDFKBYlSywmgjmy1LZfDqabUEyHTmiwnDiKvjK65G4
P2Zu/IkvEhS5BdFaBRNEKtUZd0iZFleTnI6MuWfOynQ/WLkiXcX5kbGCGj2yAeiQ
iHtliKxO/0puDyz2kUdotVUMCtUW5GZ2s5ZRgsnqFYYGTHHC18DEZEH8XazYDDSM
QD1LPfYSuCoSRfR/7oiPbgnsBDX9MBjpIVqScCtC7bF7Ef7mLVeuHnM6+24jATs6
lL1HYc0o4JO45nrKUAZEKAflGz6olB8AEyyo0SWH3qzNpsMxGm93fsoIDgmFoLSN
vWraeqnsSkt6WW7cmaYgRd9mzzu6grDnlMuN44GANPoZP8SOVwfjBx4SJIqlOYc6
SxqID1nGzopX3PwOVsSd0W+HSTopkPzq0WsQGURrxpYBpQwDG759++tirbtpWgQC
e76JWQ0BAq+pD7O4WDiwjMA4I0sKo5hH50Stvf1VaLMzuiZRMdWyQOkM8kPB5z99
Fmb9/WWz68z1EocYRA1ga1wiaIQuELHJNJfpZpCAxZFnaRgJsTylmciW92xMoC2G
nAcyAhrHs3E2cHpIRturHsa4SNj3R42pI2JoRyXBcWpPN6iYO0cPaIiFxHPCYMnC
L+WZmvgw/w9+wXjiMOyZz0QpFdloY8a+kRn1v9/ZpWjjOCJeG8JonRo6qFE1nZuJ
e/M4tZOEcCqiqmHPh3a1sWprWOOBitcl4CXCVoVecgVO5G/hwBChcYYrBgZLbIRm
7cuTvrME7vBQNU2PdNkyb8I4Cgr4oqZnusBGj/2JwEdv/8FZvOLHr8QBl3BCW/Dw
S06NxcfBHT3Hqt6K7KDSwYgPX5qkubJn3OZHdgHPP9fr1PabGBwZ5hyi8S7kNjK7
6zsVkDfEoTMJ0yMSuN74mbWnEVNy5jT4VKS16niPYCd6bHkNkhO+W9rWXllINN21
YW2iV80RKu1Qs5b9OnDFJsKfL60DX03R+s7C40ehkYIU7Hu1Nw4kJAdntl0v/CXu
F8Xzy46ZekhfnKudzemIRERSwUCkFUOfl8MFeDjE7ui/cbDG3DC4q5pe9j4H9jfp
XAR5uDxywkhdmBVJUy1ayKk15UVnUDf1SbrmH3z2bmPDjraUqdnt/JoOGx5ldYSe
pcYijdmp9bGBCFnJQQeUnIOuKfDsrP9T6i5Gmp35PG5fcfRTSFeaq9ZjNxXzZkTr
VJTBC9Q+ZRsYw/CQqQmVc7bCCTXf4D+HA693c7pgq79p1TUCQX3FlaqpXLBCSzKf
cjSZQSbTHK+EZyheV9fTAa3x0sgMw6LyReYhIOQqMmy2fbkqgj49KyKkLFWeRfFY
NLKEyHy35IbGnGxQUmF51yY7et+q+xBVWuBFHJakWjybzH/B6KHb/yc+gFZEgbsj
1VwKOrqgiDlw2Sp8UOed84wvpfMCwK2tHPqGwmr2w72zAQ4c9p4T8y+Djc8Ds3Vi
dGiLzESQ18HvmFApc7CTF2SAoW9AIRj1I6igtL0xW9zkyndNsIyQiM2+vX0gyLtL
LLMEolR8uw19+jbq17WLDEojrDplaOINWxqG7l9uj9WI9hXbAhw8Ft36npxzujc/
cX/TwXlCtYRCxEJAbxuqMOjG16ZkBhvxR1nFy7xmzYUV0o88bXMCjZh0yvV3wDng
zis/lJyoqhRlTe8ZSo5qUMn+O6RAw/m2Mm2jSWo+JAWXb+GvkCm2lMa4rII7Nk6R
qmnLZwCxQA2fwrH/a6oT55DJgkfPXy1tg6HGNEgDEgajp/NaMROj2VR7Obe6txI0
VgsqLrLMEm45Lhplxoib+unUvBP///laFU5yagONkp0mgTE5GbX+8p+APOTSX7C6
h2u1Wx01Koz+237sm0enTKuxIq1Urfpn7VooS1H7SLJ4dqas8QxZQpjt1ZwPEdqW
/45meWiEygS7K80eVkbGwN8tN/B0uiBSz3yF+oe1WisHhgO/c6Je8Crg/ImpoqW5
Q4xF99LGqIY/dQun7SoJXsPOCDlCwKZMSXNvxhU7ddSnLO/Wz6NGkbduB0VGSb8R
x5cVY8mQTbFxTMonRrox7LL6kKRoakKwZWvHlk9I1Lyb/w3HpJMefeH/d1p+uOJ+
6e4gf0UqYHH//5ZvYSy/0s8uKJihzu2qvdxOHG1e4i4XZGDUiEMCeCN2Ip2H+BVD
YmvyfsWcBmc/wOeG5l7Ta0a8QF5QzNIG6zTNXAd943pHR7X/m/Vh5uSjCsSWJ6lt
+Teol2gI9o0OjWlMG8QszRwVEuB6ZU8IhQB64Q2mjiKVn4cUy+Ikjt43oBRgoi0D
n+wiB5sG+kn4EuY15bzdEkG/nGj4DstfwD9oGS8PlEfNbaG0xcfPVHyA58q0IyKn
3GjhsQAJc/+eOAp/+a/E1IYy4r9EiHhbyDsdCkUotPoHBpckyxyvxeMFsz2f7sIJ
61LQXlgVHSqRQ6WLTvda/0vAVcbRKMPHgNtpv+5qqwhoWPePQ77pBhQ3lEFQtC07
j1Yo0R9taIOGkzLLFRe98OTdqXKDySen0wnZFB286y4aC+vwjq6fKwuYnbvVAg3v
FeFFeSSTeINKZu1acktWVeQ3ngoRC1DrDO9aQ+ABpWwFOphjacAsnvEwAjbWxNYE
i39l/teK9kMEIeK0WJ12f+jiti0NCN5cBMU0z1ZZwW4WeDLHkvbqwYy0JSxTaMXm
GXX2k1siF7iBy6+bMocC5AsqdL38qtCg3x4VEa/hcS9wEn/bEcWCIQIuLemlJARC
Bl20hzJQJdjHBDopGRHm2z7O09dEqFaseS7lKAsGqG7aD9DT+Xxx8Msq0gSKyHfL
mNzpYk5ft/tIh5FK1Hv01JJTXadj7/yWWJlWXh6kmjGAN3f8mbQZVlTKyTBzXEZD
4wQ7Xul20NmvWd9xE8LSVr0B4ed8VvskUNKeq15U+/vha5NLW4krrAcLlzoDiXDW
PBb7CmGYM+IFiWxi1KPHuhFZfMjsFP63o66VO3RW+3CbzNOuL53Hsdyy7Xgr7qTP
HGLNNHweNaOb0K/olW3MhJEi0y9R7rAD3JOB2eNE0aeiSSnrPFiOcifIQlPMZJ+3
KRWmXe0TEOBG+10NcJs5rsCLb7XTi1DpLR0Fdat266Lj7Ps401K5XbPPjCaYUzoG
LqGqA2fRe+ng+O1kgV1nq8wiv9yU7EFsKvuKxHVNvl/oIlS0i30Y/dtFW9Mqqm0D
jlY0c4gBxvtMGKDG5nnG4sBpbsco1iC417KHGxSTCWoE/GJdtnacwnCsixAbhU6S
Jn6lBlzb939F/XrCa2IjShUndjrIeic2rQBcfyFvYxevdTkZQMxB/6BV4TQk9VA5
WLFFCCNGJ1ulhDdFJRCMUacCQsqe0ykB8e+wqgVNS/gtmHNWNCyDqSnwQSUVr33e
B2QcA7DyCAcJ1kyj8eVX6+vLyfjFRLo6f/u0eBcpG8ZP2l6WoYG3onLYNqoDd14S
52BKom4A/PRB4sozSvOgHlALigNXAt/kGEiaioNeKrbkN8tWRLqY5DBCBC+Y05Wx
Amw0Zqyn/POIifyqUtz8jZx22oRH+SmWVgMpcjidGzd2GaZT7Ea8p4w4tuCJPOLE
HetgS9va0Bg2of8DnutWckxEHQwYJ4rF8Ixxn/8FRpd2yLxtzhcJFfWV+GvYQWD7
NrhXXrNZW6bY3IEqruWEAAyS1GOZKh1sjL9CSyyef/b8hyvMa+JbwyN1HHd22vSM
FYiKbC1KLMKrYoDOWLQyp3wgIDqmZJ5Nu61zZhe671j6bCt+XZt8vIfFzEJrSd8e
unL/xApil49pXRfGed7QFCzJZ9ANMUDxXK+YTqwrcL4JZLg1CL6FpdWDyjnxvBOR
q6zElI5pg4BB8cCUVU3hkcFFbEZoVCduzWvHySKNHIOeJpPBYiC7tMVgx2KVMI8O
pQKjFcB3YG2dDqIOyzQxRmrP/3qu42Wq7sjaqcueOSSuh7aN9P+36gTl1NvGwwVO
TGAX/nCrr8BWlGYlRDTPEfY00oBcbz3RpQrzyY681Z3zFaYy/79bi8dllAFflenr
jrqJ2avfSb0zgNGrDYCiZqnhab+pfaDTCJXquYsL0gIi8vQQMHfSM2QKG/nOqdmR
NNTd8vYC4qwIjgK7r2pwbVLuUnIyo/4p2ThuNGpqdW+hn6StUaeKjybRW0OXuMqF
awDUhyRj8M6jlf9uBtrNnUg8RGiM9tx49qpbCxwS9R90eSvoKtzMzE4l1r8VPYEb
9mRGkffdEKzsTAIQBxeUQtMDZWwsqGfodiDeV9VnfyjjdREMED0ncHvgaIxZ5LTJ
5tXx97V+EnMp/W1/yZY4A1XS2nCFl87sKETfVAvFojmSpvc8Rec1SQL91MG9+2UF
QEuHG0ngON4u1LRWdGCu63PLZ6lBGa8RsCFDTOrs45k5k8zAYdz3k0FV4i4NulPK
JzliaB1BlEGr4ksVKh0GB7L/yMePBHP0xkuSaadCufChrAn++xNzqe4EmofQzOdQ
TC9Y0DPItCa+TsS/tb8vlAHuIII3m7IPOd+e5GAFqE5pldvvwyFgttxbr0nr/v7n
N07YSNCQMgtTzXV2caOSlYnNNjen5mCjz+ZnbDP518DYqGe9pufDPQWrg31RfDUJ
oLxxOTQ5yEY3M74tQhnHEnjIARfOcz4QNfxCLAga1cu6ORMQbl1MPaEbDyQzXQ/y
JPDhLBfi1cEq8XXW7X4cxg6CFKPz+QXSyb3hfniWP+no8dQq5gjm9t6A2uU44xdM
3qhzMiPa8VtuNfGg+aZLKf7DW+DlHlT6XsXRo3HQcPQogERQJ5bpku95AfB9hNuh
FBHxs1vRkcF0lbmvbBeyRhB3Q4PBILNTHrnVzIqNFmCLzH7mlhRNkt2GiOBArKXU
l8vnc05uPiKCRePVr4BMvJ+CDGG5/RpqWv695XhFEAOW7D4qENrizWsDLIC6VcvV
rUT6cJu2BJxLJvR14ABXwB4GpR4ZeC7x69dFyLvOyPpw96y45tiKzG37TYjhqraM
K0KHylhGO5ZUzKfOTtcBQqRtcASaLTfp4cajtg0fkx6ihAI2lXWJ8qUCRuzPkfHr
2CcQtHwbocatF1Nl0OLx86EKnCT2xURqf8JGI46G+UbdwwXJn4IytyCXD5JDNIJ5
ADGn+4Q3lT8AIfcgcBgI7cIwqto0rgA+EP2grj2EK2ntPXymqSJxcNDyBo/DmEKP
TQczRr2cG1lubjEiXHStA9/zCJPzsgyMQBqzLyILtTEa3JZQLi3rHeqoHX8dNIpp
Ah+yGb4DoLyw91pruTotUNA1Wz2mbbuuZLG71YMrfmKnTjTlNzJP/y3LzyqBWXNv
oEmDLLpqTImWj/t7xQdDh1AZqBeUdidfMFZibk93swZsr65/UlnsJBpe9w6/aUWo
KBdHL5EciXtt34jeT+AGoY3yMNDHoc009vWNv8HGx31PpkSIQnr8DpHucXocJxzy
eKs78CZIxwUM6v96/AFmVWm5zO4OtwjkD4s8GMmHbz5j/esSif0LHD0VPDGTOKag
JLtwHb2VJ0odh9u2J3HN9uXahUQbThH8j+jKSbtEBUIe57zVUD1//ABIHIliGON9
rwuykAxe2s7RbWjS+aqnhrFP+lu/IfCIXMZU5RrrdS+m5khTaAH8oJ5/jHCfO4Ug
wnzU1+CgnR4UwslCKgX0FeK2t6qeY4JcxM+QqCfVT6Hi0dtXof6+45Txpj9Bjo7/
sfjmqwRBQAHgCGetb7hfo4zakQRknqHXY0vVBOKOt47eg8ZFEsRkG6tSHqYLrer1
VqdL1h+0Jbm/eAjUxDZe1G8g/IdgT1OzeFuBbE0ZKJzPeS475JGo5pVInp181cvN
tCRUCsuk2jXHT6qgod6LqUT+hsB+PMs0gzKgSptB/zeVuI0KlIEuYZdBLhnj4AD+
ndZy2zhOKflh5QDa0EvwITzdrTlB0GcIo5NeVjeeBW21sVZVrqE4gLhUTkJJ/u0d
L0rm5PjYjLHWuxsnZ8okuxjB0+Va0UT05qm3YP4so+5U9SKCejKwbjZpxK9F9z0x
Ku7tGL1H3HljVVgriQfVQ+VmwFGn0eYnsJ7x2/ytH+TAe9opOo1nT9O06JEsThCR
k9D/Ia5IW/KRd0YM1VmA/JkKs4zb4xosocqaeUewK4x3d1o96WC+gD9iMpAIBYd9
4qoXam9elulppz+ZtsshAN/SwKBPUbU2I6NrBvM2XrwI4Xvv4WyPH9gERYE9vXcK
AinK2zJNvLrO/3Z+I7nFjSSHLNAblWKAfLxS0n5EuHq0MuF1N29NtmzFusg7LObs
teufiOgudOxBXnYy5ZyO8LpoogyVKV0LvJ0brbakmTs2qHVlYMvdzodwyKqw8UHG
KO+F25LprIz4RIdLQLEpC7BCIm/8DqO/EXXidwQiaBSYLfPnKEazelSoQ/jOjjhZ
2VNd/pkHrd+99yW8UPWPccTP+00poUViOabAL84fzJEk1wnMv/JZOJjXNKN8/6vt
ac3eDsO3I5AqiZFVLlJrdkPGFzOwacC44JyyU8QC7J48AlayIGShpirNGmkEDeCm
aPHNgc8x2gAz3SB2yV65CxFa6jZ9PXcpZbuIncfnwBc2zUn/fIZeNNMtb6IRB5Pu
IbjlrjXpgghHys3cDj6n+KcQZa4aMnTOfVfwv5OE1bBoMGY+k00Gnwft+ackKn2c
JHImmYoE5L3tUdYE0kNJhYEYmainDxOV2DKBirJe/hBDta9TB4+a+s87KDZ95cLK
ZnpI5xl+//vnx3Y1E2n1XxBLkei5/lCG0kUNKTEHz6/+00SFv2iNVA054OCUWSeT
6W0ZkzQZXXuiruskyNijJwIOFiaGY7L0plzCyQd+y/5NoY7u+WTXWCL81IXlMtpi
vkM3Dgkc3GuaFqgoLVlsPH/pGhOIoFl3C+NyTrlCo+GTS4FOCkXQML/EVd/+XeuY
j7JPvVLbO4+1bm46in5qtLsK2z3Rv85zI4ckQevR0vBRrUuGGbrf2tQg/rjkYmeL
s0Dm2Q9awG/oXwamdf3hrR8GNnRLq8IG3EowJRjt/QyM9f8/NoelIElFJlFXQ47G
sMHo+TYWXFN9ncfNGHF3XPngulxUBAcnZJhq5NpER6ZzQR7W+STPS4J3Kf8ysG/z
Krko0AQ+xDZJ8pUfYUe3/QacPMgy2ssg+6Q1vaxU2ARGqpYvBKgaGwi5mM+r1KjK
IGOoU45VYaEH60IaRxZoFnB10cGroovx8SKVQOr4N4p3ef/KHqLHTnwc8AmvHuF7
B8XYJyvptfQOpc/Jx9S2Fxy+If5lJhO1rGU6D8B3rIh3ElK7gcBwvQ5c+gN9gHQ9
Z/oCMVfbP6pCDKSvh1QSA/iIE37z/znkUW4TWNiGQEJ59Hu9GW5cFWI1/w1yYIhP
C0obgnxS4wzVSNK9owzXakOuqhD0gd28LPH9JaGXeYafmtcb66JBnEfkmHVb7u+z
GqYPL65KEkPX8lgxX0XVX7RRhYsh68ymxFxjfrjMKXXrRKOrsdjldyl1Q+1PMMYk
tazZDUihRXCPEQ6HFqOTVSafu6jFhPiuWh51kF0JBbaBVHdgEjmRC7/Jpfd7Ow7k
yTBquBOjmcEtmPGIVUf8vBRZGbmxtNImmxK/7Wb3NhyOoKYBjdMJNCYSa104J/gG
ZPOF/p+P6o0bgWouuPujQn1BMMEX3/Uiat8+G7tpZO9q4F1hkbPYIK7IxhrwWmHM
Y1lFPoV+KA+Oaw3xPbhh8VFScGk/cf6Gc01kBypzda/J249WlnZ55TqFrckABjcF
ZFCIZFcSd6v2GHfeUGDcoHSJRM53mbDnkOIgmnaWe/eE+VOzAP8fDofz63bjy3N4
VWal1Z0w5K8WmnrmXnLq6I4KmkAGpIIEmJnz4eCi07UHOWmc/mKWuZx6fMVmkooS
jqXxlrV1Qx+CeMcw8XHVEJvcjC+VaaQm5vwnHxkMQn/u+gT5Fm9diQLUPx8eYWIX
B/39lMw6a4PbMIcnTjUfog7Ki+oKrnaP7oXS7jNVITxwS/UvXVWYkX0kATZi9ZYO
A5FLHIAHvJXKvXRG2mCDkFCGhSKxPEzuL2lUGrZFIIgrcfx1XdjIAs/pf3lth2LF
g+B/g8+iyP8GTOL0L+4K3fu76c4qeyc9pSuwsV/Lodpi6IPbnCHf/mXcnt03LM1V
OdRzT6HEqGV6ieOSTADU9Itr57Qml+HoQvCRNX8CiZnF7naVDoLU8aiMXLJKnHDC
oZiUz6f52572GI/gVSPiYsDLofHpSBpRR9+SKfNm7MUg7cnwxL2MRgmF0WVaZ08W
eUP2IfjODHt1ENadwsU7dPGX4scBpCDp6HC0Jk8NYh5055TCVDWumBNPLKz3aczM
kHMuTWiVs9rotSVkB8iR1nbibkMl5G1MCglabuJC8sGG/3ukr/5hlYU8eXB+RpGs
5eyvK4vne+kE0tnom65c/liEHsDzAM4r2l58FSh3jEBkpeLCTJDAiJ4IKi2z7Xss
c/hhqax9z5ZwTvwY7fhSjsI7fvTO6tAVu7tKJk3GYTK4wF0DtJm/99vPokG9de2F
DP5W3cyMjCpsp9qGODmAcxeElELWXnGThgnx04yMzc+rYtd/8ZWkDhmhVWorOoKw
UNcNkHc4h3QaWjNeK9xGPmYrGtafspTZ32rEanB6LoKXa4em+kEz2iSyi5E9HSgm
FpGe4+ehWm7yKEolxsSknqCciZllgo0qyCuiL4C03dHu5dTrLSuEUFUbJGNVwFyB
68vAZdiMEadCrgJq1KJ8mf7uIklU4SncYHVF2TiKOIHoY6z3jAJpa7aAls8dCGLv
lwlF87meB4+V4H1u/W9SNAaJKVxfFXER8PT0gGMdSvG48tz3hw7Rp4vYQoXvqWzo
aCN4WaqqyZ77UhwsWHaWa7dTZVDbsud+2R5DCb/6hk49HshoKdrvp7CpH1tEspk1
/arJSJf1zUr2g9zxjydwefxjs5n5roSLE/6Aqv1MlV+ZwDHWQ0rYSyzd3cCRnVxx
PkxPxA3WnbFVzmjTnTeXJtAOSJSb3V04TzKUKpaQdY+Q5I5giGdZ1rsSwsvUVPip
E90rAe7+eItKWJacP1yGdfRCqfvEkGDiKXr6MuKwo8oA5rTnnCrPi5T/RILCTQ3U
bggRjg+wdDzkcAXYAWm2/5uPgyy1ZaWwA3QFmqPHLF5EbINRCuHPMCiqnZY50iS0
QvFki8STseaJZ/R2eHiOt2tfKtnI1CW/xx9ITI/mVigGekEgE4Ys1Qj1DQidgEDt
bEgtO+mM4Rqy1Bu779g9HaufxLDSZHm4ik9DgXMaVRntKv6DuilPSRww9ZfE80XL
p8UpmowYsd0jqvEXzqAiQVGoaqCqcEUYFF625ttdIQ8KgJ8JOAc1hSzh5oyRCNqO
Zv83XdL6je625Mr/y7MVXBz5zl5Z+vL089/bM2H4IBTmmUE+ijUPD/2O2vkexpWM
xE/DTle9RUvNVmAgHdsDWoMPBpoG21S/si/fVNQuIr/LZTywa5sDcN7SJM8WAtDO
4v6Nxq0muwzF4lwOb9NgGDnZQC/Vr2fev2wmVBVFS7zTRhBf6Q9sq9Dmy7WgDeY5
rXSIoYVdQ39dAn6RM0HFBxRIJS9k1BZmCKMiw35NjeiSAXCJkbWlU6DOD4ayodMy
OA459SYut+Xdt3/NKjtNyf3sYYPwciKQQSb5TsdJse8asHfBqETlSyiBoOGozNz3
0sT3c28Fc1jkcs9kp3IG7DOSCCPlZOJ05LUOHG3aFSTtFo3Cw/t0oMblyCo+case
4ap45x7ZGt8kaDEJeI8v0lrIT3mmoXC0j+geYhua3Q2LajhbH1Ofoi0uY0k2tVCN
yrK2jm6isr2nMq3WtRKdiKLPWyldBuU8LnLwvbDI+BZD2YdfcHDiPaTX6LrawWhX
vGbUz3Yl2PoHYZCxlErBXnbvI2AmJkNYC1yfFqUBaX4cdGQbxmRUHNP70umUm5Ze
TBxD1P3Lng+ppj9fTrKTVQzkmZEwU9u3U11vgbFbItodfjoYOG/3oxUgQY/9vPJT
ZY5LkBH5JmrMF+POYsSQ2h+l3SWbjAIsQw5TXF+JJ9OT7geEayMKmU6GBS70w1U6
aIPxwYRT9oi6EXy48N5Gxd3Uq6SaMf63aiiGcAgz06Qsj0jJDAwrtZHZT7AlrKcw
I1eM4DiYbiL2a40RpQNXpcLAfafNeGbzg5J+oENMBZURl5/e8FFyi1K2MxffBt+K
RY0KURZgN3OCVPHzDICTfIvN3Gsw61J7JPpmZe4zF/u0kOmYhkeZUCEE47QXSIIn
bMLMvtaGY0YcMeSwp9gQtHjRa4vn6GBmFDHamvejSReOym+0GpC86Br1ZsWfruRD
GtuJKuDc24n8n51ouagfwv3a2+gn+7Ck8ERWQ4kgmw7VGoxha+HTKtKKyDyB883C
szdKYzeaM82XTWpjSNPnxmzcFoy6jtyJqlxMgS46/I+euSmbTuBikrVhUB+Plhbs
rhsLCHpz7JgdGgz/Xri8iQVXx9EmTSb03HSgXieZ2NpXVx77uKeUJpmd2hPT7HZW
y2C355p8eKMSDnYc38tlsm9BeKDFurLRvjNpGbdH5TjAqb0YvOk/7FTBF5xr21a6
7LhW8nizYUu+OSZWT8SCCK9t96B9xAZiOoMfg7MuD6mL5ZXr+xptoBi+AAsfq6bc
tpo1KT+XLmywkGB0TsoF6k2qnKR1aMPu2wHIhE7G0MQyELBx3w4KV/6DzRHWPYkK
FK9KtQWe/5/IzC0BPtv0lxKSHRWc9KbzhkxLkKTrydIg4v0tNVkXtrlsSyb+JBbb
Yj/fqxJDbOaOFqRDvVi9B/u2r/YHLE3pXcw/hVdOEqwTuFmzUP7Za4lEED/Y4ZPv
LnaKNPwRNQVM61Z7l1ubw3IOCPFQi207WAZET4IJ1AvlqPEgot/o/Re1INNe6Scf
o3+MPC8iwJ39BC0YgsHmZbMISxe0qwXb3QXVpSf0SK/omcQrNVarVIZN2M7dchKX
FRCBCVeHLgWS4J8/Dqjam5LJkWz1EsGTBrskckzEYg/cmhlMvKYa7J+qX9KWUlhr
7vUxo9j9IvXT8hiZfrSawwsuBjQqGachrT4YjVgBqtl9Gh6OchwwEUofMQyGzpvM
43jKqH0IJV79StJlQIefznuBjY9dRVI2gUaNOMTB0HlGMLMHWb9xWxFmToCYLLMh
x51nauqVSNqNgUEaq9tGQ0D6Ez78VY+qcD7jqyZ0KDKYc+ooIuAQYxhmj4oRebBx
Wj6RSMqitQKWTTygYbsm/wYHsmbdLrK3TYLd7Zw0Mz3nhwlmMOsQL9UajUoJ3c6D
Ku/JUnyclXubpADuYa8p0PMDUsPeUSxaJcMhRAR1T2khPjlA+5G7s3FC+PbJkLNs
S9LiTYHMS+o5YLVW5/MApnify4a4jhio+m9pWbkVoqh96b1lMIDZli+izV67vqI7
4pfMCHYZpnahOSmq+XJi85L+WQ2exejBmYGGal108J3kawD5xsRUSKz8K9+XpfG9
pvpQSYRciITXaJ1BjM+4QyMx95L5i1JLMBwKZ2mpm8tUdxd3yuAQ4azjC9vV5k7w
QY65Rt6yXlAIz9AeXNwyifckui564jdw6ZasFOP/L/N4iRgHrPJDkplDqQe+bPJZ
FheKsx4nElHkyZL/kznqoHXDLi+AzhL0wbCLmO5Mx6w1c+gtYlLQ4/Tx/5mBG0Wk
NGTGSx7ITDiXq6OvDahEzWq3agYNeZ9O9/A4qqTdFt+hvs1DljJd0pCClK1FvLqN
NONW/IYU++hyHVEUvNt3+ADMnALMZMy2+3x7ZORZBB359dUzwgr0pMS0pjuMNZAt
0UDPizfbKw5oLfjJ6NBvWRrKtfkYR+ULGcwuv+RReZJah+2OJxh+OO00NummHEkj
kAsQecqR9gAxRyxuszi3bX2l23nsqCHL2pc4jRa46RMXWh2xUsmq5TtjJVlwAs7B
zsGLVwY8PWYXUZDl5YkyCWY3BoSdKYl6dLzRLebHaqZKH5kDScWG3XRlvDtBMVfL
EQyUTFsmE7CXIXY6T6UCTxRMiCFGsgnbna4yn/D2Tf07YOl37YhdIvAyfrJHjmob
/UAheEw8w2Z6mN6OS8eGGJzRp0RsWMoWg14OyQ43l4q76ytiXnBtdOm6M7YUqZG+
TGd8n34Lixrim4ZEv3CLFdYV+xhB3guzePPqRUbK71znTJtcjkt32C3No/UKEzT4
r88W52sat8zNTS+3vuJ3G+zbsnw5AorFlsPXkVvRXAsVjl1fD8aeQqFWl4wa6tfm
6dt8HNevu/CmNaMDR/Rugtawlk2bucrFW8qUcHRHVDV29FRFC1orc/kS2GLibrJ6
7h+gMCI0VH1J1a1tC2fe7w/rWi+LsdqY8klwm2/pgEBixZrVWPk4KMsUeOZr0f5Q
dD7Ll6I43B7HxMtM+CvdSjopndZRNIf8eW8anidxosXLBLuXmy7cXwqi9x8oL/d1
a24EN93Zm5e755O2l0addc5Bg01kgny+mL22aaRhD1upWLzd0TdKirMk9Ltwnr1t
tihwnTumFVEiLzbbvSpDHXgNmYrsmo3GtqRrIQ3mk8LF8vpC9PDBqhcz8Vcoasni
rHDKFy61KZc7mH0WwoWl1SJvSbEao+iOj8aWA48x8TwQm+q/kOB8R3yS1IPVGtQ4
T6XzAKOebFlkf4U4s4D7NFwE2AyvqGeIgqVxea6L1PXHQrIu/vUg0b+PhOLDQvL/
fcaG3ydcEAiyp8A9Y69DAMvVA0yI4zj85ZvjwH4sxv+DwvII4PdUQjCXysUAN5F0
3y1a4lAgrl6w0k8SfJp/5ngpovwwpWnrLsvyo7to9iCHwGeu1yz1dNiftzrIKIAP
kff8EV5rBmwru+VPicKdBbSFRqsy9na+MAuX/0mKrJva/kO/MjYslLd9g8u8QlKe
dCyorZsCRlm7NwZ4anHdgGwTuiCpuyBhyMhmd3XHm5yUXoElXbZb4VUlB5Vd1He8
u3lNIw67tmPqAz8L2YgXZuhibyjZAjyQHfwKanlc1YOBvMbA2d9HI7hqFuYGJnhq
G2EbjSiSf+UMBfYBeb+OXq0RSugbi6vIl6fAsC4NxoxW4eKewJgMVNlkKBVFJKAa
RKNLrw/9UelABZixvAbVaZpghke6hqWP3XKoOSVVO0OALmgQfQNIBHzlPTw//RMu
4VA7ch7hGmxr2GbrAWIr63C/SuFFfyZyTtAMcFxcGS1K15dGqVS4RrfGG5VwK4d3
S0gRPfoSeQzpSphAQHHnO1XZ+kB/SsLPvpjE1DpPgC5quGOYhuJoYzLbJD6nO7s9
//oGRkxQ5XixkIEwvnmarXzQiBBQC87PWIdRvnfdfMeFygush0WSqwQxQSrAa6Xa
J8gxDx2DQY8yAa63ZyeVu72MGLsy6dtp2yGKrN4XUPugfYYmwTySiB/7OoQbvc+H
VBW6RLMVM0ibWLIwDcV3eyrCAwI4p+NSuivkLNqnf1YhaI8HZ/1LRmkkUVYiLvEs
Bm1HLkjH4WTG1BS8A73BQC3IEGgoiUvwC1dlV1zmAP80EWRPZbSxLXtdBTvtxfdO
yRnkJ9rGYGY5Gc4bx7+8W8WN/dDeT56f/8Gz1oCNFss6bso0XTu4kQrRu/RJY1Vq
Ip7ZSaV8zhzgJoITR1WFwzefXBktOPKREbbVYgkcEK0qhyIqXADFS8ayJuCsSuUa
XPUTq1gRB5Yewt2PEeiddhQwa2Tj2oX+85SYGwM4gedVgN9r8DY3N8VHwft6fjim
qR3xVQ5PupljZhHGn1fyi43QmPC86nxYgySq5EwOpS/s37V+McoYDpRqjf1cYCQK
IysQZcvvMrRDAAyAm5ExnRee60PfXk/nhq/UFr17BQi+5CWl2an3cfuWcpvtnGWX
wHv6zeODuCitBrLxSUiwA6vOYhKcge6Z28bullaGLbhHDNYGyRhGp3BR172ASLAq
MKoxvjsiUPan/VJOJfva9XL2g0I4pLXJkCg3CCqV7p8lrjesTcK0nk1AEH5cRXj4
ccAG/qGbDK0Hp01YD9160qnfZ+421X+xZpdXbBaWUpm6b8mJMdEmRhZMVcrKvrHf
GRwSnUb8qF67WnNtZ8ZdVKABqChfLGEKFBj7mpim30I6wdL4WJ+7pn4A05sUcyHL
DRKxmNV9JAKQlNaWZilpxa6CGVQVJsNTJyV08acHrI/HZ3eVvkCpHAEFNUP7U+EV
tURYFjNDBtPCcae+JTPBsUg0LYPIR31jPxIKMzaUwyoE6RJg91Y9SnD5u3RwUOsj
Bryp+/isCyfLULoAjTqvuNiWPmSdkQD2pmHGuoppML+keI5SkOJGEhuLs9xAu2V+
Ssaqlqk84dJzJ+Og6COmORbSL+R5aUPwtzLtO5gdOTgaegdxi5fckZKNUGqCjx9g
Gj3UK2u/Y9Ckzj9CjOp/vehb2rgC9S4C1DnqHpTiqVHQFXEOTgq9+AdZvtFVc+Fn
o5/198LCSXuNHrZ5nhjX6Ha3nVh+dFs1ulzXH8Ox+DExm6KZZRnr6lGp+pGUVslt
E9/yCNVqGU7Gu0XFzp3xL+52ZS2Pj5YzTnd5fLwtzIwodlEK0X8ZwNPqlGobhXr8
yEfXAnsksALbLOZ9yP1uBmjN02FNosW1lSwiiv+6sszB/v+jYktiZXF9yErPLVF2
j3KN6YeOWc6g/GPmK15RQmmWow6/gI2lOOeUcavN9uZu1Ypt0IaJH0BeC2JZOrhu
jNZHfGSs+M3cZb3NvisMebepSckAoLLgUeDpyktdrB+d9cRS4x53rHjTkR04u3ov
zsTOT5sYKjYjTLpLNuLkz3CX6WcUTeZJ5TxOYG02Kpcb8w911hys6IhspsvEcm7g
ISUNTgE8J+V6eYrcWSjQepWWSbD37TfAYZJ6qct6WBdTnst6KMPMDgQF/N3GSLED
0RVd9wNZ3tjzguQplnEFbKBcNsxPVZK8DeBaYDmTH99Ov0TyD9eKU7oO/Q2HzOiI
L9JSICaAyqnRD5wtlgm4w6E85GChtuhVCk02O6/hf+5/A91droHl+rLJfVA+ZUz9
ENG5nFEsTB3PHv1P5CBOSxxwoCTZAInk9T8J7ig04OfvUtgtQYEvh+FQCUYtEcr5
nXhNqQ5Ok1eRROs3JJh8cgzYz4sfLzE+kkIExU+OG+8QGlE67v9Tvg3Kuizcs+Be
qo/alfCgK/JQ8+tBCT2zYo2E8HqDTsoiedBuHM+Iev2aQFd7MIDa5pzrF6gz5BL/
EwVKdfip5BqD7DY8WsJ69zQhP0gDxjtqbrnfK3WGv/LZm06mrJuIiHrUpSiE0UrA
0Qz343CAczINZ2rFAfv50svpPnDFWbvqaaQM16A+u/K1oNhlruL98SP9wupp6WCN
6ehSqEDaITJrIWbSKbwQQ0qVRLA5CVo7CfDmYMPaCEUPB8Se/9Is9AaXMy41uSMZ
QjluqULNuW030kzz5MVqPQU1paXSr2T4YxHUegFb/vo6xUrtmyyN0FQVTR4QSFoE
45T63eLhRQ+Dqkgul4xJqwveRDShSr8FscKPJgJ8IXnn3g1yBBp5EtgX82alifjE
Z45pM51e19mXB5we0REmBgfv7A9YH2ziwa77X28VnIaiBjMzZY8jT77w5xmoSJXN
RZkE77HCkQPBFpN5YYSDBjqrPCLV4FZlNkpLWdN+V9pRqOXGTDI1wUePlGDeRE7S
JXNy7+vHsmw2YuaPKNsGJVZeCMIdMKukC2G1rFlIDQoSIJh0YP4XmWfaJk2Ke1+2
g3aN/LHWsDwX+GXzxTQ7KJSVxX6noF2DhL8ueMCXKqudjmB+5b5NJZeCqjqAL4Gn
yv2KmMOLu9puMdt//LQCNtNk5sQxcgMQ4nkFRM9sfDNIHqB7yle16jlQao3L3qCj
/+6M3+zlUhhXcADZTKaTH0Oti1GCn4HpdccIiSGBf6zNuo1BfVclfQgYBRGD1g/W
sV1UG5FmaQFVu8KSJ1//LWM7YClyNzP55kWyuzKejOT+8Uu1S0N+Rh+O8mhKWFvQ
EOwH2SkOhEIR2FL1oy6/NLo8T3nFJesiapjJLOYR6ku3OQgvXeHjAZQgxZE9IxA2
sKo3PVl5KusA6kCbYHAMpZ7pKZW+CRuYBnTcaPyu5OuwQdpwxWbBtaCsC1HU5qrw
MgnkJwmjcLjpzFdBtwgdAZl4y8fvUPK8tcuNBPAtj3UAKKRSEq4zU6NqpKOAFV0d
fuixSoeypZGZFu3exSgf/RESHAlsRZj75EKqiRIvVcLrIZSb+k5qZoqj/XrMeCUU
abUesIqu03XTw1t/DJGdrr009hzmIbVRY/YtUUb0kInzaXihuWuMSZ7c9UpMIbrU
4O21ZsvYJ4Xtko5jyEfLaze4/HX5MGTA3be+A5TfbzC353j9StRaWr1gSCBvmYxg
1OO9mXMw2GWMX5tdpIRSVWD5/MqQseF9USHWS58Ovu/jJBtL2QWe++5UCb5ZMost
lYSpmx5i1WZaYUhEZZQAoj0/AZrJzZPkHUFGjdCwUrBGVYEG7y6whm1w1X5redm0
AcKzukNh38JV0DQUfsAQ007OtR0aaeYQmQD3Tb8kXdwY1KL9P9c537i7RcSwel6Q
/mvR/8yiHTJVjdMHU/kd5EbYpdyiL9DwJw7As0taC4AFibbC0cyD0ta8n6ahsF6Z
Nn6DxOL/uU/RyjB4jeAIpB1v6T1VoXSyYTmIPOr5Ejmpwcwuxglq803rb7F7e9S2
PFrkRDwtKSa0Sem1FfRHq13YsKBua/1JH/qyS+2DZ2DODyunEqqSX3Pu8Ux2P10u
BXLIBaMxHUv3PGZV8sKLpt2A/iK2BGCSLHepc+zKyySFkjth8NwDH7LqNzmSoDrd
YrzQ5vLh1jGBC19piHHQ6X46SlWgUJUBvwBzwVKWvNx4SVZ5tFMywuieuK23mEn0
Loe1ai5nM6PPcCbHMpQ7jykwRNtqXLdL4BWSt0SGXEcAamO6Qxfv8xa7UNjX1gUO
3iWu4k1GSvU1vWsTM5eaAO7iB2hQJImmKUYeBkTyAT/7U3s4CAKyr47lcM6UUVec
d0rmSZjw7sr2b+JgYpYObvMX6/U/BP+sW80giN3Xk8X+ckAksLtDXAHEvFyX/YJC
NuSFyRcRziR7/ivrAuzxxb4rPrV9WBW1LHAGbn1msAvlcMDMmAkf2+TpM5Ff8WLy
g/VbrQqRoMBnnLCCvynJlKeZb39kcA4wmAv3VB1u+e5WBSpyQsIrqB2XOBUdDsa/
QQT9z+9C6m6EkMn7zGAhr0ynsZlGDGQVRCsQyXVXlebGAxR7yTVu8UI8IHCY+q+k
BMXkKVV4clKvJ4oL0JyXcs8i7sg6GWuO/ryUJPQoOUtGoo8cC9odMu0zJ5Z58W4F
1rmdlgVpS3olksY/6fZLuYoq2YFzzBJNNe0HmhV9YT7CF1hKrHE/Dkv22l2iduJS
nsklHL502cTBYK/83qJU5KIeDFoxkHjt6rPjYAbveRjt8M/CcPzk32hZSTsbm1PB
ZJEigZ/ffWYuE9wtfKXmcHJ51d2tm3PPJ2hVETvGQ+m2HARaiuf6bw1AZihnL/2W
g1u1DjObn07I3hwP56CGCZP05OM7fPiAZet5IjR8VWTKXsq5KYcf1NHdFynW5LDg
7sNWgoYXJo59T/JZ0Mt2Snr+atv7231hkIOs9s5rhSSFznS5NspM+PkN+IRNKnha
H/3ccPjbvXyukQH5sj+qul7ei28wuuwaxkk/N0Fp9RcQesgFzAz8v9Ynet9SOehP
5e8oFb2YllvwpDjUVeyN02hPrcttxYmuVxFwBqZv5AY8WNzCRFan7tADJkziQpB1
ihsrIyN2MatRJgdMKMhw08j4JWj3YL/VdDdWvnrsa+CGabZtCOdonmJgdJpTunqG
5EHa5WSmXQnS690bJeQj8EqrqAuVz7ewTiKI47I+VqWUgWs80H0io81yOb5saqtU
4O7cRid1j2Gzjr/n8AeuzCoFU/bua2i0gd8pHZHB4g2K0x7LTW18XuPQ8Q1AZeIZ
JhQVK5AIrOW2zEJ0kNfhF0bbN4039TbbKhV4/3gMDTrDXbxZQAkvJZC+wf4I6n5r
z2VLIBM8UNW0GwQRuTAFKcRmoXB9Xp36zxbrMszUY55oIykGZilm4aOLRgt+RgIw
GqUynou8oBcdSfVlQ0ZFtALMARml9lQuKb+mL1xx8lU5bF/h280K/o5K0fsC+0s/
+eQQ4cqP6SLMhO9My5ZRc7XOeT3e3ZzKopt9v57WAAUq7BEEI/3otLMVpcMFGKUf
irQIv6TTCbUCj9BKk2BpMsdtq5CkzJ/0RT4jfGXi6ab+Ru98DQdtidXTpcLkVElV
v3R1jvvbyHhcIDrq+shix9zFj0zjVHZb1V1pVycgrPQjUrJHCzERKPADF04Qpa1Y
TUI1K2NvfLsRd1CwTYdmyhYHfc5WRPFiu1WRRBih4VpyaQCk6jYbrUfHdYPswgUM
+04wvSbc5ReGsnx3Nhkh17gIfaJO97uqB5yOiahRm4VQKrmgax624jheCEC4MeV0
qppX5VCkHsSINi7GROVMNsQ/Eg0rrrTRxdqHtWVcogNEKFhZ02dv8QcHcinixzcD
/8KQ4IH6/0cbzZOVcZhdEHQIXcgyClmkdHH9vxoiA/Aej9ZQpEGtAjV74xXRbBwi
TrRI2B3gEJRvuzZRcxVtD/ITlRkrlOa3yQKojt0AIEsI42SlO3TMAmCrb2cbltBu
M/wjw2YTR9vxG7YQ8yngdQpYaEJTZl7xoRYof9A/JvFojUOiwi/4JN4hkNpvFLfm
WG1+8mAZE6Ccc/EUE7mETlsgV04qhyqDGTOQZuAnrwm8Z52ghciA2zQDi2N1zUd7
y3VzNFdYSk+rAAgy7HA+3BNIFmPT+YPRD26bmo97q2xQcmI2oZ3RwuxP96PFzU7y
eHt9/fc2VMPtyoNHVFkEq0BLjIms097YmKCWKTgZHFuMReWmmg3PZxta9B+57udt
tKWB8jAy4Y66VLKzUiJaE3cHno8PqwzvO0+H8nWxoYSwbUtngXaZPSZpDqrNXhES
SFvtriRNrUp3YNaxoInG088Pzg72aA8ZYnvsIg9xofgrCGRy55zc/b9LKCZnFjSX
9Kf25Qx2I/5Oux04uXNbmTe8AHctHuzmeN7qeLXtPYHKD6cu0EVXksaE0x6Po+MB
9TnhVTfcfr0131UVdBCox26SMGnRR6ybL0Q/cjPDn6WKFLYlkswYO4zpAKBnkhFu
+/1/dcEXw/5mcp4ltyIHTFKK7zPRE94FSr+86knlGBhBscI8iIu/9Dz7UediFgET
AMhoCUf4iOkzuddeSWFYfSmnuPqtBvebjF8W4x5a+OibCaKxKI1DLUGL8t1B1Vhh
DevZvE3k/Laz/Juk+A8/4dIH/gI83ZWt2Dybo/y9XUFfaDwOcSVKqTiRsXwKpIJv
8nfFpe8Tsgq4iF1v5pxN4Zzetc4Vd+5Jd3VDk3fgGZ55G0exJRFESPt9aeRX14Nu
udUfVH5VnsLs/fBR+h7l8HCeakZ1PSqCtYA7QuDbXyQP5ku9AwfMBcLRpbwS1DvZ
FEfgBaodVsFWY+33GfQla0cAxtfwWGVcy2BiAwe3pG3+tX5S3W+cZdObnSJ/Ard2
Z9ZsR5EiLnx62jpYjQ44FJTtEH6d3UxrnFxqr54vL4D+TKotv92a8hl76a69FmWS
cWV2J1mYGau7KsONnvHHvx+GOSZtvIXNv57LW2aSQlGsmfVa2iArpP8CYtRPyVXj
FL5mbzbpNspHsQ1KsWeP3mQNuaXzUc75WA7BfcuGz1dq3R+Qja4Yxf82C4mwVnru
+oW0cc7u6tsWacEVr6QZIumkuKvk963+eozkcWEWeRamtapfEalDWQKmN/gRrhgi
g8mzMI8vmxUoYXM2R12HbQNdGBMOpBji7keCHUCkYf/Z7qzCtMjX+Eo3BImVM8xE
nxLGTGUcWLCZbz+6NuLOi0V7Nl9JLb5VRy+6sJO5MU+0f6ZOW6z4xfJ03l/3g/mE
DcpggQir7j9//apFCyKe7OjmmV73ekeNX5N+wkN5ePD+k8Ja3ohmPr/TaxkIGCxj
UTY4OwYYMiYPTc2N9bPnE7kD39mHbl12xhNIIOe2udZF9pZzxs9fpazx1GthpVzL
kL99UKMp/rw3N4kbTBCIsJa18qX/1bP9T7W1vESdGjh55t6RA62eM5Ea52n9yi5M
HufQa+rQzZ6+stsXJkTQTTsuHD0Uv/QH0L/f9Zr6aW47ZguT+iXGuh66fDOu+knn
qzB1WGxoC4giFj8zgizWIwjcLtpTrGNLhvjfqTXb2c4lTxQ6rnsIfifiB5X4tUt7
KfRmV+vWbey52rOOhrPKsnN5EnZGJppDit9bIpUjBhxpKjnUS66GcKw/iR2bRx9f
N66Stpp/EbpjdeMsDf5t0gu4Gts2KIigyHH5/50uw8MYUxF9rssQmJndMrKmI1VG
6+Hvc+QD6PlA2vC23aCMulQTVFVBtfmaPD7sEHyrOpBwOs7JSN39pfdXA/UN3VRm
/RT5ZHrGnn78dfaf0Rv1V6A18xsFjFFiDrcYn8ASlCt8rM+ouQrhZ4cgelcI+WtM
1SXleZr/cwXxYhbAmYhIZ3JXBZyUv/6o6QPrUCZGGAKxHJ3pyNPZET/hScbetmH4
QvPd7LYnI8DisrjZWPhHDuMWho8cyo2nuRNWtDib/kVy09q0DeT/pq7H6edH+w+X
vriJo17Aqi1/jPj4B1VlgsZMqHn5ahen5NrljET6CEAYd0rM1b6Itp8p5TsY9XFD
nZfWvGdgwxdHYRkKFZoJrkiWE8P14Jh1VTdqyI6aNe8cYgmAcsxtAlC7ZcR+v3x5
D2xvz7vRf/Da2w2kTiclUCpKsXRUvzQ/M4UDxwYkBgFH95+JKdEeVFGzZF+2jAkf
DGaIGy9G83Ym+HIUGL6EwshW1Dbx6qMq1EOy2YAuN4r7/kQWjPI0Erbx1XnSDlM5
wrROIhSVvIegUZpLn33iCSY9uggdTdbULLomRiL3i+OzY4DubBMIHhNjOHyPlX5i
tCfJjwjtGJKnymPupjXgYAaVcxTGBhZJqm1af7cnR+dSvBn9QLNznlEnIdIFaH93
gO6owmJul9MiGqimfki/iZ23KG/Oh3kb7iLwz8zxCVetyo9h3DTKDekws3hmOnz0
czhivRmHwEwe3zgn6MYbzAmwuKvXKwG0hlFcrTkSM8WWL3pUeEs1wtqsEwRDgWtL
2YPER4yX9HCB5eAFyKgcr/bPyApF51vTNhLk7wZVZO8CUk+JdMzJhWLtRvwexdRj
h7Fx6AyXRDI/S4w2+K5GpyjYpTQYZ8aZlWgbyPFY2fIEpPZcYdKoHpNuKN9CQysM
3xDGgDsPHHRkdGunXPhs9G3WvZl8oe+7SWrT7X1R/eb4ZSGE+IC54xJn/0NLQVqh
2EtKjmWi6KW0OGe+ohtL8Ch6ejPXEH42AZLZwJBZ2sOcR4OhGxHnXR9s87kwso6k
a5GZQPJ9TCwAbNRNGo/0MGvfI32+BxhTZdnoM1kUai8s0zsnPIcJzevPPfuOQu+D
KldfmftN9vpdSsnCiuU3BQBCHf5dM8ehYwRR/n4z8wd9uwjNWMQz+trKKtPT8R2d
ib9ota5dsFdYFd7yx2rhCJ6bHnKGu/jputpGng0orl8N4AR+pcF1Z5n2FROjMtxz
v1NtPhl7rHsvy/soufbuuq7ItJkIHYHQSblUIvkIVxqpZIScinTFQ50JnKkBBGhk
vtL/D5RkqzR3sUUR9/m09ag7lvyQi4Fh24dN6Kgjq7ztKgbBfpazI0CwdmXVXRB8
nWquvy+PEaKnvqFBoY+sgDzSS5HrGTQ1a1INAD2OLYvZ29e6H4WjS78IZfSnBaIi
NHS8jmVZp52xre1guc6ims1RYP45x2UP6CE5uE4W2ZLJCKKejNR1JMdZgNot3lyE
VOZJtheDZRZsVhWMm0c3e5f44fwLjlWMggbBzvLvVJkX27HMJmfr+BdtNA/zOgr/
+cHRGhfVrO0n0RfKMkfzQRSNUqbMJ4hw88M4LlIVFy8g0IXr07PUyvsRsEs2AxHd
+LvViX0yCTUY0PMnb5k4UlR3d7sYbsgemuyl2wz+NelGSVS5Aoq9wTxdN8VK8iCu
lRXhQvFKYdiLRxFhUJJrs2VJGX3MA4lr7sgAN97sOAvJwOsDPySMhMJ0tWTZ6y9i
9hyIh+J5fE5JoBkrFNmoF7gEw+5s9qRbSlgxV7mzjSWdKsycbGl8qamdbOZu2hdK
kpwuVrs3gzxLTScodh7xtL7tfWbp5VrvIi0eoV3NvM9PDqcx32LjqnRXJCcpqc+G
MMqeHDWPVDRDAQYTah5pxiaGv+WnZkMQ+ywZBl5/af4o/kqH+v5Nqf5QxuKEOF2+
FgwVpNXCvQhi+pDa1dcOjyjp3C9YW43obmdJzmSsptlENG+NDX1M/YnEI4xKq8NW
lIhtIx2P4HFgg4/Dmh0uKP0dC2+CoaS7rsGdlMoHIabBlZMlauLCmSLCYNC97g0e
TCOtdDS3jhsXZ/u6uofMnGiR+/4S8vA7p/POZ/yQvgaSfkwKXUQAGbGZTQvw+kE/
MROe+utVRw0p/9u7wAF5/hX3K6m7kwX8UXPN58WDuqFC/YvcYIhz4dCmva91weve
4czRQluH15HUfLp+HgpkH1AKcsSI01wiLuNikhEXwvqo3qU+z+Z7ulmSbseM9WjV
U3Vu0E2Ax/jOSB6HR6VjeWcNvK1XFY48hWGDBSDGA1FKErURdFasig9e0vuK9xXu
MzICPWcmj1qqMRFSef5/L7O7EKHq3ZFlEWhkBEtQeLdz+1nOkiv3geKvPRYv9K7a
kKn8RJXKtUCjRYnhRwK4/RBqjNIWAeCXS1qOldgQGEN9vuka2VCq2SwHWPUkXxsn
kMGSvrw8qmnc9yyMj4U8w2GvjXfhj8ABtuu/DZ9K/Ei7KM8WfbYkHdFzQpqW780w
yg2PzWUOvaxbhFUbylisJwgio0cDbM6fyHykUDycKey2PwN8HqBX4Rdcz3QHRuNi
EI0mvdlGmBaY70eJdLzrbG4tQ8JdlQXvEgel6/G5n6U9e4ypkw9BsuhF9sOTE7Hu
7zR7PUwNHOfCpmHdcbCJ3jUXtEl+yPzLWxehaYxU98X/4XhThjt666vSAEn9mnyB
qrv8fptAt85SSK2dTe9IndESqF82gkWjC3NKAKrQnfmE8UOCZaA77Z5xsb73vgBv
3iU8gjw5UPFaAZlTY0SPtrMiCI1hueP2WwCq+16rltx+T2zZcrm79eVSJc9+Oan3
e3NqUo4VU84jN2IdHA7eXOX6vXGBqe4rvFnG+fKUPpp4QNKeBBwX+pj45jP0wSne
n4M5yugPi4RYBCj931E08pJUtuBinMTo6PyN14N1zN3S7GIqUV+ecIKnYFJmR37i
y9X2ZDL0SXSiVVvmXwN1FJjeBD9bPsyZ8U8jM4lzKM3YpAbgey3Dae+BkJlraXjA
3EdUxerDSBvdDuGilXnU3z+Z5uUx5k8P1daiVa20XyzdpDipgO3LuPGdc3uORSEo
GyttPsvY2XaHGaq5O/C1QiU+tO/FM3zezgm6c7VdSwR4lP9RlGPH/60HhjgVdG5N
0tU919+dX3YjwRmN9D+dOTWdxnwa9gQO5xFOikB8tKreyV0NtqT2pMRT/NeN/qKn
cZcwpn0Msx1FPCGW16CKKqlPakxUKzBqg6VeXE0aQ+sWxbZinq71l/09wRjTRYbu
qENH+3nGPTKVShsggbV5WL0zvdmXnuYenZuHejjhV/I14k+40FUeXoVMm39etEp3
DAavDMAxgtGyMfOvkxbLJ6yLqrdHwW7z/eg989cVnQg0ogqVH3JR8n13GTLX+/i0
NgE3tkkFqZXRYV7MzGKXTPgpKBp+wzyJm7jNuX4pN0aG8fN9xV05/P9NC1pxCpaN
R3LOJ/TtAQ3SyBG15e2vQd30BpgCpv/1aANmNdRv/FYJveqNstAFYx+HJtveKD21
DxqUx1IfiKruFe6gMB5cyW51hpNUUHMpJ+IcCdXCnlhQ1/OYN5AHjlpZiPNBgz2u
PL9uHCtvU3WcrXuhadI8p66odWMU7AKW9iBq8yK7gsbiUbBwWPVbceOOJyaKG6O4
yIbYyIk3qoyNks2VGHE/AM/fFg2J1O1cYUgl0rr039YswtbhZtdMk4ymkZbJB1UK
5sVXgoTZub6pNOq9ORFsxinNlfo9+YbHKEg35XnwY2HFr4jtcr5N3tOkMN96S95x
gxx80BYKXsOjZyZiZXWrTCMz4HwVHsUmCvvL5ggrQxCtURr09vmL/1IegR03+WYP
uBkxzdAFMsZ2dKcYcPqZlWueFjXPrUZ745bTnOV9w9UzFSZBJM0iAZhb4IcW5yz8
wnFRAUJQWuYWhIO3bMQZIybwRz7fvbfqqRQoXW2z6fyMXodmRCSG6x6wr4AxBwK3
SSXaJak0DhwjYL7sXttbLAR8yT+PsJBklJJUtvy2fpYclx9h3yckHnqxJGcbSMgv
FanQVva/KXqteV3plurNLiwUDm7nP3cCERi33GdnAYkLrmHXhhTl4Wgjzz3XANft
098FHBE+4kWRHiLlXzvapJmPHSdMvZ1sb6AmeYSTbYoGMQnO7R5S69S97hMCb/52
TYC4RaTKpIFDpL36D+ZME346cAJtnwTvnJvX55V26OCQr5xn9iulp5pPxiJkSoay
8osKo/KfyFsrBDk36WkYUYH39df7nxEOJUSZRKgEgoP7GeScDkSlgDWq7G+GVri8
35I9LMMMAdS9A8t8lyGQq6uz5qZJgpEXbEv3WZn7vmxyw7bmcLEQjgrq8VCrzIhr
Oxv4GU6xUShfGA9U4ZYx2IA8sG8dGBdd+wOUrR3qObq4EvzXWry+Tw/s9gG/9DpF
oITGEdo7YiSU5DjPStjGBXNTPh35ETBTX542f7q+L8Dy5dXqzBumgpdFpJtSXTHE
K1WzSzdlBQULG6upLRUr0qmj+ZGVxIcTD+OcjlBsH4HIqFuQrbgkOgOirm+vBNlQ
OrOs1ZzlhSZUKDbWk3/NT7urIZ8pATk2EfbolPCcunSGIEMv5yXGxT3GqGzXaKiq
JcTMPf5QNIlpX43VSIJArGBJSHG0rfOdz1223fPgYc8dNB+/A8JnUm0Jcj/PWi7r
peQUZDXM8Ih1ixIF7vniQhh49FxMwlVXIBYfqBCrf8gl/YvN/IBsWH2x1MdxRElV
26CMbmFUUU863FPKh6+dnlVUDxljwB+G6aGYKK9fX429Szu/JHq3GKYkUu744Ffl
P4nJNqHPJ3ACvGb62jsPRYebi3pwvDJGGEOy3egJak7wcSrnbbWcpkzhd//syGxI
OP5/KIk8jwj9ymkw/v+eifcFdXw/ugyF7ur7XiUofoYiSPBqyNuMzo35Q9er4Q5J
ylo4Iv9SrV+B9bnOiHdKMQtwZywUz5r4078ia6AChZ4s6+EdxaOsxfoX0NdKRmfB
qjjYKGPncOgnbteb+Nv/2jzXRdZR4rHYrGs1mzeQmCOfFfrFJmIt+CCQ7zk1Q+4g
fzEmqwXtqRc1IEj2Lu7M6Wcl6hFwyjEQH+ddN35iLL/LpjOr2f2f2Qeh+1NZJoZV
3/SMyNEkhltIPd1b4iECioFIvyaXAhbWRJB/GT1/tZsZaUIOOyGnr5b8EMtx8k3y
ejqW5LvKSqE4miytNPqxb209cBy3pV85Ws1Wt3z3ULukEUHK0MQiFXs+9FvHD6YT
se5s3ZUN4U8GyieL87wqS90hWRfbGsBl9vCs+Cl+ikPhHwJ474epY3FVBPt+OY42
w0NIfdoTen8M/qvPaKaH8XHHJp/RnhKBVlQBqzMzu16FllSVn1USg3Omre+RgjTl
3Yg25Dq6krSlirnrNCoi0GGYNlAlw1cUPSe4Jp2p63ugkL4YZB/se16Fs4mXvSvk
U4LP1iChClJOHMHX9HbvaAzZOmDczszOk7GlUQBvKIGiRUrafWym5ZIUGy5iKJLy
nvsazmqbhAejRuQPusluZx4hetA+ScBFqLlj8/mBis/ONkuq5XMsPpiRnx95pzEy
GGWHZJX6FnOEfcdZW2e3kGQN4oMhs2/yVa168J9G96Eyjfg2AbgtLmO1e1A3q/Kw
rNr1ADyNBpz3hN8J02Nipl1rGmLiwrAvXWcQZtGVXJTeMWN2dB9jHgfNh+myNNPj
C7DIafSjIuc2WyRefgJgo1C4sNuN8DYW9aE8wbhVV58Gbfpc30k96w2UjfzhK5Wh
ZXEH04VdGXE809i5FIoM9NgBgDetykdXlxV42FPPnxqCN1SKdISRKz8W5dbYSW85
ps84DY+8yapDVab/yy4pC2YiOHXjDOf+OonrxmAw2ofusFJ98EqgaCKRWqhgx0C4
veHaI+y/7rZY71TBDMyoxXShnPlD6D1JKSMneBwNCDwtINUMQ2Osd3JxlKbT2LW6
9ZSoWgAV4y6yuC5G8WMea77gtU1lBLJlVRsVR99PVuS8P/5bq54AQ2WASwi5Qi0T
x1B1CkneaeV1uowUn9W1eLvn49VzUM6ePWjPUkgVr7vlTYz+7bF+wJFAdg4i04X0
u2GJ+GQf1TcDvD1T2vXaDAebLC2tP3KcfCDaD3fwv60zoOAuTfd4GKvl+tIwoWR1
ZqYdIPzVlrXgcTVpRAvH0ojIypSuFIe7i2JJNqPuSipfhwWVCf4yog9gL+/PRdYT
MQc0OPxAWDgOmmC7O4Pt7KICSxwEq+js1d3sr5+08hVv4Qfm1p0DD4ewqv4Xe6FT
x6NhQ3RvwE3HfndlSpKK50z8EaVPPLYmYC0c69RLHE9smTUrrfKrDH/7tRPMYSHC
e8NCyZN3HBgFfxrbEiMPfHasvTEvgJVwU9UbOASzO0bSYOw1YwgLK3nspcU8ZajV
YMFVO0TGV47KgBaDkb3dVb8u25kVCDrFTE0cuWhotzcaKGj418lLA5OkIvX/sq8Y
ZKKPliCuYz0WjnfZ2UA0tGv4TszcskY1JXHTZkBL9ebPdtlW9tEzKSjMWivHrCF9
niAgwtOZ+nUeCGIfdSwzcBdhhytNtQ7NvdPgodtamHdl7GIByJEefejcN76ENO5B
sIfc020yAwYgdlO5/hnfhDhCHad74JGl4p4Qqwwv2ICMMvlQru8eIygESMQTWW70
aq0hBMdBlon8QgzFc3q1leQPAV5Y6YG9VAfF8V7vluF1NHefhhVjCaQy16gFjBNE
AUayti3/dgOw++QhJs29GHc+JX6XfCnmZZJHpIgsQVSVprK38JQYEKG/S80FzbIS
aSZz5C5EG4XtMi1Co90OgSfpTXf53plwtjO8XjVTpL8hZK1iUmoi33q3xQbSbOvx
a2Mn91teDab2ZuereTtua/Vn7irC0MFtKWX9+Psqpsq34MggHfHR7h97OW8qMVpo
7bGNky6rB5sSudI7fzmKqiE4dxFrUy7e9Yo9O3czeFTR5/XrO/FfJ02AigSWREZS
x6hhR2pBaYq7RoP8bj9bBC/7cFSwpag4GxyCKwn43PL0a9NyGDqr7ZXNznMbAox3
R6JKBe634+bLfgOmyktIauvaRkhgX9GblLRU8om9H5rAv5wZRbPNLdDDBWKAI2v5
HxozOupcW3wUB+OeYTf8aPQjrFw1lWdgyEE7Tk7E+M8ZJVhbV3jYjn2W0sZAvi0F
81vJyTDKgTNuFlRY6L/cjoWuC43FwCvTB6PnAldS4GzBSI06nGzhBXsspFsZHTuN
19UCzwVOqKUk2uaoU5HoQYI+VYwlQgMvKIRSg0NjFTMYa5YNrXhURvhwYwwexyQC
LFBJwQy0u7yUp8O2hjNkFY/tlcz0e43lCGcjIP7AeGRWtECp3O3/mDyc/RDIPMn7
K5MAMBt1H/yfqjZpdgz6b8WXcDIMT6cVz8mXlXBdoX7OYL9OMOirLS1iqtmWkCxS
A02bYIud7HrNxjmcr41ToVtY/iuMEHV9EmBng82/f+SWlH9ggnx1zbBr11zDNpsh
gi2MvAa2WxACtfSN6VOnyqFoE0ck5jG5An9jO3cNMHiFGGMR+ritqEnX8BFOpWYm
4chvct8/E/8y4BQ5oNYZYCUfvUgYfn1ZJYDmMozL+nD/R+BBuZxnb/uTo7hlEJAX
t5eh2BwALgOHIB1siNCGx4Ccu3UFynvduabCSGsLKJLS/cgxRvtjthkSJgG56CFo
MUFtu75SieXoyfdoRlc2wmZg5EWIjddAF5itxVccptGKQYAk3czdYShMaL42eebN
K/mnnzu5rt73Yusx2+gNiSmCKfI55gdcFWsVUBbwOgay2oZ3OQkoqCLXPOJE4W1R
mzN0uVUZ+qx/cC4ncd0OtmGfqiqcIqNP2pRPqmvXDE8R2Mhyt5hzWcccNqhsIyFu
eS42sr06IL/4+oocKYt/ExolVSnaF+yoVnvcjQkdIbGa3PqNMGPl6mVG7aCwN2pc
hvW7xMqrxm28ORs4gvLiTHZvGF1UMJYdd7+gLnYGjf2zTcus0aFa1tQSopLHfkkR
YwAYRjNboKDK54b5H5CkcQmhDS58NuIWR2mDl1SPRWycgMGlP2ZauZeuc+9U59/T
hqguBFCaozgS5NsLpP85BhvBkVOw4C9nq7lk942uW3E3/LSHU0EzyU6QwEeY5649
5kSS078dkbY47zwua1BghZyf/Zlg4X1OWtfmHJZqzBTRyWQnnbnY5sReMtvVYmfY
37v7D7qwzsomMLd9zGmoXuqkqO4aB8Rb8dgKOvV6ASRbdPwqFBjvIwXCYrtPbg9q
dyafe5XIeY68U5rSUtBSdGYRBiInfcuwm4rujON1h14CxFPu2BThJ36sde+5hEzy
WfhdyB7IcaQ6APqvSeIEUxjlaWVwN4GYJTiiEGJv/05zoOpnNPnkqHjZT2XMCgVW
plHZ9O+LvVTP0YnxCgMcmaBqAb9tdMmhIFNg7OsbXVwTHtNxukiWfsvQc1E/NkvU
xOvkS2NzgdIbtmwmFkQg+VWgAwWdcKDyAjmux+w+poFCTs7xfwotxieV/qWJLLZO
IJvgO0NqlxoiAb/CUqfGkyn2GV44FxmNG/AnBLF+8cQk8gEUC/jbmVnNiNBlQotg
s4cgXE0tDOSANRcqLRjf+4SHnXOrs9e4KO5FemAkGzMKFWFrU3Q8WJIwPRLpjWhS
HzYRdCbJaixHFFhjskY3hWGAdOf9uaDTJlpvdlJ2oinDrqJsey/6xuUUNMtCDVxZ
pM5gIhadYPZQ5v+gPgn6/hs5W6EWesfunaSNGa9rmf6fSqcqlvWecvptsEckIcWP
NjB5TAWKuIprkHm2SsGW6kC5Ik/w4B+OGSuVE2DBI0UZpGG516g2tpO8TE81yk7G
t65s4PYdATnPn1R3lvmDVYufPWhoCiUcknnQCGWw+9SymSccbD4Q+l/4Ux94ZQq0
TpQO2AzGIO+za/xStsKhZg==
`pragma protect end_protected
