`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hw6e2FkubiGub4UHyLgRFSVsvSw6Fe+doMPhBFWsYmBsFhTST677KQDwcN2KUmZi
p4xqqN0GsKpmO+MxD8h93+HgydNDzCBK6SUM6d8QVtq1wGIa8HqLTFobeCGDI5OQ
WYpbCZfgkYcSXxlJnTBMeeSGYwIKBe3hsMx3rTlD67k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35376)
+WgpYWgQtxvIhKiNLdof0HrP+f1TYRcFBiuuK6XPKaxCDEHDXs+5BO5+4wS70YNN
A9kr7a35P4YAbNxeKEkbx5fXo+sw6pTuMXVKZActJ4td/T1+qJdEYsWRAd3BZWnE
HzmkTd0awmK0d3lguWWJFZeS7xgPHI7VzFBwDQ7GWqmA/uepFdM0DOsmZBiWO/Iv
QrtQTyTvDiNYIsYS44qufzwHOYxWZsrZ5M51gqO0mQE/VOmLd9Cqaa/n/rBtbXZh
6XUYH52qCPCpEJKXGtRJfOQwxh6TMb+wzun8PYICkk6sq2dPzJ2UcurzaYIY3Y4w
acCUJPXzhPULnM9ohac6mI20FEwVPkHI1syoeiT0kbEc+8gx1L9D+tYbifCEFqNV
jLg0rrY2IEj1ZaUNuL6cTMnGmaFj7Sciwl+WpW/4CoInBD9Yf1usP/6wZSV/uvrM
k//eNtJW4ylI7ZHldIy2qi5Jyf74GucCZNALZaseydvylWlqpjkg5dmvcE6a3LLj
otMIQnwiaDZVHEB1Dpkw6HAa/aGPDccRiX95EqdkIT0LEufruFcXDYkAdrZ4Gvqp
MjbPlO234fb1t0Cl2xnGzKt8XNqqaGIs1FhfZ4pYdMeQzTyRaDVxvmvfu9oXDm/b
GWtUw+x7ck3d2E2MvI0XUTr9OOeBG3VJbHNWJVbgsM3E9ZzC/B+AR2QnQR+yevUz
gmxnGKtyTOypeS28Ldle58Tzrqv0oHkXepTPFt/V6dt7F8zg/pclfIfpLMhvOH/j
hxBjNsuxfs4PX1kbBIgJB03gKrhaarEj9NDjcqYbhV9JpRv79FPis9bMMCOWUR1l
ATnSqRwe8NUGYsSt3sVhq0NDNqlqdeBuKP3mTcwQe0F4og/yQC08M5SZJYqgdyVy
nJBuWyQr1suFb0zLdT6LykxW9IvfIDcupllqh7PULaBOcjZYpmPidbIueG+EHNUN
8krBeBGlqKxfftt7sRmniTB3H4aJd9TAdUp/cAx+a5ww4HlaAllgmYU8vjJr9ngl
afUqHzjYrMSQc7IJdOOtB6EObKE/54+OPwiJ43irjoq07pNThxzmv2rzNGPqKybp
ymS5+E6eVKosyOqfRD8HrU4gF4O41tNc2VRlgSjOB1qfvhNoGyP+zJtnswUJVERo
k1fHJLc4H3dRCOLY8XsrrpC+dazK1knKdP2CfaD5N9BvwcuB74gxqv58LO61dQQN
nOOLzkRJdf9JJ0GaN3CQgdhL5rPJaPmait3HDkseZbzZZ8hTQFovtyR3ehA9iEZA
9P27MJXEd7AdjyMSjJkf1295kCQqeE24xAgv6fLHgL7HDZHSvUnZEq+YugZZcx1N
XAA0jZ9OgUgfs85oDEoYTutvM/DaY6DzxbUgX/euOUsQKPftwJTx8Maxgd6vgnEz
vcXWDYH1gbtWvxLtFe4hkQ6zeiRbFvultJOYlYl9Q9acsef9SoDGp4R8JavKocp6
BxKwAEvqZme1CuuyrUqWd8+mPv4kvrrQRRTFn0bxceNeYuf7sjitC5T6AlNnAin/
Qg/wyXJWRXaEV2kFTdGMLLNu9KcKAs+qTTWPyVrUrQOibjSB7krtThNrLsntmPCk
wZX4taB8tW6YL56TyTQvvCPHV9dt8ToazlSXuC6uS92MU6EcFfRBcoewxejrfIGo
o/JpAMq5E9wxEF4Fx7j+2idabd1XgzpzyfQj6YHyS8OMpMnGU/rFMfKBXm5PCqFe
hR71oRSrq8LMKK1rlLEQ1MBEULOE0XL92cs8ptCRRs7G+YTViCqfVwOHpVOdZyB3
A47oiWi9QBtWCtBCzrNi8zKXjYVgyWvrvUMLCfm6wDg6y5yqv8i8qvR9zzViHWij
bQMVjlbd/yKa8XVMzNvKpMpYLRlPwOfWG4miqEWoi9lG98aUjdSc2QXlDSB0OrcW
lp61svv0zELr11lzpj5MKId1F2sfMTpQo9aCRBTJRRZoLhiLz615KaB7AZ46/WXo
QL1hJgSfLvOjLxTbR6fYMWfXhyY29vT5TA+gEq1Jfv5Aoz14KNufbgIV9YQQnl6f
kHq7Oy6RBwJ3JPcIiuB0x7rtIYMOVBc91XkBrXIxcrB0TPQq8/fTN6FLm4dLu1bm
ws94PSpl5f9dDHAkGXNvucgtf7F7qcHkKtQ9MwXxipAuIjvA/UXfcC1XfHrjh7Zs
mG+3gI/qEJ2l8bE7jFfs+WclUZMl8LntTk4dogQLXnbgrm/KmUsNjBQynmdH66QH
6fmytR0ZhPXLhi7QOLVt8BNYk4Haij0SB0TgvS2aTZCBMwZiMXO956btY6bDFbNL
+5bxE8I0kBFe/7VIWxWVABu1qYoInsBEjKWSVjGa2gQKwOBg4WnTRxve0nm9y2lO
/FthRK0ClREemrFCVTAaU1xyPEmPW+k6ylUXir32AjbKIrTo0YL/BL9I7K/eW6K2
InS53E9agLefj1ZetMyDMuceV0SkRCPvNWHiWZYmXFQfF43g1TTbaLZNa1s5yrKM
kbeSbgTgH/9u+DYm2gNWFNbzbWmMIxoRLmgvbUww5o1BvTGAJp7IV1aJXOyee7hT
bsHYX2dUJyUdGYGvi5BipShytpyCtxnaDF7lPwEpXVaZM+/HlGn/Rosv/cFgXszv
a8ZieFm75dam/CvayJ/RuxVK1BYldmnICsF3K5N9tGL8E/1Q0C1YXBJsJZEwORlV
X/7Wvl8vXf4spSixiAvZd/t4CCzufRDsVOenmRRFEZLm0X8q3pGU3TX9UWJ2PBlv
Ut1rmQlug0Rb5faPN2XN7zfjJ5hoCjvfV+NbZDnEj5jd1v5jj1mt7s6hgz+Pj8Yd
/nrR84uBpB+NPHASNdVwiZjffNtsRudBTFFKWd/myT6QVzGz7xAMxV+YQvNcpyJE
KmYoqbTG5tjOj2iR4DiDFtNYrEqne564DnsLb2WQYiFv7pb0EPZVbBMqBuSPfyo2
QO1COhc80H/eEmcOubyRBKXolPSug+EdTJR/aVF9CWCsmOkSZp35cC40C6OJaTNc
IFd9Ql+KF6m6AW9Ow6ErEbHO9uAfLp125UhHVY2itDVA/Gy9jglBpzxOCpOxQFz5
V+3cN9+Gbiw1tcmQr4TIi8Nm/aaDNuLU5iuN5CEgQlMViqO7qFtnmqSKFm4q5pdA
6VnrIKJNljblS2DDJe825MQ+ojpYmdGUFY6arC6PToP7BT8FqkFhcTmyCU9dsR8V
xHsFW9o3vfMWjicEPhjjUDmEi4J1og5eY5ot1LGO5HoKR4fW6nRPvgQAqYersGlk
T7Cu2WPWSm7OjpJzpZ0gkhz278FplHfB+AMM26zeBw7BLzBPMccKqLwJI1LYfaJ7
0G7Pc/Fzf83Y8RmMZymm4nZpnsNP389Af/aAjUBPuYY3nlLsAqXo8LzwxdRu8Sja
7MhfX/deyrThENraBs6TIH3RnnXgBWF7wozBEHw4I0gaQn2PUBt2QjWL2GFIKQjS
D6XrlbbGGkM9NNXcDSmXtSoiBhwUKPhdDpvxW1VH6WDNCBcc10eBfoPzG0CpQukK
u2UO2Id6LXrkxISwwCBJqpvfXOW72Xm+YYL6mLaBxURaMviCyLsJDX728leZU5Um
AFSZAjnEgB4OgtE90lbHhXXOXBpUbHzrc7lH7W3FxajaiKL+RbCbvSFYSvRZcjHf
EUbob7F2Y8DmMa7M3lMazhkjsP0rcEgIvdkbXUuMnu5Wg2EblGS/85hNupWXvAIy
WajgNo0QBa322hHJCVoDtLDMulKIjclIzVkW4aFQ6bFvsrFXmIz9EABbKqRdUhGI
W2W5kxqAUqQPT+FlxBw+RDyG3Jc1pFKBxj0Jh6l6SaQkumay1YTn+zRWyGtYgvTn
DkoZ4BIhwp6xzIyqQS7jLAsN00WGd1sZ8BRGoC8Vr5yeNWJNWxDntCaJM3JoyZSN
y6GVP+IcV7hpSYldnzBDErq2HLbPf6RapRJ2ji57latcH7TE37Hzpi7Qm5w6SE+8
X5O5ymNJL890BdQBsjmpxq0eUGREPwThSm7AOdNrTxqxWGX+ZqiGIlbi5PZoa5g9
ukIfwjT0mRGmG1oO1zXikuNzZT6pWJA2VME+pcOjEfW6eQEqLU3qxs21wM/mu2u5
jy0/JZ5jj8yXuvezz3kme3/odQC4pEfS4ei/Tn8HTCMiya91c2IGTxnPVLLWqBpg
2zXTx2acMY2lBS402gjjG2W5O65gvTZSTn8ZZ1YSod3ajbdyCIFP0Qimv8csyd0D
Nw1Pi1oLUDQJ3DCPaNhCewxCJcxtfkjarxGlzT5OPkdHN+hh2t9MJ3ZbiKjx5eQ8
oZbvO2DaZFLTbeV2lI9uNDoakwb4udyRsAMwTzePhDrgPTgpYIqYtZaJZkA0cpAg
5k7VzX+Be3iKdYliwC9manp3NY2z9bczrjRy1rOC+qH7NFVBSUq+X2nPK2tlXLEL
30NDbG7WCSrgr/3EBLdRQ4j+ee4vkkttREZsEmu4y4l94Nds6QM3At7CbCUqMK0Q
uGMiWIKPB84Iqta9bEejQLSFOYixrKnIOVKpGGavBIZlgKIKV/IPQK0vw9GjnvG8
VDBQukFK8hMet8l7MhshTCUjuGzxjV/6GHzKP5CS5iucL2zF/C/wdxywks1+mUeo
Nx/Z0UClcGEqj7ae3exCJ2G5hzM+w5nrs1Pest7TJ10IptsvG90GDzdQ1try+1Gx
Yg0n6n/ZimB054nB9aQchSaEWalctuIG8C7jicvj0i1fz0T10cPe20UlhrZ+dC+7
iTtsIILBkZtCZhxmCH5ABJHBB9VsDwZxU54dI7sB3fAAif8HigpkCoSJf3wvtsJK
qHagvpyhICKR1ABt2zykpKEOtsghgyhKBksjj4gP3Kf0eyo6K6SaF5ic6nQJRjV2
1CxgOSEPpX9eZ/CbHfMQV/Ju/aMqOwyZ9fvvqzzzIjBjIp5IQLax5e3XRRFDJMzS
UcpjR2LoCvRwf1axDn75lOiUakan1Wd7Fp8CdgzKnbDh+g/rjdxSN2DiEQYihT3K
06aen1eb/2X99vMHY2NkjEy67O5gJ2WAxrL+GMyrMxqsWEAbc8Om+5Tbk/QNFZKv
P3+QFFHRACrI20spU+aFPhIqUQkaWO1D9UeKdLZTI9XSp/DbE6KKR24cgI4GqiNz
/tbm2EYIdYOOFTOg+F6gsbNldW7LYU/WuclBT9DFWuQGCr6aF6KFtnHb7jQgkxWt
9gab7mTS0kpHojH+JmnYsPrFEWxylkKVatKcOpXT57bUQwvB/Q0fQopJIT1oOoSk
haddwUcq3YsAz1mmBe4v87PZIXn2SAkcOjx2TCVfekpqqYleSb5XsqA0QfrRbmP/
JkOH8bwbfITHeLZ9k9+0tUUxEBVEk121Y+UKia+/HDzZq5a7SIGD+jkBXFuvUx8h
ptUrt6EL2dT9SxS65rz8S9X1gMZFGYfmyawm6nNvquA2N8qdt5KutDGgM4CaZYbp
00bXuk3fPlhbnbJ34/XrApcj9kUT66OhPbq6hTlza2ADePggDRYpDFk3zovuwUhY
rLD0I1RlSHW8xePpNqVqdmv2WMbOF9BOhyT6Gfhes8OM5dzQVBsvxV5YbXGDIAUN
R55I5725YQl/aar3R+lvNw2xTAZEh94Q+Cm62CiVu9vn98SVuFXVasQJ+eTePdgh
yDcuFbwYKbbMibOFBhOXN3KTRHNfyWXaL7tOceu5gRdjJQbNnKUiWss3TNqfyBq8
968PkJMvNCPTSBIFIONFsYEFTRFNQoNXIZv99Mc+V7WKtc72xoss63rNuHKJ+1bi
wlt2UnewIoMOZMpRKa93+uXb8xlhnvDL1MdgcO5NmmhyRCtL/LpUL5LWSvQ6vgU7
v0u86gd5aBw5i4koN5Tag22oK1PFaH6wM4xpTut2+vJ0QiWJQufXqldy5Berb9EY
y3UbgI7EFmSp4gMQu3hS22eoON8yH+oDVo9k5kWiS6om63YXY3p2/lN/O5Rg0B+V
KaJ4yPEuw71+AMaQIXMXfVdc4KiZEu4TCP34E3vLh92AcLOfHIfC9K97vzVE0hBE
+a1ec8MBnHlo5QH3yjYRnJGNnIfRDGk1FkVxgyJwC6x6mSnTM88UcBBgG8HjEc/p
OEXuCFJfJtdg3KJzXwQ3TrviwJDlaPNKL+cE2Z7K8ZDkN2MVthU1jQva2EmQrh6Z
pAxNlNqqyWW1bhlMj1kWlRaExIU5JQyB3GqZS52KxYJRN63xDoRROQZqg7g3uYrQ
jSgik2Na7w8Mnmbfhk98WNkRhmGUbaVC2X13WRw284IMAyWPvzAGUUo8vB7DKgc1
5I44tN48igw8jMn5c7ozs8SgfTyHpd9hUpptBeYKouGqB/fXk2T0MIMQNnVFFdvb
8e6lsRA7M67rRNMpQ86pNXFIfeD+5tR2lkDmZrSKHdA5/OqolQHZnMoQRkm6Lzc/
0DYD7X4+x8IhLL8cFgzEyjGfsyewoykxf5WgF5ZYIMXqhpoX1mLM5BQE6NXjB19+
UaorDBxkEG7q/Nz/5P0XxDviAFQtoCnQDjwiRUgFUY0MjsMuwHuPvi3ewBX/Txqc
mnTX2zCwZXGy58MwyZco/A0J+3wDSusgi4qyEc8ssfPfRFxX/2En3V5bgOYePzdr
8hi0QY8zRYL2X3CjE4C0ke3cEhJNTJkh2M1K1wmYq6/Cacf+Ss/67Luvap6nAiXC
fJHpRwhPgBkM+yv13qJCW2sJebLmmN+zwJjCx+TeCUY9FiVzxY5G1lsR7DLaXGZ2
me4AIrKsqUpe3xqtm5XOCw00JPQ45cumcjqzQQldU1o5yigeJb6bi0r1enJyWRij
gPLUetOEZugo1qKBTZT/PkPnE26kCDsaVRB97KvloKuT5s8I3tU7MImYUtnFDhpu
wGbOvPiFZx/EGK/2g7JE5AK6SfVNrb759tY2kMekwd00SfVFZtq67VBEoSO2ZW+L
u5UoLgvzR62lZacHY+YrIqTRbRjSwpdx9vQVikw3Jlqlg5UjEqy/h6NBl4A/dmdC
LOAsl8RB/ABGRB08jGHR2847ZlP141lAYNC9YFLbEHK+15f4GwArdfxPDJgJSktU
NbFdHD2e7fhx8UOJtaEZlslfdOkf5O0xljDroTWzhHFd3uGIE5l148JGx7yBHvtX
E8bzxQq69cAtKKM0P7QqLHp7ZBvf4Gyh1iUbkk2GXc+MJLzuhbtrNyBEFKyvHMFI
P+aGxlubCS79snQR7edyQhHt2KG9r1dgmnlxraqosSNvpyrAboJe0lqEpaSYwCQR
oGcKcvpaZo0lJaa3FY1ygkWy+G/xYEHoigYHFVaiulWRbUBvf2x0dwe+r7SQghYT
0mCaEGT+EJ6XdVsfldjoRBOsgSvPQ/znPodiX1aCIDvSVWDfRVi0tBYptmJccVKH
4sTIR4CIGM894Y3ItVj7r854D7dW5tOeMK5MTxiRfqcRIVkO255VvVQBV0xRRLAi
7tPgvEVZhUEVQbnL0f3LwgGAeZfg1O9RQBbP8oY9+dbegevHjdtANZPiAmswA/DA
cnU1Fsijp+tmVl67S8kDzWBM3/Lr5DXxSfMv/zPgeD9RGAiNv9dHhkU7uaYHwMMu
VD0f+k9YJxBpZfQ/MTpNt1B7V3q3vr5J09db6Fq1RADrw7Ky5kAQYdFcOdZUCTbV
mpm0Kgv+qXAunCiQ8ruzNhGOJA7p8hzZouSUCxeDKUa298yJPI9gZHmJrU80/9e8
QPJmn7EH6/qyGVvOH96UQZQr7DY1+6H++Pa/j+xlCLrfdQowP1EV10OApgEy1DQE
f6R/LG8y6t/wxzyg1zdCjDDZHuU0rTFEnx+2RvH1PTaH5J0BXy5Hid8kTOOD+rqb
TxlrH2en3QiIsx6f1OafZO/tsPnkJATJN7vEj700M8S/rhy11MOGGM6kT4N91VK4
dPSfAi44058qdNid4Cb8I2zAVJnF67KvL+KVOHoZTwlSdjURNSkLEIR12/YstOrV
DlpS86XhN36cU7iowcDf/FBK3u8CBnIn65GqjGjk5p0Nqdo7fdmh6bQnW2Cx8rHb
vHTIle4ziEDO6lBNSfiWd/lLtukm3N4ZLfz1X8dkH7KuMF+DLXTY3oinfjNZ5H3S
yNNEVMoKBlDT8imoDy9VfBupqPVmGpxLLufd6J+AolCxsGY3IsIX7Enpn20pqeVp
S3vXpkgODu12PV+PRjBVKfmt+1hMsSeot4IC3oefu3tKuCzCarVcxTrM2IzlPgwt
zDG23u4UKmKWTQcRlE//vamoJXCG4znChlyghb247/A4sI7THykw8kddTqP4ha87
VGeFrHMAeomKEOSk4itPW33NDnYzBsgD0EpHgY0fA4UCdw/fkqyf6FamI7gKCgLb
m2U6KUxahMEKZyK8EQnOki9zRVzecp6Mlt5IcaLWABWf7UXuD+Aat3sYZY2m6VnJ
AVq432ZdYYBUOAsjsJaMIhx96XCYMUtxvGXUy4MtvePYSPsQw/+4cSBUcJhPHDnl
L0ukiSxzFLMZf0dEi1DszNU9j3Dff/LfKBRZFzeZ9sMJl5GoXy7FmcEFqboleOGD
ONdwCmMZXAA5MQJ6gaV+XxOAJGHcmyP/i7Rh6MwlIUVb4a6al0QgL4P/+u5/PYTu
dFnQ+hsn2GnD5GkITH8QKpNpnFgjl/Z6pO7+h3nMABDDzeAEuYW80cCn8tKQcwL1
eS8MGo5/Vyoz+exVPW0flthOYCoD0zY1fFo/zbAaf3Hf4tMR6srJquDFENpFlsO9
hwab6kiLCf0smV0uESZhVSMmYyTgD29yVhw7IkcSubBSMaM59WtpFJ03GQ9QUNDc
vMLYHprYGl1u+lC1f9h+g7K60tnzv0Y1YNBJaGwNud7AXBbJJjTFxWhpJAogtMZE
eZ+ch/NQsPHMwDn4y27+ii2hpiTR/+Ffh3R3ghBnptffprmkP+zUylpWfCWYFhw6
fncKzwvZ8S0MFGo5oEIXxLVvvp475FeXGtwqcxu9ysj6c7x5zrVeNSVqMYt+GwWP
rm0zHHf+8T5FO24leEORwZDTrgs92lnHwN0mx8YW3hMaEBKRUzWXf4OHyL4n6wvq
lfgADhJouinf0cLhxDVZkkMyfJL+6m29aGpWP8TwpPF6SkkjRsOhMHgWZWY0zE9I
S+oRLpCBObkdfgV0AFlBoAtK160JlB6uo9jL03PHuYnoIn3PgyKg5meHTY3HaS8M
NthvuBoaJgYe1vDmUMpzeo5iHxVxPybeajuiPnkpKmoU6DkTUFlFoDXRJ9sGVWUy
oUjMSNMXW14qEaorATRaCOgah6gom6Z6VUVfC0DIEEMsWUsgoWRXTMRKeSoKmW1S
KGBjFA2tvDoPPn2UUxaA9Ga7s0uUWvJqljkX9hU+UNdSMjQDhMzY3J5Uu8a8pIiW
76MQR1wXNkmB2PwIyG/tfDwfLEswErkMbrsPgobjSCj+leteIjc++8Nh2UoS49yk
WMnd+AG8QFMyagLz5VNjKypOMVSu2Xm0aNn5CwHH75J5pvTy9w52ezlpBv3gK+l9
yYaH3inHupSyDzN6V7KB4Xgn6y/PGBeE793hCLIlkFjqGTLn8LtNjhg3tNYG06I7
gsfKLg2MODgPbrAHBQZhdwCTThD7DWHe9RSWrVDicPna1qoXxysKgUZumvfSnS6V
guh6yIni12VXwWMJPmw0dFpJzGLzyp3J5+uBRRAkbc6/KgNtlklE7xs9S/KqLqrQ
lmyO0Xm2mN2gOv+YsuPmj1qCzFodcYPxjVO9r08Q+csbw5FWpd09o7hBBn/6RpmL
dG38JbW3nK0+zIDeFytCnbi1oYc4y8aWt5f8J8h4ermq/sGLmZ644BDAhMujuU9r
6I9BsFFzW14fU/6gaogq0ok3NCx/saCJ5C62s/SLxOl5+rkB9BWiROLNI9UVWiRl
80Rne0M1wNaXMCrHHDgHanQmdpCoW35YqWKkZJQSg9SZNIpC+GJauyxBqN+HYbo1
uWttIGpj8zUQT9ejJqhQl9CkfpQQNpVX0NBBYEI0yT7mwOt8ru8LoUbCKXQQw7BX
cXE7jb45GoAVcMD+o/PW41vX6cOApS9cYmOIKf12qa/yQGfPVig6pMJqI3Hd59gU
wC24FHhdsZNZcddd4i3dFC7jUJUDMaQ7OLzS7UNN8oSw+g++KagPm+Aj/Wdb+8/A
I49GV3QYKHlUqVMHH0QVdwDvwHDk9xInE3B22Joe69KisD+8Xs9hPYBpapx1rc0L
gKrdT9ecD3s6B0iL8zNnlryzKmZF0d5llpyEksiehPco6sNDPdETuIco0igxWOHh
RJbfx46phJTVsYoVLk6AxfG0bLBhAcsr2vRzNIIU7rjIijTjQaYxfa1jRiNKKvG3
sD7HCIfD/7fCVdcWjGlqvHBJBi8kCpDRyV9vVLYde8VsFnihjZxleE4s+VPiYsUe
8JZbf+l5N6kxnTFREDum4EYOy49uw6ynTJrg/NTVBy5z4SNG6RyG+8JXdK7+UhrE
kN0IPuGWBzZbaJXyHGt7CxfYAKQZFxO0+bLwKyhuXNVu3kZxpkK7ItDnUJOfpxL8
p8ZG6V7tlk1Boy0fmMzBkl3cCrOXvi0IctEtqBEXmNr9tJ52wLqcb/K1X/QfpvmO
Lv7/Cma1k7X/G4R5q1YPBtX9Hk2GNVA3FIo2XlU/ZksgUNoax+lhzvdTxIxDoete
LCKIgfWYUwBLKAXVMS0mvEQaE5y/M5SpIvp6Vq3GmGeWK8bu4Uo8ribLpZpFdegd
RMkYZ63PtcbURiwsrqG/tsTPznmu7PoyD24FpbQFrvld+L5OPqsN1EyBnEPDPb2G
xmqTCS0BybjwZDRhwDtwnFvj3g1yMQjKwPlrnqJp4pfuDGnzMrjdKWHOSTE3Q/DD
EYWDZSM72gbgKlr+DIhO+cZh4czKcyeOOV++B2VoGcI144e7kjPsI8XFft0R5Q6k
dzw1SxlQeLwiPBHvFgeaxM9X5zDI9jN27KqCTZ3RmK1khl4pm92rgBhwxPnIk2uU
soSMjRZH4VPLfTQAvMqctg8n/iwK4N5x/rH1mry0inaZIbSZDZ0KXtk9/4IXHDdT
w5oy6bnETqsKKtJLkcCrs1K/WK6PjPf5Npz6iBtx0ScieyWa7pX7Z3wvrnzDPsPV
3EzGmWE/uT6Ts7OEIMP3jSj3YbjwLgk0PFOfMDTNZ309a4JhtHII5FVUl9sBjVv/
hE4CB5CejHFVCdk522lnc1RZz2j3wDw886an8MXxy5J2iJ67faRFcxmeEIt+dUfE
cKrfNniFEylaikBUnzpLNBoBAOZWTL/bO/2pqAumIauH3Th01taTTfK4cjlqx3qb
TJ4a+BNl3Sxe5Eq6g95RT9uWrVJBdFJDeuZY7jYsyySUm1C+BBHaKg1Y20xZ0MRc
n/UjMOt8BGqrKS8h8HCFspdBcn6d/t8R20Rh0rmS5Gcd4Epi2pJ1JJ3vPOUq8F+e
1t7qW0VfHQDUNFho5tzjO+dpK/zeR085d8mCpkChY9SynQB43slDyBYDe2NPi6iT
2ktB7XSSYxtwWu12Hc8r4yTO3O1sZkZnVo3TtF8sf4/nnnrG4j/xIzDRKrxpJyri
9HCERA9F2zwV3zdrwtQwVS5JWnuOsFc6t4BWmbTlvPVZOs68h5BCk/xqvvjO1lWI
eTO5OVGT5if0kg+KDqpYtOsEiv7Fixr6e6ZbafUcso1Ri0Xe6NGZ509MVo+tNCTq
vqt+J0oeRj0yy5Y1AyFZTln7kG2ceFyYUx7ryy1hSvYPwPbXSicYnxs/aOBAhGMe
1jl1MjmmCt8FCG/4yulZsSM2SGu5L55JKnu7mmbmraMkQqY41v8qGV/4czuTN3tC
kRmXPEXBRcYwWeFSgaGeiRPcLsmYwOdvnTlg/QdumkIW8WYSwM2CXOKzu1leVT/d
m+IlUsocPLwwXz5cXUCBqS9GzfTxtIfKUUGQ48Myu+I8b8aLCiMhun6Xs/s+b2p1
RLl+9Q05QPDGjdo0sFfMBbGDrl9o4X+0A/uEKEyG72K+xo+oN2xsqyd0p+cAuRyk
90inSGL72kwFj6fWsjrG+VcMCaTVhjfJEiR886/yRDNVFcilhT+FA71PRvhem9o3
guFRDVIgZ+bUwtQYXXeDo93LLNEZBvifGl6zRgOEY3rMHWmP8SpQTyQ0HP2yrZSV
CGPpB/T27akIPmgJpnyGbGmHgniI+viSVwZ9ypcm+ricHHs/YaI489IY7OAEGCnE
M9UVaabRBFyo0VCqhEznjz8jao+Udj+p/aQDL2UoHbt8IYww17bIBkVbMFenh5h9
aFzgYcdbMsCCFJmg+Kjmb4+2X2qXSaXWOFRSlAgD5BfuXQ/IVjoCJMV+Dm89gkO+
rJ8f3UFpT2a71zXSRwOJl4lhih816FEaAoZ583dbhOTT5qIpUY/RaIjhMpnd18sc
1OJ/hOT8zta45q4e2dAMcfB3msToKfpM7k7SEeTb8RAKvy7Zt6p5AtOHvzueDTf1
xEBWh/pkdpUAr4iE2vkwo8cQxJYujxYszRAREq4FzaBW+bRUufHRwWf8eGXZ0IQ6
f1AAAhBAdHN72DR1W91jzzyVlWUa7acPxuu4AYX15BX0Vet0ODvIpTMDJSvVTnFe
ZX1P4yJNtBUZ67zy3vRC2MpY+OrE7rJJtTBgpD+r0MuBouU0bKr/XhQ8+P0f7Wqf
vNAR9mwOCReaoow3RvJSrCEYqYISHF+H1OctdETCq64BT2Soga+iwFVBYe2xTZ67
YPPdlGZjH7BQF8fEu0UeO3AaT3C7Sl2sqbHyroB+V7HjKacgZQZV2RxelCz6ybQX
0yKs9jBLOSl8Bg+MZdxhzubbWdmfKcSMGNWI3U4vlUYJ3h1kaFOMHMkoO49EVh3p
IZWexRKop/vDeey/JK+i1B0uvQK443UuxsC4ku1HnHpdl9v087ivzYKRGQ1DPYsz
DkiieEtKvr/Bd11AzsPWRB0xeY/kY2MQvXCyM+a1m+rKN/BIglJ+hj1W9SsrwT8c
8i55reFdsNrj/U/ku/tvxdXLjz3g3JNca8VK0/LJOM1NvVPWnaJ9nl/9zv4EfZxn
sGnz4DNbEkhW67Wb1yv354kvxTCSL/a/Zk3RMRa/kK4yPpOVp5GgYyetiVmehPxt
cmAkZtkYXJqS2Cjpx1NARqydFLTb5yQ2GezkBpvGc7awUwYDToJSzUePOd0uHgLF
Y+mRbzwXJttpjMMGw6FK8NC+apYS7ywlTTIKpy9n1DayQvR5LgnxT1vy5hoDIMTJ
K7FtwRXk4fiGPYp7NdMZZgcgGg6tyJ8HDBQZ96HMf3cRpD6KFvpeBiCUxGzMp9UL
8DcA7yofjd8gHGCfSg5un1ll9Lw2GzUpFlZwnnc1ylvcrH0jXX8w+THl4XXxJ/rt
XGQLr+dFrXvBm4uNqtnRfVMUSWmHvG08Tsu4WMbVSWFK48N6rM6+C1Za9KwVf6gQ
eF+js2G52bCAnxF/uhwtovPUxLjrbEVWdlhsUkNuwhBni2vRapSj/bXknE4f3mim
mecOc4VQ2a894ibo0XjACeClHdor8cSrJZCXTVhMMHmBenk3S5SWda73gPDsdxP6
ZbdsIjEorcCk/F78jz5dZkKD1859R3jOhzccauUXwXFe29IksDpKuIktWi0sYneT
GHZAk1RSdRygqQn8Ixb32E03ApTKlCVy6C1cC7INWPg4a9vLDvP/BR5U8VXvy7fJ
DMqOVsJ0I01yUMLlVqfpRd2Y+euKxLh2Cjbzioes/k4XR33lxJ/9hQT2v7LMF5JC
6Nj0hldEbjMnwVjrLsRkWEo8lcBtnAv1Nmy1GuJHsjHKsIxsnibx7P/zvMZHKJeE
0OAcCuB+4EW1iPKz9MpbF+j35jKA2kI+mLNuOTPvSHVdfQt8KbS7LxeqCL7wjUZU
By8iyF4KgeVFXq3LuZNo5JgcCCbuiIvCfFjkD/Bp9uX9JxoGPBiS+rHk7+7qC/eI
zwrUKZDakFycZLB3wvozSkKMYA8EANjUkD58FA8SWlJE4U5S17+x3UJqvokxp9ta
iyYmbBUqYCVG7Mv1xaWhz+xnxNLqqqxHO2ZowhKo775e07dTQtTAT14dv29ulOKh
sF3Mv7KpD4yr4BR5U14SqXFfWMYG8CYPhRBJPvXdv28rFearTKTnlBOxGjA+6D8G
STG4jIg7Gc5t0DVjUgL/Wdhj9PoVIIGm8K27AkWAOptd4xzsj3mX5dnvxLYwCOQk
ui7PBiNmvarrCxNJ4/STIP95Y16MGfmvdgzHRcG2XjbTedBPsdWoui/nY3huyl7W
GPJrlo9dkbVmr5ce3eiba2R9sO4CSKJuXFxAaIKYujhJ+r+4X49Zw8lMvsbSAXVx
XDsa0JOkCkYVXQdkYZvKXljHvZWBDG5HE+1q25VI88qlq4S6iEhwfius4K1Gh5n2
py1CfmrmnIHd8I3KXrInURBezB+8M0PS0cjBsuSvQO8mTsfsz+vk15TBpndQU1xU
J6xle8dWwxmfGwTeNH7n1P4NuSa81lKGSAfnSV0KXA07Ms5ifFUQPfiyt5y7yhZ0
1eMCaZlmk8ywpP6SH/ZgQquS3tg+h0JrHrXAaiUCBsaOTrY4iMSQlvVP6IWpzSg1
0Ipks5jpuuLlMuujAjlTDz20cM+YItM2bq12F9k7MGmkGjZ/U0ik9eLvA/WBZLa5
SrxdWYVGgjuZQcixkByZwsW9dXzNO9FOz9ILAewE7mOldaQewRdBikzjwj00UigH
qq2olHYNkqrBnlvC84Oy8eqsVE/BwmeAImO39n/h4LA0wZMWdU9tW9dT30TJ1xcV
7NdjQySfi6nKtqAW5uRNCM8JK88jG5evXVjdGlqikLCdD/Vz5x+a1AxUhHnJ1EVI
qyvm5CfNLQVz0JhC4dPL95eSczsay0iK+Eynei918dD6Yb/IBvk8EcrIDVZdzAah
rn22lkNMrbzaL8c23yKQllEUZ/cOzNh4OM+o+LRgUUz1YT/ii4qSsT982wTZ3T8D
8Clcl9vbkZ323cz65qHek9KYB4W626t/nXKSIP8dWgNCGcDEtgFPCWkAhD/yx9b/
TcN8Fh6kJGpY7rV5eM3AXWa8vSaSimC2evA9WylYx1f3E1NWaKbWfQTAIAvT49tk
F09l+ha9U7cepJlHYH2T3NqWEiffzFAeP+pDO9ZalTX4B0f35rivMtsSTGkaTBCx
MY2NW4DXDhYEKZhLMTcjiL26kv0UraVsomfOWO0LpKSsIalXrcTw1PSgiQU8hH8O
vfdYjJKUTevY85+U5W4aFv5wJDTfodzuSjpJJnnIzBdzwwPBpTaOgPwkyAz0rlRx
lPIGf47xqLXI6wK6IiP5w77ORXE1SaFpB8jpPWExKBVtPsWANke9uzhqpKPVHP3c
LaWoNHH6xlt3K3HUKkv1NyIrXk50wm1E7vq367Gnz97sQDEadErbCd0Ec0gOTiqA
f2qJoAVnB2ElptDEpGMFVQBmFt9b4exbpjpwrxyXXcDZ5eE8QJlxFkmSZcNLteXv
pX5ttA0lcoTVTfa1wXMV6UroQQMmWE6yvDHqYZuzUC5dgXW1G7SIr0YHCoJFy+l+
Uqr+UYZZ4DJuxmEckc1kRRcRcNXqZHhkXv+rd+yKMysQvuhwzXAovEiEk78HJc/I
KdQ4saWRsEMnQZYrLphQbYgnrhovxWUWNfjZ+AFVmXTkYLKBuVw2HyFn/80zT6C2
HFPftLo6/YTRyjxJ1VMqPDy0ZAtuO2d0W2hbHA5td/LWFWUY4XuR85a8FypDsnvo
OuWyIYJolM4zFuNzMzbAlxbOFDXcgSF8JOc6H2z4FxzRNTNDkxm+ivy6MRsDCkJC
vLYVSX6njUyfuTvC+GvBBgLWVwAgT4eAfVpSGK53ypBOBsn/2/BYfVcLOkTRXf4y
g4NAhfdbSN2jTXl/jeV8igTqCuM11liqpCMLS11x5fJ3PTfCUtCi+UCW2zIma+L6
S6lcfLN6g4zYnOh+GK5Ffrm7EhM0z9GG0JcI6HsGIL5vwiIAhReOk4+DG5eX7coc
GMteA1tVxLhioyEPjAA1Vg6Y+wf0DmaggpiMpKRK/IKjnsN7KhEHDruH0GqnvfaP
RiGbGeeg+9kzCDpD71KhHQi+enN+duHbeGKcxByqJkl5pqeicpeeF9qaMTD9kO12
L4hBQEa+OvOEKwSjTlI3y/uTf3NvfU2+GvdmdBtUC3+Pepza41PqA4DMLs3i1hyZ
WLA0URlyNji4BJPhLGEneoBBJjE1VMK400gngaoI8Xj+20Dflg89bM6rrfF1VfbH
mvgRyyF7z5c0ntClCBbqYXiFzayVgMXHmyO/HliHcbB7IyqPqYeHfxFSOn7hz7rN
cW4KfRub59aywVGRNsX8olO6lFZnEg4GvD7SF7DVahvO7YPJ0kKH/OhGW8FAv5qE
ENsBq5Y072C0vdRyHxaAZkf3awzY3pvvt8RRBEhtc2vUd48N/x5piwNV42l/Izsl
c2XIhJuF4vBIn+Ub0VF0UtyHJmOJfYumTgpfm6NoEit11yKmrUJSG+calBJhK0+A
RHQVOut44MqEb8wW1cIWfErFsewJXu2PaRrX2BfsbMEF34nc9jjyg9b7t0lXrErL
8bRDgfG6FE/9bKwsRRSlw7Gb5pESWQErBINcKVmFoWVInQQvGCaQAESqA+X4SNJ+
F0XbBBSunHhIb/8UQHXn0jDKEKYddrgi5xO9BsuGOz7nobSiKM/jtDyfwgcb1mq7
5T0FPBSlJw7+h0X8pOYuAzWUKMabmEPxWCfaYgl93xNtc1zZaFD3zTz5TF0H1mPx
gjwz/pNvSUukhm2rm7W5kCUCLWbYHqyGAG/PRkCr55IOyhRWBG3Laq41OuLDDBmf
2FCavr3L5grEsAH2qw7Nr9wGN5LE5U1YSmZHF9BOgSOIR6XS3TQas8ajNRDdLjg1
FuOSEaBB2CnP9xa5pawk6BGyGcZAHVrenvXFNWP9SO9kMex8aEogSYnhpLTozShL
dip/L1j+U4bW46abJLTXhT8kOH4A+6raqCkBtx3UChbTPMbAiE5OZKFl8DlFot0D
hogTM38Qn7w6J/nDml1yzV/v6oDJkw+/guXpmL/q/tVeZHt0jBcPp7nyuAAFEDUo
LpFtcIGbqc7WAgBB8+gyL9RT22tr/2z0bC4SULUzTKeWJizvwoiQcI8fon35cGRh
ALxh6tqKkmCxkcBwvcH5tR+/UsMNN+a3OeaSKrQt9rQvZMlHRmR9BSPzv8ImoQqS
3eIKzBTve/o9+PKN/hF8JGJIhSII7xrow4pFae4iG4i4jlwh4k59z5JXMiKGI0Ao
nD2Opw1P0kPFoCAmVkFsrLtFbyyzl6OFyDGfUg4ady1D3d7/IdwAHYa8RPwhX4JM
nsEx0BTDOb3D++tmKYJd3eSct5yglH8TZd4uj/lfULkGE/PMnO9IuDIGqIxwwMiF
Or0aTtLt0echTKHq+3skbE86BZ2a/CnfApY7EUnqKAHfYhZ5GlJWccn02idzYfkk
dJ4D2FwzbJwz9ykdC/wu+0A/ibGKs4RsZcM/NpqNSymrMNEVd0tne4h9ugPcT28g
LgktCJDbGYSmsJBI34FeDWavFi7kqlT31srMOSLRU7/oJDNKWxO7L6TDYUeRtuoV
+bW7N0LKR1DAxwJjXmvflclRTeCLcnRGVHHjVYuekmrtcfdYibnjEQpoqJBUk0L2
EuUzOaF5QCoyuZaZXpRBXIqDox+d/9WWWx8fKLO7oAO6S1cbrD0UuCQcShNuTGBB
EqsykhqIe15id5a1nS3IANBJaXyJqMgBQioJ49Ts+tAWPyXceRC0a99T7yYwvoM2
c1gj5ZIwwJaKdUZWeNQUHhYq+sPLfKdTcJkc3XbZHxa2q975adYyW6rh+owd0Wdm
6vHNBKDkEtd68vfeNG4j0h/l9sx/hWjHXmpeMhKCs5GnI+3QyXQ9HlA3y+qPPNDp
lLI6a1sKcWPwSSL3PzS9QqqQD8MbmzDlbfnaKQ/w+8R+l/+rZbJp3BVn7fQUvQVb
+7o2GNYrlZ+19QSnATB4iP1+srpGGqF+CXaEKz2V5fDg8GucbrjQ5wOAuTnVrx+O
TnMxHcbvwhp4CLuzLAnyrJNTMa7E6eRqr+p9bHEy1zF2Yp7635AYP7OspI/71H2T
q5SssIPyszXX1WiSU2/PlrCEzZ0qDXKO3O1lH/Wq5Omwe4h69MAEzqRBYA2c7xfs
dKI5tJ3a8wfxsca0vXiumw5BsHRRcIZ5EhtHGwIYFDii14vzYfq+HBFTd9YGbgRg
je3EcmQzGVKSLR+cXoQhHMIyGuKr098nCbzAL5IvfsKcpzpxZkjE8RWOrn9Sl3H7
CW8MKBW4wWDMswwcOsklrn/zoUCVUK/w65u2fPn5jTLpZgdiMyZLF2XtMjYNh8g4
3LzGy/XdMkA8Sk+x3bWAvM8EHOO7U1UWj0bja6e6uqBuQ3m1r5h15dzZHzMl1quq
phqgrYcoSD7xD73yF/yiz40SAG2kPuFYj+lzigrp8qpgdS0/4N8knKV3LKEdxn2q
F00O4uaSsrfnpJ754+o4oEIwvAXqYjaykykl16TDCng18M6eFiRhKfK3f7LCCa4V
JzG+/rHYK8cxmC6DzpJMu9nDHae4J230q5gU31Ae70Z4hFE++5AieCRm10XHAzfI
4TxcBI1NJDSL91G5/LYxjvuavqz6DSnSxAe+9jk6CUzOhB0huJvGi/RL7Wj0y5lB
TgKZagdQt5rHqyYhtB0SoZIz6yhmctfMsymasGM8DVEFvjFKgdyXeFTVyur2cR0F
pIwBS+hyAStpbFDQeypoIjBf9hnTFTxf5ZQZbO5ycat8xe0e143+j+4PyQ08UvJB
inOFGrD6BUFyVeRe4u2tvTrDXLd56j+M1S83wVd81lBYAW/MBBS/zD8Xdu4my7ND
OjX8pWPR4JQGgukEuATy6yH0CbX3I5hfJr1VtxF3dQcNGv0s52Y4nWSFmrbh6zgS
1QDVQKZiNSJ5uXX3bR9l1ys1LF8MGwSXJWzdjZtnL3DYenO7dCuMeKq+RdZ9em0c
75H56XFcghEECBdrFwrYX8pOQgx5vurkzQewtbQW09lMeZdpEzb1qs8X2rWKkcvv
IbjFeaXLHhUde87aKzyRovjMLLeUa+4okIogMbue1TAXBfyUVxK/hrggzeBmLYrN
/cwvfN7alofbvO68FRxolyNe9Y2Wmve1TEtoaS1WdFy64vmn09d+cts/zX20pQVV
6cCm8BqBiDsqA1/lgczQ7ZBiyowraXxsjeumG4xitQ94GpTO1X1sWB1oApyqrP8B
kFThs382mcL+AfQOkyCliSVgg2r+IK0O5BHmwmcrLHtYi6Qe/P3lbwfLCqxeE5K7
yUJySXg47MAzxYds6bwyrHZ4th8osM22glMS2THA44E5ieoyhl0i9x53yVhS0KpI
HS1RDVUQIO+pWpbGCVB+rYpsAltHgkBit/TmDw5bFwuKaa6TxGT3BXmfOkafXhFb
gOOTB89IOR6bs9jYhGs8AJKw7MGNSxOKtcn9rGFBMLjQ1etW1xK/fQhWV/y2770S
hgqZdQuXo5BHDgWGYtHqkk2mr0Z4/wH6DBKVF0CzBcGpAi3ySkBc0JSWLxn7YR5u
PjKziXUPEMvgwj/CYRxT5k0rWtyc00UOdRIV0J4IrRsLueNzB6ysgss9OdKIoDtf
QFv8VshF78lDkFFYLLSi9hEXudD27ShsBwcGyKNCSDHvThVcVgqP1C0/cfHOYEYg
EABlexh7eYHGSsIO/JFHod4etgzMkB1xLSTaCUjzHKRscl45FAmuWbjxwp6q9Lrj
ZBL3+4S2gOPUVxkyREgDDpnKIYP1km4mGOvz28cImuf0GuaPqEtp5lUJR6Q4ooTx
DSzARNaBh4F8+Ybg8tbpAxwUm0P+td6/IC/iG1OzRvpEUHLtwdTTyk4MccGbn4PD
WthhmMoDXVWx2bp8KLAIshMtMlbRIzEufe267P0uiKS+tFYGHPBtnrwq6sJevr55
P2SYv3qXyA+i0Qr/h/MBLqh1jgoadzS3UG84MUlKxdpPU9TGl22oNEzWS6EEtOxy
VUaTXIs8p9MUHt4rWfGnCFn+4ZSxCr265LJQEMM/kTaFPD+jfOFCLqaC/F4KejgL
Szt3V3SrDIfHs8Gz0veaND3+IHzVIP9x+ttGXfXhy4JMiRZEIzKGC/0VFbwe5F06
zPng5AsheMW0FftM4pDVkEVqSxJ/JIae9iAzop8p++YsqCMni57UxHZF8MoT0E8T
viw5H8bgcSa5et3m+ArpVynwhBBrLol8+rVdjpOReIIH0X23chX62XG6tJr3FioT
14qmCdnUfGdi98jmkVmIFfakFGsDbrRfpgZevPtBBwgA9ZEdm1DEn8VGhMT9boty
osjH3rtxDS4pEvkcdLJScALLMuSOgTUZHR5vNfAZhaNOlZQCfS859Ibf/xsLD1wG
fVomIsIZsIub8Wr61EXiT+NA2BIa7g+NCTmFwaAEAn0WmzO7Wx1b4tx4Sq6xNcgp
o+xWVAAtZqu0y8PO5r8G6QYZnpfeEKmanErvHzQ3f4u9vC47CH7hXNW+866S3k8Q
WqPBUdyUACg/iUI4RH/ONvZHLO3NE+4VS8qclYSNY41jaXkJZodsk1hFBiX8zWtU
Na6p6CbZKTvRBuagD3Uva7+VN9TKo61Txb9cmwjrsQ6/tnIG3qwbd1dQbd0jaXLo
SI4BjFovPjN9xv5u7oHwIExUHpzZMuoHe8KJnyeZc+sKstEMInbJRjuL2no7MzvW
+1yzWEu5okgTG54+WtsrEdQ6NLVvt/4YXW9HiRQv4H2+MYJ0g5orzRmHLzJXbzN9
w4pZFxT3jyAftXlaYx0ab8we+42ZZR49Ps/R11MORYOO5S1iiPcCtX010TlSw/6c
TtPwdtw1o3ey+TX+AOHmBwODd9Y8ELiwjU1KRjAmi8kKtNB6F7Ug/fcR4/HgwJka
VSp8gsZAelmAXQ29fIjRbF0XghGlGhuQoyQnLT2yv6Sxjs9r7MeCa9icJSmmHyq2
j6JVtG37Y1bnRTmRT83Ul40Y0s4ZSF93IQMhB8TOelM8gK1LIB9FLi+YXijSIbrM
o4psJkzOaqb5OGjhk9XfvZaOygZRH3FxzkUQvJqGe62MsN0p/Mr0aCyN2LO54Ou9
mLiFnakZPwMxYagPZPazDhEDesYcsSUBpfCM7gqdOQiQFzNLR+HH8KHgzjWApZTy
LUwWd/c7too/TC4Ouhbc/H5C4ftUJh6HzBchIEhIL+mep+fU3hnOV6GoriHda66F
GJ/u6D4BIWBIb8QXOIfYyorMhHDh1YCFgEhZmkQC9QSzFGRGrRHGMDbQXesHokou
NJTPdqONqOljdBZJ64ZGEdZCoDaBckS/Kmhs5FlOabqTV2uOa6oeSh48atP+FatH
qhWvz0DHkOQUAbBt6bhUItdk27X3whSYVqOX7e0A8EaLPwj0b8q2Bpi9Q9Y9Nf98
IHS0VgQ3A309tKQ2sU/LpZcKmD72Vy+BELly89fnrG7iEDztY9E4RDPrVbH3OK5o
0LmZBP8Wp4deG6TCbwvJd+2hPdufCsQj3QUmT+3MJpp7b07L4z+m18t1lohr+rxk
muNIx5ur2ydnCuNz1yoUJdrU/iD78YsfB0jYxP73PVciaDBFcXawcs9z5A/w4Phk
YOd4lY7Jp+mfBTY8ep+PAFbee/LlKiO2wx8eu1+Z7YvfUOsvZWahrbaVC+uMRx+w
Jkzv7RK114W2WWUSlbgRG9dDzE0qvp9UaijXMfXGHLF8NZPQxoKU0FX/5DUlrMGB
daubSoSZ2K9/diVyMBy1p93PEfNtWzgIx8AEzjc2KFHGS9gzdd8qYLMwit/MaQKC
7kkfmYHGZthWEnhjy0oaIcC8kRBDuNwQFAPhOqJFwxaFNxIp6FSVkOyi2Njm+156
HLPPaU6dzHcEjYorEXgyDWdd1ntZpElnj36yKhAUY/uJC9rpeNso74A6yknWicyn
p3UxftamhzTBOD+sQBl+2npvkvMcsp29HidKXh7n2jrjdXVWwIw+KEkercnlZ9H3
SNMqRkQoXxDhfi/ePaQJ3X855HNMnF+Viqk81BmDgnfKiHtji8u8WJ9mBnM/NPWg
oM3zd+7bOjrh4xUfZdb9yGibb3bqObTeJ4TnU4SazuJaAZJoVuNMA6vb128iRZSG
ynMthqpODfKOBf/IxAl4WZMsr/ZiWKRXsezu2/MJw+ex6CtcnxYR5pVzIU/IKnbi
1ghBaqX3WpsJz3m+E3RnkwEgqJyGkmhoiU8qFvKCnb1vWOD9CbyjH7xe5HueSWqm
mQjJiQzqPzXB4u5YylqGNgTXJczDROgYiNelTBKlB6KrTblJrP9Th3pZGfKZAfGv
iw1Sm3A0XLMLrxAgH2Q7obUWqImTlXfZVAA0mdwIy27iv7EDTj0Bo4Ysi9CZOvWn
diKgQF1A3TKDSW2nRSKfZE0keHj8hDgd/U47f6C/BBOxYaxtf6uUN4thN5Zsvjj0
qidV5uO+l12tgHmgfaxtuDMIGkXrC5tyqI2Vf1cx5bwiR/Q0/TY6k1vjI/0jVzXA
F6YiXeNcY4yT6esR9ebzKiIFm5uQc1d/vm3A5rsSCs4cK67+eF8NNaCB79rTbDQ9
X7x6uJGv3Wv0l7EcK2gv7cwuQu8YWHZMt3lYOv3t+BjsnIetvqatr/qefSZ54EUM
eidQavSdLiFAPUKhYPFPnhPVAT2FF0pVsjr4mqICnDtbztKPfjX/pSiE3oDlNnXv
r0c7gPIR0suxBQFVbHYIxZolbRn6uxVjqIsU+j+gYbxdQ6g4I0fwaHIyzvG7ZUzJ
SG3IsU9lU4s9JMSkwuV7dP3gTVkW2DglJk0fqhJonru72Q+6LiUOoMZV56f21BEC
FRzkSrgh/3Aj5MUt7/2SvrmaH18/Obxd0p1c1oPWqqVFtPbMMQaJLxujho7kDWpx
4OcsDM9fGja/LW7rnOL/t5j3LbH4ieIH7CxGwC7KHMehJlklDD/aN8sXTPeOiilr
hyPPzzYV2Y/6WOURdE0DKIX3HK2wecSXu28c7tRhwqiIu0lStE+wh4PLipHR2uGL
JkHOaKYSQphKuLa1CaMDazIRTJIZg3nKJ+Qf9JrLkRRBDqeOF8VLNzeoSNFKjRsp
orklTQ3xz0TRkB6yZoz29JL9KYaIWjPYy3n2vgaVKROZWkmwq1k0z/sQUF7G1K75
cquFBdGW/eqxlOgTJwDZAWmuNmrcwdmTqJ7xbMzU9bIuoU2xmkiiGCCiDelAVJ9h
wZC6pJQJ25IJmuTkQSA5EJirD1ghdZXLEj/eqReqPALofY/TAocNFmURMR7Emm0X
0SBuxxy58Bo5ZYB7rdZNaSJWtvKY1FgtQSJ9OzQYO04+mbbY9ohUGWoEXxMw8pYb
98hvFOqH9OgvUrDERt4SoakIIqEnTI0UIbKaPOJdfoBx1Ao/KqTfW9Q5qpRZcG+S
ty9c2064+RgYm/1hn490pMCSP792XWV5R8ktDY9H9PIbYVIHUdEODk0lS/rL1acC
bIONZY96LQhJqLMjdAMuZLDZSXi5oEreAMM5MnEpINS7Vw+eeCAn+f0ZH5Tn+7nW
EqeDo1JuxBS5lcUf/8YVivsl2V36oA7qppIsbSbcT3Btv8tJxQRhgjBPY1jRJt95
BFyYkMouw+O/Twmq19zh6tEidPTLY9RT0wzqf6RRW5dattqtUUmk/BJlssh3OjfN
ox4dq33IVzqXJDUEmc6u7UrgADvF4zMWi62UrkLJmPl2XbYvF0/CAK2SVWSkgK3v
PGHZAtDXfdbzzJbVM3m1BHWX7HgtTS3zL07pD7pFL6N4s9yN1Qztd7TEQxkz5BjT
kFowVxNxcAnKTEZ82tV9TW6JY81eHbEzSs4vqhbTej8KrsJYAtukpEHXDT6S8Hxk
S7aeUsEKRc9gK56LfnfqyrJTUIrM2YoTrigpu4yqn/Y5+lntTdp5Q3GYe7VHXrxA
Nob3nA5Ag7q0kLi+Dy/oHr/bypI8cb6HXnp0w+nSdVNi6XqyyWDACsgCOXuA99cV
AdMVUbDk4zzpJoFzGv6HfWwW5HCkQdizb8Y0/h0cccSSwcMenL184dQFns5f02FF
DkoxdDUfT4bl8AhabMtgs+Fsckve/eyYrf/eehXZV9/igIpcmr2QLYxDjk6s68CX
xmCsccIK64+1ONHnk6IwJyYXQH5D6bbsiyulfN9dLgpRmL6Q+FrIxG0MgCDHq3Vj
pxuZrfgbEg7YcLqOJGr+dKLLnYGAc75YMWpqJaB+KjF+F1h/YGBsyaIgwRY6eu1J
eFyVXPemFyAajRUKiShmzySsk8DAcGPhue4WIl3d4M2wngrUir677Tz1x5+co7Kk
a3bP4vd9f9uccF4NhVCZA4/DrrwPnW7sQgVxQ2NTsOMwUKUDdqEItN/tbuu6aQss
h7DDTKsfsfuXxUCk1bcak0x8C/CkJvcThNRY51KtcslEKmRPZvhoKMTfCPbz6HqL
9/It46lJxp4M0mcTr9m+f/9MWQb4SwhKyHFhExsTa+oA3TyF3UDczkTM93ydnqy3
Cv3xjipdda2PcY3cLW6IvOFyBJ77XzbGLAfhQxwbFBC/1401+yrO0MVa9gfnN3Lz
GFRZe/SYpnDNOQ2xnr/4ccBFcimeI4r0cBo93RsJTeu+/K2UNXNBhJAfDaShYkAj
U66MiRNF9JFk2G7OMg5h5Mak8ggTiHGkit9JKkinwOIVTRcSQmF2bZNTx6c+2jk9
EoFVAczcv8fzntL8dEpIV2mgiOnOObJMz3/kmiKpd2flOuu06FJPKaJ2bUhsQC2z
ivgYgDPMgode4KWfrmHDmdH2JVs+aLzzz0BGi4OfjWQ9O9iwYF7zdBTXuLdN8qMh
maBWq+/C3+2+6Teg4uuqMljZWVSMYqu7mfyCR7VBvB9JNWepyOLK9S4q/U7VyEqu
mlTGpyqEVAzNwiLE3piwgG2WVmiLH3sC/OHICx6zbP4V9U/eMn4ucgHiGFNp2riV
wT3XqnjRfpz+kt+0CQbpYLCrMSSxpYxldj2+qvlUDgN41ahvd+fuQ32MzLeDypyH
0TsauO68pkGYlC8GRjuzZddcvhAbVq3/eQ1CEYySxPZvaYCb7YOoPxsXqhwqbE3L
KQQJnzJuDVo/1yt5YQoGZsIQ9LcQTnHLMNv2cTiiivjpvSPcS/eX/FXkXClny8fg
aDqcpxwJWqHoh1a7iC7YO6meAsJMsLVKByhNFowdOUtp5ZJZqSEHcBJbSRizu1Q/
3mpNs84D6xCdiZpQIYBaFsdkeh08gtaWiQJHAh19b1Tyg1DixdSDPRRZpHbnNHW2
5WJzq9iD85s88mVcNhDTmg1+rO9soT18R4CT04HQ0ifjXMypK79qwdFkE31ruvCM
az4EwCOJrTcBkyC1EHeQUZ52CnIoojJ9shDu66VAQfpUTmy+ry6U1inmgcc26Ppq
Z3BXPlOlTT8/fDAhxPs7u6Gi9WrVIXPH41+k0bOeyIXWfqGwhGatuIcKjpXUPmhY
yBOtf8Kvkj4Ylz82w5zCf/OvjZJ6CqF7Ir3I6Ob+YtqvGPEUq5tCJDPbtlkJtdad
kmwL66oodIEFSDzJuXgoDUxoIjbV5DbBFUlCYgum3SKWrFqLeSwbmDN4UYuxZMYW
kxCBCw6kBU09VJ8kMsH93uwZU31UACQr5Jd9WGbtstBK5/lssrp3iejKtJl/Vdgg
zb49kHt/cn3Vd6slyF/t8z98cvC+runPiUW8XVBDBkI+E+3ujiwOmujnUHduQv/1
Pp4NGsqQ10uO38qy88BzrJml1iC/G5gvhACjPG0y6ry+d2MbBHxe+jxdZP5SYVAG
7NBGfrdPQs1B/3wL4HAJWk2+ck1uxrPu32+lEpxCBMKgNsazliYsak5APt25bjT7
oDVwbze2TI/OsKTTypaVNHar9CdhmpsDrUTguOGO1K5AFaoce0PNLRjGeAmi1T5M
40CsTZFyKsT6VLzekDrM4RB+gzMw2Hf4J4PhxLcdqP9TXlFCzkU5hy2jM/1mZHV5
f0uhH3i6bn2EphQlI7ctRLb+WmO1QiJ2KL18Ow/dAKPhUC6belU+HfAc8OjEP2Q5
BtlpFAasZlv7fQgY7a2MuKbRj1gHk90BpScHwlg6Gnl7dtpXR5xAQ8qsjVJ3QKKX
m6SIAG8saJ9VuF4sVypExNLr+ytXJ+a+1rwomBfgXvnm5C7gNONc3NtcFBtAx6BW
rFdlgTK7hfX9BQEUpduKhLgvBpMt4b07fcHakneAqtwGWIn+HfmwlMccqQ2Y2H/A
Uc/e7E47QkWZjcFazZWbyd/c3lRYY/V6mriJ2WjWRUvcLsZJR56mmVYn/JmftJQZ
aYQ96OD0QCmoMqSXcNmJUHkYHt07B4Y1TJoysFD5SBgRmdR7osrkzAIAi/Mgdg/e
Uj7ZPcD14BdtEPrg0JG3/IEjdV69OB0gADkpbsTiE4+elFGn368G6GSZK38RnWuV
FKudGuAaaq1c7svPDOf3/CYTP+Vfu8MISrzXFgdiOWs9QFPTAqfDF/oC4efV+dua
n/D0T1JAc/dbzS/SiLzmkcacQ8Q7NDKo/5uvfcz12hLEofCjEJDERzTnBzKllo2D
++5Fdfm5PVZIaBn99VRxANBsVgCvYS9NYaTD43fx9cnveV5bcJxjussk8ZomAAJt
/7a9DqG/0lpmttJOr32BZjgUfxi3LS+uUcS/6FV/PLYAgUaMGvqO5Le9rhF+b7Go
v2SXmxOIdRl4wktF8rqng48fq7laXENuuK74fLnwj1ehgLS/PUYt3sJeJXXqRcUS
Tp4ZocXdMU/qsN0D4jU0dywNbs9kUnt0OEWFJsDCHKpflGfxzUK2sKMzeEes8qQ/
xB/E9rxQb+LH3tsyUS0Sp9PX/olSN6xMoKLrXhxmY5LlYd/Y6zWefuYd9oOMyl0I
0gnGz/HRAcEQVTrUuE4y/UHAMYD51N2LNZv1TBSMVq9bkYhoSPzLZtytO4oJIy47
Guo3AThoXJyVYnKc7aWU3PasvixDP2Alimm+5YiEfzIzuBkAG7V6DnqJaeBmIID3
lK5HsmNaKMObom5zIT1j7TmzaGoK5VueBjgjVcQ1Z2zoXGPZwUSxWkfoQufgZYDe
uHTr6KlSG58HGYcl6MKE6tduSy1ckqZv+D5p06/0NEmPaUkEpdyMeNOh+idW3f9B
5XiVdN9NqY4rM4bg71z/nEVt2EZSdDWQLM/w1hokAb5dg5toqudDbKly2qDXDxfl
2KiwCVKBTbO4vm0kO68slgO33lPMZxP6H8n+gJNhuHSo2lQDv5KZfVyVtFYV3BHx
nBO8Kqw7vjKYhk8yXFVPntAI2unBurYws/hcZ0DaC2fJx4kZn3lIgoBsNEGSQWbk
hkuvS1SQur+acW45QRAVnvzlhbhoLGBnu2FwEYI12ALOPOWWAzk41cNsuYTt9UOd
7NlnJzB1Am9A1Lruhj3KWK3ca9gN6WomoxFxq+QMNAs9xNoIayR+MoHuLVCI/7Ky
r2SigbSgHoa/qY5RmJPAa2+xXk/CkJCUybl5cc97mVTzErxhyMa8kkb8LWnMEwZZ
90fnxDJ1+xVB1I8Zsd7YEi8YTW5faQq4t7SMmi6y2I1/fHS6MDTLHVUZ7RFa07us
fW6zoQ9zVO/3qd/WxtT+O34ChTqFJrDTJFMEcQCeB7dsxq7JMs7GU/NhIktpLbKH
A+F465rS7w2uZiK2D09TP1DXSjKz8VhK0tqLO7S8Li0t7jLiGtlYBgXZoLNAGilX
xRzDwwTEhXKbk7dwX2pxWeHWe4719c9oRYJYqBV7kU6wov5uBtSuatzzq4P9+IM+
TpdDwF0DFotiNh9fm/tvnrIbx3truPYry8ZiV5q7oaCGaxI7VJqEXZcwQUtTfee5
F4W/+Chvv9V1sjDtplq1wVeipy0+w/nd1TxVVYxFlh/00Wetd+GxqiJ8OPUGwchi
+DVPk+NS3weFlIHMQWh7rsxMKXLiN6dz0vJhTLz6IzAkL9whva2p83jIzLN4/u8S
atlGCTF3CalpDMYJQddDhvRsLaHfxqyMd2jK1p9D4plmp44ha1XTpMImnqYANSzP
8WvOtNorxSNY1CPkx5+MATdkNe26VfZm9KTpQk4o8yVzHmzuDS9Mdt45cTwS2mac
HMg8jwQIsg0bWG4GmY4MNHeTcL4lpMEubDrBe6HNlndPGkpxZEWBieOBo7a103IL
L0LaRcmLisM3bzyMw6CaJDI/kZq812qAHQNCK6b0AvgucYRBGUcuI5tudunEmTqk
Tl/U9Itppt5MjSztkTQalPImgocBQi9pIPZehAP6FjB01vvHw3uF4tLFGV+sRbr+
962O6D68wysM957BdB7m9xcEUKUTgVeruIDrSSrDDD7h4C0/oSLXBk+wigklZPEV
zZCO1pKY6/3IM5B8CMHZvYPQZSjraBlG1wdJH2JYIfohFlTT1No1srJs/96tQhcB
SS/brdzanYkyPYdad3wB3sCrunq0txACVlbkiqYl1/GsskS/rSR9k7o/iQLbE8le
RKD6ikCgYeGt6JnqJsvKrDrgV/bRyPwAZZWMN/LFs8/i0tOZbNDZS1p5ZDd2IND0
1otjH1wp7FplAIEq13osWov9dXixmvI3DF20gSiAd2Vp7pWHnnghOqQwbxOlfTlA
XmmRihypkN99a4xXG9rrUCw9FY3oImMd0OzDZbZbKvpnoQNNacbo+Oq7HgRLYc1i
M8FZGGyGn3q+Ldr/7e3QSbyZ7M/Qd6WR09lemhheR/I/NWg/hSHbaCsQt2tYLd1y
8S4cu6+zQV5cbcT+3vK2YNeu4j10AcHXHI6H9hiGtwx+NoewXoSXcalijbfne9r8
f70GxvC8z3n0EUat0alQrCWWe9aKS98/Rdau8JwbBZuZPPudFKEIYcGArPvzjUyA
9D16YN59mk3OBvjhJMqmzxtTdKs0/VfzJ2wy8NyHNv1dGcXxVrFO03MD9l66xwYO
1z9TDN3mSLKVzGwDuCHBjgcB7UByNlOYnW0nBmxXF0IYr6W3SsGZVNSttwc7ZLzf
ZXB+asbjMGctc2zLTcavbs80XD0i0UowCvs1U/RQ7Y3vsaefliBvDTdm5JQ3IOXI
+lyXcJFYysUEqkMWoyZGK43Obyd1/UIGWa6EYqw1SGZys3WnqziqqOOZfuTNbybw
seaKNvJJEIHZhd7pAIgvzaqTKs+wxP2TOjvl5MyxRIMQLMwaqqS24USpimKxZw54
2SH8MgF+qTB/+INIK2F14bSiAVC/ScMaj3os1exmESYAY3LrjLtGyJ+QrUfbJjny
SwmNWp/dRDuka6YK1OA5++A5C1oJ7Udc/21nkTRJtXYJRirWGXHG+A3mTI2tccP8
ULCl2UgxhLKkxxRuYR9rm4qojs107WFCeTjqRZXCfA15siPmHlcKY5lzEtBSOCsA
giQzLTFDgkb1IJPgKKIkEXTT0U79qI/XFgZOYHIWmDizgi/0EyjuL0kAO0E0za+R
euLUnrlhL9GSBWrNA2JcdIvgMRsWv/OfNuajlj32GVqw79WuF5eZ2cUNKVblxLqp
5mlcIynSHpC9af2Wr/6TPdZRALRLoA8ChPMyHLHXRr+qI2BdYurVU6uYOGpy7QsW
vokw/aKzlj6IXKzuHkj5/DFwZgzeWeGE8OW6zT+8GVgREA/EGahXFanZJEnvCMyX
cry973Gh/VWEissLV5z6PI/+HeNfysO8cs4CjDoH2QYter5SRC9Bu0YQ/hkuBmcn
11hGYE9FEkHHPAosS3BuNagj66UjJCQYn6fQqX5obxuwhkWXndoSyaUBntPfI46H
EG++ZHePRRS68eF7BOokOtzwYPjwn6BLHS0dWADaGT2kM/CTJt3nfRAXBWSy3X34
kMiHnMaS47xzC5qyPe4FWUQ0sd6z3VLSg1qLfYSw8aidph5Z9SCw7EPkluq2e/BZ
WdR0UHhNnt0Pocvv/tHDodN3Gr64NHxoq46O04N7fNckU4khwB5liMeMPT84zNuT
yhrXD0PnZX6RtyiTxHS8kUL/YsRRVrMbQ66cZHjo68LLFiypnf9OSUnq4TxKbF6r
Ws4ReA0DCt51TRB6c2OBxMC7JGOKD1DR05vVCu5k6X5EhAeKsHLLRUcKJx0qi9n8
DQrhIwE98sWEh4Y8E0aYyVSB+pSVE8kZtZF54t75Gjpk+5+heamaNMG7cBQPozRa
sZI/AaI9Sm3XIynXwAXktrgH90V2M0sHTRM7+SlBt7gK3Bg2Wm8mlPuIiDuYi3/G
GGi3kuRAEw0+v4XbNRnV28hMaxmisPEFm1Q6WS4RHCuiHwQVjzJiVHJ+XCSfiRFR
wmtn5nPY5fz158FGFL3w5AOVRYfRPCyFi13OmtD8oPMUI3V/rcY3X2lHsckN05Ec
6KrGnl08stNW5185FMh14IXTYqFsqkRjvppvY94XNb/wfmw/dHdXOtIq5fZI0PpO
SCOGwZ16cmeDwQsJvKq+kDYLR76MRtEvp9TOqyXWVhGYTg7FTFIU3O6bfwoSX2m8
0aPFXt+mcmYIRuolvPt97aTdsMGT21d2aXFf9wXA1kEPrLFXuD/bPsitIVguURj5
F0m3Vedm6kAbP0eF0g0vrkGtotrYRkOCTH+BP4HL7YaA0rWBTa4CfNdqgDx5iHTF
1bMf8GR+pAJEsg+Rosx7q7tjC4C9dP6NU567RS+oKGMIhB/NcG9GcY8K5YJMqjC5
gMBcdZyc7Gb4BRR/VZU5C0NX+YeRzByzZcMBYK4SJXkFx2mWfa0IwHBlbTU2lhjB
oTxW4308QRa4lu1j9zvRmuJKdboDxlzwEaodSiEh/LeXUbhC9J9zcY6PiGwIi7AX
eLnu+nNYZjx9H8UD5FBOcdxnNrCjxwrhyInMCEa+QVtuN0GQM9l3tKBmaxVyEdEi
UceK1Vq2abIl9KLfbzvWV7OVF1jUN6H6eeEDWCBfv6AlSpc1kSfQybE/Rs7BlX6X
5BTxXFm7EeEM5Y5+V7Dp14gBvSyxzomSGc/RIuHne1jMDvMwRd2yLc57zGy+HHTY
GjR6Sx+Cwr1Nj46LuTlSKQfi8VfLi8JQ5p9hj2EvuPnxt+D4w+nZB4FkBZgNiqaW
Z14aHHplQAnUdNOZy2oTrMZiKq3eC1F3KLztKocbMMTB3FsuC4/l0+1x4hZ7pDas
O108yVVjFy3FNV1KNIk7ZpnZquGEjHCyT9Ohg/x+QPNGXk/Q2TY0o0iacO9JNoOa
xScT/D56bG7IEIzSkSK7XL76OO/h7EjwVh/r8iPCxYYP3bDWgqGKsFTrhmpAfIL2
d4UE3slhyySvNDmQV8XwYjVaIYSxis2c1nOn/LRjATXla8ahrjBW96lWYDNM3pzF
36sqox0PK9DMtdBAO2uGgoXQ89mUTfyBeWgtuoVLa/3RsqDh1TJi3Niui272POwH
9JXYHq30IdhedOoT35Y4qZlFMBcy8CKaB9LWZPpLH138krFhDH67vbElHGj5y1IN
XoHCyQsyUMb9hdw0ukB7j1ihysPKEvfoXgUcgFuLheMZaXWzNFN0hobUCKdI6D3v
6ejwTzJWgSQGIXAmMFzn6c3LCYkxdePicGXSGwIgvwy1EkVjM8u19WeYed+nHuEf
Bvvuuy1jzn76Gp6Ha1a2Fo8ECWQTUISyu6R8k8EiahU7uEOvZtqxV3ivB+LLk2a2
2g3F/PBaOSoNN3eimJQke1n6jk95O3V1kdr/+cr8aBTmKfIbi5w+eREB3eaR1KYf
+K63a77Kgu+Tl3Yr/S3+8eVgT7JApBxKFz++SlPUx+ZsJ3mfDJgSeKbkULqhoXew
2dyV8yRpJPU6Y1aTuYAwqwj06K+HeCjsYKGOkcFrl4fmafAZyfMoppOW83MLjXQ2
ku3JoIku0vsGA7Q9k2/mZUPFPYrfsDK8cj2dey6Gpj2il2bbY2vpcBPRQcS/Tkxm
pc1g2JJ2+7QQm6j8g/T8ZXx6zy/7ju5JjiHH5dUzfEIXnMmtEhq57bk68lkw6ZI9
lVS62BdzqAACrgVCcwDvzJXp1nAIvL4e8YhzJTzaLZFD0bYdy2dlKLvP7tzsuf+n
yUPcmAH0P1IdAC9qal7AjxI70gmOzLopsJPfDRBsc2wsu3tuM+4uj7MEXymanjDU
0sLtlYv9ZoOKUPhQ8VExrABcSSfjngtjR+JfQ4QAe3uqPlyp7cpEpkVYLrLJL2bR
NbyFcvB/yvS2XSdTbSi3aL1ND7AW63xS3a0U53gcNppdiSqfAIQ125QN+Ap5iNbf
a4mMtK94Q3E+sBjQ0ST5kHXqkLw4iBBL8DR7xqkqW+UPn2kJacf8A73XX5mnrtuU
hy6ywbQg/8yOumT1kAEaYZzHL8VGFDMWrOvZGJ3B7r5EDq+gFWYgweaezIE5H3Aa
lUjwY1nhYvTRrEN9Cykm39ffc/mLt2pjl/UKma3V51WJrIqz6exUVg5yhifBHEj5
yz+DdBO9tiflHNF5Pa54by0Z6+dOd0tbzYEHBITNXgijls9CBExeHrMvM9bzVc4M
cDv4daZr3JdoRRv1Em3mfXtjdua75oWFceKzAnOLfDZsfFLpOdtN7WVFZiUJiI26
0yaN2/ANwBNZr3W8PsWSkIFsSHMV0r6pO6H1sX3wF6KXP4IOfPT/ir4brs0L5v5N
rdLmpxCVsHXvBEopboNg6CD7+c7z38uEXyj6YPcF6+/KgjVnMDblPfC5Lv02NVZu
QfIUX8KufH1wG5TXPL92KQrCUseA3kV4zyXcFz5Qh6I/R95xLl/2aWLOegNdf2ln
Atrw0xkt/z7TjWzBhUgXPZRJ0T3W/LG/XkZFJ11ErqifbAD1pOkIIhy1CrHPtoPk
oziuzktfvN/3KuLdBjVgCo1aesZI+Kq6nmuG4YwmkfQH1krinHqbT5QFDCeOgtqF
/Wl50L5keGN3ZSMqykh+mO5Nt9koSdbJIqoN2QVWpKsDeQeYSYZ0Is4VMfguZfnB
FK4H2HojM7TbnhwPF6yeImZFUhNamNAE5WjK5EPow/kXEuD7dkd/CzpDkUhT9Dj6
PCrOSD1yAJDGSq0sovDQNzaRz93brYIW1M16+ARGKwMcpIBq7QiyNJbN7pGbK0sp
IzIwN/Qz7Ej06yQBzRmRybau6xo1hwaxjkPRym65uugurAhui5n5GBsEWM9hPZle
d2+448qxw6sHZdjprqeWlM1Ql+qe3XOwAsV2pFvzeqLio34Ul/2NMdhXGTh3BFaT
bc4g0OF+oERbVMT0BSB6hbglOOO80LJL5o+fbPVDJnehemmKEg/kaPw4l0CzrWPm
tDSJaqwYrPDWbfwhj3No+5MeelCfz0tE90Yc3CitZ+DTect2MS89w3z7CDZl2ooF
Ty1iZIE3wkOXsbDnZoQf70yxF4dX7ZcKWTXkbc1ftsOcKyOb6TdJaXAo48nwRK1H
G3I+ZNGQVvfuDJqV6QzIh0IoTHQUB1y6MGDvcWdmu9rxHEZ0BbnBCwyGP1Brw4Gc
JmMnu5fhMps/3wDVFRdxVbRI20fuvVUZVOTJm3nnxYMaPPkG2xKQfxYwMX/XxT5f
lE4b2KCGvcUrBEms/ZDWADtz5vjPCC+cwNmWOOO0T10B7JdTMPmSqol47gd/oRpj
9lTQJK/neHXywm838qIERdt9ahnjz18ZoSEHrRM+aY0vIMUSnVcbpAal+PYKY077
EaynQLe559bUGuaMjGmRUJQ/UT0ELOuU/hn9oYTy67o8KTP1PdDMnpGMEBFderP5
hYCkd0VhuzaYPl0/blbJfapqGkzsIkxhXtCAs0ijo6p1sOYxtNr5iV38VeWVmZlS
FzBkdl00vJaeTHITy8JsHcnn9/ocqHkBq/TVNnSevwRyCchIKC17N4e8/1Pr0eDV
gHtXDDWbHEW/ZaU296XwDWhs5HLhgYfgUBtYFK6r+KuxkiVMOWNlIZNNaurWyKVu
lVwyaryPcOG8OnPNz67nD/hCbXDsWNktB7ll1BJrBSXC325Alo/ji1ZgWJcWriVh
wHMu/dBx5+Gm+sP58zZt7vB1CTGTQ/P6x1kiURAklqmmnYYBmPNEOIgsyG3q5o3T
ZukrNLgWArQAWk8jABnUW/5BNuOG3NCUp/66lrGR4O/HSGXUfYjDALOoJ5YgzfoN
t8M+g3idccGPkaKTSnLkDTIAjSsB2fPX/KF6Q5qkFhLF6NMqyjRqs0pjblAhbgSc
OMLmKrX9pkTnZeBb/398SH8cJkzP21DPH0+a0M5hM1QG6yg0/TOeudZNS6jmDOM2
1dlcDwDaZJaEzkL87Sp+SLB3hT72bLipgZCd+tQ+pUVKKpG1diQ9lfJsyn+z75Wy
fVaCYN+uLDZSziZOTyBRw33Q4WB00J4e9LIw4jSHO5ODZWUVhbHOc39k77AD8uOw
X6/ubZFTpaow3KQGgX9U56FUZdTscZDN8pZap+MG7g5Hre56UhxsxuXJIWizzBF0
tWuFE7mjMDqp/fIR4dpKJd4V9N4cTUWxYsA+zJ/xYOIpUwfNTvsi05xU638hKAYL
/UhAHKwKa+UAZyapS4HvLLHE6g1tJLS9cS0J7aUnBqkIyI6uMKQ8FA8KC9+3bshM
xAwX+qMkBRbDxEJPwVqDv3Ujl8xuJI+YOwz12i7rCFrs9qgZMo/88++aeUCE/74S
rxaFT0RmS5wcUHeZe4ep9P2mVaq1zshXnXPoWlp8uM1+42V/KT+0ySHtT24wENtp
qbx6St7+D9xFy0Bwp7weENz6AZR2ii8OU9eT2cUtAU5xiz3cE1eFTtenNW4f9cnp
U2XIO4z87nmvpqMp9bjthKo+olHhEU5VJ7d3EUcgkZHGv8ijQi/G+I7pM24FdWAM
q3Oido09JpzVrZusPKIkPpfsPXS7GXafLvO69h90swB4+CjC7nZbozermDZhH2N0
17BB6k55CsoC72JpTWZokHWu+kUyGH/gtvxWYtXdmcUyGjT/kZgIocO85dAGCoJ8
GFHRJ+SlAStGxXRlDxBcuu1uk3om+6yOidUU4k+QLfmlqRqSDe/ndKvA4BRO3O3i
yZlnK/YGRutj9WEdQPSQ6QJSm/lPYle5g71IoAsjCusa4LDLKp5dc9aMTPWVW9aA
yyalSFs5JeuYEGRyuLGaskFU6nsnDKjgWjNI/zmnBNkGg4k8S0F7XNR8EkNuChQj
60aF6MGaUl44dJJqwi19P0DYIqwce9UVUvP3tKglXVqJxML/6dXFl6rb+KEYCw0F
MYBXRtTTAMbQ060PPSw6MNnr9HseMDKz3dVbAMx7KenZXzpXVMJKsklMvz2ej0BM
+Yq8pIJidkx/SyZMhqpKw8ZXJxjlPye0FkpLFAPqJla1/53ZAHez15zsT2uX0QV9
oyStJW6Hz8NQYDpZEISqlLVK52ORbfWxFY6LDv90wus8yD8g/9IVvyHZF6Vpiv+2
QyhaeacQhKO7lRuW6eykP+1mtHkihukHXXZUqYbUZEGE4lsfuwTeYxGE+l5TYrsy
iBS30qvJBM5IthXjBopkANZSbpxNv7w41xPbaNKYrYCoNdYtHzv0Ql4g6K588uF+
1VXOeKIVG3h3HH+dT/xI6lEiJyCd4TCdO2Nuan6E70YbCTtjGE/OddufwCP70+/+
YFWylbb1pZpkUy4fEE98oyQo+5tYGvE7bdhz0ctJUPm3pay/zJVqoTFrcSYLU4V8
oGLg/1VhO9a5WXafildz6I6uozA5QcMS/TmDP1bV0plK1Y1IX00nDtkB91LF1asN
vy96hYIMBRRSaU4MCi3JJLPUYxYrixjrCcqcMo4so3MNqybCwjYTQhbRwAEXTKOE
UOcSDJfS76pMhPMvVwjGaFIqLOCO4LIgSBVcJ+ioKyajmbimWtRPFzXVASdX5opz
LC2P6oNDiLD6EUwEl1dKqOR6DvYGyvPdqZtP45ddpv0l431w8N2RIoICEvwFQoce
2OS/5CZEhzHGzKNTcLhw72WRKDpLBt6E+vuCB8/MIOWSHB+0BjChT6NT69nYOApY
PZfBMaUK6Jo6hhW0yLwfgs7IKCkxZDmfL39WfGuTqslWv9PKegGCu6KirTssh1NE
agNLaX8zLaAYesr866s8bO3rZdA/NZKKy0R7rp0jgg2YNYaAdoN9VqACm+ppojvS
YxzDOFlfS58nqmWG64d45oi9RJfd1Hgp+HflkUDly1/Xn9/THkF39Tgq90PXt9F6
NBtxcfYgnr8P87i+OiH44bDNlMG8SfmzRam79mFk4Wvt8A+VlcAsNxsVI7wp0/YQ
Xj/SBjIYjdu7k0rQtrRnaq0HOCXdPlAdXV7DPfyn4BFcsH2DUEv10HEV/IH7XZn5
DSoFnQ2qndBfpeFQKygc+QNyW2VuUYKmNWSVulzMJe1CF51A6VrrdFxwKZh1lvrJ
huqYO2TX8QC1/rZGKcU9GPIDp04NNJ19ONFoIK0zOTS17zyO3+ohG+WbtOcxZqFl
UGzmBjZAc3CKnWd83molZ6AWt0nGPrqMGSYaYDhKcDBwcOflSi5ocHLiFcomlQrB
tRWl9QvfESOrCGXts2RNiRM/kJBRySshESCVcE6+5z9vF97qoMS06wldmD82NI7V
Njfi97uMxNcgsexdhA19sqrcWDNBd6+yUwYrwwPjgac6dFocLBpin5SCmfFSfOgL
802WTMMEq2HOkldzpz6LBBZkkE3waPd26CbaxRlO2Sr9WJeMfIS5hOJQtLBIJR53
v29qhACVNHCvcqQVcdq6/q8FRjmaxt/l2WzWBAtQRhti1uiE2nVRS0BE9aLXit9s
pGw3l4cBplI5UhLRG42xjI8dBBoSEz1spKiSQ6LhV5JTpFGM8NjxXrnKlBjLXPIy
sMMpX0mVOQL+gYHVNZ0xuv52KqUT8zBDCJt6fchcexI2o5JYn0D1NI85oTskrPKQ
i8eDO8uiebDbblTZn/XJFDubbohiUepwkr0QBb1YdAVOn1dKm8q/XbT1de3kbEZy
0UYmWAY/QOY6qmNEJ3VAgpPmtAg7dN2P8BktnbT28iLWJzB2EIhMUJ0a9K2hPRH8
eGqYyYi43ua6yEnWRzC6SaKOHEQddyeusMfyP1gz4P0clUG5cc07hXllDKZJZ+Qk
HfRHdo0kGry+iJRpoG+wx3bnEVhk+H6TONowCfoPeubktfl1Yjrx1fvrnY/P2Vs3
dAWGiDLIX3at4AVzgeDOkKGv4MDYBMTXVkuc9vxh51FssB4gZ9aLmuOmtoXKU9iX
RD8r6sbEiFJd74TyJfGgXlW9pMdFdVzfX6E+G2pcAS7UlWURrMP9nLEeTvwkaQJE
pZmXICh0EV14RY3+broZWqhgCKtct5XgQlo4gQUxztdkJ35ektqmT8KYQyZ5/Jla
SR8StItalOlIZD+WVMc3d5hUYP8ZILwEx1b+5YJEoYuDXEl2AvEkDSnn68vmO8Ot
QyJAl/GVjimuBi2gxpyhBJdYrlRW8yMhYakdpK7ByrH2EaN02uWWLD+mGLScRTK1
kDJ/U6n/zgAgdCvIpBt/5hNbyy4a625Hs38BHoYG5w+LV9N2B3xog+koG8hG9A1J
i3pYqVQ3TkUdOMt9IBx1sagv3nOXaSH1erdPQwRMVu14VBfAJlSOfYVUNK5mkbUx
GKxxpXKVW6wKQB9PT+1t2Zy3V+yiuY8iMTXDDQmJnVRamIxmJ8XFsqGqIH4pDWll
OQg+LNHHJMyoZX3CvUJG+6OjrfJplCwTtu45nYin/K7oioVZSdWQFoKYxqEWfoUF
IcsvPveHwOICDiekLXE3pEAUyio7Ddtmssz80+pCjxZN29uuczUHbDo1oy+nPHTT
os1OA0NuzY0bhEQUNqJ+PGx8UTwlvEjAccHZBbc+wLLakDUAqh5mKI1Xug5Aqf0U
SgM6bWlt1yy4cfaLW5qJ8kaA2TjYGLgDjdu6GOLhFKfpnTu0DPfBsr9J+v8X8csn
Sk/ovhkPteTmm6J9t2amo1vqFJVrPi6dDATb3fjl4/4LZLhoKWRd22NeDq7h8lCH
avYwbwhUJffvd1FTljVI27YzTQuBB0HWjlWzT2ebGNJi0qTrboRc6MulsrD5nAqA
3gxHcQKDLXfpCR60Rc3SKXSMfZ1haHuc/1VQhYjeNWUroeorRQwd7qSJF8AallzS
9PE52Cf/fYafNTF9FD7D+a+skyJgSKYDOL3b/dUx14o/kN/9pSmvrB2svGzqTY5+
v6vExm2JXZviNFmdZcFZjolhVpWaDVM7K/GgBuOySCHPrP0fOS6BPL44jZ1UReam
HBhyNdJWfR8aV5TKBPzw/7IjXa6p0xiGFyzpvtmS/qKIyssVAxWaklMtEV9pPiIW
t+H19VP2mHPjv1AXxG1x/pEYVlS3V5b47weT5RPXQ21uzGdMDDuKUqIQAH7xDNxd
q02oIGy0kmlHtv2mi/NTtjRK5c9P5r/EvLXCfDXk+5aK6DArA66Z+DyrMgahZjkv
ngr4KDD/TQLMX57pIRQJC1njAXhZ7VfUFiNuuMaA2QeoqTjswkWJ/Zq2a43HDNQu
v89v1/QImmPxLb9YO+ikazdvutwur3M0Um5IgcS/qskiczfzSlofCwGx/ksO3nhd
aMaBGgDUHPIKn1+8gMpal8E2LCyLFAjffiHFU0unKMqfwwdOQ1PQjjiA3L9Qdldn
SuzPI+OuYsGw4dZUfP4vOJ2ZgY85nGWHCpuGM4s7JfzrmpuKFDzkIsqeiBnkx7sc
BLT7c/fmluvm01J8SUTFCn1ITLUmcvSzxuo1rGIImcKsOkycPG0DKst2s7rYKMOy
p9KHFuSALOrIl+g5J9l/fxLxjCBfsYurgvHYyZ5ysVRcXfNx16vuM4WxifCVljwV
ra9W4rYAGymPyCS2ifynJ6B14mzfDKGryh0w3mOiCv57T1lPO3R7TtTZLX8T98YL
jdZa+2EyZ6Khss632jttgnNNNQVfgOwaoCyMPNGokCrANnBeytOKv6PpIYSZVrUG
6bTlQOzz3QuDaAOqbj06l62456JXaWYyLisuDfTjqc0RhHCW0BpwFAM/8TpL2no/
pAZeyq34W3jgYuQgMggqAGzTv0gF3zgnTsosev+Kvb5laxrWUGOjl2j/yY7MoLDD
SUCrgISpYO6va6QpD/+AtY9bb34aI1uv4OXKfOWDexd8hux1/sMJ0Lv+SALEPO7T
0fAMfpVhZSgIxDDtZKf4VG/xA3RY5wm3FwIyVzYagigV/8chzIfy8DgvbOewes8X
Ilrrfiy4hlJDBpLqlR4qmpP1hzQGagz5a8To4ZVEl2zE3F6LUKeugik6lzHkxKoC
g3bl1+YeYn1nuEUB7JI6buE+qxQYuBYhPSTCyX8ladOUWdZdayvEcTGBZZf6WXKD
yXw3Of4/gUt+4Hq2EG9wTv3Bct7N61bGeX5m1Tvikrt/6k3Xzkirf2pprt+tbDHY
Qd4IPUQiphHW7nc/MpVFm0hI4hzG/Q6w+cP7fRW9iCg6plfPNSBdt9rLR564MHFF
51kLqU4BZSo1gTwfOO4vmInSR2gpHykTp6RyEyXaDMYvu7+CNoRHbNWWbua3blnE
Id1jRpJqgX9wJLUwEkkXp9abtGudCg06rMCv/GpSr3X/G63DS0ZEkWLP90wQcNn3
z66LBv6jbzX39zzvu3RBvBQQSSvk9rwneJ6FQWrh6HIY5sHpfSJkTNZoj15KnbZ2
IeAXKyS0CGzxxemrXOFC7A1vByOLY/EdSoiEqkJUD1hbqQpLSaHldVmqbIZcS+qm
Pz9qHiPIodQHt21XWbeGSwwV9XZTK7BnGRiRaJ1mzAx1DbDXRgAAQzp5ZN2VVVyR
KQ6r3tWTfhtygrQi+bfrT+JsTpN2pnkdBSxe4GXpXCfIrgzLaPmmVAIog7bnx4tU
loSxSsp/TLjdXupJsI2FXlP+dfDh49mF9lKCBpXry35m0jFiTLQeR9oYgUdRZyrT
oN2ZLD5GQqNV2qiiAaJ374cDGQWK61eYs6TRnF4c9OHKjomyJZKOhfaTlRk1YrBL
j+P6ub7TDYFp6bL3JPOZiJeAYdr18mFqLKYesCQgcbnY4asAfzrQ4DeaGlf2Gjpf
6wNam7cz1frVLrk6GAlQqxKJ6COvajh4wwcVujQCgMbanuxgdoCexsKOOEloCSH6
oe9syLlcUddOhR9yOBnecxtRcASdMY3x3vpcEuiyBp9vnocRG/wLsigqd6slHGuf
LTavo7J6cX7ttw5NeWNHmitH1SCt4+ACHBJ3YU+AafM5O9b6XMn9F+60+WLaE4xF
XKjYV84jNTe9hChkwnPU7nscBai5wSJWtK7vQZxIyIrW3NDRntgzx8dbnMPkMwBN
zFFn7FnErHxSXXma/1QZZg/VbK+Ep0UyAkspb5CxHHsXdDBqb79CP29n6ZfPlz40
72fap2YyIs+QgTy+fkK+OheZ+xeOwsiyB/rfUoQgErof69rL+HEwO5OAMpJDZWfc
N785kvjAD3JLFKjsC/hLBX7b4ccOAkR1p+GURjCxIFpeangs7kMB8y1QNfC6cBvq
Ktn8s6Ns19ikYa867Kj1IH04f7qdCIe61BfubpBz+KfprHa8aXsg/UL1g3W2XZjr
s0WG+ZO5JmQUTK8I7/tUjfjvR7U3v/3FugcA/gZ3qNinROys+p++zFmGtexvDt39
TAgBjMV4GHbt7SfxCjfUfJtJoIGtfn8+rY+yK/Xj9xZMC/dDRNJiyjB3yEmD9JqZ
KyB2WG45LGUwOBJHm8wMkJgb5d1uvTMDqhikzk5eqaY2FBvBc+0HVAVvMN4mC+0X
UhokejZfSX8jDwirhs/55q1rSUURZxYqikktY1mXFTjWWdQ+IOCZrxOa3vt6qusa
pmArkWnzHOQeGfj8Dzf1nnPFyesFnYyFnr9oWIPvTpgljV2mtw5d8ztzVZ7OG0rX
r1cY4XmC9qW5axLS6+vgvo5OJbHF4eOZaTpHz01eITfR0lDSf+DW3QfT03aWEfmZ
InhvF20lxh8lm4BgYYzmViY4r8qg5wXfIBkhORdJqt3isej2vD//ipIaUzIpF/mq
f0aGhD/c34rTgP6JgkHczYeE1MNE1XhbSZpPesNxTBpDTOD7EmL4UunBolkywcwI
iIEaKKyBqZAML1J6g9dXfnongb5YuV9jBLUzoKaGe8ZSOPZ1mCr3+g/W0H2meSje
f14h3wXHtbtaaIymmw5nsx9hoeaAsoE8JvApLl4JxzUqnJj5/1RPptPQl0zWwPDY
2astvvWiIyg4FItmEt+lW0hdJst8z6WlHhgbk13sHIy2YmpwvIUdMDoVymfNzP66
WtG/4YNOHGLpzEQKmwevRMnBuJXS8yWCySdecmIKhmLcXzz0PBI3LWjt2oAvYjqh
2HCDytYbzaLPgGiXOpl99tlojf2dA8EkQuyGic663yk9DOY/jbvt/PellfpzuDqV
FkuuAhzZT1m5dLJoqIPfqrdRVyT1WBYd8r8sPYVAaRMzSEgp0f8f75Ex9ynRqbXm
++5CaRY/dyyZcGbUyLjdvgLXamhOhfwOyucsLZEFa6KD4Em4+naHasgriumucAUs
XlPyXbsq6gIJ1to5jvt/puqGVcpyhi6at8mvXz0UNRej9SBFr/AHdTo0+Q4X5sfT
YHIDQ2TFwciE1CaMUd4ahebNWsMLXKlS2kz+tI2Gd1qzrLuxZq2Lurn7gZAJcYVw
WUE2UVbqNhvQ60ocySN3kqqSa36E3HKgCKVCZfOIIjdsDZRjZePWUY5VtvL/905t
7YxeJU3u0uauJxwEpeqKDTIR6ZBFRPDyOuxpwGbZSANq9mQxG8/weeY8ytJJO3E3
/7lPyYxUaVMIRcZiOzU939Thr4uS58sWD4DqVNGRNmbVMDsO1I++NtremYqo/L5T
WwyVM9qyaZ6f7HL8ochhTauPelXL2ukr4JCAih5T+XGpn8HfFx6ihcKr6PI73hvf
rGtQqPH7Du+1ic4HAZujr3O35/ea4BJX5+uvh5sMliKBHN+V/A7ZWmzaj3TK2zyF
EcMuBApj69u1ajbKy//A58iOFAaOpLltbFvdTosbaDud2Tpi0/+iTzEJY3beocc7
Klnn56VqOooAEDo+RKABG9Q2UQROMp44I878mw/+Fk4n5aV4FwU8jXW27sL6hgGk
hi0w0siNTiv9Ryb1DymHv3sP5n+cO1nflECG3CbeOIUxEgnTN7lol2MQi+j3Z4+m
Jq6UL89LtuhnRTwI7pOybKWqvYCyk2/djAKuiT6s3CYv9D853Uf7DcMCrzU8hjpj
h44UiyZlVzlExea/AZCYaLeGNv2+fu/FfAUpuvG6CsmOVzqevcWpoBz4NbL3EZb/
QYAMGJgrm0eU0h3cZPxPBBss4Ib3oTFuu1Gb4BRN9559T8JD+2kvtpN39Y0UXwwY
IxfSBa/v4UMZ5jJluWAdUvQ35SpX5wEtJDC0X/B2s1AO2Ni2I35w903m9UCgo+vH
PKYy0a0ZgAZTv1W/7OXmj8MOckTkWAQ6L4XF0nNLhw/PKu8mms+yBDcDstJZD0C6
ZTG8V9RLLTlsx9rLa4kGrQKFXJ5y51pMUXZ6S1sT4D96wgSknfdlC13p8MCV3srn
AMQLdk5FT+E83TQce/Ymnl1EQEHtvdz5e31BlzUGTSiUBGRMsFYjDeBB+Dp1X531
fmaTBpYqvGjMGu3Gucvtv3JuS3VfHVpfIjwIuBfiIVmZKnrlUE54ITO8pONd3CHM
b8PTpjVE54HGr6TWRMw+Sj8KCWOcdBrm/iIZsXV486g2dIRce/u1LbJKQI4jKVFZ
QT2vivPrPRFdqtE3e4kirAVbKRMupiEajRrcbfQAU1EVUBi9Q9Od7rMPvWps9jRs
Xpp5+q486DQemW9YN98y7KP8xdJoIw0BD631im22XsTycdboQQiMuzBtXu+mCeI+
wmlxwueUh8zGfgucGu5yWvwNhlFVDEN2A5M+T2NV29XHqrQr7/N0UaSZpZGfBJYM
z+3W6otSqdAQUMv+mrOhqM9S+fjuMERSoeRYRE0oLRiZCHK2x66EcIUYk2pde0I7
zKqfYp61O7+dVDUaSg2zGoZr2HSRopd5i/1JTvwcS6rOjdPB8o/KIaFcZw71InOk
T8OL9hPy78ZeS4ZvsVlk3H0TVIa4Re18NtaZo9bRQns8Aq1fESfnAEoawogNc9RN
iufqCf2ZUhY/iqHN9u/I1JKVWaGY5Y0A0syRzWjI0vApAieKyVExkMdJcjCSZFTh
9j/WFUNR/hKR4Ikde3/G14/R8l2t4sCG+3+UxbPTuR0Xau33kzDJrYL08wstwU7v
aGvOrSicou3CPXeHQarsdnMLSeFaqTfGs25cSRU3da8XFJFGaC4WL1Bdsy+ScB5D
5vqpb6eoPXLczoKL4zZnLEWiO/ss3YQiHHGv/0/viPpuT0saFkq9HHgAmFQZiLDq
ReyQSiz0vbRPtLtT6wJL7+YyuUNks81iLwuijzjlSklVCIoHFhDhF4G71du6okul
PNegCBR2p3a2d9qecd2eVyruj7y/G8ic7k5QRuv6krXTdI58y2YfF9DQkeDuPsgB
Bpl6jlQZUXkUUEZYvwuef39oJMNFtNLM+ubagTq0S8YgsOsOdLndAdaeKBZB4A1A
ldWfg9aRafQSyZMA9LRrZC360iqtZ61KMl2XaaEid5hN04tARu+hVNGiuCPGjVP6
FKZflf7+PVeEHnmweu6tOz9CyQN80mD4QuJ/tQ9Qvz/I2bSwHsAw9PD6Xnecth7l
GnEFyxGWFZ045154p8HIJ2pU16tGD3hfc6tKlecYGmrWHIQQT3qX4Drtgz8LMrXt
v2LMf4TZiXrczfH00hl8RUSS8RPvaDNi3HskuTUfbGdOSo9IsZSDPvzZVwNSwRm3
iEFKFIoNQ3THSNNJYvRX0WMeIkarJ/m5WJlY50l2pg4WjZnmsAK0uZRnl0ABhPZL
3XiQpA+XcTEA94vGRJmsdAdHzXadkVB9J+wEnQhHVdt0u4u1J1PmnypMp1eVBsv0
eyWExUxeKywr/nCL1dRG50JCkGgwHY39VhY60k721Hmr1Sy594TRaLg1r2Ge3qq/
VO0QhoWDFQ1gp3NXZjTsFI9nJKlAz5oWuZjBx3SXKdq11gY63OQCpnIYa/AWTlLh
6E7KyOHr0yan0WyITTEViSWdWAClpl9/6OrCjPvzKYnUc6aaHGTgW83qOMwOAtHX
uyJGeRrKgWJAn14yN7DOn5ORtMF/0Y9x6yQz01NhEviAkiqdaG5RNpdJXx8sz9Cw
igmEK5iUSPEtH08x0MrOKnxzbiEXQzsSjVxsWIgM3fW/WA4gCo9wq4FvEGZeXvnz
H5jljNdwQJLOAJzZqtLaO/S8EFnG903sgEQ8q76IvzTM3WAkEQGy/dUctgt7+vwa
NXKlf0du/j8KdI/1bh+asSfnlXmpzbtVdnuTH0PyI4xacchZkFyqilSJaBo9j9sF
fdq9iC2i6RhIP/0w5dnnpRMfOacwV4ezaTAvwP/9vH0Yklj1q0hYlbc80+jRw8Ho
UrFzv6SYz8FDzYm7DKnOLvICzOF0RjhUi0c2anAJRGdrOccwSGJkzEaISnkokR+O
llqlLxBYArc/X6Vqh27Vd41sggEVY79sVb8SHFlgn2TA8KvCPiD+H9bakIW88RDU
Vw+n9ccDhBnDGbi6JeNxVZOGFWiDApJjTUqjjaRk9Om61OOQJDyuZMIMunFxYJqR
wv9AtdVrkKy0Kq0UBLUuXDuttQ8M32kiI1inOQ4Zh0dMwiUB+MLgJxTuRT276nnt
1SDCVdCyXAm/pRgCZUQfgC8x0NIrfF/5s9Y455c0sh0ZxGF7//easelCMCYpo8bv
6a64r8HLI5fy0WbrWbXoSjJTBpa8c9u4yKdQvxR5O94VUBgFJgZdR9VLYXpx07i2
aqmbhxpULM8UrlPKS7Ad0CGYlS5cK7bWoBUU3Br9Ggyuae0y4a90qJzoqHta5z1n
YVWGp5cAzzA4SL7HF2E2u0FI3a3DdW6XhNuvnI36l0rJ/QM8w8T+0A6FSUpN4KCJ
J+SZ3Jvuj1NIAc2G+16qPvU1z9QfazmFm+NmWnTHoFwV36YfHaQd7FPgtwy7QQuD
P/zLaiTJA03lFQYC8ydanRKIbM7PR9rztKklo7l9EehUxX1w3UaKMUPzSr6RB5+Y
lsjBJxpxz1D+zt9GcrSvlfWIOwEJLqFTnE98qkX7uUyk2cjZzpO5jSP2l0Jt4z91
4nVTU7ocVi0zDfQXMG5SoZLN0C+/Sv3hKID/YUKeKIokKux7qjM5kBSOw+mNUyJL
9jGNXb+EC7wLapC4zG9RYIM8P19D3pCSfKM89RlMva3RjDM3t98tflS76VCLKTnF
vj+T2JQsD/XvAjOxhAYFCpOUbfuwROu/AWyECdoPm/+5TE2XtbYcAV90Dfppm8kO
EAsEIfRwDPf5TB+c+a1tegj1fTwd0N3Mjp3J4dtUYX7ZL7PZBa1Ik8z6DiSuY2UO
WwRFzcC+gJZhYniu2OG5F092vYVtqYQahWsUNz3j6STnk+zxynBoym6ICJmnqZYr
116hYtDeTp4T1VlMYqosIT3DhE05P/6gKqwgsFxD6kKxRR1yJ8e00f9kziRV2U3+
A3Cl+n41O4rnaDDCruZbVl3Z9F1IDupqJWs/+ESSutGRPtIiZo1uuJ2ScQFRKbgd
COomnBdIw3iOa8AFfq8S+0CFSJ+5Ko/K/DNV/UfnS8YPXVQHgX5+tItZLsLKj4mf
r327RGb98449PXkVaAtICM1MnUt2gPJC88gflCMhvDDY0vHznKdK077bKORQWLF4
wan9S+O4DnVU3FYHpkAxNxwrmvIcuGG7Xj+BeRd1qVVuey3+ytNWzwvfpafPehZR
RJ/fDQAJvUQRn43mLJHqEm/feqkU5aR/20BFcKhyDRWXtN6G1QrEKJ56xDtBm/vo
jaa557Nq9uxv4XTaMno7OnVLdFtMsXvd0KJLKXXkAG2IVJq/tV5BWR6PphTvJl95
wVScTzGgdIAwY8+tZ+Idhwc573MHWzWLqKtII15Tdbibp4kJYVIGFjy3XPDLGvlB
PFUwAThB1bof1+YbBo9nkBBUXe4MlbUYtjdonWuXiFc6T66hnZIeYbmnRCEurur/
wbhfg0GkFRd6LI8TR99jT6M/IgrPA8eh7XNVgs5n7jDoBYPlWnxiRpQGz/MBBluf
/WRli+D9SVAN6QIvSqPmV4Gc71Zj+IQRiavS/8pu+HcIdxnHyX438a8MhSm3XV8L
VqvCGvlAAQP5+7usdTXDuhrtQ2iX2yg9X1SAwOuFbamxxABbPBEuOLW9O0HibalE
4q1Z3FKzyfeVkmlFAozKrPFdPyuPRu73e/VIywCDmPzkptv0F05lteYhnBpHYRZG
bunTIFLXoohrJbijYwbXgTtMhTMFtC2mtR1WeVYHLPz/2j3TSzH9vHk0vbOZFHbK
c4Xkw9AlhRnTa54cRoIrqxvvRWbE434kovVAO/PRboMfQTjQ7WsQbjS9NunE6+Il
R8/vfcm3jjMQqqbVvTu6iQm29UDIl9m44QHcTioDU7ERJ7nkutql7BaPR2OaDvqs
/tDeOpLS5khs164j7LhwymYHsfiCSGZliN184JlEL0CXISutxlSLpf1gleQW/rfW
EYpXgby+8RTLuo/c1Es0yg5CLP+ZphYVsslpWp5tMc3FgwmePot4ambNNlcphvCq
PZK6WFctD+MwyadcqaC2fNmDQHKax0VrrZjD4pEqiuwwvWfASP+7iskOlVoMXuOl
E6AP+T6HCMeWorM+awivptH3vZ3sY/T0FfNGuYtW0n238dkdX/4CnngbteagQrPn
a6yN9eMMxc/4Q6s7xA909p0RAgfhtI0QP8bnsMskU4EJw7HihYk1R2D3x1r4Ld6Y
qaatIGf++ou00IFe/NO7Ybi05nQHmY6rDs0uTumnAJ0J7sT7msk+zHGCcDci8PYK
KTrwC/eatAnFdGWqL/qbCxfX5iNdfjwUZ5GoMNLCH29+oOfNCv0DZLf8FDbTwl3N
phecRJAdTbjx/yegr+Wt17roddjH82RZm1l3vrBEKy/vRET8h88lwqkS1klzPGmY
YJdVQJGdbpleMX8yAdn3Lt+LHfZguxYvXpFDs3B2VNiVBvGO8kBnQzEM2MMPW8we
VtntD/kKaq13n6ussWv/oJA+QIsNsHVWJZJYLn0PuEzT1XTxiTgfSN5TGMF9sT2K
Crh676TEDdY/a+jvMgoy3KPhmhkTCHk3eeSE7wwAWnMVrJ5/5nZuu/dgv1nxSyoX
7f+MXZs1f5xTXuHDhWncgiinhlM1ee2Vgs7qWMfO9cnordxR7cDBxuJhaXd0G2mH
j7ACL0Ca/LpPINqwDGzwhWzu2lpfcE2txa5zHaNF9EoG14wAVfyBkcB8N9M4Jdg4
`pragma protect end_protected
