`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hPNWqETS6NGxn1+fd3GqNpA9GroTFg3/KYxpAVjDJFvjtDbeMWhXbOsEm+Bs6NBc
FP1hZlcl5td9hn0TQB2NF1qE6a6bjfmKgZkElABqgHQShTRUDUXF81whWBMMMz/j
B4hH1IrjkBg9w0q9ExbYSLV+K7cQsu8iFifyuEx5DLU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
Obo1Kz7TGSVRxx5QbIYqKlcIlRHSiSW5tH1mX4gaTetZs7HTqVQBpd65zHUM35uW
U+c77iUdWL7R5xowDBCK0ywjSL+Ye6d0EJqUtZX/d+7SF+eiKABGGGxCkhdJiEf8
yqO4md9EYUfmOu+l2CHaXDZn/sMNwhxVxmDOT9TrwIm+auV/Tzl2+Pp8QORyq2Xx
VlyNR9AidGsM30RGxMyc2FXaXn8uCT+ffnIuXQRqCBGP1MQEmhCoIRMwWTLa6MH7
hv8Cfun6i3QdA94XqSrmuo81oF9JFnafeEBxyfnlI2aTMJ21aur11AfTmT/kDhCn
EIyWFkWqgt6f0RQAbrMyPMB2nclKcT+Wydksk1vwae9mO4E/lXqxH0oSQ7aSu7Gr
88e6NIvBNxu31Gq9eY+OXRzXC5VA2iIsz9k46gnnjD6Pqpb1D610nQsJJo62aMRy
QFbiPxvMbQcIHsC9t3EZp54XPcFu+Y1PB6Rr5xUGJEnyTFnqXk4aHqc8rb5xRBxg
BM+liyavqfaGt8AG5UyTb4iIl77ZBbyWyFnxPZ6P9tzZxJtDVazCuNRHKBlR1QKa
IoHuQo5odVhPsdXjVhicC3kbkfv1Rv4FBcKDLeTszPiIyL0LEDBODSIgqmRLkYlR
t++YCJ3MRJ3I+p4x7T8NZUkBp8/T+qcoQDTUBU517uiejNgEFTucLtebKSZqTwif
Me2av0p9RHdRsgGO8TDo44CiI5uJ3E/Q/kTrR4HAzQp5gm+A0CvhBQvmCQpXknbz
wIxwby7RVncxTYMJN7/drF3knxm7GJMjhUbTZ3cqhds5ufAS87QzaWA68p1e6vMc
a2xydjMS25qLPLTtKtUXZm/1MGnrmrtwEFFFhJ1guYOht4QvaIMX/HmZTacE9kE5
Kh2hHmRMJqQ4iz3TFCG2x44ZqKnm+ljnnEZYi5thyLeg8GqbpeJlCYAxRtI76toG
jeRhsD+Cda9IKiLuQ8cXC5CMCMedK761sxdzIoeeApNp7N+s6+M+cSXaJBE5j+bM
sg8URU0TVrXoVq5/T4fnP4utTgUH/MpX88/jCtMbOMeaPEgHMeLVv9mp68glfYyZ
WYU52avpi9dAuJk0lfYVkAmN2rqQTki3HyiOLo4yQzg7lwwM+REyAHwzLo0FUzdD
QNrSWHLWhGbsaQ1o4ciFs8F0F1S4oCO/roUZUq2lylx5ycjpfPLq9a9Ps6PKWIyt
N/zIsNKBieyFbtnGJdei3C6VslfV5J5oH/BlZAbJntXCHjoXvoqRqnF2nkPX7Knf
hDQmT0UgjchxErTjPRWFy6hNJ6r7Qd5aEwW6KW8PyirbyksUfOsk8fGXMBUYlYdn
LNIg0MAQDgB29IA5vYH+lQZYGi+Wx0WMtZ0aN91K/Dytt0LHfiKeV2KfLt8+EL/d
QBPYKILFSVewIsEjD5f/t3PSxubFNoexCPXjK3NNWLVkQOvrZvW+f4NU28lcsDZo
IUuErrd+d98/noWs0XgLLJXG0cIdibr93uj1o9EBfbt4bOHoWjv9GlgMUJqj4W/K
QIkRrEfXlsqi8AiXvz+G7ouY+vt4PZ5Cblh+yiYH9/yYIFX0vYO6WcAaDZgXxEP0
E1AjcjKOri0eU+Lo789WUjpwhQaJeyLPEcjzbzcMsrRzLlMF+vmKxWlOtYjRCNeY
XcUQS7x34xNGUP9OHITIID6Npuq1EwhyTJfGDYUVxK77OqDn9CL14RxjPBwzOU9/
IOLWtsdGloLPP47pVuB3KtuwED3c2jotpUDm5nyVG2LswgqVB5mfOpO/nVP63u4A
RFLK6Ve5x0nR9djGZwVNAorEvTyr57iGeOKj3SMAKvvEYjpmiQL0FHaVnVtppd15
+NIklOXzoBHJiQyNgeuxv33b3+aETmzUVJrhcNrfrt5ZABPiBi7hmolerIaVkKM9
AQDO0eqhNeJL7/1YqmwOYSABaayudPNWxAEZMQjVtBb+TnA978W4fdNzgzoGY4ub
aXod7ZdHR99mORHtVIXzeglySNUNQ98jqzr11v4/oS9PMrjNzNrGpShZ/7fKPQfh
pPlDugO0X6h6q6oA4BKtnR5qoE8NamAGgcuiGDao88YODj0S74XIiGZXW3YwZvWI
SNi77lT+2SamvHLZoLi0AKstHaXCr5mMoz/X6YkWVjIrStU4D41vjB6hU3Jl5MC7
M157f1eFAhf2r5TvEahi++Yykl6rtpF9QxWzoB0aBRpgybyjPeYjX/ZXrKduicSH
W+gKTvFNrjFrqrbh3tt2frKBXtoSQOPBTidVDsFN9/xvpvK6uOy90SEnvVsEFZGd
t5XFhiffp8OWNpAd+1sjguOPDaAG5Q8e5aeOdAzIoaVWJMs3iOA9ECLf2X+u6+gx
/88ksv4V8U/eil2+palRYPI0wcpzA0lQKNm9HcOgs/E9OVn9K2rIl8L0Gi38/2Ve
IDTp7JI52ffY0+3uHBrknbTKHtJwltccp428uoyun8MQ10fHJYB3dqOE4XhMaDqI
Aw+a6/0UO01u770kn6Yd0fbkiryvIVrG7hv6ohY590opKpWIqsnMH2CqOpNstl+y
coppk8YfAglQlwIASsL7YBAshrtRNb+m7Y67Uvn5w7jfJlVmRfloHZu+KbMuNaWp
e+ecZZ+2atbbLPxUf+ypyfey1On3xq+Rg/idGwiGInRvLqrFYCHLY/cQ0ORcsYKk
FJZSvtMuv9L0rokhXN0w9IjhMPu1rB4ByjC5XuSwnSza3DW8qj0oxwJb0qH3zD3e
Yuo8eS2cIIqIraoBLdN4mZNbhApdAChkCBKJ+zjfT6EUbwZ9FjF6c1qT3+XRDTWQ
YuTyDzMyN9bVfKoWmChDIOPOwiAAuoNiQQz9CEeNCO8//oNQfew3voQNH05NiGx7
LQyAauiynEdy3chuUmHICVkUtMUQEiC/qgaq+i4SPsGrajwNasoga+2asJ9oFmV+
wBX7AcpRDiE/afxQnFL12yrmLCoPKA2Ji5jvsjWPs3qCXip81950Pdhvve5c7PVG
08x5Bshxml+OWGe8SawCAtJA1FdVFcLyV+D8U6qGrhLzO/bJt4U5kwCzHLc4tJ8f
QvQ8jsYHBVvwgLQDPpemTXFnebBJNp8eWsbLYSY3+0yEowwkHpKBeREVN5H53xtL
vINNvACJIi9xMpFbfj50An/0fQvy1Wb5JUAbc7vQKIe201GZvPLmrHV32Tj9sA1y
VmbwX8l8svv5IuYENq8fhWUku6bepoD7RwD8EI+QaSDYze6n0gNul58LDWdaFao8
h0g7hLZRGtedv5o9M3cPqBSuIDbtsCFgqsS51fo5sAKN4y/zOsyvQJGR3uiDd/pw
TOCFTXd5EIKZAyDB10cEKHlgjy4JQmq5FKtb/MNeeG+H3j9zCYiGiOrtnqvBen05
Y75bPjB4xIQo9IkvLv1xxn8v2ZBkCYREIQTr0AzENU1hB9YA6tzw4ZGgfg07/sW1
aaPrqgZ7IAKhASv52N4qhabY0iKY9Dr07gQjF5M3TWWheOp4VlFNUjHujpMhjNk0
U5XY+LtIlD5VUT1VScb1AaR7ggkdY+pAfqwxmwa/wMp1Ty8PvBCpADbn1rYa4RGl
FpNHZM0xfny/W2FDE2QBkpk3w5jnnrqEgPm3PHHfCxNDo3/Zuxnp7GXvkylLyxse
82TAnoDj4mrlsSECk3xDJp5u7rTHIiaKlE1Emh9E5wbw3DF2x0ewzR6NpFmMNJ8D
1krhxFMnKhv7FG1xI/TjmfgEtMjfU/UzI2THaZ1ZiizTl3IaSNqLhpaiDNv5uI1P
8uWCQyNJ9vUd8CRsLrhGd8ol2C62F0rB81TVkx7jzDMAKtraR7V/4z+5N/V9qGc3
mcbqtxxscp4GETymenK9Frin7wAn4D4Cf8YHds0hR0gLOAPiJUAl0ouUJaiLnVDf
Dk/ZoHzg8seFyk8AUU1cWGsww0EV4xZZcU9OkgxT2m5JwAZZPJYMQnrKtfVD8F8C
Lth3yAM9W5rLYoOzJEIqAIcitgZTBVM1LYw5ffmdh31VNjjNC1/WzAoRIKPZcYHF
IHn2ghvro/BG2gKcrizcm1raOW/mV2MVhDOd+/Op1vCIZyg2Nizi1bSYsO5gqPnn
SkT4/gB4N++9peIAasIHJRsdvuONPob1LWJ5wFKCDGTdRw1bD9+F9sLDIup92oH0
69smQXQyCb97ATIYrMw77sluOa8qhCZY4onHmpdQlpCr8LAGGiXrAnK7euQRxvoU
qpAtHeo5xW40RDJhMHFh+1ako/pHudJoyog6kRV2R0qrWtSUAy17qN1cTt3W2Apw
L1dfmXnaJKSRPYWv4sOllz/XIERUUfeDKLmgtwIBZvn3WW4vl8HQd0+qm6db66D8
ywhOn5Rah/lyeKqLmkSlpD71H51K71p2jR9imLB66+Y6ib1MHkypGTY7f/DAYaTp
qtg9EBOqwHblne/luKm9C53NCxq0oTsJejyA7K2sUzA4O2wbL8vF4KySlYkztNkO
pGOBERvCtXjIP4DJsBf7CvrOH32DKPCZHvxMZVtCULEPwlhPa4kxPS85GROvZXYA
pvBUPG6BClSB5+kDLiQhgKwjmkcc6kOLWQS7kTAq42Hk8JgBTIOtqNtSxRPEKiYq
q27TL/a+KA0SoiAkU4km236ww1oxHz5jMthewNRM1G/9KCKfKHdiA6z+3n1Vj1VI
U69tmKkCIuEXQFAIRB/z6idgIPb9MnNZbrqmH/+KGSt6Ie3NLZX3Zyet1Ze0wqr7
jybqmMWmwDpivRZ1fKQsddpsvQ/7FtSLk7JkKFK0vaQkSC4nUOTwlusoGAPfE/1R
3vGWbNvLMXhBRGNnLVUV2TOyzkX7LneesFMfFvMxNk5PYvV3GCDZSQI0CaThzpyi
pJeo5O7rSN1iPI8X5GIOKMS1KC3NY3WR8BeSXXCneOjEgqcRAc+cLNEDDs6Dae9r
6gwy1sGrOe9lRPISUllayT+S6YrbiPO6fOom8S+DaSAuGSoqnDoY2GBNDvAlh/VG
72ToQbj54lx48Ds6QiN6BSoR/JIjcYkM1/b1Rj3j/Zq9IwACAoYVe8fan8eIaoXx
PadxCKHBS0qtVULx5NmXfmqzlBqWD74iiJFjpQn2Xfdf7oBoLLNB4S0ArsDNVVLf
hQ2g5w77X6JhXNfjfVM03Eelt6t8D/W7dYo2bJRBUJ2DN1VGiFgGfuOqoT3Vn0nR
++8FVwrX1XthYq6YHr0c0BlsQ8B2lX3A3E8q3WLqVDo3Pdt+wJ2IihwWIb8ULY7Z
DC/7SOEJdNiX1YSuH4Q1vvix1zeVHHTg/SyhoX0KCt0myq+kB5z8nF86wdv5NIAc
ELOhz9BXnSo/k4sQHMpT8SMMhssBjKwvx6NgAv7PV+x+LkMwruJwTaEQ2ZXkYD9g
RMmwPNZ42Pn8ATFWt8CueFoh0dakQv8yPm7pOK1v7+USv2bxzUu7B8ms3mHvWvqa
0YMQ89HwxEVF8WozmWQYVAQKmUVG4qaGlrF+7mhEV3EWMtB7EZz9uYB29PyHIYLc
tSU6FkjVOrZAVtd9L5eXG614yYIqEMgTxLiA2uupH3Fkomkd07WVzMqDaGAX4eZr
bihNFPpWL97mUWgkyqLk73QqMXDe6xwnovU8u2bVLa5x6Kk7PXyqzid1G+s270gL
j3AH3LfOS8u/ofXnx0XYWbh+1L2QQjKechoU9U+2sNU4eVpo/rpxNXgX/pC+Kfot
gE8t3oC6AfrGPY5zHsSzTLXVWS5i9IEriiasGU3lRQcEv4SeAzs1QKDx/suAw9bG
OX7Oj6o97l9D1LBJZvTcX3BSc2QMuOLgMmp/UwqiDOg+Ot05dfe+dydg0NnTZPh1
VPNR0XO7fMw3LgAAOu3KRZcrQV9YwN8bZml4LjnIoMHqvQ2tiAtfC/fl7tnVt0x7
awaWmauPlmzap7OWqmWIzqzMLswAFihMS9oWToZ6l4M7HeubvrZMoBwdXSU2lIII
1pVF/F79+YXSQv7p3k70ehei6K+J2+tDBo7Pp/pWsuSqecqO5TUX/U895Pzw7igl
J6m9a9oJM7Do4jp5veS5/fT0zTBg9lE44SazF1Ftxrdok7dRPMlX8bSXrSMfytlY
jsHd1v8igQQE5sNy8MQSJ2l5rcKboP62VChV9QVcQPqCwk7AJayk4lM7nVKpTINw
R/pfJ+Rv1u9e4pyjqIbOnYWsLYQKqNFWnzG9q965mhWAbP69qD2V4k4XRWut2dVG
A5G2quLvexeCPGZoqtwhVwwpdq8+qUg9P7oltud+KwSNsOI2tByDUvdGL05GDw8I
igp5Gz2LARMGUBrvafQ1md3dGdQnZ5EGo/Hv+qk+StEJkWgWI5etmUmL22H+in3Y
GHXYd79aU99GI3RHMt/d5jeUTZ2HZuFaYXRlgYDXy75ZOrilkpPz1Q7Xxsdqrn4V
VUkcuvWq1q+wvaY7V3bH4+GOSWgG+g04uOSIWUXZ78dvlPH6+Ppe0uDOl2Jp2r75
U2phv+LVf2/2ZkK4kVfYjGgCgC3pM3YNZIkxQ4VWQWxM0x17hDhkZ45FDcda0oTP
bL79OkXwVuP+gB0kMTbQtXwTJMHh6X7YYxG8AS8OGDNZp/BcE3xjup+eIZ16u0Yd
sA61y2FG1Uy7+OfgKn0yczG93I5JKK+fr5i6xdOnnR9J0BPwInjxDLocAVdXhB8u
wDhq5LlQttN2rCQFXbALr/HnWFOdIN5Tlna/TEmyHRLHpSXVpVaKDPBIBdINERjg
+4FbIg0tbxDHEwpM6zpLRFCrqMZSsIsHFOeB0KC3qW1j79Ji6h1qMeKmkVpr/rW8
UO2EjRWoh8F642UG1yynrBqB7ys9NY77Y9FPPZikBwzCBsqyIEfrdXEtRLxhqLKF
MPLpUz7iPbzP1YU7WKXZMAS2swMNDt8CHiwHgd1Y68Dl7VyDcAez2TB8s75E9yPX
vRK80XzWX5OQA23EFo6sdmwLHh14bltfXUA62Is8RayvIlXAET0wSosr7NgSGJhW
xIX6bKmlRX9p98gHLuhH6f5DvNFqCJFot2JM1b25nBYt8qrbzaffbdUXwvYYYXn8
uEPPqPyxspJrkf1JujMzT+DUS146TNERoWyq2iy60GHGniOr78pVIEcAQGiTdktA
7uMScur76Ht6BhOz5sIAk5Y1dltoLTM/tUfLp7X8bJnDKVOEAyLvwbvdvbULfFjW
tDB4PROmP9YXc7M5blP/Rj/9vJlUHUOrFnj0hQJG8DLdXh/S0r0t124wnkIgUOHL
paJAJtBfT3KBwfURhymwT7V1+u9bylZV4jVXffSACN8yjYANVrWQAqYy4BLGKT6g
AriiQyKghx1q+R5tou1rh2CNNYdo0NJ0hme4sbEeX0X0tBAEBKspBZst2AyTWjBZ
9wiPQXnKD+5j02BiEvVGsPXzDCLZkr1bFW9oymTygnC0A8M+vJsiyWprS8a1i6gQ
OqUeMG7hrevNGxwInwgtvw==
`pragma protect end_protected
