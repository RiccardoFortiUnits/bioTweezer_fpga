// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
EnvJ6tDaMhTLRvbVlYEdxFMTLh4FoTINihIvq5S7Pk729aRxPZGwlcllv/RtcfmBAMM+tYqE83RO
MmZSO2l+7izT+/MLPite5g4/0rd85X7Gc0HK1Nu2DvSB8+iC+tFa8gIqv5AIl5/gt1svwHbB9znJ
bTbjplrE+08rSZKFjtCb7kcMvYklWMfjZh5vxXqzDcjASv6GsioPED8lr0DzfdbvLXPoCyppNrdr
+ES3vkobJcYiJqICjw28WnXIP72UONc1We6OCu0QnPCWYsnrksuZlOlz/iqofJeoPRxmvjJl/Ewn
yLiyYUkS4vu6kAX6AoSNHMi6+VDSxrABdGPUXQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24432)
bClk/uRMQ5Pa32EzlOgIXqcE8i6I4JqQbA+sAcqSRlHe5tcJVYT1hK+Silh45OWuBlCaFZ7+sD/O
P3jxBM9ZNzn353iHk6bnISNUdcwpf3eLnpNC97KfvX56X+oqM4VwlaN+VRWkHX528uXiz0A4X82R
Y6lMLQmxw/kxFqtgIcSWUA2KS1bjzhQqWMWZqzRZVPx+ZqVNuC8ieAITmi/+vWE29EPpFDZaMNOv
EQjN3sc4I61tvQyxMTJMhWS05JrDhH9zKksEmivbEFmaAVKvqhIAHSZyKOopMimlLvWJzfEkiRA3
Ie3+jgvvZlC0kG41ES/OpY+ofLRUj9D3TxB66/Yi3d9GfDPzlKKqtY2XweChGJS3m0GRvIBAZkgN
3cJqYBXvv1OtllsOsTicRhBA/0/GjXppsPhCIrcXjegOY1bRMN4c1Rnzu/Wl9PIqSn4afmNRNe3V
E3ckW4fRZSDjGXeYciVBbQGoPl/80z439mtJuExS2HzqKFzgFHncD/VQnc3JTV7HY26r/8RpvakY
+4V3Wm6i/fsvMbdt6blMoTc7CJOBSwA0M/F/vzBvVw8jPaQdypx38G2NYtjGXg2it805fOiL7I2V
Ha0DgxMBYIl1joxtXdRpGovzxs+GpF9EL00Si/znjj4JQuExlftmk0wZbBQD5rVm/NozsJIEgGTL
yMnrz29UxyKX0h5xGM2fWBjr4aO/n4of8rQ+XxzQtEn0j28GsJxIzonPz/yIVBhLG3BDDezrMOtQ
Ccn5Wv3zZw4Lic/zAusgyQmGbEPgSgsRrzN6961Uz4ZBxSAK3Ki+mrd32y070GNItjb23M7IbWV3
Q4Hbn6JhgQgDOjXaHQIyiQwOPgGAu3NBY6kEsx/xRNBwXniEcaM21PFAswxu8WLshwvHcT/TZzgz
sCYr6oKniHw8DKzENMXuMRxARoHkrihp1OcUAv0ICYt29YR870xilNht93Dqb7clyQnu5fHvHLbM
p8eS7LjeeWFI6Nbl22ivy/oqqjQTBTC0flNpk2RrfQTQLHbVy1xCGtvQuURtbz+kzNWOZKUKLxDa
z9wwHOxJKCcls9+Ofx+etc9AFK95HMzit/WL5ajhu7af14fEfQFGu9I27+n/xDjqUGdzbWEYb+xp
gJ5wtXfG7XfPqL0sat6r2hKb0xff39iCTnq1G9qd26ljlvEOEoQAHiid4klLu14q9TN7Dj1Ob+GT
W6UqfOpIYoMIP+hZC7OqW81M1Of9WCiAhQhhyequ7LI3ci4cUYDKvWiHvwd6863JzTUxZrHRg6C/
UKw+YNL91OPBFY2oWdza9QdP1ETBqYylPZZ+65fHNlwVYRemN27JYISfSLiFIqQNQjPAXE2FJkIk
Nk/G73OKTkDhDolWON6R1V0ve9n3usqkO55bnJD4pTC9xCsuFDNIjyF5gHSJyO/arG6TelKVV7F7
FXBtMOtbnkoMwpJIPMdXjhX7OuSCFI7g9jrQ/k5ckBmyvsZAw1eXvfrB6c6LaAlhPUyBMor6kWfp
oNBKQ72FupvlSLbnr/VGO5R8/GgAEYxZsrgbZUZMyiU9Vm2jq5RZlTtNLROyQgw78j5nQa7kmW8y
P4ZrVrCsT/ixU5UfxwXUpAXIs5+IeQW8fgBMLzjDjfyAxrUyAOl59ZXy4pmuTFM65V6PKLY7MxZ/
hRJh3exa/C+i3iQaX1xgERgI+e2qXmxiWhwsJltarTAzdbO/gOGpalfjzNDzAbQShE/aPtch2FZX
nzttp44/lKYqXhApPDfE0a8NU0nAeBzOAN8+9xc9QTLMG76pc3YYC2/hlM06ITMowm6vMPb7aJOU
tp1b+nqrntsOi6cGSvX2+BQmteO1yUK4ddmIxy4JGEcPpHrfbylDutPiNIZesRHiuBpPhr3tLH/p
lRZcmU4slXfdrINoUla64CBZ5DzLBXFGzMNAmMxi6LQE0T6CigkpnQ37WA46DYYAXW2bvk5ODZ7q
1HAwaM4J+Pkjzyfns4m/cnQLYEzK5/e0eFBgFlHqMbqFNTJNXALXO6Q8Cne28aCnRefY0ZWrTjo0
Ju//Ft5bEw5gwkMV7sXHWbXH8pA4FEjtuf0MWihb+f2n9GO/MZvwsIaE9865p385DSCaWuthOfWN
def1gNWRsu9SVkeMh35lY+Wb7VVYUUey1Waad6sgdk467qc/XKzOf9T3geRwzri+3odPql1SHG9H
oZSG3Zvl4Jd9+EW8lUDorxsY9QAEHdSw5kYk9QizerwL+7LN8/1T9i+lpQolLJTt5ba7FNpLD6/K
rSKDaUike6RHqYUm5pZUS5ZNsLbeh1k/67ADiu3PMro0RoWUOEtpP0LplTOtlvj2LAeMfaSyAat4
kqj5IYOj0wYSJYo1NOJT/TVbuBg678sa81qXb12xvYyQvJUn5Hi1jFJVnuGC6RuxWjw/IGln+PGV
liVEEuUlJSnmcN6CF03pweGq0vzcBjZ+ERRWUuonVh5ognSQnLUV8qP/n2pVGR5oBauoGEytUU4S
MlAhCLLy8sdqnOq8ikLZImYyLr64AA4622aIk7EfXhSbIQsMpupEcf7ifKbw1mrMePxIOT/RBS4o
pE2mTyYRnoHGwkfOyQpd7dRipweu4p0s/BMGDUSR77rvnafJWThdSXxW3XAgmvFAWUosUSajnQCX
i7XbmIzlYwMoLq0IOsTDsYU+6t/mGeojzWE8+B3ijlVXJLk8wd7Rj6FQuy+NXE/5sUeVReuXVWar
8YxNwmxI+3DOmW2koxhlSaD2YnvGumj/0UrVJtgKIu4DeG5hNjrGTwCYETF1/8eMBpeNdOezEiN+
i1oYUm6cVVu2aggVT0fYHF534ZhSXTF26a+ot0jKNsfrZ3c9hJvK2Khh30mzTmT4le0eHgRtoTkX
lVEtL/KB2AY5GDz57FBkRKs4Qpc44VmLmots7n3xQWU/q8cwcaDDaD5IfQGNADBn9ZidnUCGaHSG
R6r/Puy91hFr3/CwSrlSW7fc3Ei2ECFG7B2NRCIp5l7QFUt6RbrS6Z0AcsQVxf7JZAGFnhIUJyx3
2fyxtLc7kqbyHnzQWce+K09n9mqcQdH/l3mFFYGmGizaFkfIQ8Jkrnu6lcCsWeo+jm+BeVqtUXD0
zPPh3TUbMt02b5A7zQtJpTftt/49psG5d4CtjK0sDe04CasXqELMEliQUzRe5Af+KoHi3v6bmNZJ
ttkn5Z7gK/IMRkT3zNo9azLuthRI+3Xer9Bwb7vhR0NGJQ/nFklqfs5pKr9lF/k2Pwz1fbPbEm6z
t4FWNVIv13g/j/T1XWFEbQ+EdjfzkIGh73GTDv/NlT52I8qcp3KVBrmpL4R1CX6/WKVJCpDe1Al7
oaAwEPXr2eZaRcXevTv/W+RVrztqMn61Bbos0lCXBTEpr5MBSrUKEwKQd6D37LWC8U7GM7aGAUrq
OwlXtlHEgLyLMuJU7WJArJz/1fiSdRcvnwDZzNguTdGLS7EiPi7C8cDrgtIA83UxrG5amoVs4i3D
aWeTMQPIP6tLWjMEEO5krprqvoc0xVC2Nf4gsWOSPoq8gZTnMQszlzVPq32CK+EpriWrQNK1HNiI
zLXm5DZ17dL8y27tx2kbwm+LpEqXqYrNuFg0mdcau5t/KGEKYu+JpG1nRmrnt0MSBEKuiYdiT1Ed
R4hAlOlmlsPiG8y9G54MlCbj5M42FoQhmkjJ0k1b97ojggm9o3G5n6++tMIS4Fd3xylNXB1zSeH3
qFMP/epD+rywMBkxV3G+6BJ7XthvWdCGjPbeWeDyM67kNusUEqhgmBLs6tjsJ9RmHv0R4vDx6jek
UaJl1RkbEo0XiVlA6io3ALsXLIKq7Tl5hTf0YH5Bk4XjYhbRNOM4TuGTKMuOEpnkIsU++XZPx8gv
aUSXcy0jNE2LsxhR31bH6WRS67FZqBDwTM3W6gETqt9hP8gSnK4R9tL6ccS6MCgdtTo6Ye66pNJ8
WhTOIy1e5YQF7uBVRlgb/EVkA15MZODvlNK+pSNgsXD0hmgATHdA3g6fRKtdmGcBfDNHfRgvJkEH
JRZhAMPJQH8N3L0IWUA/gKbht/tE5U+2TH+2PkILrE9sEfuqNwP8JFOrLncS5/J08IyooNU96qDd
JwlbQA0Z7iQjdVmVF2qVKDCPSpOwRx0J8RAWodh8LLD7BYlYLad24k38wooys5IrLka+gKTBeuid
1JfdFBcJeNMDr5p54XssiesnMso8o4JDR7PaUXDREhbLgtnhHviWY32eKC7cG9jq85qLqz7wYzpU
puVbwNvQuIev1FyO7hwIBFmZcXcBx16rAIkwbtanryAkjh18xvJIeirpJXTXSKaj9hwAynC1BEaX
Swp5UfCp5SOHZ8JaKrIHjXnAGiWilzECSOy9gICVFSQ5TBtIyew7FByQQTBXRPbGa6X2Tn81Au/X
gWQDx3F4/NDjr/hwIS1p/2s/ZA8TEP95k+n8/f0fEYVWBzVrp5WYTc4BnNgfW2vma9+ZGszeiNtK
4UbpBvoMofyf/XlsSpfj3JHJSDD0hcIE9p3kgNayeahAFOM0holnV1HoLvXcVgoQesIscb5e2Wsg
VZ4Vrmf8WyUL1r8gsF1ums1MkY7hGc/i8Q65la/L72tgxnJPn7u9Seb4YQrKgAEnaVY360VoFFsq
lBUMtFGPPDzVAiotV/2ddA5hF9jsLjw4C7+kvdkneKPCTSUUQnXWbHHnJxLPt5JxQS0SO1w5ct+p
CsRACiEsQ54UZpoX6XFJsnpCPtjI/PCFVnUV8Ynm503m8ahdlpHLkD0KxWfsfSduGhLT4dwYLzoW
YJNAs1BshuRcAejwQUVwQjN3U2cX4C4teNvylOKX2k7Llb3kz+LpyqE+vmHi8OOCigaZ7J51PfCN
O/oNCreMrffGvXM61ALh4DMa26SMN7scQysKib2f4n/zGtYScYMk6MQDio14dV4WKFe98C1XaCbP
3rOOMesN9R3oj9AeiM6+qBIPYI+F78rLF9dzZgmudMC7caAmPFJPPyqZFIgbBcxB+XS+xO40a/2q
m/l4nrABBLOVOu3qFowfBcnVNv5MMYaLXBpUZ1mMyYA8oLxFXw9+HUHhHbtEaRL/MeKqIogIfFHb
sp4wjSQtEH5BYTJ4p2XBmjPE+kW9dtykWT3knGZVNfGPywrVLcfO61a02ZY2r8riO5Qn1zj3fOMr
XUl127wmMwrsuFB7K9FheDB1WPmLKDbZTsjwJVHQxLLPCo9wTpSX+gaDoqUn7JqlQEKz5tKMx1YW
FauoN0O1lLiAmjfRKxpdAyntPwHMULbhuFhK0Fwgx8brhRj9HmrSn5M8r7xDQlhEB3HTFbVYJFw6
WF0L272YYbqRH4Fjl5ak60Zy/0nE2MS4IptzG4/SnNRKy4teLvSDfHJBPxs408YlLILBJblf+k82
3Yfinqs/sxVaIRox6/L35qa87brpNIKuwP2DvfMB49nscH/R90xBhzgJWHAzLW6/UnM5Y5GBhU3F
tlpyNtD2eORSECxMNGMiPwjiA2vTWZJdEEDZdcwEsbXXKojOkjyiKTeL6deYJsRT8twxhyEwzHRk
Kzs6sA98KZJ0GkUXZCJS5M57OSevwYvf2wveGCtxwDUoNnLRJrVbyD/jN6AokQl+jfNzvgML3lK8
nk1WCXIG76gN+UzvSBSIYq/R4ggylJFIzChXPZU9NnEG4k91bmC5xjE3RHdUqp4nYuazfuTQlMl7
qXyclF0MOwzqbodEttRmTQZWywyhDKY3rlUkRVl1x4h3d2ZffwM34ovAs0efUlVdH7cjqFB3a6nv
bSSF6YE3R27OcDiwm8rf7YuM+omMb5Syrm1ve848r/RAuB7zbQctT8AprPufurPvPbP4O/b89tsY
JfCiJhcgeW/1zraGa0C9DpIQxuOgaTQV7AG1vfiPC0GdOk/ofIFY7ew/gGqak0bB9a5R2E3wB0RB
VmvGdmnt7TwCERhZMzHw/3o5CyGJYMrbXFt06S6skX1OiFIYlnJauDECqUQWkaHXjpiYRxmkfYOK
68tGNvhDshcmKlrmTClOmbSyHyEWuAERzCo6dSfytwjLaF4ImSQZmGXcxswvWO2s90IMvQHGYo2Q
45jwcss5im3Lh+svOvmR17JFyjZkKkWZB1/D2MrElGfH1HfR21cM+JE2YgEXZGIttywAijpfuiQz
1ampWPGVRcZS0zGZ81tr7FX0LM+78dNx3rFGWk3ZBRxweSMaUyryXjKUYgtTFvbOKDlSPfZfQOMG
CX3j3ya9f22VJeTsH8OUKSGtwr0msI0ShojQwcZWrP7ZEM/Yq4ksDzVOYD7AK6zJl62qLAo0NxI3
FFFs4VKqfC8aa+huM/8HZniDuheV69P7Ucbpjf94UyzMoapmwk7bZYOYA1HeaKZKETwia9q8gYTo
K+KoRMxOLtXSSXpHMtokHx3Hh0WsdXTa4mMaLXUl0HQ996ALlQAOlKNW1y/WVPDgrZ+RIwAbpcY1
MPTGR6xOmzwcrhTPPfUHHh7I3hSqsELMoc6cCTheztypbG7+oQN1Ro+knqrbMSugXLL40CGoCNGE
JvHtynAldoaEsPXFzJqdqU/1iy4sy1RNGnfEEj5ilaRiDn9CLuandfF3HFpGeuVLCZl+0xCVvBRI
qpcvFwie+j1eSmfzIF5VHugIDpupl64CwsWG0ntwfm+W+63ianfRyxojv6el+K7wLrExgEeEWqFG
c0N4DB+9LyNKk0d+kn6HYa9xqDXSVbbuVEgN7C/HAjG+F4NNTPuPhGj6ww2cMRyixU2kbmgx9TDa
gic5zxrZka0UnZjWLQs2olLA8/XBjgMUjrjTpXMuY5OzSYurZaJPJ3+ATy/F2MUkhCEgNYzbqw0t
ADk+VQSCoSPgloxqGF+wkq4WiopDbjF1kF+xQD9XJQCNgftaB3br9Qis91waQyU+8Qdl4dAcdIvq
bn7Sh2Xo6xR9OFBsNI1hyxtvvWeT2MkUS9Q9rbn39RKoROFcD+fHDppnQ1In/KX/iVEEG3FTlDhn
lPlwc3WivgBWD6LIYiI7brrHLMBhdjidL/7aeas9nJ+sEPac2eBJGM4gkSJC7racZ3L2IlrtAFm2
2ad3mr6BY7gbTkuAbUM7aZukmPgT8Ayhfzy3QGy5YNYqBZuL5Jj0xOKIhBwUh2YLJ1pXbiexHjdM
pOrdMqxphbYk7SJisHeuP5vO56drhaKMF3BSjc1+l0fxH4iOz2DphfR2uYFyqGbC4fxPzEiRbAxC
QRjkDEhlDt3dEk76tYtVMsl48o8xgU7IPuv7G4ntjK1Th0M712dwSIQ4Iocb5kfFYzigdQwaHW7A
rcRV2scFIQ/kZlcRgvD6sOEFiR+Xhga2oQoNk35vXrPh9n7opKhgw8htOpqc3JMQXQjl4kPShqv/
qltiKPsaRzD8DXdgk6tW+gBxdLnRXF+C4gqRykOK/DfKVmF4uZGLusGGfVN0ld8bD9QDeUWEJOG9
N28lOTMelORWq39rTw+47PSXE2XKlwzYf1JJTUZVV9Fxm1VGJrwkPQzrEVyTOY/zt1VNNwhq4Nz8
b3tk9aXEHxDJCI9Ndc2S1JiwmU7urFngXBFjMiLfHMgomERUUwsY9PQbdR9VimRQq3xdqQcUkC/X
SkxcAYJRIUPOnekPN+mvqcD2LNBsdzxele569G95wT9dXpGOVkxFLhymx4I5S9mSqjRKtOAc3Fja
NAjixqfiiPx8FWZ8KA/3oBFRQ99U/bib3/vlbzTybsS5+JRI9rVkaRSxqUICCOIQZ7p6keoyznU6
8SeuVQhKJ/9vCC9EyLxybLHYFHhKr4TNhYmv7vzHNuDT0TjPymw3SJh1CEXIqJnbjJ5D1nG8Wm4l
ACxmjWne7VA6eJw5CqnbfxYn6M2w3GGWDwTEnVXBmZnWrurJLj0DxuNE2n6sNmQyyX7D8CExCIS7
am1/+NKeI+jkjs8uBSZm1kFzS/uXn8AvC580s4MBSDwMo+eOVozaQDuzWDXfK12F+DNE8x5CegOP
L0rbtl05efPi10XZp5OyoX4Lm7ZXlvcMpTwKeT21TMP1CCbCyJZS/+wnjt9Jw80O6GNBapL3rfi+
pVqMtVYsHBED87I7ov0ra3CNO7DxeTPKz1Oj9Vsj35USJpVpiHiuzwOmom9ZOv4cXm7bh/RzPrQL
9d+UIl3L7GBfFoefE+CXiHk4/HBL5RcLZpiNNl0pu0AYpVAITJKb8QmQXRso8uam3XUPxQS0M3D5
WeyWCBVzxVpe7BB4JvHXqZEp8yaW0FEnkHSi2/zFBU2A1ojh0qJk3BSbcO1bJ1c07Fg4x9JHdwXW
JJqM5Uql/plt+O+sSzKycC2fmr839FlxrCMOVBnQziP3U7xm1B/ZUQaNNgh9AmXmOfuG4AUkOpZG
3GbiTg3zPK2irjCE7Oj2OwoCUwcZH1JdwnhZK6bZDQmHLHZPf+JfvrruKyu2Xx9eiA55OKjjXGW5
14NbXMXCup0ibymPCZv/BCFsnObhksIDXtd93ejSVzHf9edodWhUsSkRgxDRCMGJbN+wABausis/
G13NyZlqFw2iDI9BcZm0weXPQ563A/4eZQcPo9y4hCop2N5nh2k4kPMpGkO2mevfqgRBAsBp8xB2
12CqRncjlb81+ucp0bi3vsQp2V1hbFxtZF48sto4i7AYvBmEU4KWM87+g1BHZOH68iDGwP+v0oYR
4sDdOOm+GczpO4evXg9uyuNY3PSRKhdb7zmdqJfh968Oioxx9RZwUl8aA8kE1jH6KO2ywzD0Xgmh
V2qOFaUjhRoA9lCcjdFHYjvXDn/nzvbfiwCt7UV3cjJTLZUjvbseIHinKXKCNpMVrpOgEoc9DPF+
rcVrqEkn2lAi73TWW9a64QJDPOJZx1LfoZ8oSXt/ELg6S13bK+NQOH1QwOvkRnMddi9brtrlu1Vu
hfeg6s58xUQnFBytjx3NgPOvcz/5/S5vFVc5+Uvvhm27uKIoJmE/yjDwmLpIgODr+BGuXa8qlmW/
v7MtYvNVizPVpeiTVL6tc62Un5rRpKcgZ1pfDVyd9+WxnS5zUhHpIUSl/F5IAsOHoCQuS8+xWWpd
DxWpeiyO3SEKcnSaa4npq1eSc4BVKPX27BO4NF9oRiQux0dLP6QhYtVwVroW+6vEoEg467iy1XS5
Hpdr/FnK9SuNjOcDaAb0l3g6sdraDBg7uE+U1W9exzHwFfUhwPB3GkBTRl7nQtEu2w9mqD6AbJrc
OIre1Z1Df7sCZqm+r4egFOFdeHbgVJOu9sQo2ps0bD17gQO4xaYK4iveXzCVFDb8OwIG70/boF70
wQtVp1Vs4RMXCFUBjxoib4VoOY6Go/V4Extk6Yn25Dwq86wThNV028XYIZUT3TdJTQDn7H2StXkO
557TDLxcxdo8AZToyX5kanQQADdhcQvpPAr+0wM72WYyAJAbUKd12rGRtoiW51dtpj1ujsoRyF61
zsJ07mErjKe0J1ZLomPX92jl9riUdtxo0Gj1W2uZCvqrwonvkXll8mkJLzFEMOWmnOZ4B3sEzdcA
X0yO0y6Q9+3/SPNiEoe/TmQ3sNl+fe+Z6dZqhuLzVG+GTyczgqX0egaQMoARAyjsGdT1FW/wgKHV
rdKPTMbqE5h9LKkcDaYvIYNQuxLFmPy6+v6MFmtSHziCwrgfdg0cJACYxo9WjtCUiRgw3B1w+tyl
38PiI3L9SNynKrsUy21xf5D/CzCwjvSEkWZCA+POSIfaA/Vd/fnMkGCIZ9GKv9xS6cUVLNjzDxgV
ZV6cPiK3s5x+0UAHZ2pu4CZdfHEu2c+KxxqRcKlArC+MXvO56Lo489h8YN7sldRw/OtXk83EAltF
TJ00CHUQeog0lp5XaT6KKxtR9t/eG4T4R5aoDsSDqR01NMm8r0Z5u5uVGwYBdtZUimWWz67/0TKX
mJ5S7MQc1NGRm8KFsdO5zOAZIibZfYKr2aT4nxoK64eYii6EWj7tIOgP7stT84CRAFXnwUF60SKG
u68UKO9zGftUsQvW0uv2w3yTwQIPCZy4l+igzqzB79wFuBS7/m6C5yk2q/9TDcyB79LlNoZo/YAV
TuzXdEI+YrKSe6BaQIEzdMEHxMyBjPdHzGY0GSpMC65qjKxSea2bJo6YqRkaqUi7SJ4sTgtlAhrF
Vf8C4IeP2MfOSU//77DC3L6gzNtfIKKorUGHy7KeM2zmU2RuhbbrxChDKVna19UC+AhO3trVm8xP
1yDk6Sf3vS1Y1bUjHphP7tapaXd5IrCVb78+w90HuspxB1xM4X6qz0jjrNf+41UQFuYgGu9VG6Ag
AQ2e2oFSGTbyBNnWKsbGwu9qTCMJVG4tBrEqA7fSou51FEZmE6aE24pxDJgwxDBSLEYFvjw6uVWD
N2eua8jJpL8Ev1JITrGd1sZwhpRBzc6FDxE9afKKrMdwlkyXqaASlMG5kgiUAGPugHPX1FZamp90
JWG52BYoTpwicGGNoa9O9rAwuW9ZXNf0ADbA/jWeu9Vm2JrGubPZBtlDD3rDYo4CFeasXASWadfg
qUFPxnx4/DRQUShwQjLHdT/aEdOq6gBXYm2IMx4lxu6bInVsxU/S7iDlWYA9zcLcIWQVSBBWnk6X
UrdBu5GQXLPwKnYnF77/+LIIFpROpgLwFv7LCb4yXOGLIeSXU9+LG3+Hl2zgL2qLYJrjzgHVjDCv
kIPnrrxzzQI7QQfrQ8Wthped5+LGeyCFe2WiIqZbtZdlXS09sKoFpTbN3MnC/iyz4fgGuWNHjqKe
RO/VUE6+bWPEtS8PUsviShAdjOXcJR+J+errGfuO2nh9CyoOoXk6seXn1x7cYyDAMjRJeCK/W7qb
gm5+9vWovHUJrAzwSNJjxdenWqmypR+nNDYcKGPwRNyb82uXmusP7DVq3lyOWPIw+l/xHAlZqbDg
Z/wMuQL74M9m3YvPQAPcFH3IfSJg91cuS2emgFxdbWjt2+gUsdpruBxW9P+bLkcN54LNZgYsGZp5
Rps+ordd2dREjlQnJwIXkZK4KS/x7qZ6SAM1YGNBncvYco2upjltp+ZpV+mXk2xcPRI7teoZ3p4F
Vz9r85nhvJ3lrb2vfmdx/PsynUXkEv1/lVa75MQVX0CqQNMO/FMHakokP3c3QyKsJQXTDunEvO6N
40J/7OmFnDXqG8+B/zOE9UpZd/040OwSp5zw8XbXpf30G1LD0OXdroroJQspfnm7BjKnCJ5ZS7PI
iOE30wAvgdgqiE6yDG2UhUnPz8QQJRt3GO4LmgvBKDjaBV+EgMX0j7upbO2k5gCUE+mcCoOxOM46
TZjIUa+dQjo4rVyaww3wPfq3STfYzbpWnvTGqUVqjV/FKvRtVcMc0KBsAorXE5AT+186S/8hTdpV
G9vRRwh4dF4kPkXk8d46BQqfc/zar8qctbv7cDKxrJBQWfXY811eET5iAqQFSc0qxChComce8gFH
GtPDf6EG91OOg6QPCy7u6fUsn5UpnSbwDlrEOOXzpG5PKBrYtR3u6kmcE8eVe1rATg0+mv45a4QG
tSjfebfDjj53faGjNCO1jStjcdBdG2/LzdxaejVOGECQ1OpfMi0QaYP+WguILNo2oNXwzpEw7AWz
9YrzhSks43hIfp/eOIUuZ/tzdrCkXBd/aroKczbz/PS4VCNRiDdRTE2KIufmLujiB/T3UpGDDScC
bsKbGJKnys9Pkbw2HTXh6ilsge3ARMuPrzZv4mXpM8KdWTa5bHUpieyKqr7cu/3jZvP3CkkJD//D
xk4xWPAGeuODhBjwB3MdiA8jMd6tsVWLXinCqZzfeeBk2rZJ8fMGOJo6T4oqT477YaI34pGjITpL
62xQQbU9UQMZ1ZlmgaCJKCjkzjVxpobqNRkFiC9WuDMvZvEZeYrY4dhi+9DGA3IjLqZhraMW9D4g
+eQ3cERpMZempjdq/0KNWfpnv7xBv0+/2HT0A+wqRdoeeKSWRfYeKi0maRfEKH5W0T+ntxu69Tuq
E9Vz19tOEmeqKezDM1LsX7nsvPkOLirWcf9T1rW11HzMkuleHKBkT39ZPJbrF3kkc/tmEkOXunHU
yugyOBKzTOkqrQtFxL+iVL/G2QZsks3PvAKfsfY0kBA73CD2MoEGhF/SOb42azgsU+OvWmMhYGvt
HbaxB0+sA1Pv+5vGel6UNKQHrDXfIoM2ZPudxM04/ogdUD8tueg/k0AtDnkkxmJXxdaPB1uiJcxO
Fjowv2ZxJbm3atL2si/rzxq7am8yotXFRgXfr9YkU8wnXu/ExZsvD3Jkmsyz2yudC0QOzv7E2Osh
Sn/0pm5Fmz9uMKKP2DHd02sLVD51/pZY2/zApsPJYy8XyHzrCezU+ucbFaSI/F63JB79uQlg31IF
dqCWxmOUENHl9/BVWkSCkjDzlpIrrH2UZm6FZA7eaEPzQToV35Eop2wUwYAkHQT41jB3G/irh4fN
8KuUzc3Wb9lmzl8FtplYx5NnRvtCIE8CWESedcnxBLoP8qr1Z8Xx8cf7XBTSC2KTIk1hrkH/MTTF
2hl4dqwAyIsURbfQYU2K82u6oEtEMdbY4xbWOhyds4dAAPcx2wFtcICRDFWsHLngMH6soLVVfi8a
RcfzAtGqrWFxYALKbk0p8aXVlijTLSr5IAsVkA/fXQVEmFleFpHJCVglj49pfNLGuHYBoRTs5fih
9/jfCQ6FQyiEpMBNd7G8p6KXQIKxztkMPfLWq6mPwKFqQIm5k9pZDAWeTSf24o+KJTdCvE3bKvpN
Tf00C/sEd1OmYabcyR4TAZ1kX0tcptn93dHNCuzoZedji7FcuFFd714Jp3EvdFDZEzr/Unxsa2Y/
shc7ISMVIf2nLeE5ypSp0HdvxlWpRWTiUPTy8akAuSvriAvKUo0RF3mq7nmvRcAjDGADateqa8dt
RBeUjfaH/8fVnPEYZizuQvneqDj9u6yMaAqM5Q3f4WUY2BdvTvmeaDMKzFNM0dHiaa9CeVh/pQme
aDy19iq52ssjFUXcmwlfq7G6ksffnYrZiD0BlLDnOAt7AuiMuio0g2xHKkjq9E+hg8Qq3xDy2Fdo
Vc9v05ESOHOI5zmnQoOinGiYNK86faBpCKFUcVtHAS1qTyoHeoeoaSFiTxr5rEJAb4aeoYPEAEpN
TnEzgWyyGMawFWM/Zzne8UOcPYNycsX2q2xz3/j8SOzlrwCpcaCSAancFCCL4QT2wf1HseBovPNN
d2iAXEY9YgDBTZS4MPiKQG3162AVgO3N0jYOy2jwN4xtMGZp42uVm9dFPGlNMW3X7Xlwml4cBkDX
IHBB58JfOq5PqT1hEIdw8Ih3ywjRi96yPnSdFRI9Cu1JHRs4xznbVTZjqzoO8wVdU25PxI7fHRt7
YlBvOgtf/ZBXU3afWl3gKUFEAYCvtygCjr4ZHATDE44ua3N7iqiZSXZ2JNaEQtanjedl8iH7czrE
sHrsakVI/Ks5ctvbxwOun0JvjkCyKHUjN6TKvvDlUDl/oovGur/R9Y9tx5n05pcuzORCGJIpKH/p
Hgbn6k++UFCP8p/jY4gycUFpJWw+BAgJXn26TfaVfPi5X7ZCTRfYEmDjW66/jWi+CnBpEM548fZx
7mvymlszmn4dRKmlMFifnf7jpIEHi9t74MjHGc4P21VxtVphz6msItxmQptQGPxzo1CbsOJExUPc
8qUZEQXceG5J6NOLONFz2UbQpSzmGij8VB8TuFOPA2G3mFMGecArPlITm5/EB3yXpWH3CnI5OM5o
ZO00AWaVDBFDzqVZwLFpU68L288f2ge5dqwBFtg0ESBn6SFFbCySQDXKpdLyNZiVX1HyXc/fzp65
p2mffDPkfd9UA/Ufr8NT1uVGTtUpRg/YDGZzyTQFiT1j/3hZe3j0rhY0yTBFWeRA4N9qRXe/WrK8
ibnJHQYmS1I+ujLWRnINZuM7HOTq6jXnEY9cqRgXCuBxfmqyCYgHuFsDTRZmLtcYwbGP2Z3ge9ri
hrapsZj2qSG4T7Wl8L3v2WiI098hVZgdkMQWi81v5KLwSbUCQbCYWMaGWkULmxSgSSZXRzme2oHr
/9uuzSDS/qSOve5qbgRdkKDh8cLHcPFcjT0dRgiizIizLBRX9y0x+pNsnlHs1RahTterBhFBR02W
1GU6/U4meCb7WrrKUe34933L9RQlfNF30Cc8DrIB2XplyomQBfWVT79tECMGW8DJc/mML+Ww3ljY
D37lZkYXF+lZS0YjMdlrXDeS2q61kn7cHgT/rTfE1YOsYaDtxNZzfRUd+airzsuDKYTzuRCJbSgv
l14cHoOlrrLCUiGQU5T7rIN4SoSmcUd7+an/8+4g7GTKq0XEeHJ/N0Y1xSFgjzOpZQ8YOm2ceI2Y
9dVhSpix4GA01f1dFpp+VBaAotlgTlCXEcEws+VrPsnNrQ9j79XYLdcI3y30p58lRH+yas8kvfs5
Ktk1U0SyrB+PahBaGAmeR+aTfcFQ79ZOgW5/oXABSukXozOlj2PSPijdKZWNiJbH7705fVdtBAoV
UCgorRWJqgg4Zao2ekXKgu/S5Ue2IdnMNDYyjDjnB4PiuVqfL7BIqsF6rMIC5cVa1YohdXlSkC60
UBA1gU4PbtnGXfAr+4HXxaXN14KPLD1U6U0Qohn0b5pQxQTMbgXCNI8rC9nKrhAraklk4Ulhl7WQ
VWPGHHbbCjr7FYBPSMzsHo+MjlVZ69LBy3lndFSqsbJVq+RhAjd2yy/3iqb5BUJagHsK6wBdBvbj
cJgLSa2PU9d7sSU8srpcU7abIvbF/8ODz+NJcarGuhzYsa1qIRgiD5gZq8+AIeibz+XxRC/jdgjD
BgRuMPkT4XXbvQJ1fl7StKy2geqEG03s+TgQbBg8PL0aE9oB01K8hNswLyhPpzDAE/Ha9/1+T5qQ
Avlik3FwlV47kKKFdhzG6f/oSIZM8zO1HCMNQuWOhtVpJFZKSluzX5HuJKN8AZsoqIXbMEjQukVA
zlOFRa9z2p80Tf5Oc07SmrZilnxpDGlVYB2qHHjfYk8IrpxmvXOmkKuOQKl3DNKJvQg+S7hDPsTi
PBovimafnYtMChKJtKDZammpdYvY0mDzu1jKNXKcspfLXWttbUqz6AB4TNHTYxIY6PPfkQ5UjoNK
gQJIv528qEFxtmpMRVK9jpYiSWAzVe61lo6OEcOSFlDYBQX1ujJSUusmw8KZVOmqRH9MUaTgui71
Lh68/hX7YcfAGu9ML6OhGtFazYFLCvT0a056y6GBnZeOpfQrVO3M3n7epEGvlXCybtr6LyZ9z/oJ
/dfsxDPlLnS55GzVTtKrKNVtMRvBEmz1H7ujsT/e0KE3LVYOp4dbTRzrvEcYQB8usPMxcmd+MdT5
tYryfMv2SX97zxvvxljbzNByskB6itSa8kU9IznhDWINx1V2bnW0uLNw2A1x8o++cTMAsUfr9sfT
INpWP2LC9+/ahzX1mAL2KeORzE4Sl8BujhUaaXdWN/lUZwdqAw70s/MoMrT0TjsRaSCklYa2DCoW
3wF1IXs0yj4MZao0AmvrCQgHt1dGX1f6hPJ+l1POcm1cXrRNpHBxbCqr9QkN6PL02Bj6TPe3/lg3
WNhfp6pFYte1/NZxgYuJNbWmq7SrQD2hWuq6ca4S84GKLD9/4dixMHWnF3BDbOgrZaLZyH6mO1uF
RMR93uPofSUQyblCM0m02YdEqlCQe8A0wGqyV1089qws75RxbysX/VeZf/zLdsLG5TptB/ATj84U
MEH9mN9yXNPnkIjspbr1ZSC9gykaxCot2315a7CeSxpw9p1BlOewspXkgugFHSYjsE7RLntkY98A
YUzzLOC0ZJ6zzDvQt4qGi8ToRsS30ydshaF8NPhVAtmdvA8TdQ00nUUR9CG6FTU+IqHz7HZDf0LV
Da8ULKQOyQAfQXY7JSqyr3KoqA63eWuv1SLIkmdb4QKpTkxc+wBnK4r9cltYcPoFUSG2c5z0X9Aq
hbYydA8bCg85eoB8LXnEo1mOa8nVOmnLvnYFxxehRQrHAxCxYYwvUL0qChgNslErC/2EKoQOghQI
V0iRRBetnOYiGmX0XRsChj8z0mdUKTuWJMUHLEGG3+W0JHgrFURVK62PwhazgQFqirJLJPG9VL7j
skKnHcRR5G/lfxw66NhpeO32AaTZ0o+90L/1uW+OTBVGNB8CDn2sMdud0ZEcbeUD2JVpyE85GQyS
pG/1nhQ2mC2Oc7EeRNhuzSAyt1C00ym0NRByitvlDtjXwzHJlcBTmEGupg25CQmgKr3J3V5vP/Fd
dRRScvSLy7AHcnPuc9q53eeKr1IbRvx0kqVXW55EbLrbxfSfKczLpsG81TXLSoymkuVr4J+yZcKv
1UZlc1TV6lqfhL2Z3V7krMq+9LZ4n7PfvZufkYTjY40zIlAetU14sbOot+b8G6OVhZeOFZHT3u5A
2WU2ahZ5MGO78fgKPySs41mLByA/UJR8cqK6U9cP2xqd3r+jKeFMPAxK5j4b35/nhXiJV8WsVHe8
IxqbjGE1AMmst9tpyc/wS3HmFyUWQuzwUSX0UmzfrthSrYhZjigBaIiTNALhzlVGGR1ZBtF45HlW
chpIS6XdoIrY5Nd1esePJ9smtBB4+GYjkyAXYEXLdh6usUMhAcUhayI40m3xbVUfYaDuERsgS0Ds
3xBqj4xN63Fc3tJFvfv6F0/T3IqgW889sZamRyrITvqsKKaOvGxTXBDs+jepQBK48R6OXVPZL+6i
AKBKTguTAdT6yaKVydNJryxk9jZ6DZyHjYsLili27utugVgDbYbKHF4i2xmAnlWOdlKHwnCxV2W8
4DjCA13cpQzysmoLCc4USBoWmPFcto7nmy7jlovCHz4a9c+RBbswEpG881DPA2O1geMqVHe7VkiB
FfQIO/MSctq12hUj9dQKYXBmV3uJ02zeVYBbUkCjR5kAnrkC95EBCvQAdR+mnBxeA0Cor6k1453l
VVURY8kIuSMFv62zpomD0eI2GgOaQiO63BXH3BNgsH75uUzR4O78Kj6fKzp9d2cLGm2VU1lczCs2
X03d90RFyr+XfwZhZlRD/hjFBIGtf8afdOdxLwbEdvp5uDFSGu2+l4tNrZjqHUVMPOFkVyVng2XA
OOh58DdYwdtarpFjrkgjghQVHB7DEn8OqSIkWTf3pr2OFGeQsJ8ny9mVg2Ygx1w9xwhKtNmF7k0F
CYgEr4rFKfoa5qLHCEaBKJ/tmu5+AHDHMI2XdC3d51c+Tp+EzenkBREzH6wEAPLWXXoUyIv/hjFG
BV+aLfiSxxNS747GX+esHesn3CPNUfQNU6/kC4uzgeRkGgFQTFGlv6kXy7G2RfnqSy3Desrxr+88
YApRNeWlvxBZ0hbKrtQ3PjJCoF8YyT4LjoQDYCMEFVLqlIZw2i14gu6nXtDP++l5GZ5XOkkBXd5w
I40E5y7sIDrPIMMfZNQu5bifyt1XuquHKEthvvqYmNNXta8SK4L/J/KjcJ/pVydmvBzkDqyKgx5R
6cPMxawvnxqViFrkkQzgdrqF/tPrYB6p5PPlb8q+1frmwqRmaRcXaZk5WsBtRX88dODI+W4+UCER
n7evPJF+2GyCy4IE/QPwcctqvuc5rXQG21b3wc49klJTKrBzeHbheDAAF2Y3LxKTktbBsJcMKaFN
DXlxnoYhPOMb2C76eG7js9tQDROwApeHbO3PHl6IaEH4A26uCD/voBrhok7P+AKvI63psGDZO+vx
N4fdHX4v1x89OsvBaPX0vVZHdyV8BOMWgJdq9ypdiYb9qaP1eUvJcFdT6ClYp4WEy8xDxTqFAaAd
ID+IRIxJgsz9Uv9rH7Gej0VUuuUkBtFoM9sXQuazdfBHGkVoNcaC2jjaZrh0cSnant7ODCT4Mhs/
Nq5l11raG9dCO8eRmL9QxZK6ZyIGJSbN5Cl2BAXfM/vJexZhjKJ84mGk6cCDKUth0/6tE3oX3oTU
ivMxQZikEv7IrdBaUxb5cEWW1XKFZ8UKNy3F+Ia/aXh3yaGMKlFReU/0/9OGyW1xdVtfo2rm1T2L
BKBmGvduUrUAtnA367Kdoet0W9Ht7iyO6XBXLJBKmcsQXVH9RN5rLmWbSXfiko0O4FuaQShupiin
s2aUzR39DnmnzbvxXYzx9o133GSjOKXCtqhrivn6MjW5S4GNhsfPB42iDt6IylFdfVyA1Ub9YqSt
0UJtTdf+wuKLfJquWcBU0+qL64Ho6xDLGPV3kQ9wF+ZBl2MT5T5g4pWRyU+4+/z/wFJOcVeExrrn
FrgBz3dJHkPd4hSW00vHTYz5ZM2sZEkeasIK9A+oGzltWhQLicqwlM7XnKdmoJgOL+g4tV1/sM/Z
tMyg7sT5QQwllcLc+7fRJMTMVKyiDdEsUoeSajkqzB3JZ+C8L5I1VVtKivHAV0GnBBR3HP7dktfn
+EpbgVdGNazCIyJruaBhfA/iy0hW+LGrh91VbsUe3DCWr4MOTiW4yLzmzJ54cq4n4yRkXgho3NmY
SLsmiVtLtIXTu6JIyYls6j7cD/jtZb5Xlwu06w7o6IJoS4JVyr92zvTDRcnDk7jKsb5U1+XGyaQK
gegNROiqlwMMaweMUvrGy2z7UZtIpHvsV5lJLEWuwpAkDqdQPXi8jzwthzZXALI56bTJC50J8mfl
sVDcb1/tVZmA0CaDV62L8RxkOo0qX1Rw1AV/EHHVdFvmWMu6rKMhJ/7QYbeEPvs/uuaOYUY58Ln1
uZ0fYfEhIRJrswJ2mPj3DjYjO7b8yFkB5HyB+ND1+YVjPSNk0xl5PJzKQrwVGjI68Hcmsi4ckyrB
iwtwWP/27+R2gBUWcMsM/7wZlJUDA3KD+4TVd9fa8Cf71CGHFBXe6FU9xySTADUPLXCq/S2Zx1iw
Fxle6Dq48xccqcRf8HGF42fj+GBvvBz2IUssk9stUKVPvtVr8HI3ubJEmGp4IAd5EB2RCzbc1j6P
6KdQd/pL3UY7BMBejbwArG5UlFLrQMGcygn5hK75Fiv4G+yZPVuOvaJgvT/WhaBkxWSQo6+KnBk+
qiwHi+jIqo2fO4wYbCgr7cqf7fquhjFYMMTedYLYxZr5Ki6yd0Yexg6mOUEy5IpU/fJG80/eLRYd
eZryzJ0KIOWpzkee1eq5MyOIEGZYgxuxPgxA93tntJA/beCwfpIJFT4C1y1xoPgoUzC/hBGkrdeS
TaBE+j3Cgo/jo90LWePr7pvqlbM2vzLB8D3WpJkVymylvIFKb87LyuJ8+6wgr/IWyolHuiBvOwp0
hq/EyPy/q25dYyUusp0tqjEzk4gkpywhGhiqLlHaDOeiEZC+deexSi4rQ1SfXnhMHDUqvaPs8Yt4
hX2q2KEbIhaZKgOBOzsNnGEuOmVdqkEfzfRAHHI0vGoIkjZf7z8R6kTIkGIp2uT0sVNBPik+gk9u
NJoerFF8u1rrsTnd6TpqGEo1+pnEnUYGDc7Os6mMAH/S3N6SBvBxHEpYRSCou9h8nKBjzaNgB2iQ
w9szapsg95yhw6RTZozDAMTROqAx80H6/qlYp2Lz2WqF2n+YaZw6I/eKQoVCa3Q59yy/EhMHri3H
00/oF0k1O7tJv8VaxOjogjOxtmerkoNz1l3Nn0/UYNStQYLqyEjIm5+8vAFkiYl9X2IqePwUj6D2
+NSMGhfQABTMgSwvKTFkWKLYhGw/9kYp2llNOzcEmB5HNEXysxoaFvUnQltPBEscJxc7Jub/jGlF
SbCczfoI9i7Ewb2Fhmlh19V7+d2WI5F54z8C6ztP1aZzKkh/8UN2bQQM4pC4Inmf3Ua1DDTKIUBi
Mz8S8hXmO+RYfddGHi6mth9afsvmwbgHXW45Y7T5yyBidD+DXBxTnT3Pd/AqmueaucXvXDWq6AE6
5azBScvdO2Vc2aAM5rg7B2IVF7VYUSABrUtRf87kjJ5Og4h3tOkl5mzH+Nqy/mtqHk/maC/JnTIa
xtH85ZIqlSgGjvxfwox76DmO+riUkV0zWmMV3ndtcOXMl10QVKZadqBwGtYu+GBGcx3j58ccC2ML
ho3wCV+g0L5kRXa2ZQxWmkhR4oAh54jVQMPkC1QzfJcgAXI8RD9q/GRE9vnce+KaxN7u5Q32KHWS
O0xQWwYkAMzs7KFHs5JIfnntZWxaZpkfCqJz48RYcIHnEC9CfC8T6ZuCpIzuB8OU1dU4VpcGfeuA
oRqP8EroQcMGYphXUDmZX0YwNXWlhCGNY9nO0VSVB8HgNDoEdGcu1y3G5lNuggo7aTHqsqC7HfhS
aXjn2s5jxIQ56CRGZGFaZr5uyYUadEAORPwPAcegb8FP313jmk4PZEDXUWECASEtyBUQKWiDj2bo
io2RV+k5NwrwVBRjOKc2MgP9iKrhyem6IV7Is2VtddvNI4aBnf+cE3YzC5Xm31Qw79w0HXQjEwIP
/lCHbDSRKN2IB9hCKg+KlIj/HOwwCppz0YsflukwoSf6s1DqJJZ+Ug999wdPuExRjdZVlZAAJt/p
LyuJXjuKGXndT+tfylSmmcGHQjI57hLksdqxGnE6Z9wwlP7ZhGcaY0VybuEE0ZnPXyIu4+5dXktv
CB8t+KdjgCyA50gaxzSmdamNcSRxv2kwVzcsYtuho0UJWZNuYOtBE1ANcbV4C/rjHXDMyBfwybbT
uz1F61/mZbe30t20UYsK/aSiF6yM4AE8/yCPy3Rx0cX/H67XKC08K81O4uvoxrI5oxfD5+wuy7Dg
85eT0nJcOnD/OOdl0BjGSzm8iV7EISu172kA5cddd64q5xuc1t9QzyxByGO6iVIuAEogTraVjMdF
sEO9yYDXhXu8cLBmeom2zv83VgcnNH3/gGYxSkkB09KkfqtjZ4VXoPkl5DknDOIKi6WIvj3DPR3S
PBSxFu1IpBw6ajVxNCca6IlzeDxid194Yj0jZMRS3g/zcqjNUFrrcpmaqd6ukGiSBuNbkkfn8vFG
A04xVgwqGVeYjNehZkDSc2w5l9at7H/WVv9WmlQPCTcDjxXA9AVstmN9oM4bxg2wKM3mus2qVMTr
qEJ/s7hpOr4X7Ety4/QfG2oAytRzsmcb2SZvU0kXVgPCdeincVGQ1N0ZH2zPD4/XsoUXHLFyXPuR
92a/Y1G7LBR6JHiPCLHg0w56CU7pH5HmO1FzXuYBiTQGphnLzCO9cXQQukGpC9dJDU+Q/rTbQv3p
QhNJXs5+zxWVKv/SJZXeijDXnsITkJj/V1+0Gz5eanJ8qf9Kui6dXHzXXntGC1nCQqciosexOJ6f
9etOi6ZaQHdDTh/BtFDTaSdRHL8p3Acht/h5rxIF787kaAbhDJhRaucANNCJ+WUMWQclGQF3reTU
UwJAnIPoP0dE0fcDB+Ca+ys6R37tHn9TrXIMe3+W6O3iLiwQHXOcJpYY5D/Yu89IkOipYT+Yv+OX
sq2s1cVAvhZk8XvckGKr1nhJ38as6LxeOC2yFdKzXJEabJmstENl38uccaP7/zHkRDS2Q2jUeaR0
pWq5uk9vCQaoqSmTFk63i3kF/NjovCCuITbuyJfayCOeiMv36kUwSJo4anQ+j7SsehBzuTZoaC2y
JWFPRh7TNpV7gnDpPfJO9bdfWyCKa0bXUc4KZzl6VJF4b6I5bW5Qp6naslU0du6ejW5ek8s5/eaE
zvZRR60AFe15hXc5av++lrL9pBXe4kecQCxD3B98xwg1kd2sYHRzkeBgRsEi/oHzX6ao/ZxKNgBD
DTryGx0p0eFG/EeXeyeP8A7dDiwFhvC3DWUhsVXXGSbbWsGjLBwykUgyEW84GIm6Vh/zcT6RBkVQ
jY3hSNENCo9c/sP/sGto0s/FohGK/vE796FixHNH4qPcwNoVxY6ebibWNFxqu6/5mpo7UmMkd0cf
WM5S/5WAfgK35JtlphlEl8zGnrzjGp4B8wS87DMLg18BOLOArDJp0GGO9KMwp6w/GGUz8AGdgD3y
M9HzYYCFaHNvg+Yj7FFIUq5nlM5Hjra3y/xOan7+mjqVtxiRkfD0OwhdlMKUa7wHbpRck0wnaijI
k9KXHjH4uWFa4idZZfop3p9eWr+Ye/E+P5XkFq4ZB7BXn89lxBUbkmIf1fUrW3zxVZ6R6RCR0N+I
HoZYjBySPj93yEWZUHPP/9I52UdLdwW2hp57Y/J7xedJQ//d3oVkbmL76RGPOMSi81eDSPSJmrKI
hTMc+sEePodsgEUVt1Orm4BE5b6SFZS8lMMeYuGD8q+2wnnR1YsfTXNRqvHEY5ulppPC5hxOTBVS
P8ClKYFhYd05Jh2Jh05iIZrPnGh9uYB6nHDbq2kPg7Ov8GOXPQmIyhfT+rVOyi0M+bx3GVrQzVX9
wrlGET/XFQoEw5FkI2y3HJnYXU+XvII8qUY7cDsBJIKKEEWaWfuS+oBlCgiuVtrtqjvA60SMkwQJ
86+f/QeD3WdWAORAviv6gQnzO0fruPONzYFdnFY+7vQLP6jyLTxu6vnHG3zEshkJ3hjpwA4f2pDf
ASCzkouxSwtFpWwZsjnX+Y0L4EUfryzaRJUZTUFRSuXxD1e25MDjoaX4mg2F4e9Ru18B9wV24OPz
Prx886NJQkVjEcWhZIOUZi+hW5B9CEmvIG634JAkapUdX2aK8Ir82twiZjVF7NBnP5D0jOupkTDe
QPgVkMka1tnJyN7C0nua52CHPlxhHOVnIDaFIBZVRoJ2j135Qv3x2iItVzJLrp6F30izQzXX1vdu
iKjdiXg13vRDpKDAMZBnqg5/YrcKRYMTvuTzWRt/nXKadA5nn5ZbM1nCjddMq5DjWZTUcIMfxPbE
LPngkbSfMmH4dOGGGxDRkgWCEItTYbbXXsXsJVmXTWTjSUASug5DiM0OcAAPiXQCVh37BbVEdFaP
7dhovYhFaCtO4w7svIy2lz6CnMMT4yXKTnxqUlv2G+jyduTpJJw6SkJVPEz7dHSkhbkmSvErP0ii
9Hy8HLNkx1nSjazXcLY+UMw24QGeLE1LOQrJnNOm/XI7tQR8sBA3/vMVh/Omg8cs5S6WLQTwUBI4
dqP0YXR4q+ow6mnS1GAF+FXkLtNLxzBEYwUpxdDGt4wSN6MXWIbwc7Xo6G93DDT5cOb/qX70gaaz
AmLnnVwOvgF4XHGRmVW1bVgSFPA5W2/bgXOlvl1VsQHsDMMzvZ0mBdy/PThndyHlK0cRY19IVOxO
hewb8wVcnMXYGr+xxLEjaSww83rPePt2tjTlptSdFRWHyLlXe2UOtGCmP7t8TcwpUyrIDMOe85Wx
2BS16+6Glj6nZgNymIvKVzebg8x8/VHJQtsjd/AwSRARDhAqvltJpdnLP3BvpcsqKQ5p2fmrahcC
sbhwFgawgAAS87+TAviDLe/olqNqIypmlo5Ug3bCDnPosaTZLFJE9LOuN2wPKU1JzTfiIyvqNPwr
0ANH1s7DifNjN7uz2fBaA6i3kj81Yxxjb8q4SejPplZEY5qfzCfEtAEVCZunQ3gvS/3XK7GTlwu8
4dHvtA26Ndr0/SXCC/dNA3DqtiprIS+i1ROVfOMhySshuLmug1DlTyYcDEw4h8aMrmN4sdxL7FTT
foXwclIx5AaKTGSZ/d3AbEJS/yzdJiSUTYri85D8Srw0jb8vC1OlridO2mX/NllpX00qvnBV+BMo
L2wc9+H9kZXnvWdj80tgCyEyRNSTu64jKE20yKNMbaL1sQWpHrFsN+e4jdgXHB6/Q1b6VuWIZvD1
PgbwZ53AbCYRuEpTjzAQY+k2P9RKv+vtOloPDWhPFnj58sIJAO3TDJDrC92MeaMkOTOtCuesmHx3
n8E00b6G8TzKKrFdSoL/OnXbYLOqW//NDtZfABOtfqQZyRTqbDm+aKMiWbP1N0bJgFhPgutjFmob
c/4UyxND3KRxC5KIh97MQJbXv66pJOVu279Jr2w/LkwXk2kTOIUR1vGHIivoxkUxm6P7P6QZ5w5y
NhG3cQM88/sAK3gBS3HPQ+7OjstmdQr5EfAAiRcYHr/niW6pagpMG3TFSeexYwJzLUxfGlaQsQda
pcUi9DhAj1nvC29Mlxvfn/dwkJLVmSOOV1r5QFv8luC8ddjekiX+xnHgEDmS196jOQe7iXkkVNQ/
x1D3uDo3lklv87+pevgKvor4HW4xFgByrGkZ4dVOYHZw01uYls46Vgc4+3oTHgzPxS2742sglQvl
or/QPFkHSTpNdQIZQfkA6V1fqF/zPXkwXygddVu/ApQ3RHJDCUYH7GqHWoZ5I0qKrpjuobNgNmMO
E+jwLcFJK7FscFouivMbiBby/mElXctNgf3O1ZtSpGC/zq8Idu1q4D9DOFye8tGhQmTs5LEvaA5g
+RxWTNvb+SsCZaQ3zl05R7EfMhYxuGTkpPzY7VKuf/0BtBsqAPNSvGmy9i+4p9LpopYlRIrcE5wp
Hm43SLLMhvJR4/jNUXzbu5tokH+cEaWx4DFipEMat/YCTHFx7ibLyztSCqr9lAYDDicaTfsZESD4
84RNlNGYzkX7sWRLdVoaR8OAnijjrPUDAJ5ou2VQl0fA5wg38iS4/a2ivz2B/GD5ATSvSpH0G/N1
3+/c1M173TeK49z3uxnaGLXoD5egiQr/2qPnG7aTRcTAO0AZ0ao1Bfc7aSjpYT8kGd3jUOTl7Agv
cCpua+LODfQLVDmp9n2SCUoMqGcxSNqDYJRMMSwSXq1/m4bRUVYjsogJv0Bdzps0xHB1r9+mHHTT
ll0T7KHPqCrQNLg5gkLL47mHAY8RQMAagSBef59O374yteLuSK9vQ9keiCj+A+1rxD1u6ret9AYP
/nu7sURW+hXYWKVAt3V33avaA023WVaA67ii4Hwb/6Ope3y4xBc0BxOOeKPdlggWFVTYNiklj+12
71Vfb2CknhCQbZjBc10rrgg5T8rGDtPCGq7+pHVCPxscgPpbFJQ1jn3wB9miRWLneucsbI9eOnTA
lPYO8zf7hvWONdH4dJr3mFv9OD0180YufYT8CAitjrJEi0FSkupqFC9D0qKP6YkBn6wpcRLCY2/0
JTscjoBO1/L6J6G4Njd4jqACDGxFeppcLuHP6/EE3FJSFQVMdhKzASXGMJo2mMbiFhb28JU9OwdU
HMnugiaJycReLiJ/XEj/xCmsGob47NWhhelojeVFGvPPB2bSV//uutedTGgajyd0YVuXGW/ZkZNc
37xxhVSh3K2u9vuKsflCjTZIyfVc4OP5lLRrbiPH31VnmR17/0nUlEC47d7h9xmjqsitg6fOClQy
NVobZJAmDVxVerxCbY4KoOlk6T9LjsWKpQD2bPy7t+4bHw5Zg720hG2xNr6WBsoPqE6CglSyqp4Z
2QPnojbb0hKM1NZQoMdIJQiVETW7vyuiD2Vx/jdbKpx8E/ZWljsnq0Bw2AdViYctRxwhdh/bp7C1
BeeugtuGJqIhK+B5UzsnllH5z/s4MePY+5yBK1oxskzXaI8rUPfl3TmtJHHLzX8E7xZZlGEfVzks
wrm/pxkOoePQrOcalQvxU5HoP3hZgGwGSMArnA7RX+P8RWLfvvGp+ejBBK2p242vcDjbcWrAMvXb
CrQCFQxq2kBjQ+8blSmA3XIx3XVNSVB/AorcIDvsTw4XHd28i9hN9TkfbYzwpEFx14NyJMPypBMh
WsUEqfsQpMYw+tDbZS6KSRagEfKribHWeenvkPJKyRbieRurghcFaDaR0tK8MrOB3cIjrdXL9cEp
hxHjpKodo+mTXwecOfwgJIQQIhjwl8wFfrcKvQDQoVN7bw3B/KNMNKzZ2lxMz6a5c+UPRSjbX46U
7Wqck+HlrC/uETzzJP+/8w++JcEUi2b6xhFvzhMCfyrb8FJjk2IiGBQ2FmP3TccHrgPsO/0DLr3X
5r9/ponhGVdu5/AFhafcqeWxPDCk16DXVFcfMDof12+IRsYJxBqDHZvnAuEDzwZ6qx6fD9V2QjcG
fFTQbuxfOCpAdz2A2i3ypmZPV7RUJGEJH+wd1ry54IJt8LhXCmcx5Yv+2/m6HTCgTTJLT06+2vxG
BgKRqpgAAINu/34N5urBAb0uOLA7FPVme5k/fESPP6UFP0mB+RfP0Y+htvNRy93GP6lwyTFQuzFz
Betw14pQG7NRJ304Uln0tthO1nX9ca9515oirxTpSH3rCNmZWTnGhnKMpr8JuJeCdcqlBuBt0QVn
Dx6HCmfDGm+1SJ2ia2C6wVdMuQH4opTZl3SUl0Hu0+1gVEYhZxsR7CceMA3+L/+a7vfwFL+0l3Vj
2bCllEx65LMpqtsjygysIfVrRSpgLR3KdnkrvtV3snJDfpb+GKlyWYmqynFD2bdeilQapzvgMkNq
9lFty+66QqghMrYIsyaPQjyyy3fBHxIf4rWeQERTem8YNA6gTCL2Oq4tBqDUTkmQlFSHGn/zMTWv
WIPBbDILQmW4NjEge0Y4xl+vxpZXWBYuz7MgIrzjos+XFdEzFWw9svWpU/pQ7P0x64/ebs07Feh+
v+WSHEY1JId3nRMR+G1cq5Ezo746QeInJDZNKh289wb9O/pLi9cscFk2WmY7NBq70jMRLSauhtc6
fZpbAQY3yVYEt0lzCnTbIaZa+Hg8Fh5taujDtTHDxR9mjueq9y5Zv66eWfEzdNcNxbgf+/8ZCwKK
aZHP6PfloEr2/dFQEHk0ItJ+hsp6M7frdfckpdNLKNxrIiTQWIuolp2zAX5v0iDmPvVFFzHCJMaU
CdiDstV+/YIXMkJTpqi0/kNVZtFCTwSSAVN/aMCZbVZRNkNCvIhdb8DQMRcBVy8eyqoa66Ah0r03
AJQhKytQJpG6AAue86oPS1hHlE1aIRvXG0Jah7bWbp/QU8mLfxhPzYzNMnitMAVOthuleQcgoPY+
aaVlfrh3g+de8U/Ckb3lWuTs973qsKGz3pTsGEXt6NGeGHZIzxftKSX0fyiznN23W1d+T7x857bH
MAsx9RMgJ/We4hQ9Mr3kXihQuGR+aB8j7BrD/a2DHf/jmsH80FSoAlAO25ENo20CekggQsEHFCGr
MFKjWHoCB+SpbzO7KskZCsKPrOMiij+bx/OKNeCe7EFtAEeuLICtz8UimG5kZsmeeRLHfIalWZM7
9XCbIWBB5Ln+AVS+iMNNdIfcSSEEqPn8k4P4cAr0S5AZgEYM2nlMd4DTVXiMcdbhFhXRhon290BL
Md6xp03+OdPulYtHOReDT45Xl2gJNAWwfsvmLGUFD9pICDGt9Q6Z2LEvmF4gFUwlJpkXNEr2fytX
/2F9V7bjfqBNjqQrPPMGBB5zqL8IzaUo58u6lR5YWIczM9lv6i5vXvmhm+8/CWcZ2zID9nzOO5n9
kiYxlohv7KXWES9U6GW4iDPB1M9CYzMVSX8umNWcamItPYmNwFX2CuxIESybGEDLaqpAZbchhk9u
FJqgtZcSlc5fPn9VRwswCnsR5YIg2Ur8sfQAmxTG8VK1Y8Tlax2BGsFrUYKQWobK2bhUKZMojfXo
1ypYRIhXpHF2E8EGtn/Yyv72slRS6cKHJHA7bKI7/d5hQSibdFszwQ/xrzZ8UZUWjw+5M9bXjFrC
FBlUiMy4z0wkWzUtsDiOVwKsJTL6iL+WuC/S3+R7eSxpW0hbCmrXH77aiScJYzHlaH4Fqu2bfL5I
9LzvBqbhTd0j9HbUqo3WZ0HUF2u7sMCNMl3viLrEZ136tii20v8+ACTqCemV4/d79jOZACi0mokK
uXAi4TtVrAhL8L3ZDFKl93q4pjInCEXsf8Isci3hpqJHTvBTBxzlTZlwZ983ZaSk8+rrv0WiyfBb
1DsXUlv2fYhqgQ8Gd+TixDZQMxPz2NV+r2lHW9WTb7vuVm+RkY8xo7vMqiy+xJw8LK1A8lUnuyrq
bnEkMXEEkG+FKenBAq9VlvgqTe8widhiycsvpzNdhLmYguz3yyRZLC59XF8fbtflaLBx/Njecrsh
jfq0y6D0jOZpcLYnqvu+PpMyZgUuoNpxgc5uwSdTElljgB1VeE5of395SWPY4Sbhy2R/kti644kw
ccwvheaV6jzqh6TByfene8KkMGMe3FUcMoJuVyNZE3ii8S5MNONix+n8faUvwb6cr6G7TL2Y6J/O
ESbc0Im82r1QyPLBhSkc3uODgf9rPTadnq06fmsvbkwQK+bOeVmK3jT1gg/RfLr5r/psKd5oEhja
yBMUa/fxoFiMFl0ts4mAHUi1i3kJ0QbMcI8dfGPfjsMtYdTqzlAQYcEbc/AA+AQPA89WULNl2sBB
gTeKNcLd9jCWdFJBZLUX99YG4eggJhIgf2sxFryyPqUf6WAv6+CCzF893YqiPHwg9YV9trAcmSxl
ILNtYgCfnrQTGHhXbz/XRrhi/rZHwMwHGkhVC78F1ECgBV2TVgsi+3XrX9uZDGtLBGyE/ie2ZCL+
DFHzVLA5jqR3/EWGRLdU3lHnQKNjcuNfN3wcTb62nt0gI/T3SWIY0DLZgk8qJGZ+6LgeS/bqPuiq
sN6eQ7brIu6Z/uBJyRa4OrPU0wVKZ2PnhrUOIKK7fdkV0jtzqA5XlT25gRgf1ZQ15mGR4hVWVusg
cpCNJqNqolbQruQn9cnVJHNnere+P12hJLlmx4Anfz7m/nx6PwOmCTF94/OAdd6RAA0mtZ1JXo5u
tCSoJWEfBA/anTqu/G7Qlwv6Rh9pyFCvR8jdSIjl/cZu3sxHMxooiCb0M2y5oAcVelhgI4YUgk+o
jQsbZkjTLeq/EebTlz/hTU4vxMEhD//NyKfsYDYiplWRU2NeQok6Y7GI2FnE921eGUxhaB/F0E50
CY+CrHtJkuF2Uv2yMH5p4yYJJ+qEeeUEM42g/XBBr1dw2Ngkh+8TeAgavLqhnvtOhBybSiITe2Pm
MiYFnSbWGVlgOCMAJC9kDdHk3LUdU+xcpFoykt0K4dXK2VDIjyOsskVl2REu7MqmGRyWM+VWrAfJ
CdeNQ2vdo2r72PwjW0lBc4hIJZjPg8eDm2dWVRT1MySYsXn98KHBfndTZiC1FpORFedIjvJahRkE
MmpUbyAxrx6E1rRvUARoOmEKlWqrWMA+2x7jPNaVsp7k8Xt8wZQs+IfYg9vRexDz/qRYCvW3MaOM
/bBoAUMkp1cwmmpHTCLkJ9qFYMY64YB2RmeRArlAiJsqOXN2ZbXTW4Qr0k6DGiFuD6eRPwl7WwFg
47bUaktUFB+3rdfH1QSrvp1U9ZFdyXysmVkVjoKfhsvEb5+tUy05qf5kGai6k919i/XofZu6eqCY
IqiUg2QsJIismRBI+HaqgM/di+0d6I1yB0eXHjRBXfbY74icI68xJ/a9RNtB6cALOyvrqpicleAf
ZKupt9gNiEGt3CZ60djvilwEOTt0lQMk8UAPeljECJRpnE/pdSfyk5C9lEaSG+NkRmSsirvda3Nt
bDzXS/cYk5mB/kwfy+QGy74pSsk6tmgzR7cnd/htqI7I08h1UPJtJPqa0LqlGa9gQB1W/030R28/
5W7VUxQ3sBzn3lZBTZyB9MtSgiUiLtMSr1PFwjd1hs+JklJMJ/8aFNGnBSpsqp9VmzcjHcWQSkxc
G4pRsABeLWCqJfzyP4M52biD8iNbibEPyp1b7aGKsIiP1bzECiQazyRKDTwzy3ZrXssmgyjv92JT
/pL2QC/H6wzUx1U5M/1WoSrbtO71rooqPUISm/XHuEgnQnbeHp86swSaNS2oudUuf6+CQynQwGI0
aMySxDv+LtwKD6N/Epb/Wr9tBEAACJeyuAMCqCGTkSKhSjKaXAzQY+/rIqBYwzIfrX4NI8vpOegR
u+u6oI5HkFT3s5yHddhcXwW5iLHRRtQ5FlhUqgIOu/Vphlep3eX1qrFtNnaODJCocpABdta1B4ZX
4qYK99Ryv7kY13d9FirFHVrAisPScbomVDPyVX3g1fCzFHJH2UT+d3QThIuJilwktQxJ2UqJ3tvf
NsmlnTlDavHGfXPgiR/MjijMFwTooN+YzG65/SuGePXN/qW9u+5Wc9jm4GOIZVNJ9yVH+DgvmqMy
E09omTlY3e+J1iaOOax4HjwnTZn29jf1+nSKY2tFoKaGdJI91qOgEHf8I1yTXlnvfno55NuN6S0G
Vv/tYT38rq9H4RtENpurhlpTneo3JQTGltRkgGpVvcswMU/YgWEhRkYM6qeZ63Zh8TJ+Ra4OdGLO
V6bMZyxnpQTbCYyQPh6QNaxWkTOwQSrs0DkuwWykA2wY52DPdTnU41XNDrsqNdJfyqPGXbWIoWIy
hiUWsplf9QY20iEyeuppul0MIco5T5FajQl8ybUscv+SaeRzVwt+uzrBbpRvjJCiZI+b02j0ObQO
A89v704pyUKT2ozockhn5Bq2x1JdGmhkr8qcL1eTxol2NC8EpzzBtuTbCShqTXHOtW7+Yxxsr0va
6JrkE7gljGjHqM8w5T/22FcAfdBPvWZaKIYHsRak43Ctw33ZWSU+jCrbDbrM66/TScMmwMERGeJp
iMkhSK7J7d08Wktb9sJmTsb5wqiJ19Brj8i0Zf+XWEPlAYbuJ1qZiD0Hn3lJaEX+3C1C3bb3SFQu
0+HgfXeM4TYW2m3+Ro8lHZgVr3JNlyiwxNdV5Xm7osawhqtSlqc6COxV2QRy8ne2baiu5YI8kE/A
hTV31DQGqBclExbwkZKSw2nBFKopLwA5K6jwfHjjRTuNZQzkeODTJfUimFZqq5R2ad8bzz2JyRKv
fsabgSXCjoWM6zwl0lXNO+XMi2fUGAXCuM5mifGBWdDOnXyL2HsEabr5SzVzZ5G2mdBD1Vtrd0ZB
rDSFq1T1peE3YbeQXD6EZTkuZF5bB8Vu/Zq0cPI/8PAxUAbiy9HqZ9lyTOm/2unc4WeAYLyJDWgn
mteY/qZGvh4p+rV1PxjjD3TOlMitO4sp2Ptp6/MOrXB3wlR1RMthc0P/vA3pQWmVvVo+DfFzKeVW
0rxlMIuj+y1sKkpdN16YtcK62tEPRi+UBZIoPZ0YGU2/jJatzlYvPxIsSSjOIfjfTZIRHYWi+F+f
cKS2UpmeLWxkYvYL71pSX9bTQOX5JmtOIhkBu0aGBis7URVG3uovKmo4JzA4o9RlZr/dDbg0y7Jr
6/YVtSahdUFngn7AWx+s1yM+fblouKmN9s+DJ+iAZ/JpjShMDREHWn9rgn8K0I4ItjTT2fzeH1Lk
fSNX/gOdbHZ/GckVDvGJKuBcZWKkDkT5zWNNcCrfwEXMT9icfyX3VDUF60rCUPOgH0FlkAipEsgD
Pxdbyd3JMPc/zLdEn5nCMHrftFB+IxIMHKDToo7cy2ZA4PTw8vc1AleMglsSvLVb6Lz9xbFa5GO/
Hxp4lR65DQcrSxJ/A8iBj7qiKB3ZPmi5VUftakGXnyU2FfEmCJ1WTOfrIM6AyojZB2ItrpwwO+FR
ZrjvIIKGyIcvShYtvAkBQ9TaQ8JZom4BFnjW1ah+qdJ9f5iYoD2tos0230NKpD5Qf7eF2NFkS6Q8
TBucUMqdOHR/lFXSV1rBan8EKqSv0qRcXNBjxejLUf0dHDc2Is2d3wnkBw+6eo6KHXqXalhnly2H
HXfZ6WKN4/ClJJsqGYY6BEZztMRPqETLnY4ENUhikgRi8vUC4tQE89VrAaOkVkRwaXP2QJWqbmtK
PunlT8qmgzdzOxzvOcJ0aOG6DKmPWW6gNn3AMpjQ6/cF4emwQnwbnLdzxVt5nyoTyUdSigDyiOzl
mmnMWRF8MRhNU5NiolA5asFgqJFeAqGHDIi2Eokv0cRKJTYSG0dkg3Y2JnakQcWEHNW/JuIMPFv7
L2HuGPUw/wN0dsBaNM4wMhVB6hFMosWm+UV8IiK77Xaq/6gAUKA7jqQminxp3SH9iqyO45uUnMoR
ahUyqEniL1KCP2Uhe65KTrHUFtjPl4eefl0FcRfmtIIeHYGt3j3q7gmHA9Twf2cuwABe/5vxym4N
kZZRM7fdCDL3w6nSgoiQjUa+2MqdxW6pt9FXQnD4chQmeyqJeI5xzJAiD4dfjowF1GNqVb2j2mBx
61lBac5TvYASZmVR3IhP5pF3o40sy3aAQ8h28+/KVYa19tB2ZD2Hs21IF8Kh9Z/1zXv0xsCSPrev
YYUdeSgaOP4mze/E9O860Ueb+/8HJfhmWIgyU8PAHfBc2pTXuoP9dU3swB2AEa0livqROo1V6YNL
P/8OW6cRF9ba/EtsaxkDYzQ91uOX0qNHh1b1iQU58FD29L+kH8zWJ09kr54SA7JurJvJAQ7TdeNO
NuEjYzGF5kZSe14EJyjYzEgrri3N5dD/oVAioQGZdKBrBFevuQHDmOTbkInbsr/vp5DlNOiiBD7r
fjL+GCJxVbKPI3kyVoT0ny4pRsRmH+mBbhmGFVHQgpM91jEgWe2Rgrpe4LQVyqzYyiAJslr0TFQF
hTOs1Qz8wsHestieYrNK7pp9cP8lARwVdUAWmTRu75A0p6j+AOmu/jaWDlSsCYBLiBh9cULXXSoZ
g4mkH3ybmULdsi8rd6pzdCENZh7ya64v/YxyNEVsNQipvGBGQnombsyM1rEj72VnC0HRQMctJKF3
KpQw3mNsSUkikEjQjvrq48Z1AAklUJfRxB31ki2Z5+ibO+/W88tvxnTCofUZlv8OwdNYCRY14j3K
QIStnwB2HlZLkt2D5Hxic0u3YTVzgru5Sc9qxE/tiZYwOz9VMkNIJYFfbtnD7w2u5Bk8YE8tG+vn
WYM/t8JviZv9VHDz6AHsI1kyvXKK4Y5aUNC1Bk0ter8JsMjwQVcbxV32++CC59bea7LvOIvet/Hm
kzFzNt8SXSnwYrIWvy/h0HzgKUIGpcVSMsB6/dfZVQ9WvMyi
`pragma protect end_protected
