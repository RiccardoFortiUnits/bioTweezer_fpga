`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jZxb3NFCUgKEmoTjxkfUA3zkuZL7VENVcgI5LeszoGXAtWAIztLWwlEdwhfTTeDq
2X8Q5P57vpLNmopzBamrk1PLdd7GDhsgAOM00H2e08rJgPCSQtMv7K4XLA6AEXMR
YBf/W+/861g9u/r7qQDjWLeSLqYHO68wCyYr1EYR198=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22608)
VuPmQJ2lMC3SYBnUd8hG9u37VCAV5KQY0yVnN28CMSpdHp3RRjG0o1EQtiehvxSo
3IrZzgWHXdMo/FDTIJfYV49iBj2LcowX/HUuZOzw1pN/jB4diapXvzLR936smFen
olQuJyWUWbu68mKgwSr2QciSCVoWrwW8IEzxwJY7NOOAr2a6TEJP6EfV4ew7nuWa
pIS+TA55OJgohHmwx1CA8Rq9YorIcZYF7k9PsfMdQlCV07G2fR6iUATwRY8num4Y
qgGKU6My3+7sk50Jgq3yC0ACrO5FRoFlIuJj5m6qLRX/qnd9Jegs1cSSTT1yJg41
26DJWz/U0IlWuRXy3V+JSMMmDJcRvzlco73PxbL0asEFTjrbrwlu3sm12UuV/xl+
XBTS6g2Hde/Nmqug5kM966y9IQNWedCm03Sv7v2G687Ea5Ebif5l+zzqL+xOCGj4
ht+GSSRFu+sCb4MrwJtK1/uNHOKgabHmyX2a3LqLKNsB9/86ytN0OZWkYZyQhHvc
/MpDNx3vI4Ept/ZbHZcoCxIwuik0IYiG+66h/JZqABuzhIbmgehCJGnmujVo8Yyo
6IJyLKkv5Drc8buc31TRxx2pJA7oR5I4/8ju/XM7q/1czc6K67VEODSQbeHYs5QJ
+earK/1ajSw3yJo1OJtHCUrbfjTlmpWZn9QsY03oUttPkhB4uOFDFiqg5JFhSkZA
5gwg0szUaEDkEQlP8+/mQc2N3SyKHrr+vclmqO7a4KeW1Gnsy3r20j8Zbfx25il2
hpJ1LpmmqE/ZrZQk9rkVVJD90dt08tyC5EHHyqszCzQfYMffyRek1A0HAyyiHVCX
Ya28c+j7Tit0y8tDXiYCjVO6GIBlwwfYuoG44oPMusO0nwOJBYLKb2pNYnjmqq1H
hFaKMNKbc91tftzEkGbDv/03icRlNDfrLQvLMYS4iLQcG9RFnyZBVvUxx97q+Hq/
vwLggW/rvZ+DCYGcIcxygZXMvKeJ3ai/lZ7xdECcSsXLgsOrirX3mHLZcB2u+c9E
zWtIgKMGTx9RyEsABKiefmjST+q5nRHMrGrig9halMX360ziy+ENbldsyYXGkEHq
mkxJ5PaaDg+xrdkQmjrAaShYYVgaENkNYBCLQugXFzMVhvf7uu8kNegbifJj6qk2
0izxCdltmawRobY95+CLhx0et422TptDARglZQQ5ZAgC4xmbhwcvbgbehZEkJsj1
QXlGZfRsGfJUnl1yBic1cNdOJlk7DqTJe8QA48EwDoJ2LDANLjDF5P4yDQfrykXT
aGo08oeum+I7s0XUFO028vmn8uuNxxYrvDuDk7RqtLuSEJawx2dVHGjltC7hdLLR
8Om+IEX2lt0714SRX1l+hzCZb2a6f8uYN9HXUXDJcIiiGSMtQCPfAsNmeCYk9fDH
4zgZx9Puk5jA9ur5yxmOjLgTiDASKzKengiNxReNjGtL7dWkxV614AVz6p6CjblL
/esv1/zbkSUBqCbqcxV0f1//Ad8nurECuioN/hmk15j6cYorWPwk4AbHcl8Z5VO3
A/aBkZVj/EU496AeXGIUUcVM4VZ8WXxto6v4zoXwMNhK3ykkNxNDY7LD31zcG1p7
0tAxV1eXzQZfGIhY9vi9DugUtYbXLqwlQ5iwR+Q4kfDGCDaADDMmI2/pqPEvCoYm
Uu8bkzdW8K5ha+i4Ek49sDednjHUfM3h7TU6b7JU1PBzGvLcCZEN3vPJFbk/UJqD
4Hx13mfGR1lT9QpxA0FB7h4Gg3WciD/QgZSXiooZnmhOnZMMS4sShvjylgPV4AIh
wNWPB9Sz915wIC94HLFeOfm4YgVGW2kU8XGWyzocpCi0L/26g/uSSPNJC6ZxHjWJ
BZURkBj3jPkEynhlMzA6rLfoygmEd1t+f7k42WJj+VEd/l7u8gyXCI5DujXbT+NC
jUiMSYqNa26XuTCnVfTYre+6Tl167G5Kglfk8LH95ROLfp62LdsSIs334z1XvWO9
xHKfXAoIOwuX2yPJUNhH/i3ruXjzkz52fpdgm9/Eg/HtrguqUPwgmPX9dfcKYKJy
Z7/+sRxeBLGcsuct3NpFkDTyvbD7xDCenq0ixLa1G61BNJbRKDqTe1kqZdl879cK
xe2ThE2lFNmTcgFEElNNka9ae/ILOYmB6h1CR/swciu8vuclmZ0RM0Q+7tHDlvxl
QIU85HmFR73R0YZMF3pVm73PpCirYnunhfoeXzn1oVpj265241q7WNNcYmDW2q4S
ONZ2A4zQDY9V97If2SQ2gLFWZcfMDvABKLWSSK7+KVbOjS56PDxpfKThreDZN8dM
s6Do16hf+D9na3ZW56+2G3hhiEDxZLT9yqz614Sse2BaCZ+qVKCEcKP9ztTW4nuA
F7UlvobnP0p/yRzeUv6MAs2EtjIXePJZclzUuphAX9SZ8itoXu9Bom85uAGWuNua
cLq+mF+KB+Qh7ID513zZdb9MpJfdrN2WaSwKpT07ej6+to8O+WNn/d0A7u/dyYxv
NHLWltw5kX1HHN9pcbxUimt/+0aivSvgDgJs9RoJXlbtZMo3OCA1YVTb9Pf7jvFH
98EaUHapX1IVwQrS7xZhjk07TTjeueB88V+Gdu2KY5E+AkPRX60Pk98LoToumLV1
KdIHH72QfPct7Ew1fnMQQ+BdRMGN00v00/QK7VWDbYmdx2YQGUJcIIOK4PFveqBR
mC/P5A4Lmn5PglXBKvqc6NQkk7yLJF6ADL0SGNEc147ao3lY+axEBqeTM0b+N/VN
m3jkOshRs+UsmsLAqczpypv5XdNTkAeulr/f4yOMCamTPatSWzi1QniK0bbtodqV
wtsssJxZb17Fzq4gNQMYsfH2K7pap4NxJwS48J52lITkUhNedtAJWx7adIWCoYg/
qzohKCDvlSICB8ERLZxsbpenw/rs20KOLdpYuLcL+PdNQRPItOOtqR6A8pnNK3D+
b9rQhIctem7Cd1k5y5FNr4ZQkqtB66chG7tItrsnklldKuTHpAFmww8Gp2/TKC2h
PU0z4cr2pglkg+Z1MJcK+6DSfsF5mKYUqqntnaBE9NBOSxcphxw/ZazAPsuYgM9a
sQNTv2xV446OMc5I6GxOGts138yZAPwv8yiUpU38mPTmC+zST4SNEnoy3yvxkZPs
xlVJ51hwA73tJk108bgRMegRgfcayBtV7EXiMXNBpFVTNXq523wrUlp2h/Ha1+73
DmFMYfYYUsMXmbqWjJveQoJhx+nkB4ODRFlNfSMGJxUbi3iPZ3hz+a0tCEh0LrH4
I+EMBmAxxzyi0hOCawzHv/XJlVj6e+QDRgFbIDZe1qFl38eLmQaouuxMLEzu+J1q
Wnhx6YiR5LpOor+gsL6Emc90PDVOmZgAnGbCLEH6SbkYndWw1HukOY9+SdJqzapc
zEB4sq36vqaR6L0g0i2pEs5NYdbDBjIe4p/uY8MP788aJDd6+27EPW2SF8vhIGai
RF1/WeRSQarPBM6eQho0vtjMLy2hgik/nfWSolTUl7jp3TXQa7KMErOne1AHDKEc
6gtNujTPNNmyCu0aq7RxvmxJM8dIrOTTZm0f7176pzLkZjnzsPEdTj8xw3qfjTDb
395ZSOajZobVgOpvkVIKlt7LWNfPwp2XahH/b5c9cKI5gkMS8UAjND208eToDrqh
ui/bYfzwFII+3GrxmioHMj3OpNH6xp032nEBz8ekAU3LCUzuOQfsOaz1kXZaZLGq
HDhrZ/cFTRZT4kSBiPdvI7wqOZac72GkyrV9RHlcJQ7osaiuAmar57p5Ko7OXyR/
Uv4BjSwydBkRtJ4xSpNix9AhDokOHbrZWzDt9MVuOQcCtOff+t6zwXyUMCo2c8NW
qzUXhJBZ9/xTRDXv93WSCkLbfORLBEivw73ZwF4cZs8ieqbLX+57ubeWQ98UAiXB
wiwIsspGRxc0nj7vygn1byUWH8/ZQWKNML1xi1XafPDuBE1vCwEd6EGsaOQ4n1n1
Maf8eWt1P1MKCT2+MZ9zZbEZSbuh7HuQJgq8iYVpqoS6D0ylo4F8r6LOuH91DvTr
eFs+KKlDLzS6RzpYLXxz1Z+oGW633d8OJraP9F/COU/x0CcZ6NnbRV7b0xyCNRny
03yJFjEo8bZTN6ymf9A/kbLEL3gyYqTNnH3DkRP5ByrvyZ8CZv1/Qm0CI7DdKnGH
nwL+d64CPo57CxfcPZPME0zx7n3H7scj5NlO/sPSnmAQmb7nsS//GDOfFW7SL2mv
1VwLMsR7PYUwn84PdCueZdCGbyryIbGEtFF/OIEiikYSDrFUd39z0dVG87OEctG1
7+NKNrnK97OQ7XBjs6hO67MEbaiSrDdb2h02MS8FnaRCcR9bDKI8mmanWcMHlER7
aNDG5Cl1iQmASQdMMD7IkdhD3kGDnkz0hIxaSv3hF7VbDxRqx0Z24TbzGT0PQkN5
M3L3nHjxRyMxjJVBW8FtM83SdzPo/lg/kd9luZNL6OV89Z745RZuXQJPqMm4Yxvx
quP8Q90/o5YnLBxvUm69Kt9yHoX0Enkpfd9Kc/SUq0ij7v4ZW8kPgsRNTjm+2OvV
PtGxqMzYojlT/ct1dzaGoyWu5hCZQHCdVPMArp6GTXtEodhVJKTReFE4+yMOzJK0
uMFIOD66CjWRSCwjN0X89bcpSKwoiK0ZnMXsUTK4iDicb9qJVrPp0HlQud+HEksv
fSwskaqyxjgfwoPlOLjJA4z4VnI105hJnsfr30TbOvlIZBRcG0gis23jg2aHGFJw
H9N3Pnq4B9e5pf5QwQ4MKYsWTSj1jvUs7228YeV7B2BVXjHUMymN1Jp7JQzL5tcY
79wGPT+ockR/AVDvXtLW3z+ekFj92fVvXOhR9HiI+q8sPaYMwbJOfkNju4bUA6v3
bE8MwIiHjHrI4lUKyQbVvN7DloOuMdEAQCk3ACEGl5jcm1/VfIw/ECSz02l1Gx5N
fziGtwPt7o7wqUwWxjCvob7s9l9DYD69PbTS8cRpErZVeez2oAqH7VJ7NL5gi7B+
sNJPPILl4TeAFyd2QMn8AhjItZn5cA6FgdeNglw1UHNi1fbgmKG1rAj+IdUnWaMo
DQQAsEyvFZ1UcT3w4noP8d+hD5Ekb/6DmbfqxOw8Y3o5NA54ldgAVXM1Wyjx2let
2eyxjzyorFyu8fxAnQQu5jCYfkkTvY++HQTHOH1Q2geayF0Hna/dJeFMhRUDJ3Wm
b5aB9nwdD2GA9kAp0ZbNbdJrMw+YU7XbHUIyVhRMYnKYqlM3mIzEr8FE2DJ7vvp8
A+rKdnyO7mN9SaW5kGRg25YPTEZsIpA8yXCig6rvVQoulzSsw8UiQLNcSshO+zFA
sw7SPfG1WRzyfGmnu4zr5o3HDHWcPsMqnKTFWsj9CvkJnIyJ9448i8s7sEHLO7tm
XjW/WsUKN8VgOCtk+O4xWAu/SFHKPxpqKsZqN9lGX/IivbE/ztR8ZkMrK3SR8ngV
J7xZYeLXNTpgfRUYxf4ox0QHyKNwGKWhr0OawN8PfMUQ3TCS3iy2NLO8WOxjp+n7
hrt8oulTrw1DM4ukVETVflXar7I0hFHcC3exv2/weo8NidOOqHkBR05eQQF44bJu
sBkR5wo+VtSc7jd38yU8tFbQ5vXiVBFc3nlAvl6dOY64aOIMNJk1esg5BXayGRM9
g0/zlhjN4u8jkIoJlwtEW58jtJepanR54jSHSucq1+ZK0jIh2FnzIapFIUFS6wDr
MnuBq6dzeEkFLNf/EawQowwtXqzM/iMKHOYehy6H5EbCZX+AYkD8Rc37vw5F33k2
d1dIaen2PzUJfEqYZqkYq3YQ/4iQ+z7IX3BBmxgZn4iNFGw59YgfYwwB+u5tJRUc
riOYwzsNO5TpMFDnmyE3RSer7QH/D6niMeHXbGTdJiGRM2DswsegN/okXYlzZSR6
M2VzG6cr4S+5+Yx1sYAXLdAOddY7VlQhIdH39QfMMrodWT0/iXA1s8MzKQlk0lql
t/AcTOyU5vebOdFdYHuX9WvDcjJE9MHDdWNf09cSIzsrQDeJLueU/ipV6TR166wP
rHD6m/dL2vPZTY//xBavajyeASa93qltKjNCTJxhuS81tRb5P4tH4ZjNgYxZnXsd
dYJHPQo9YVRKO1Nl3ykMhNQi7x+tOUqsEQggl3d/hdipa5wrl5jp086EdHa5sB8q
VZnErCqdq2S2dIMWIFoAC/hzR9ZBDYCKcArLIiuquQTcScqCSpXx94ffT9udCT+k
v4we24k6tBwbJi53a5F29DB1byTSHc8L0EVPLwCA+VELD2lsZVeZVT0t9zpx00lB
qVcEzbFSHelpU56GAIwrqklkYYMUrjckewT7W/jg4GOd975LqU3we02vhJUbRB5q
sQIgyo2wUiwCbZqVcw1zw6RpoDoEk/BjwqesuIM8KhcRyxoANsGsR0eIx6E0lkts
YZBnYewy1WX4rdKDTSnf7tZpJvVf92frYqagtERjtxSD5F9XMR3xzPArwiSElC6J
8y9cVgEnsFXU8JmStEghFpXGrLgetFqplIH3E381qxQO2HKesWFIIo0KcRa7FRVU
hrVXDMbjYCcToquulXZX9X3oLMC9gtxItDseJ56fVhIzejvgd3VjUDj0BX/6mAmF
rnFlg2HO9x+yBhRpJpGugsQMqI/Ig3QyDiPUNz8F34FT6DCfzyajlwqky0yh36Hn
mdd4J8C+DXJ6piLNALHIyAe32siFuwNS3yur+9WXCFV5lNSAIh02qpU5vKqyP0fi
r719T9IXXqoI/Lgc9UTRx6aMI9489eW1k8uaOZKbXBlBbmbuaP2oOPM3h9McD/MV
a1SzbZg3gpW2RoV0h9jNt5C2z+FXra2a7mTM0JluYjDS6mGb3DTnXw35501c9yt+
R5OZruk5xprDnfo8NvE4YlY1Yw+pMcwX54AORgfkbHPRxmkW5W/VUIae5Cz7JvAW
kL7wAxQ/3OIbYYhP2QkADCMgggNgH444Kw0SWxhLTPoh0ZwnNu0qMVR093k0NnzS
jRVyUMWdljcvawf3NHi6a4SrRvHHurHpftVaJem5NrJCuR1b/ukDfH8KKRinbKHA
Iyk3eIXXMfwA1r/ub7QBuuoRGXqPU4bufzXDBkDvjrQRK7/htldvx7QwzqjOOalc
k+WhktZzGUOaQ0N43nldUt6+keVRWaSDCYBk99v3R8eFzxC7IOFxsG20TgH40O9y
hRFj8SGbF8e7L/tQ9TuhNJOYOf7Z4UGwuYeOaTJ0PGZ33D7K9L58BQpXWhgZrRtb
A+xiFCKvKIJaRcBrWQuQE1t8dyLGc5Itz9xRHBL7zpmZbCWECvub1iXNHT5DG+SS
+y9cWrKsd5HEGWzP7XRS9RPRiN000aTWtl9N8l1TR74HB1NFA9yADP3sqbV7cqvV
MoLFtmNRlrhHPLYa7fugyFEZUNGputhQa9ia+XTRlcDfLxgnjzbza/WEmCOszTfo
bMelGYxfxxxuMRNbnchbhWbu+jespBZcPvgUYsHtyow845qGtFXvlM3vG+64ZoFP
63BKJ1gX5R/65dsfzJP5XIQ42MLdWtV1Re0NOQsqaA7ckHa4i1jcmIYYCUogEl9Y
aCWVtcmPd4eChGyKz7ayJSDn46kfcqMNdHns6gcnq3Ok4yPxCpXZj//NwsiIKIRI
2oEOp9psuOx2RpOPN92gcmo9OgRqqOTkyMUXYVy9qUThrwWFCZCl1raiftyEDrQx
iQHN5VkLZIhhlEn3wNnZNaJw1ufljvWJdmOez92piP50D3T9j2Nr91fy452i/Vh0
VIdfBEaIM3blh8sXKuavsZMTV2yTrqQEC9hswhh9mm4REo18B9q0XSNPBjrZs+vv
fqjJkR5GBxDEX6Qdoqr+n7dofT5TAEic96e+fCP6Dlw1IJgYLrPLrKWAmvfw8OfQ
XQgX+rFm2vOIy+MKDe8GwGwa18cASWY+B4/V/PSLP8DKgJkwrmvFQDvtDUch6gH6
UZuJmzhJd4OE+sBF5Q1pVh2ZtlzhTvdreRqRMZva87Gk+dOfAHVCqtR5tw3SoP9P
xfpV1KnONnwepx9zUkix2YNRFTJFWwK+NzcGbKMg6dNBxfQ4ddC0uyA4X/Eujyrq
DUCMw4nTfb2Kp5eaprGW/AV/D9qLTqS7e78HbwzTDxYFpdXuqlSUVjPo7qPjN3ri
Xs8h02H4QWM5TdUEKn8D/6eRmiExE/JsDVKawOP/789rl47i80XTaW/ddVrWQMWt
Whr1Z8cMLqi4sO/eyDeDFEAKfqyVXcePpdRNYjWPe7SHig7MEDQ/+fF23rSBdCrb
taw66kzCNCO4tr1tbAyUsspTtBX3Gs6ez0yBrNIuo2u+Qs3a3ZLH/3pQRxZlrjat
tFiz7Da77/MHX6bVcmcUyxgDLtKQOW43jmKZJUgnntLy0yHGtY/8zASAAyfRXGCZ
VMOuZLnY2JzBLaABaH5GKnO3OLwM51JlsVkEa+k7qPVyOFJ0svnV5pXYtxOILGxF
GwRoTwkIRJ854MhoHTGuy5HyYsqq58/hoPiHLXeU87Ay/llvpweY8MB+diORgYoe
bEHXbwZ8qpJw4JZZ/dMcL7vDBVOcRIngGUSTilTX372vsZqrbJzOfROaAuw4s3ri
KFIWETQZlhVv3LWNmbMQBUHnnKPI19e0CjMvx0/NZDwX/08zcRu/mbIz82JO8OOB
PrI+1rD+k0o/bQmXiPtfde4+HlqJDjbgqL4nL+l0ckIjIIR2cjRxApgIjW2rQhmI
OYwleDSymGItF3hfQ78vy4XRtcZlkKnI46xprGLFY4HVFuyNBcinUyPlZcFsW32A
gwpEPt4Lu3X0DXp3DVl5knwrwVdc4jzh5uloYmsnca35vYEKMX5c/BKGRGa8i+4h
OGiiEhMFGMpBzzHymxwWLIMYjnZ4hQue+vU1WKyrwMqUWIxGMWkX9od87Lf9CWU/
BUZoUYEAQmHZohVSzmvSfyTtTs/lVLJIlbY3Sr3v7ti62YuzMGvQdgDKD5cbrjCr
w7aDBPX0NoVmB7HMMeTkWIHlfwca4LL7QkkSBaVzAG2N+EmZWppjOwrA/ikqcaBi
IERhiLpLE1m+6YTmQLxsUOAMzp+bPyKDJ8a8ZH8iazvjI043MGibkzyC3nmuUOU3
vCtzqKbUlMsosMUkwoi0mJCO7EGM03XgGp9CB0WjLUHt9kwW+CDI1AYGBgwmEK0S
rE/y25Iqz1rEFTtQREOjsUAAKKym/sZwyJbIFoHNPmMI++949JeoBBA6Yhwwp+2k
mIFLFDiqFiE30+dxJ3q6M+ZypfipllO7ypwI0WEQYZV42wtJ3q4r/+G2gjMzypMu
frLjnaVP/sw7D6XShYdZQylDCEVV4E94U5vSflPJp+31ZxnGiMVFXiCHBGY3neTH
OEXzNyLR1lKVm9wsrVwfYxpZ3/+Xv0eLoriPcrEAS8YGIR8Le1yRsBHLSaOKsJQW
SVUXvzXPuRruPx63QiVxFELi8vA+fF/uNa9F1w03ZVxKSPky0y8m2VdprDQ606G3
WYlwTMHulZC2PGkTLt1V5PK0wl02giqzJmO5f37MjING7J4MAQFGvCoa7h/LVQIg
dEV2syloUiegLc8CklkIJdiSE1DhaHJqAfXNc3YVoxCCodezg4KWFCMUT2bk/6Z6
G5ADI/CfJ9/k9QDRjUB3vouVCjMa6fjYSl8Ui5G64LKfht812HMTOH8GdXqHxI+9
pUdN1hewtLkfQcOwwuWkMA/wqBVvSduCMYk5D0gCQasWNuKJLsGyrxDlIzbqFoDt
ucgSEOAP6OQ5rVrguvNKqGGf7+h6o0Een3+XAj8U87js0JWR1Pz0K7ZN3LXebitM
8cxu5BFPOXaiCPb7y6Uddd4HbEcVmcrwOtIkLd28GE4MJGSxN/S8VEhGnfslKTDN
A6zOUasGN7FQRx4epVyUBn3JKeP9JqXjRF7MTSJEZXSJU02Obf/wuVrkKw4XtzNu
n85n2UztOt5fxix3wGyWISklOPw76mSwQA4uC6IM3X9qzsPoz0AVc4mZeqPZiE21
NPunGclPHoFheXVA9pAuqFCS5HKs7IfK4mRndxhXdASdnvUocWVdL65es9WZMgLX
BcLDuvMN8rf0EBYSKLEF/Q3UAKvjAuXQEK5fMEs5AUtbywsBNdDnL/c+5Nvxs8L3
3z3k/ioOjHkIu+837v8gm1juoEUL2ghZhomEqVMIjaxKpUMo3ewDQESGXvJBycVP
5zGi43heUtcLzL9L8r4dgGLQeQmdWZfTLLh0RzYRnHYhAuC41Gr5KvhCLfwclT7d
2ZpsHxFHFwov/v5CC5AJwVGyj8hRGLj7m8vXwseTjmLwgtUbnGUAi3e4HJD9kuBz
HKn5PMoFmp8lH+JIcIGQo735MEbsl5huv3MQHMYcdCFVsltjz5vD1MfjW7sjrInq
ZoBocbk+RrjLaor4JEMszBwIFKADptuLzGVJZs7SfFoKOsF16W4JDesDOvcZ3bEO
kegEZAvHp4yD0HeP8XlqPogs/3/ti7OdHIjf6BsjOj/gzkAGwDEeymLSiKueN2+8
GJps4MBE2QyVLUAhxeCPMRGHWPKswAT6hnmiot97IHtSqG5pP2rRYs9YsE3ZSm9+
B8BZ6Q2bj6Sh3ioIGZH2vq3jRtKvkGTy7sRD0A9KzS8ep1+XTiBilJ7RzzyZfqIk
5rDcBrQEAx9rkEgaPmrKzeL0LisZlkBcN6dnAufqMXp8xoaSNQelP7kRdqR/XqHI
nllwoBrGm0L3581N40wTg666tuEPMSXj6PBnrEwQy96/Zxw9bBhrjnXOlk6QfMqk
eV8HXgY4S1DDB2K6gY9EypV4cI7DjDVVs/OHDAR1OZqF3hk2D3DdGAVUCpe8zTVF
2aBkijDGXWxYB4as1rnFwULqlGEL996IKd2h1lYSREyiQwYbih8CH324evmr67bZ
R8KWZ1K+mk0Fy+5U5/TG5QV74D/iCyW3ih8RGegHpjWrEGTp8QQJqpcyHIoMMVU8
lEkjvBX+CR4kp1plyf97njCFiXux5xlyGzNxmhXGFWjXY7RqxMuCK1a0fdltDZNg
gW3yAQobbdbNSxMUb2PFdz01IaVhZqCZ3YqgVU/aU3SQXGvWF52t/jIg/yI/z3EM
wZCg+zZtVHeuEFgjABMobRxgChVdTC1x3mmjmloSFgpQTmiJm4pkP/Tc5COWj35u
ZbMcRd9iP6R073QJr87Mj55chS53DMVZ7ia3WbyXcQJttrTBpR7U0GLM/QTUx/BW
DrIYhwheiiLCV3jC9ag6D49fBuaZtQ85yp8L/jLwv8l7g0vaeHzGFDLkzR/c+LQD
ujNCEE92gaWXyLrkdLc9ZcdHn9GtpulO5ZIeVXepjt4yLpLVcgnaDu0rttSG3r0R
NO2TXOCpnO4bLmSEcexw6AWvWvUKIpk+OBcIp3s4WQa3KWxRUZZ+qYv+MjVoVToH
OBXGi1KX+CAO4qoFv0JSlU17poC00x7vItXvXHOJ9QJWFecztsLu/tZRAqY2yeSp
G05xO21oFwdltdvQj06NaMf5Og675tikOtoRaWPFLls3t701duIyfamKUKIg2R1G
VVEuu3weXAoHtvkbAeNerb/mHf0fFFYcTEcOEOilKixyhsftE1lLMvibRDeCEA72
v+4Pf61FbrMTeNIJuRZYxGWzafvh2atmBU80kMp92Bzsww/qhjAucFIsDEDeK5vN
Kwutv/ifGKr9TQ/WK4W2BlR7wDCtKsaeWx0sO7qmC1gdtnDxwrBXtLPLoaCU9Qtr
3By23qlFgCk5hooB1QJliyWwqmQJ8pyzsdRPQ/zPYqHt0CagbvEeKD/o12r1Y5vY
EsxDYoKreCkhh3V1i/dkasAngeCueS3aN1fwbbJvbSQ5JYNX8TX8vYsKx9bmZbbr
RfEzLEI4WJu0MyTUUvp9EABXjtY6IE1NwNgCgL2IZXx2+xVIxewe+yAQ3iWYZuj6
X9cFhAQ1LFUDyPqFOrsaFZY+/Csy9GuXuLBzG895Gpu1LfWBse/ap7OuWrnPmr+0
DdE1ecMOJBy+yRAIZak/cyr+5IhCW6zR7AOAFXwz3bEJDMoCqvYHD9LdoQTTkMf6
DtKrVrmuzcU7L70jMRtcUN8/dUfhD4Mdw07rWlExguZ0+ZpcdD9zQUmCWd5bbOKg
lv4KHFE+YzEXMkn7hvJcsSMUEVTJp0NCvvK6fCPGyJVyCyEgvfCnb/MFiI3z36j4
YBTX1wc/N+NdgcO/mtjKNXYHk3X3KdeIWR12iaeUY/Z3cFT48vwecNBUBm2K/RZ5
StAMlHwLLYHS7PVEKlyL8FVZIg3QX8c3weeQB5RlN8D5x/BLa1P/waKlpF79hNIj
faWW27L93ONlrdCLKB5U40DwkScQoX8z6mOQ2M/CG6DH5YW7ElHlHrWTfFLQWzH0
j9nPwEy5KR4FCAG7WjgIkkkBApi4cDNZbcKKlQ/qGxyCbQQhf2YqPPXFhG9DU58P
J4bJCDhAySsgzDaeTp5IU42ie7YLYDdsKlmN3lrsIxhjBCVuy1Np5tz84t0wEYu/
lYjH4jI1ja9n9nlswzmjWaiAd7gFusCbyFV59Ny//DfPzKnwS7peA5/N5VNdDXLK
F0GMQDSeY29Pm6kApZzuQpfeREWeNSw2hbtwH7SGTf5kL45Q49gRsBrWRf0tI7v1
7cpjAe2mR3CeS4s/a0wLBGsIKzvmbtIYTI5MTS7seBEIDM2TQWawY9fjXgymFgyB
eUWUbKGXmXgkcSVOsAV1F7qCYmBZctujsA6gld+SFsJWhCHfbrqjVl41AglRrEdP
zxrSU1CIc2rdCV8jWYmC/PIciL6PioSau0iTKTv8zLOMhHR67uEOuwVIOtubM1jE
RXFqkllt4ct5o11XYN5RaZDvtC3sSpDSvwQa1xqUKSAJZI9yAu10spDBgZ9fU4Bq
xDic1u6N4ivwGk1dQ3+z/K4MvJYnviSyQmZCP25/qwKv1I+EsdtrH5ImGViEQf/7
C/CB3/upvjQ8lI69P+lNPLmB4mzScAk4NwgkwCBsRR0uGWNFLv+2SZD2PgE95gID
cSAGifnAVHUb7JgcfsyQfsT0XKPWcg9AtMak2jWkQzFM03aaoa6eXbjw+A1XJKEF
CSyg8jl3IL37Q4aJyV37AmTQhTw0iY/rsY4GCvNIlU4jQFeGU91VTDqMzNmSHljw
ak8qc1zY66+c9u6SLRs9cYezcmO4bQaAY7yHDU6gf2h/ff0CBxc2vchY6NwZY5kh
NjtTjPDxjd76XOZUWAuc1kYa1v5c/2KibR10I4jsBe+3akrGRbUIGkwgioESfbJW
cAnIwH2QzxxH5S6z4UVW6+8JpFdsMfD7PZBSUv+D5ZAwUEW/DZrU7c8UwYesRG2d
LwbluObEQVsJ8dfUzBh7MSFVUoCug9mPfi35oyxGJ4OnfUdP4Xq8KkAZaISxukTZ
16dGtxwOiz2CpRKZR2YO74O/U+3iGdtDGHjRFmwN7NY5Pv/BXGC2PE227gX5M9BJ
WVgcDzQwVw9qTxbgep34Y6crOAywbu21kZlJAYSOhbY/fbx1tmZOF1r8lyF7MNzT
4+XLmf65QiczhrSTqJoalDeAo1ETQHgwVg59bgMnrLOjFNXfOsp+nl85J9mRvyzo
jmkv4jiUM1uMz5KFAUq9srHFVEM1x+v5jCWzCfc7/G3OQs4NR3AJpJgnh9hXIdG+
+f7ffb/VtPUI8wNS/fpsICx7SMmbt4xX9DBKy8HdWKm8PRSKZTNsY/v0rhzAaYFE
FjRkl3TT1HZnET4vCrVs8FLNj+5Wdht9WzM7W3CLJoaf+pzZLGlQam8IxtBOubaN
fWY3UBnlxzI81vuxCNeFAmJMsLa9zp2aidijGRvFnEZAhTCQgGAD5+YWj18x48bW
5XbAGRF1vF8kxy4c3kPjvz51sxH0zlCynMeJ+kUtYBQGD2htE6l4zWcMzXU003Rh
8oTS57ORNqLfvk12Xxv5srqaS2Mqj0aGhdOP2n/WW1TEWY89CUNFf+0X2AObzV0I
1sCnsm12ziXwo8NjeLJBjMR/1wQrGDizFGbgB7b9IxA2gBIX36+7/VGUQ8kyH9A7
7Ic6xswj+jzglNJ20giQ9Svir/MLETUAToMvCAAK1qTPUAN9OFGNc6Ovd8TK95Ea
J3nq/VmWZ9P9J08SYt88MFSFCD5217EXFQIc1B0xPUSDHtag79r6W+Z5pYeUfNMp
3VSPpwI3WEJ5YbCVooKTCqH9evf1ncTx1DjScXGF3NlrecP9Jx+hz1ZOZPhsbR7X
9DtkEOl/L0Tb8fA1vur8wMPdd5sFtbKU04lWWlmRssSqif51ueOXVpbNF+tCnYMr
Jz0whRn9jh9tvVUowN1J4Rr5mzzL16Bh6fG6QPpCXi1pJOUA6ALeDZFZo9IeWhsR
T4zz5EDFbIZbxMLwsgzJGC3NM3Qy14qUvfhtR+qYwPIq89FHBrk73fRA0/1BOeQs
KDlOArBuHWa0Q7StU2Y7Q2TMn2Q8gdXwhJOKhKNloWFkVjSkXEpFlhp+Cj9ls4Jg
se6mzDSlV8RxWHeaCCOSq4FvzFZNzZQSwd1jQ5Nfe3+XQhWEIqm+PcN/5AJ1Q6sq
bmera2KeWWiZ6IheMnXIXbg6Xfb5IJoaUayt/2yYFBB786iVxppk+USJsKDVOvPG
1SiI+Gxcu3zTxUdLmrha+XzQxNMVqajcCe5/CgmD8GZvGKfbz5yu02otWwoh5T7q
PEtyxmnBYZ8T77fi+nUzgspqnj7mApchqk/LugzyD3oGiGrBp/f8h3X/bGgPOgS6
Zpz93rrx4wo5PN0GyLmSSvFvEVR22XZ05yTgGeMNyaxi2/bB84RIHo4NR+H6fJB9
EqRdnxboGtbLx3B8kD7WOtQKxH6S+fWKxeyCsjmCft11QXyax3h2FoNysE+E0IFC
DZrTPc5/HmSZSq2zBoSFxyzTSPoUXrpH0yPjIrU5aEHTSZkVAwVNPESomo7MOnvD
d6RJ0EtGsq52IMvadGnwfVg6CewCFFVZk2RkH/Jah/LonapKTYrKf8osNhbJZ5AY
UBxMhW6z/CJcNgeR27nLOhyqCH62gb0f0KqPxZU7QpxjAgPHMIxhVMjjkGZz+RsI
kK/4KPUhMAjTKGiQiFlB9Hvn8Biy7N4AIRC1w+Ldvde4acuO+uQB9amvOV3J9R//
mpZmQQxFBkApvV+Nz5TjsdmtvuPr/urRyp7cO20uiv+2vXVXis2KFZxBSy4dzjuo
lk6iLr3oOi3YeLGy7ynI+grfK2YYyhkOPclXzugw1B3GyzweL3b35r3LO+H8tUPb
Oy6OuC7l5+z43ASJ5hAhyD7KgV7WarEvgeagRWCnLHPgoRIB7Bctd9VLC32FP/if
zgQzvtTJ3UxhnYJ7dKhe1/xKLj+vk8AJmM+cQb0yhqw0xpzuJRwrU7VhB7ngsDOi
IzK7lpO/FaoJlJli4yJDEJdIa2a/4Xs66nSn9Z9UzSNt/QlncNzpolCMiFPfUozH
QU917PAK28jGTZPUD4YSWHLgwEr5K09YiUbbKhC+SwS/LsMQO90Sxt1k9FciN8W5
nl6TTgJhBr5vPRf5krKIf7cSyOW0KMPnNrfbqxwYK9DyQTzWHwIO5YgzT1UBmufb
ZGC1jmREPUV78TA0XfOvbBFHoNLUrLL75C6syHhBkJu3jFcHO0M6HZ1DrW67msZ6
VfuE9x3B1zgl9mrbfT/T8K1K2CD6AaXKtnEJ6a76wq/ocOK1CspG3iY5gXloyUv/
FlyIQPLEJd3V3rkxwdTsnHUMT6ilKa7caBejBQybriDcqZoozFbg71GhJcF9lFWN
XDX4jndchbuxG08m+G1r4S2YAaJG6DE0DnmJYA0ozJVOu27q+Ee5y7dZJhIuJ0aR
0yz54ctkDdIfCL9MO1Lv6tBzMlM3E2EbJu+IS8dAyP4GW7cpB/62+xnnqZTHskPk
BfVVoqLkyfzvWurNRs5DKxL15NS5Lfq2dBdSc97PyfEp4o0Um0FIguQOqQylM7Dw
2i0LBA5BdmVcdXJY4eIsS1bHyH5rrjlrfkSsW6YRJwKBTpTSAfnyccBOBDLbbwv5
OA9pUyz6zAyPLwPPEsHZgQzimjjzIFIBB4fuX4/p1hgsP37KdIuYcR4aNdVXd65/
nTGA/EYJlU+haM4SWDaKYfBbcDopXH73IowkzKHk2lmN5ps2Wk/3c5AhCfr1q5d4
GcpvJ6gyWfh9DJFJi6Z8YRUKTsPa8oIynW2iZl8c6IgnGKIdabnIGjR+8Gvly+6F
EKtCJQr/8OPsN991QhoG16dLrSciFlsD1EBMUnI2MYRLuoaGUAnVrdNuyAogsQdz
uKC9L3mlZ04NZxeOE3KVu/U+4pn/XJQSaanfMOksRyScCOktDixViKqmnyvfkR74
QecFgbq9FO6dN5lA2MLPJH6tq1eacuzQ7jGdSIIyjzqYdudsekJVnwZQy4lMov0z
5xTKwK3my54PpdutwPOyAai8Iro37TEwZWBNGVYoUPAtiKXJYPFqqnnSiLvmaT4u
1UNDDNhExuYbRmrczDsqj61V9EC5cffroPBAs7ZeNIHLT9rqRean3ZryAEAAntHE
ERMCPqJjuKzkXl1gw4dytk2FjPBcCEsxRHPbHCRL67GQ95kQ41pOEHbiS5iqzQdK
Q6zc7mLLlVXas/s34oaCvwHq2Wl16pO7EWYJMwZXoB/Ox/m5FJxhOId2imna3smb
kcPD5IT3rZZBIb+uvhHNQtMzrDyB2p+/iZBInWqq1VmlbxDH4E0DWk4Z1ei0KwvW
UenkzYJcgo3ghP7tkDCxPeyTwrf2xIIaAXszomaidqwn676RcqHwp7rbGdyEXq3L
11qQ9LReRXH4pKaSIDRQw6xAaDT9vcHEo7ftaKRy1Vih6FmPB54MgS9Za3dLs/Re
9zw7rS01VyoFk3C+2U0DKu3KhvFcrZJUeoKxK7XffeyPw5Bv+IV9Zsp6S6bXdQm+
iOYL8lHbTejjwQJyQN87ZOzkg83zTtYW3vE8wWOp8NgV1pCkjB9mvlYcz8h9vbVq
sOyd9AYYbOoW1lv/G1sRxVjMxydiXKgci8m+WT8wNXlxz6xwl7yK9Cu1UoB3N2u0
xWYM/nddIOfixtsQ9eRhy9LGAYgg/wlG2RxuXtJmK1BIKcFaw+gn1oWqDQoaEDa1
XdetUZP/yyrH2P/jtk9SzGD2Y2OvbB1NUsDlFEbJKGghwt8BTyZMZ66J342WQ2o5
oFNhnJe1M660ciKH0dzjJqxtmClrw4HmxoTqQX0e2UckAVKbnnGbrhLFlVhASI3r
/YL7r8hqU5Uz4c/1MMwEH26uezIZZvEnLAyD91bo+htSIn6KO91c0WGdcZkAL308
Hb8bEg3lHg5zLHmjYlO6OR3SrfZwsV8rAZNy/crX/Ut684gmNz/P2mOAT3I7SR+W
NPt/OsvlYWZ/sWh74FuT0+soA1Lece9D2J+nSWdx8VrrDXqqpSOhbB7kpM1MYauZ
VbFfNXmFH1fRSUK9rdRZZG0U8vKj8ebsOMxbZUYgl8kKSV9rmd0S7BCR1a7C9ZCW
hwYzryupYttKHEKHto1vnsJL1jey63b4M7fMQUTYcNX1S9DogPmiabEiXXU5Dujg
Y0tGg4zaBBXv3r2CxM/plHdqyfQ+iqAlg9oSzSt4gEQjTG7GiK3mc0lSVeKuDTTV
Es2GAh7cCnojbQ58bcPf6+y/M9RTpYb8LoiGIu2SF4vgH44/9cD7ZFXF+KlgwF1x
qzbsY5jqAtYX2aaxtJ8naV9Q8hXeoHoBSTCTtv8FW5XZnEhPCOdqz0dd567lKx90
XbLfbWWuYYHEmHsRChhiWPWK2W0ems1j2AYh6hZzhYMZCAUvZvrKTqSEg0MkJhwn
NLn9WVpRlCnPFt+TWH7UdeeKBa9VX3KXINOylgzY+CH2jcmiULNFucRnD8pq0/m8
sLDQVIwbWxA1uo1zCT8O7rsk2ik9aKp7OsY4gBH+7kTOAKntTNlyHCBw7lMVhs5L
h3fEihqSITbtsoJCPvn2Hp+i/755uEBS8weEKm2OsUM3V7pjT6Sjf1TFsuhYTf1A
/zBcqXsuAfw35ytA4KaPW7C7hAsbXnpSHcFaHm0LgaSOA6r9YH/Lvm33Ir8+wWHi
EAvQZ34PNiMpMsAEjjrriqOCZoLJKdn/1MkNet+FH+8srFWL9xt7IDzJBlHVQknM
EKSkUo7HqT6pdWBXtAhbjHRUQ2tu0CMNVtoaHvSMRgtWsULYiLOM5hZKp0p+5n5d
2RQRHrjYB2HKAZnWxA7hhyWoia0gm1xMvItMTWvQPpwL9UDdGV031o7Zw3YzQzpv
OVoHqWx2a1Tc0/2M8V5kdo8E/CDw0GSuAAkxN1jX40B8qLJpUhrokUj8ivvXw5fS
CYZ0tyc0h+UAxvQClpR4XbpMjI7fK55Zjnq+C43kg9cZQExeCLwwk4jiuLz3OJUt
Y+38Vh3Yhb01tpeqZijr3AazPc8PTl8E4zyZCyZXnRn6+bw5ZHB05vLl+tKPKr+Q
yM/YxaRbNQkXrbYf1HU5ojq3QESxwqxbEdN4/s1QlseX53Xf6gw6u7JgwNOfhK9t
yNjg4v8YTVk99zyRfV1Z/xlzEoPRnYTpWLL2fe71OYvIC9V0+3+FVe3O6qEIwGFA
3Iwx0Ov4d837gd82637oekgYw7CaXcrsd0SmRHlXgbu0IMEc6WrnbR7PG+1mO2ym
FCMxg1mD/rMAt2+pRzrsfcqRa7JiUX/BULE2yaXQeXjOvUbqi0UnfKQZYzEfEhoa
ceCxtOzXVeK7YCywLiyI9pyuVokxLoF++O67fvVRPUANGr0NXnYUSVXnaHpih1gV
bj/uJFYQ/v70x8qJTdEwqwqQSevEGGfrtEEexEUBucRPbekSGHsLxM6PUvCINdif
hcdT26Swn8TiEFQzbvLA2kzYnFI4ID9M6BNqnsC328rHiWt76cQSycN7IN/pZBJf
gX/R7wHi/U5LipF9V2haizUnZmZyG/JwOO3icPZNzTKcFHXBscBI/bTmZuCMPVhk
mto74r+puiAYNfErK/neXO43W0ef0a3EMZQZAnBM2maqrgxU+KVezqBTLxLFnVS6
KzNcaDUDGwFz4bA+iKi3r90flqasuX07WNtGk+e6Zmce4NAd9V9AGmN7sZqtAElN
P+6d9HmWBqgfmzrDDXreo7L+fk83vcsgOGrtV37r3dV+iB3XNWocbRgVUI5/e6l3
a2Qybjub5QRTszSIdJCRn/AnBHfmsHbbsr9s/hXctoZTdMe/b1p83F/7upcNYms5
5dHhh5uM0p1b6vMKkVgt+nNvM/usk6xZLIjqs2Gnvs0EVu60tOYkFd/JJ/ca59zO
lqYPyAViLeHLX9H4b3bt2MQ6dciyUhMnXrb1ernaYSDlUWsUmu4auFUUEEmCF/x4
WHXoo8Vk7/PFOpFZZPbqS389z18A9BPjjKEdHUa3WxUJQJH6DDCUr9wo+Ol2qKHW
dbhckpI34RdLTzibn8rWZSAzMWdvNnecczOKOFDKZ+AJ72nbfNDX/iKZrpxmz4lb
dLHQHphBxOLE6ZsHYgEW5LYEk5x5ccA5b0aFVHPfARVazBxlXwiOubl/85LZNBg5
wi6RU4oG9lLMnizng0k/Qv8OX1J9r82eShh26kkrg3HlV6kKa7mbe3+YGOFW1Eqs
3k9II8VlBLmpD1+tWQLbY31AHoiAQypNIoG1ak+Rg8sPh/uEOEP3Ph8XMdWjnHCv
+KJo4nE9vDnJPZOwlqpkTlcbMerPzwPHAvVyvM2/pOHFrd3KjEPN94OCTK87PAwc
ZAnozHM+L4XM9JrdllpIqPYT/IVxniBqpjKi20x0rAYErARMXXkIEMMDhmi7rA+T
pZdqp+u+l+T9fJnBkE6iQkeG24HB1Rr8NAuq4ojJuNunJfzuzMMUFDQ1+6DWgz/X
HwMgkoUX7ASRwzeDTszFCAPJ8PxrNaGsHXbkMu2UPs1R6JNl711353vRZ49/5U/V
eu1QGa+Bex22ry4ovtVsPVWQkV8igs2yxK+rwPfFbrQKLul3G6lolvgYt8/tDi6H
IocU80TlIGrj71Tmlj/iaVac8gjxJcVNWTZOmG13+SYB0Lz8KoKMxmOqoCntjZHY
UEZCwLjBXUf/G8IHhgVRMgMPUVyJ7UMogCuAAK9XjOuLUeGtw8asuKCvsaSl+YBi
28MfN69a4aXD1GV4CUC5oKcy5LuLPzfA1ZayLnZBXrrGbPVU3MmGf8nGsS/AfQFU
9JMBDaTraQ8RnFSt95V0fPjZOa9HUtOJmwK7vSb7teetne0iSoLlQ8SpMONML3g9
s47dRuts8S+31+Juk7LurvPWwglXRQxGvbbfltRBUYfz/U/GYrttXIUtPvOA9ev6
Wja3WQ9ZGTHZbZFBFZT+eNzfiasmV141UUYxN1MjUPBldGmbBJpXdQ9smB3u5Q+6
ujtNUpa9zq5KvPDYtD+uhFyslpVKB6icwbbnQEQle+/4ZeaOhbekSRD+00HmIQJ8
IlL+hiU7o6ne9xrSqjD2+dnfgmcU1sNHc18XIkZMxjCrljy+6QT+7OUfBsZBjlRP
bc2HsmJ/mPWQrpWrvMBPArcF8LWyWF8dJ4BBs7tFF5UXDcg4Rfx5jDXWV8ZmWin1
nRGmScT80g7WmqnLqeKhUuBXJcOYmRkJz6+JyJcNFmtrZhfSUvcJ9r9sFOJl4f3j
ReIaA+9AoAQloYgHSj98U7detcIHFBn3GEWK9H19vGCTq6A5iuivnBzjgfGJOobM
Gfvv5XZjwL75UEZP/bQVecc9FgM7iXtVfkZthdy1NuFGVD/62SMeV0kEHDsL5O3L
U1+MbW/qW0nZe1/3ZK1etO0GRg2iawcBjwuQz/HB42tSAg39zVjG0eUELARAyCbA
ocjnQdnGLqZc5Hx7qkPguHnE6LRA7k98aAxn0UUJCcXiJA+pAMKiDA4rfNVBscn/
BDK6ZwUkr+0JjJZr91uc0NwNDf/L5yIgyu23ThW8mwYh13+WwYjzoX8mkQXq2ogP
Rz5syPe5Eg/Qh6xSp7cleqW96JaSOakL1Z+KT1HzaN/kF/rE6k1wXzXF+ti7JSwk
x273NFwh1lelEx7JCQQLufkaoPXc6XTva1tT2YZdV+SJdhgeEbt9ad56viMGL9W2
azkWRBQC8A8ux5gaT7qGT0I3FhzxrjB6ea5ER7mFVSRCCC0+f3/DYeqgIo0yv9zP
/9RZre6j60CUBgU2+qf8V699sKOuHErrUPUQEB+SsQXr5m/BdK2DsvdWfhZYaxUc
unXLO3o1tTyVx5Ty3m9cUREQje9VJvHjAVHVLmdMaQqGSNfj2ah7Y5Wis9dcB8O4
clP2yKoiq/Nnr3FRdcgfcDDOMIQ+ss76RFUi9Fwbvv2YoYgy5Us153716weqv7yr
EcAulRM7DMJVgcH+WjmMJKDINbxMJVQF4dlA+jCJ15orsi8c1BdP0WuO8/L16txe
TXS471xWT7J2h/1Xi/YhrFI36+Na7Mr8eHbA2hQUa607y0G5KQtUpsQ9my32Qu3o
qi39roGushxf8nBxXgMSM9sypdLhOccGRukTIPsWTH6i6zWnuRuKe5kIdmAYkoAD
7vGxdsFGomck4659KPNI5RJG8ymEkqid2dW/y4yY6f2ry1bUjr6YXG7233O0I37V
7c+skNWIdbhWtSmRVA9kqo2rzAPpVfUKf2YH5ynI5AXUuYB0wC1dwme1UJjCUQnD
ApXRnCXzjLFEJRkqAbGkMWNEPrLHVsONK7SDmpduSa+Oqbka7YB1EX+09gspYkUz
eNa3DwD9mxX+gzezGFdITuXVsZY0XAyaFwGdKLRWv89ebu4x5Y0Z8NpmAlNDIXmn
K5yPI/zXH/hnjw5cM5k/ZeyhEsepCMaYltSmkh7Kg7ufd+B27VlwmgxArcyr+Smf
dMbjyuX9Tmplj1z3CsvmwR394p6g7IVydSL3BDh7TEbjdhWVy4gNuUk72BMbojDi
tT9Jqe8L6HaG+KwNkW/fGWjq+J6XakNEU0UtPd6ut4TC1NX7GbjfjLMYinWSdzPF
b8v46UobrPMFdVrqu+1UlJXp4ZknES+w7mCgLFENEPr9EsflocT0P+Knb2Ume8O7
xDDEKxDF+TvuwC+bZYdF7GUHqnsPcM4aKtfJozqcku/klQOIJwgrEtkAGcW7dY9M
nYruyGKZWtDgIZu3FzKYg/X4XR4yHZHOBM5c6auIJZvyH8wGpLb0ORZUBvJr79wh
SrFU6F2+l6ZI3IkEHkCIRLOHI4zGJF2ME07q5wqLb5eC7OfeZ032pp08RnexeIDm
1o4aBB/5jJWQfySNxuuCwzg6Fm+gzIIKCrcPAxYfCX7b+z1InbD7tfX/pXmI91fv
Nyys0w6BsLmfGBpYaGSGzoFYJncNjJedtxwtrfZxHyFcbfGFN2TsDZ1Q/fBZ0RBv
Pr1O9TuyJ1cnSkf7GybCaErrJzBgPqwFHmbakB97DN6BJVNhiXfykn3XijSZhfz4
wlQdezHA6T/JTN+856JF1k6o0nbzHuCv8w0+wpbgYU5lUrjL1wR9O4kjQ5XZBtoq
2JnCWGS76r9na4tmGe8gEit3Ct8GS4Q7jo8QIgEM+qUdcVBCIVdTZLfcphkxuay1
QPn/UINOBNi9Ljqmck6xoMNukDUrfA3sYReRqVsWitHQ6wviCSrHLUrHQHfsfYFh
4S1yb4CMNSpwHnOLNOmoy+cz7ocCs1zGhcdeXREiSGfHu+au9Ee7+Lc29o0YkB7M
RNj3njIzUbYG7XegvyZaNa9df1czhMYyB/saL0I+6rkrkCfVXEvLab0IvKBFtUZ1
7K6TTGLx2NCRm4MKgM+RZoFBqm7ZoOqQ8k4kwMr9HJB1su256kkycps8glrrBneW
xNKr7REslZ7LwIOPkYK87Kj9/Bh9/jmr0ryhdsTV6L6yg96gWUqxqSd6eKBad3q5
tG/pXX5STLoSblrfIzeXXi4UPEji7bdPh7E2gXNo34vEqFBD+HdKFPW518PECM+5
4tt5yQYysJTBiKUfOD2nbGQNno5rwSeHAfcMPjgfZcXr809kkLejCW1vBUlK+/IP
QKbXADNC9f+qSyIQR/OWLHcbYy1jltsP24x9DqhCTDE9USTJP/NW8FPPhZz9dYFR
6+ORWhgjxNYcoJ/ldkzRqoHTye2Z6q37mvvyrjna6E/1qsw9dRXIHurQgtnCNXMG
IWlir196pILL8E/AsV8fJ1yi/LrIVxLnFF5/1cGaN/wLRPbjcjuhBilsbHlxLPX3
KQVuNiqryDMIbKR7h1IdhR1RTPFGsgijYPoOZSsuiNUd7nQ2Qfqs9A8Qan48cL8Z
ctYnF1QDmYrsmRER5v6x0j/h7x4CHsQHYa9ckWrvhCAhk2BGRk7kDeyIxrEwbQU+
bjUPYUwSxKxH91Qt/IejAGZ+wqRcGacxNCOe/Llfb9iChPgbJLedy3kA9RmLObVa
lbHHIIOZ54etad7QMvLze96rFHQHHgTx/nlizpI8zd3UktFoxhTupTeuQFjgEMxu
H/mBnsbH2raPUbXnaBeesAEJA+v0s9dy/hsIYQrhQI7uVw7D1jsdpLKJbSh0FCkr
KCblEOltpv6KioYIsqiMKBYDd7GD43db+CXIm/yrVElkb9ZUNlrox+IkudAQRgpq
RkPxHPFMApLos8jhDr2EviLERr/XFDKsNOV3hsM4fl0Cl/oGBJHB/0GyZQ3dKxvp
+kDqpFWXCnW00ybtW3FzPHxe0OZmQhvHqCSQS6LcAZJ2b1qHbXf5Mmn7BG3EQFBs
FIzcXkJkV27bkMp2/z6vv5IgbxMX7fS6cxG5ndPII1jVGIFarKQL9AEl6CRcJCJE
IVeALn9MxJxgkn+ZH3T/R9OhanyWQVwP5jk9IWvp7X4u80BySNTkE8nHfP4t6RRQ
SSgxhV0slymiw4feQ3iTx5DY55fXUhVBG4j/QGw39pKSmxShfranyTdoEIAXaCD1
rtZAJFrgx+/PSVsPSfCAjg5SVD4PlQwuUi6s+WlqP86Kw1YBAFrJlz03uPO3N996
nhLMDiYjZjfH0umHGQSq+r4W0zEcIOnPVhRqfXMXylQUBOg5ko459+uT3uAci8DT
wmpvQr8Hawr5wGP0I9mh0TwCaPC0Jlf0Wbt5ZrnYCRBKua1j7UBjyCFXHmmZPulb
zoGedHgWq4DKXAY/mmooRtCrlJEjsSR/lumag4XYjPD4UbAlbpwN+f/khpaTVIIu
VBgV6SG0VFTLWMBfasw8j0xhw5TXgdWQ8FUJHE2lc4HVTdB+WxFFNKBam4GPuqxe
9PytC5fXOAHVXvBeaxY0vWvgP17fH6EvAC6ZY8cJC75WWPss7fKzQmzt2JlDyevD
llnUIhMW6k7G8esVhnKfzzZ7HWDe/7XLkcHjvuhvufjJ0ctZtWqa4jtlW/TvJrwj
C4cKHaBugu+VOMa9pMGPaEAHqHlROm+pVAqsYBthKfvt22elQ7DXfKQYxnuY76ns
gXQM2eKZPGWAzTOstftc3FRq6duO52cIawmKumIxQze5V6yiNcqVHiKBj9TwXbOc
Zmt222DZtMDwVOkVd+AnwEfxGhma4L7hQARIFgvoxJAyLDs2CCYt09h6852gNCiF
9X7RE3OhrRa75xPegTFWDslbO1l2kkKalgHvlMVh7fofiD7NkPGKBDWsslL639pJ
OZqSexOY/zdeXZmf+lHOQ84ikkQBpdSKpj1q774WgdTn9NXYaf3ZUn6MDrX6FerC
JS6wkHf24EtaARcU63YRWSanZ3PMcf1APZchI5261NjmX5VpZs6So/kEYepVbHLN
zw+bTS9drtZS/mobJ3DqCacr7PT/m2x6tKNBRJjYkb5CGQtRN28XP3wQtVfz//aY
kMR46kwo9co1RiPOjO4X3bQVpineaDHz+eeKPe0vKQ614McCQodMisr0H5cihyAe
CA0RXXKQZGXTzpyFMrsUM8WJznmTp6lUEkyPk/kPHqEkz47y8tnlrVEygEk445/8
28qiFV1E+eEVHCq+NVaLrF8TOAdJP6FQOk4rpd2ce2NPVDrQ3br288nl1DsLgfeO
PWagPe6VapDZfb/p3j3GnyYHTgocCl9UNgEpEWNhKUgAH89QC1kduPyia0AbSzTY
ESucEGhILcs9DdFwShBR6wg1gNqHNKFOPbsgJ54o5RYh1sfjl0X3ew1RFOZoWAEj
/eT5YdKu74osUD/dZfLGw6fX68k6KQ8u1esiGSm5Kif/sP5PLtniCBhXw8PRwKfM
gq1MwQX5hCopSKBMNyigut8BI9eenuidV6weCiKmUdidHVJmVpuPbS5bQR7gxKmB
0C2cdoimHlj/6pokMpfMRqYSa6mwgjN6ICuOxd259aGP4rqEjTG4wgsHoNKsTYTz
Bc0Kkr5IyoeJhF9hmc8215bnXy1REwbKJft2XycZC6r+XDM+NdFvqE2tYsJicUku
ktJ+HehQVVa5bJWKnWT0w9sgdjS15sBc50y5/CCWUjedjjaGgslCyRpcybD0v7gk
L9XITRiI3pyuNDI2/9gbidQERXtmMOlN6niG1/WTaK1F+HWumGHNLW8hyIaLJGKs
jiFyhXyKL4exYz5J/rLAKCysjwQTzGt0BKpz8neZnXacUPka1quayy1Q4R8etwAT
66vmttsKpiiWHCmSaJJEaKtTA6vMWtvC+qvI0hs9MIFFwKdE9gMQiNaf/X/OO4GN
IrFN5bIGoQTWfnn6IcGQTV4moCAZnw0znA1YMrLzPoIDfZJXnrUaILEkWFBt62IL
xVH/RvdAwjR4/cS1rZjsLeGAFa9S657S2ijOnnKVh4UVTWMJgKQ9mg5/i96+NyfK
szWtfE4x1/3MV5D6IgFa1kVCIE6COS3Mev+DVFmmrTWEQb9cDLhbjOyMOouU/Ecw
frQFuQbfWW/c8e2HFMmyMhMJfLaORhic475QT49qbFAyl6TrF1rV4sK00lQrXj9x
Zl4Ae9RJenq6ghIZiT2rPwxDrjNRPr8aEZ2Fily8wpAXBp/yRipgNKBxwTg0Qvsd
QGQgW9Nz31RZhDzqrR5asc9gSoMMC12LuhUB3f9v0lr4id8gS0x9vTM1GmgAwDBH
yDV9hqbrM0RddBnH2jn80TMXo3Z0ekq9p0LsbYZRzVUq5hDALwVSNSkYb4gTDIHt
eEjjb9dL1wdcxVA0GPMMhH4X4znPRHYUTsdzXFv234JmKdbrYKzl/Yj0rFfXYC1H
w6swNsA3Stqh0/HvDZybN0rLCcGYXoTW8aXNXIAlfOKVZ9gdmsselw02mImZcEjo
MANEduR9P9fRtMVNZuW68i6D9+unO7FUeGTxvqz+U/nr/hIDwO8Om2tM+KeWW6yq
nmMgbxuFgG0XV5acwhG316CNUAqXtLVDzZ7lkXFnnsZBNyXZXID/3yjNjP8UVdpC
Vja/cAWIk66IWub9dJxvVBV5xv3anGx0P3ekidcgT33UYc3kvngxbT5vfdNMf7zy
lS9PqUggswkQDBSEnbzFIjn0rHlaQPE/8j32rNZErQRJyz2UTfbchCCaJao2bdFp
9ZXOw7ajVQmCJZcIVxlJ+U42RFSqIHWUq9QQVuspGKBhF1XfgOhrLVKT5bDUfF9f
SW/qZVw8Jhr9ghwykN7EdcfAX9l0MR0X1XYrd3HHn593F5RUiYvtQsinA1JNHdxK
q5T7Yr5PKMknCLADxeI27XXxYIBEsLql/cCg/EgaLT+HGb/qUG4QdriicAFaBLVe
a4LICDy165d5uhtfAVV1b4U9FwBnnntwHgbBxkzFGE8myLTxB1YqI8dyRz7HhMRG
m5ywQIIhjO9KvOX6MvCoRkxiQUDKv79OyQNGYx76vvLLsqwQu/SJ1dZ8bhrVBhQG
AunegEcxyJZ2Wv2RHnq6ELMWtQhnvjzWir/0HojFtvtmRIbWvBA2LaIyoiGy6yFi
3wanDGWF/OsFu1LnNBcYpcI9O7/BBpiNy48kNzChx6uMaxl9VvscDK9yNLcxf4JC
XJ0TzElo+4bAKLLnpm+piHOGM85qNcQZXlBlt4Gyj1hD0GIoUI+NTWHE+sn+wBba
SCzW0/FOOXujoFX7gCT8eN5kWv8onN7p+YXxDwnFOrEtYjz3bKmWB+geMCxTmZOJ
vRdw1PDvlGr31HIWLXlD1Hf+fKKNXhKXQVqu3eTeMj0a2MgaVzlwe5AgVPqeWiZ1
+/eCUsmxuGSP9txjIfAgpkix2TTAGIgkBvtLPvBxaijaDfNhH2HVQy9lsltm85oy
qL61mk7awho2QdqSA2GcqXecDotp+NEbWnC9CwKCmolcvz9vys2sDv3Cww87NLkv
9Ibauv5YNhY0PqDRklHlLOuw6PcllkyClpPA9AX1K1gqgRSpLVqsvtec4hWc2Qgd
GO89c9pD/LlizeNzH50HJj5w8ybhEf3qNQJPDXeTmnCX/F3J9l7zyZJHq0Ryi3t/
j4Z+sqEhH82RIonvdY6okHclBM5DbhhG1cqXMAUBDQ9Os/QWf64D60DvP8EtWXZO
Tqrp6AYUFJ/lhCUrCzSjQQUBRVMmmdtuxQ4yJNSRd2kD4Iw+8O1WkERLSP695XJR
KUHzRYjkASShF5eWWG/7mXLdrusXz2h5w1EWAf0wJi5RUx54HNyeK+JKTYwrBtw7
zVaxZGjzjTnX4hF/j2vDgG39KU/bIW/Ok9XPzwt19DwgBeezWV90N/hHN7oBg95E
jqwVk3HQFN6qPeQV9mMDkVQgdMmP+YbSusuNUGlkPVStf4PJzTFGVhiQCuOvmEfR
GHqS/544Oz8OD64Gew0T2lzEgH2b4JGJFgzF3DJFxKg6SMrztxyFkyq4oFuZUMGy
tlwSnnW3PH4dnGZKuaLN9b/bmGXjr5DN+HzhC4i6Z14mG3vhceBFJw5cHxyh80//
D06BbeiisFNGd4jp0fL3TgX8MX1N5UV7YQ8E57BvYGDXqKQ6sW63MXjHGgm7V1Mn
RMG99nQqR8JpmYlzkLOeygovlHUA4XCANQR8LEpj01DPsx1Hsuug8FsgQeayjfT1
72Y1O7grkzShfn1/VaDqMLeO8np2dcxAplIp8n2qj/oJKiMasSgvh9VBNi1OESiQ
8tjoYcN8QRl8A/0SlFegJavr703dQZOhRWyM2W8CtHWphXFluD0rZ+zz8TgVIXIh
QtPHPZyqyBVgiaE+5xbCBebD4WK7QYdpRX3avhq0if5nP5Sg4+RnythUhCEUta8H
3+fNo6CRocrt6nelQHPUHBgI6GRniR3dKQ3DM+Ae2jwCcIujXOA2a6luivkCLNuA
d1kRlyBgBBwOR5U0AvMrc8e3olFPiuvRP3MQEiFaJ8aM8EN2RFM89S4Rdq5RMHa9
qmBQZ9gDXjANw9NnLBbMF38SR0oVmIi3lFFQHoy+gCwOzsYBYT6LMdDrzmbiez79
JfecmmIYCC3mzlg/L7QBPqZmVzgBhRIf+Oll5RFWIlqQbR3+rWxGPKiJfzTrz3xb
RkO7TB1LkZ1C4vmVOoJbf4kVvZyYQAx/yDnDCBJqHyrPnLe25NdUogJ7rlatBFq3
vOJfqBIpN99aPOVeUnjMvZtQ2fpDtTnbGzkcvlJ+JJqmy/Go/V9HclM6ADcssul0
t9t7jtihQdKt9Wf6hwrjFlDQgTvdtngVQUeuI67LJi7O1pM0LIo1XZBUZIgpHDfJ
i85c1Cn/7C5BvqjEmMZ7ehJIl/f3oG4tRXQVkcAVq7aaKb6Mtin2EZClSPw+AuVG
mS0lOhg/J2kJCDQKKEygSbYqiYuuxGra9Z6P15BbZufXxJrKc3pHIl8eG1wUlU0n
SOJTyB0mudamCutxLOp8yiBnFJMquA7O5OyzRDAvtsN/8l13faC4GcZRmtsr7XrP
ai9TZrcoNe27/BfahemBdUH3d3+ZT8Tcjog7LRQ2wEjH96NYcWrif064R7nS2q5j
geBcUwo8tgykS869Rtk4mPiEI9oKbHDiTVChT9MAacbRLMVjO5KW5UslG4e+EEF9
tHvjSkZ9VnxisMZ8Pz5J6ZSw8SArtFqWaSJyyNh3xq//32Gt7l9SRTKOLRoLYYxP
7xhwjXW49hlmr99Y+1GumEhFktDDhsT9qQqKCGRB2BzOSDn32PcLPYbzoavFzPJ8
4ALAKWBUfWSGknIXTwu7eh6lq8xkSi7GmmLXVjXN6NhJPo4s5YBh0UElqIh8ETdA
cyEG7bCiz/dEDjT3mgz/wY5ZEdIgUzb8I5jQ06TcPQjju+1LG39Fu+Urm8Wn5gis
G7EOdM3CwchWjab7vQ98LJxaUXphyZSPC9Jz1pR7UH28ZNZDfko6TCIfGePd/lvY
1OejEWUjusWxWaUfcXntDuUL4vnmO+b3Hw89h92/Hp9BN4/V2IjE6ICPr1Q/DbPQ
0cEghUTE7eHZIDL1DF4vxQEnI7ywT176VAlF0eziakw4rFcmecUT06xCHn+ppeMM
9z+ZUfTsCHJwWmtrLJuofI5FtaU9CPqQoiBd4r4VWmM0yBVEepfxiU6ZxOu10lCi
/+d8SJ3nBg3cI1aa+9xYkcz8xvQvvQyf9/UZmD8BhOjfCclIiveSRfvYxQRqrcY6
LSFD9pqSdw6kwdV9BMydcPPYSBenIdualCA4Vj/muu+Tt6ckpPcBIW0bT6WzXFvi
cEov3AbjpFKwvEqOQqTO/7ZUA4UUFUfENOVrUmmgTGM6uG+4P2m+1Cnwmm/zPeAN
liJCnK/4b2xsG8aDBzKn0zSvh2nSiJ99tC0S6ZNaAp4UYbXVKxgmnWohrc8D769K
W/jpytPWHYZwwjca8PbJy05iEqspTeHU43YIG28gPTrth5BS+VaBgPPYn5CIU1sJ
gZxmH2crnngXKr8Qz1SXB7GWH4j+S9+nNr0poGrycctHJ1DmvBpDtTXOkMfSZI+T
DI/C5rygA/ZmKHidvHw8mdgQsqZb+JGoA/BJ4QVb88JMXvwQXkdv5WcUM7818Pse
FHh5V66JM7i52DhmjahoZMoXfs3VhHdAoNsLbQIUS7R4jy1kdX6MTukIgZK9/zOK
tjZy8/15M7QiANrADE9+XeTATEy0oXU5OSBp2/7YANI656WtfB7bTXb0CA7CLg1H
rkHGcdVeCqQ3erQwTkIcJpXF45Hkou1bCF6eiyLogfFEuQ00F/2/8YPGPYkzgt20
pTA6HDCmZZADQf9OIVVtb3y19pOdCByj6yRuH+Dn3t3wiKVoBssoISTU4Ioo+MpC
wlttiiKc9ysbO1FO+fx4jxRWnfGkFmo+u3FZSkA544XcCA8r30Xwrhpmdd9CSR50
`pragma protect end_protected
