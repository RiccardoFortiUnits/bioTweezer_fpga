`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F1SEgBl2fPJya2zxzAQ0fK5oWHYgInU1l991E5YUD4NmgnAvLOOhYDA6JcnjqRSg
Cn5XoMSlN80bddRTrNxD7mMwwFB6wyG7f8ULnVOvSPnUTheEHq3I1iyxwd3baLcN
WNTFX1JTj+d1tibIoSqos6ooLeR9CO/mv8SiCWiwlzQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15680)
pQRpFfbbxh+JLeM2331Nv3kgCa5VSWhlOHH5T+NgoHU1FDO5a/IhlUnRuxjD04wB
PSS2+XFZbtAda1QSislg8gRde6l9/Zomc63ChFD4OD3FONGJG3u6kp3k4BqeZ076
Cs49lIZMrsDTLJV75NaEljLQBos5BJjlU1oXzkQFNRSzR7Ro00x00ptdNo5TOwc+
ujcKJJ6DHtsf12PKNDwKv4f6/3vQbEBrz82VDE2ZqWEI60lsRh6tN27QSc+MdgAk
tgXcXLlVrQIxWl9TFQUeH6gZeLQLQjYKPJtq65CtCRQSK8svLWCdOV04w8VPuFF6
BJ+K9YBZdAHjsr+TsaBw8bxJeet1/qwGrvxUTcyz0PoWStCnc90Tan6i7hwEBkQL
1pXSOeEKtIdIAdnmNFTw3BWUyXMcufVeHJilfBa7TnqO2fSD7n8PfnnPjVEjOWz/
XeKWW/Un5c2tDH5VsKxrJKBFEE4mfYNnRhfQzl+NXr1OKiwDHsZL5HRzRYR5LF7Z
PoV2uuHR9/eRvvqFgrY70l+lVOB91n8FuFDRKW3Zva6u7j8jxpfD4LW0Q0EVKSiD
pGAflKiBDOwDpBXsaQFnODlrENAzj+nLAO12Twk0M7Qlnv62Zm7MS6GH3Bbo2NyD
IufkSR95kcEW5WTNUuyVTWlqUXLF+DMt+3+kVZ3IwSQNBRtJHQg/ctGUWCCJXXcc
91G/nPFVgFUI9TSWGdcCsxaQoH2yx8xWY7DHxVqFBlp1MadB8FvsPmJwgmxWGFNO
F9RdIjCH766hBFLPlC8yf/Kl7+6JSTSEMiCwig1IQQN4nkD6ycCv7aOOAMvvMJju
Nw+CZC9gGIyq547tfNExIZbv6PzoAS++jiV2TrqLKIuVfqDifW5Y45U3hF9BKcV7
nVnMyTu0xM7lHjK0xs2prryh0dfK2SPwS8VkgGYW6gZjfH6JjZFkbQQZhaWn42D3
SJ7JmaUE0Idd81G7K09k9+fRQCjOJwPMCNcKr4oe1VTKVSwYPIDv++c3JnVGJ4bn
aRfpeP+Q6UWmi+drRxl6YVnPoDxC0NQpUDpXKXONcwPox0ap65W0+UMGTAzl8Ji5
gYyCWEWqq+fLCwO0wN5XXiobGGYBvSuySmkF/r+IQS/UcsX8rf73+9i3rTgoxjmK
prHhQcgCIy2vJ/8dBsVQjY420rLbuooXIaNWuMovctMiue1coKthGDhciNjGf93u
K504U+atZqZLeSXeTI2/EVi+H0iaPgedqPgXwpBU0TJExclJGpre+7dWslTPG/CB
F5AL5tOMpeEHPu372gvcB21eUgbyjY0i39bQwPaSyhPh6vAbyLEtPQKXqISY3QQa
6r6LVDiWLfbNyG5mgwa1N+RoDIdrECToiBFU+3ICnNhyE/ruyC/JH8bdfRaQQm1n
VvE+mq07sB7FYsaEo9JE/cRoXqnvK0a5tZgJEv7xj64FuZRdie2MGVsivGPk2WWa
kbRi359Hd6hjoKOHUc8aLo6G99M0LaW8akiTIRnI1PUEO2wdQY6kch6wwqQI88Sq
nMkoB2bB0d6T2jHaGeFxpK6zrCd0WAjtHpa63m53vapOc0VpEJkYQaCXbTc3ZnNw
+JLL+Tr6Td8zdBiQI2IJMWMN2ly4PQmNtQ3uCNjlSMEYFIlSYlsnwOLRnHykxCnr
IEyOITbOf+xf2cFS8+yZCcjrsrAJeUZMRjnhbHnAhHBQwXjjxtqDYl0af2/bT61M
U1HLAO6oqQzL3T0Frf5p4jI+jx3mamNNkT+TcWjeaEGZ2TdN50Jj7OwJIP8DynQ6
m2XSZW8Ne8HaEDlUZkdbY41flHHfN3Cmp9DvRVhgj4Z2Dz5RB2sqwk3qSkRx+RDI
aoatFjhKhHI3Vq9oBpE/Ot4gYDBJd4jsEahuSAIykIRkwRBwSEHRkl0b6fkAalpq
9J60uiFJI2fOXTOaHN5OkRLWvcZAsjImmOho8T3+WeCbkhB1iprge207c+wsaB7q
tHSNeXOtJg6rOqcSTzOAi/usOYOS+zEmZinyhABwqOlfFPQ8OMNVpd+wOO4+/Y4a
4OFphVid7hwNtU76BcfWTpTTUld2MgvEuGhrRhh9t7d4fmolcQqyCWTCh3lz//fB
VCvQA31EIvIgY/TQghCA32t/zb9HslReRvKQbpdhSBo8MPNihPTk7+yIijwPwEEI
fWfsMokM9ZvHRYkJBHlgFlO6eqXqhWGtMNHL28e1oYY2eYt9bvn1prD0uQf+m1wS
WCDifN0xJlmbzmit7n/DTaDntNX0+4ODorPRh5dFsFyCm1yUhkQEtNdZ3s4mqGTo
TzQk7YEu2oEOO6IeEP9QlyKIctLj7oIJHVH0jfP8+OtKjA+YNolgiPP13fwLFCZ1
UmVJ9aP1FQVkhcUfHuMQyLuLsr3g0wJC1AyO/ohdT9qYSw6o4SzyVJEvm8ZYG59V
KThI5yXJXmutvuEO76Owaxh2RBI15TfdbEngHIlQcMWy0iqCRMYJL4nD2a0qW15m
Z1JW7AyciD6ZWKIuM5+m3AUmyzP3psYspzRpGpJ/WMUXXBeNwbs7rMj3ughb+kJo
qgThbnraorXBa/G4XNurgyB3siBDGDVkAQqa2HWTE8wkum56rgMFwWPImrGevEyH
u93WEFzNnVL0vYGWOh92Q1iVTBO5W8GsAg9XHQ/NYW+VllLLXfVksJQ5/W0+SU+F
5KVrGA6N1tqcEWvFERsdYoCZeTw+J4J8I8ufr/alm8L2CanQNN27Oovnamep6xVl
yRkNzu3D4+t5cdyYXhbcKerDtK+u6/KbmZ2sJelBPvCx41EZONivDWGH27xRFsQA
6ge1Tv7skBAzv1XfXRd+M3jCsVcGheCQcG9eYSbZsLq9YAOMVA5OMHHYf+hbAAqR
NMaLii4w26uez9H26yJ7Zx6epIvqeN2eL7ABgA5pnhO8h3pj8Ka5APxLBbolZA4d
yJlY7cLoTYJK5HXzZSGhRPfqOSTYcFxYiX28Zs9ryT6c0j35v1pF+b3XFqUXS1/G
oYwLvR8iHRHox7otLPw9Y4gLSRQffH0ZNFC/sEXluUS0JjL+VXKHH97iBFgAD0oz
31uA4vLwnlpmqLFluBxAGPVcp/5jhgUzQxqYjpkxNdqUgffoH8/E/1Zv93YwqV29
budUucokmWZDzDdSBMOtrF1n7tqcOBW7haMdT3+TpgNT5r8uEyUuhpQ3bu2YdnbS
WKlPZxxhhqKGeKOiN/NC6dnY/5sen6rd1QoG0WWjKV4khQ1NUpLiekP83IGEpFsG
lnL511rTWcC10PBf1oOWT0IS0f4gmWlN6HzgsgufT1GWt+ZuUvFOn6LH9bVZUyMW
pleFdyEdyVGtLKGu7x9GeX2Yn41Zg01ctTH7TdiCACPFAN/mD7BPkQoVyEoMO+z7
Um3qW5gE6Hf0POXRswcj8sYAbYPK9svlsJSkbu+WIQTMNx50l4P6m9pcOZHtdxfS
w6kY89HUhQszY/PxhGixl/kiTgZyWl7gF745csyPjDFOvCcUe8sQyH6L84HZERty
GElgAJnGTtHpAidzX5sRfMGPmpz4mqdaI43Q5CqBFreB2RJUONT0GQTRO5HrBDgn
WGdSRlXnySSux7WedNawWLdTs4oO7rNR7g/sGKh09k3lEESALD6XMA1PksQQKA9n
qKe4vggxPPiVqhnhwzyT6+Dngy6QE6om0AJe8XP+Z5BkhuQUpkkN5BJ+56A42BDR
GytQ8MZUzB7cFUJyHea2Uq1GPwvArUvn7zcvPByFqC89nvOnPaKeqwkhAvFH5ERI
yCy10t/q0ooIS9CFRvqExBo01UtWBYyoocxVpy4ekbKccwFuha8J75Yx03SsHozA
/GfiaLp4U+Yr1EPhY1w6jpXBzt71a1qHav2ZWc8rzx0Qe119Ie19qcMF8gsvX1O+
nMs2BL+A3OKtqyO/tpk1QNbAKheJ0XcaoySfUTCz4XDc3y7ak0G0fEBB0437/JOV
itIM2Z9MXGEnYtvTAbrtBbkDD/Zi6m5sr/gcsE4dCdN8vK3MbpCAlaq+LWoxUGV3
53NXqltCILILZ04NFa+KyjrMAMUwLmTme8h6dtVyRYlHFlnkGmdmK+YpJh93HXZg
rG3lkZvd4iZrYGUyO7guY4ybVMfE/QzXujvnmHM3M3E76Bq9BufEofEMpt8GAh2n
Wpy2o5kyLSHLti9tEj4tnHKWjkYsocCYaFGVNM6ZEF7eV105+DLtK2RK1jorh8na
mkZ4YygL/YKCZ3v2enVKX0cDziAev4b9FkRhtCPsou40OnEiX5uHUDf/W+t3qHJL
nJfzvOn+XmdnjYm2zNXaxqlH8xWwzOzIe/+xglqFsjEujOv65uRs0YhcyG/3ZHGM
fJildGYGjhQGsnHvkVFHRSttF7Mhi1hxklA+F1UrAth6T8D9YrSEKz+Lx6pIrLCg
aLdtzR+6J4juVt0nSCqYwqWAi3wayuvlHKobUjz64UkRMa9Z7SVn5yqvy1HHui+S
7DOCwu8B39S1Fd1s7Zanl1qPNcbeZJOf6Kis6pkH89/ZeOFG0hYA5f6zq3qiRg5R
jAHWhn65pwyiNB+gUwl2Ln589yhqIbb5ESIJ7rqLfgFIOiKnzms/7K+6sqaXea4N
5t9qIYcBx8skHvfmha4FLgmPV8XLLnnWn0YnJrzI+Pr29uzIetZdK4DlR4OfHnFB
ZbqimkzxAA5DnnJvmubSco81MMYaMtjPHTyJp2Xh+MAqx8jwJb2JQDOIV72FrySd
RZ0sByh7zmICj9q/qVcyU6qkBBCG8WdheqiIEVmZXrLD1JoeEK+f0PmeAawo18GC
3gFHajG72cKbLUNkI+6BiYGW0vOW10Rl9V6TLocmUS3sehWxMp61B0nEAwvhTfie
TlPSt5HqQn5Yod0ejsiOLKR55PGosC6zusadcBBZgHm6BP0op+E2jm4M6ja181nh
p8ouWLSWKpS+d/pbwA+jLfTAZS7SgCyvZfi8VgV5W2YhSd4yxxypEpAZZ0vYpDHX
R4yWCdbBQ3pIIqvSorbzBpTXkpS1e6PwYBqfh0ziT+zdB0JqB23ORfLV0fDVRnsT
fPstHmdEjjhRr0gcCFwgQIyNGl9wbYgRlvwsX/SqZwv1Ij0KKZOV63msVvdirExl
4cJcL+McZSg8aQiGW4JGZ9OIaPS2pTDr3MFIYgH66IPWJ7V/9nndKEqO0giHxwQO
YLml+7U93Z4kUoORvHRMctAT617rXHozCKzAwY29WGGoWSWQF7pru2viaEXaiCtt
ajF2cKASdp4/xVT3dSUTrqjXCiJc+MFZNcV3v7lZImN4CvF1ozI6Qkbp0WiI1S0B
m1YOHDqFDMLqs0Q+s4IIE04dCCV9aelRu9lA12e4ITCs4zB9yBCJiVXbQoP0/Alt
tdlN0BMH4eJ1n6hZ5wgxOIji7xSh0FAT6d/hdYtkKCzCkE0jJFJlMClZIn2mc87y
MNIusdRf/tdWH+v3xSAsXWWchWGZTonfD+YG0JYDAP8EIwnDzZac8pf6hbKtVBLW
9/24+tv0vijrJ0lYeS5gbGbzvlpNRX7rOnigy1D79HY1fWFlmiSq49VaV0TZK0ZW
+xaPsZtzsm3d2yLk+EelEfFtHpLoRQAotsIOAlA7B9sUM0ekh7Z0GyC6DEnorx3G
nWke1RI5EaUPEOulwF8SVXHGTQ/HunfERfkMyCIfEFQzhQKdtD4R6IRhkI0zyRMl
KRwgoaefVI2kzXyaOtAFgTMcNm0eqfBImNWWns03dlzsCoCgkD45HWzwborBMP5C
zBU7b/csxciJbd7RVYGj8u9u93OrTw10Y9GyrfHuY3iTW9V0ixbFJd1aSudV2PTn
kiwerg9ZdvJqxi5OUAQPN/9MqLZ1jUZOxgLVidp19GMqDZoqhmW71YtzwN5rewCu
cJ/13255mYvL4T8k+FYQhv4ZvlLrKGlbCoF9G3BXYKasJuF6vSjAorzou4YPtSkN
CTjCqRnFQV5X+Blzr8NUGSG/Q+4RuL385PgpIDGMLBV2c6iRWhe0uc/bQ+51WpXa
7lS5OnL/QIJOnmxFdLjtydq48EOAnmJSGUw1+xtduu0HZR2dPs/RkypoToh17oQY
SXrt5AOCtueuuiLn+7r/sTamOrcgIE8qjzgsfyZun6SRo6TIJ+gKlUP+ZS+qGlj/
Bm3+4m8QXBSLErhIfsiqg1X61y42jOuYum/mpxBNcphRferWbSQz/H/nhCo/QMRl
EIZ2BCl7rGf0M07xoi2Kv8lPa0QosfNezwrXA1m0Ww+jCnhJSappuGwrKRItgptJ
IhOTGG1b8u4TbelpfbzIRZfBB80yZddYseEMV9ILje+0Yf3Sxv2EXeO9UGeLBVRg
6w5SleJ2BlRRpceUlcHyjOdP5H5UUWUxA3ZBd3Bg8QzB/meyA7msV/bQ6qwJbriS
6tImMPb0vJeKmrZ9gGV21plMdgGxnqs00s3UL4XB9K2pBsuZmEWteOEG6kdigCH0
Sx9n3az6mfPh9V/QPS+nGu9SZKjG8pPQJKYpWQynWrCnHsxpssELDjHZt1jfWkze
5w1rosZeWScX3hN6wJI3yF3Ufe8se8CdXpMWSpWL83pISVWKSPKBXtqbpOMCcfLM
NSNap+QazHov1x9uv1vd9z10i29FCTRRNNNZoD7HaqglsQHHNY1yZuBQ/PA4H0B1
I3HFH1tN36GoM6vlP5meQT10E9bmAgPRDuIvSaUoY4p4cnwSe+ABpjPP/4+3qRvt
vIkhc9iH1e3sXbOIrADy/sxSWid5DeLoXYzqhTmWeh0oCvOTjJL/qHNj6ZVj4Vag
SEDiBBSYEPCaRa3GXjT/Ub8R9p8esOfYyT2J2ySyz0XqCiXuvTtuAkFvDTcbKpaK
xzLkbmlYBkfSfcOmpQHbaEo513zpL1xCz2248JA+p0AZzeInPYS7GrGY2/hnb5kL
aTwDo6RuhIFFu4EujHvJsDDkqDnq8qs58Z03wjO8pfwYLebQ9r2yZ1Szbqup0t70
hLOFWzK+zguVeeOC7H0c63IHcLYJs04aNXgMFBGqrRQ5DgdL4llpMAqugupzthWQ
dYL9lxlZh+w5+h9qWe6VmdS5xEdlj3jzFl4zKbckMcLqVCk2OaenppAEfT1TtAeJ
bwfj0EN0c2fQ128HP3GsT5F0fPnnIvrrlYxzn4YYmJsz7Nsv12MTSCS9tUBDepO5
f4car4SVNZn72usvvIRq9UuTxa0NiG4EfpBt7519NPgge5A99hlR7/9e7Xj1s1SW
Pm+C+f3cwZLjYX798JJr3bDD1XeALsSUeJNxTnK+Q824JSw8H38rkJFlY125/V34
V3gZGEBSXpehsNOQNwX6wabNMybF2ZZKpd9ahr5lueuItfGhvAGRQMSjKgg9gRP/
R5MdpLusjEL5gQSR29Vo0mdqE4gcOxyyAP8n0TXrSBXVc43bDvP5q9hJzAms3OJu
N1dHiWG7kbLxqlkdOMLDk4rEyCf1LiLIpxKvK/j2yCGk9nfzpsNLbFZztQBUTDhc
J3c9XKrldhczWrjx0E4KAoeU4Hw6yw8nlgX5URxiQYPKjJpjfbUlpmZi49HJ2WAj
tJsa1kGZCm/elynAzdo9Kl3Ycj7k4gVix0ndEeBNPKpjREaIjEWy/JX0Bwrxe/nu
fhfM6BLGKrXGfS/MIGj+zrUIknZPcGYp8uJX+ILG4u02UBkTg/PFMtCybTTxi41S
2LMk7LT/AMyg6vEN1Cz6zJqfW3McA2/OnIqrOLgRgc9wIAjCHw1TJGhserYUTOgN
EWYd1Ldrc8FyWuTZCSvVnLxmf1mF5Nht0vrlF1/gO16lyPHIhtmKJTfDhop2EG7B
FMSVyP2aGb9z0ISyzXxz4gZdkU4KuZmSP7PBK3nJB3xkJZ1OoXoqfkP5vIkbUoAi
NWhoosd5sOBc/8O71LDsajJAQ+GBIvqHJ+94Zxrau1QZKQFcuq1lzfe1zLrNHx8J
CiRmia8ZG5T7oa7H6zsNQszGw63+5q/gsBXYyqj2m+ofZRqjcRgvNn+Sd2YaI8Zr
jdDyRz6d2bEXF1tWX4J5J1e+prA0vuFNcOFsXNEVZBrpSdmm61rgzqnHfk4pkBA8
0n4dLfZP0xdv6M1WOsJSPuhBISl5XKtf3Jry/3t41SSXhkRwurFDPOImp/7FbNA5
N3vJWAsR+AYjD5rbijTvEDN1KdcsBvuaFjZUPoj0B59n6tZIGvVeA3Sqj0x7DuF6
V7V6VHOBxU2wDenhaA7SKyzX17aDJcbSC5/nNLEUQvmB3JY2ypQH1LkV+Fa6cgMS
Nrncawn6YL+TBqSdJHRY5EDtzmU8jwWRouWLumvo1oIBLxfm9fMc27Izqts1fPhC
BINv8A4/ve4NILlgHiClIlo6XWeHXtDQXkQg07Deql0Ln+SGqtEJXjcTbCPyj0Xv
Ab+za/UCCxh8hD+H5bMvH+VdfYXYL28DFPSKzoVDIgbcZGg4YTBfjFP4jkzju+tt
r4VYILngNY+cg79bEb/xIqiGflv8uJw78h8axsJz1dH0achzbeox7YWEPaD/n378
p9m/6UgbV2Oztte6PkhzEzSTiEOtH9OM2pn9mmEHdyLBG6w24rxT3Gm2rhW2usLA
Bk3ajp7Ah2uKVkVLak/3ESee5yFTwC3WOcXViCeAs9TahQnRVhGLKQME/aGb0rc8
24W1UDQtUAyaRTzytQpR4t34wpordoIMetXxdZNFJSWLs5TVHwZg71GzmB/KlVwy
QG1DlYOawPJFDOgeRzfvwKzc5HIPHQZjpCw5iAT6e/on7nzp+s7d1MxwWfmZj0ED
VVTYDH9ujmE9k5PRJaoOgXOsQ/CFG+tDrzDshWoqVHzDyzpr1qoUoii4lR/xOvRi
YwixjIYbxMh7+Qiwgqez7+LQsKTWdQCd7GuN06ARo12fQ8v6PAUN6HzLFCZ9i9JR
PNUe548oQuPFANzN/a4FFYX2Sxku9jzfd8T9TLe+spVBJXr3xyiaaGQt8Y7YuDn7
bnAj+d3szFGELrOStFSdbTCtGPq5ZmUSH52a22IHZ5WQ0bVQqBt7b6Nn2TpCupLw
zG7R1+zbKMi9cEh0H2R8eJFWWxrpzrQHI3/pTzrIvG6EUp6aeCGpuBtcwtz6i4v7
5rl5X9egxxXRsRs4y0hDJMjTvYpWzk5xH0gL6baz3uNqXZQZe6TaW5rSzHKEOM8q
73gRh4z+BIX8jI0x4PErKiZWSCagGn9ZnJ2Fhvcof1md9EU+MN3hWir9ZO8mwoeG
L4FjGL40CHXb4xkF1fklKAcIrY6PQQHZT9qs0JWVw8Fq7Z9PCzg5OqyL4ILBWSsi
ltuVt/2BB0WvcTTSeWW9yExFPQUbdDhI06ZvY6Lf/g8nfrMQU2mVK6ec/VujQFtE
alo2kajixjaH/hxaR/0jsHaN4KOj6j9prLDmRIPX25pIhVoV5hf8Xyu+57OdtCQQ
Wi4svNbQXi+iELE93dXgtGP6j7BQJv2eCKHNZV/+MN/TyKbdBwaGc3+auj7aXgnK
QEMM001wtK9o9da0DWqpkpPsm4NI5dDs5gVnuKOHEaJ4U87/S+O7S99v95Ri6RT9
W/KzKIc8mFUnNDpaEmha59uzCM+yfP42bQIkhc/GJ5yVCI5BOqcjoJ7xlNEXAvGd
lxhVvdNElMfEuTEp18QfWe7DjEG/4buHnqkSdeotuLj7thnaJ0nDC0VkB1u9pRf1
AgFBvB1p9H/wLAHi4lPRpXBiau+LAZxb36SZaraoayyOI/9kkEvC/4RtUq7RWOer
HzPsCLrhnaJ36zCqNITG+4CaaqKhZwimwbLOpzmPF4lF9tOIVoLYA9nlkRi6RKAu
lYHzRuaum5Af9OuUwN/gxXkaIz9CS7RQvbZYYJpCBfnu7r/XFZYidIpq7FMvgZ2t
8iTWUw4T0mb59ac1JUcd8Ij6cSLfnh2Z7wBmzXKFm0kNwO823Pzptt4GyJB7DVlb
QC5MIVDi02l2jGNTS2OVwLPsiX4gfNpannQ/D8zvRX185uw2ShdHE4xJP0yEXmTV
m6QMeeZaf046cKboyAa+RaiuotawDHWzaYXa6IoqYnPgmT5zdqvUEZBFqs1feq/c
ILu9RoAubTw7JY4IHg/IU6Bu2BQVdVbRoxFcOpvXnKJ8o4Jh9365wm6tZNEkYk9d
E9f1uQd2Lf2Yg0wFfSQ5mWaaVgVBe6qm8fnFq4z2OeOEhuKP9069mSfMuH5jBdFu
LSaLutMr+Wg7yC3RQMIRD+qHybGhUlxJS2YmgSL30kIDVZkhi7hxogwoIVt0f9nG
wLEcjAJ8yH5iZ9C2zMcG0yaJM2ttELnnBeDQNu4OKHDZB2gBC+tdLTjgOsK1HV6t
jQivSNRnboeeqa6sR3oK5e6gie0rwq9Vz3NJ3xm8csFcqtOnUZ4SWnnqxFdK/t7o
1RzVAnN8+n027hNXRlyP4bw3UiqbJZzjatMfQiPqhee/Yrh0K8z6CrxkEW8gdYxB
+7vWk9di/KoORqdu3tcfDwyDLy3+cm43tDAtkwGPlvsrTJDKPXPf7WV9X92c5SJm
8bmiINTFKC0+iL7J/VNQiqCJ+oaGiXFZxrMRya/bGLb6XAsh0LdM6T/DDjvUo8Li
Cd4xkJCNFPZzb7F8FfvXbfjzz84uqoJtd9/0/3d42o6l8BVFYpEPPf+RhnrrMssp
a7FXGGPDcR3iMMtLVL9ONzvstfCTUVzqI4Un9bygJM2MR+Ew1JognYEFHmjz+/o5
rvTH/yDHlp/XbDafyXXTPszT2addTLuhOSfQLaTSfzrEPG2MkAulUXiY/6s0ZrpT
Im7sv+Nwvy3EdzQFXzefKeOe0b1HZirtv9GQXufmXIkLvE8+l96b+YNFJz0yjd0z
DFt2rWh5sW+uYFM+akTc5mR3F2QUa64THfGWdPuIjkIQBdL5EU5CkkTyh6uyxmgO
qti1mRb+Ci1DNel1FpD//jzULoLoI2hvBG+WayXszAzlzQOh+z5NjRtqHKFSkMcc
d8ZJpqOcdWVn7Vy270RgDIcGgRtWhWlnbTnosyvWPNoyRsQePGhKmZCgMT7qvmLn
thQth5CyjVL4RPRNx62F+xQ2DYquStKkw6yvQphfGIjzu5AwMdcDIlFanhZdZD0A
XmJOUe5BqcEWWAE1rt/Bl11Yffp6ahP2bwgxb1AtHIXuYq8zZTrGQ0rIq4VZ8aBg
2CW6jE/mTmnf56R/izx+yL3sY4ylSaLBkXDw/8ZjqYVKPYhIxPpg1YeQ7N9TKbu+
9ytPZ+cOL6L6Qb1MjtIcjyzG+FFBmDqulbwPm4e2ff1rHPrfKgb4rrzJBNipOoxf
b0M8Ta+2a0yPA6Doygpoj7oh/SwqvF1HgrIn23MCAlpOm2/EX8sn/Geww2prNfAf
4lF9vueMLbebtvgbCmE3HbyreBT7kryu7Xq3RaonuklC6n2oGbAG+DWu/IZrDAkr
CZpJTBsMhL2Wnk7HEloiK4U88K83vIIEmrkjxSL/obksfE632ClUaWylq1b9rSEk
dPwiVNc+ZiwILgbgrQlvEfrqSGLaa3+xPOa9Z9ghOSV1MIAxow8xJo/0CjhC+IGv
zF6H8K53xm8JLcTUTuxoNWXY88IhayM4Hn8VvTLngIY36P4kvM5EYSqCTC7YPALT
zXgB+Sn1AGRXXBN5KMCySy21tudSWgC+R2siA7FKx13aRhXN/wRMlwMBsiqstqkj
08uDL9YBJq36jqc3IHrXUmgL3RaXI8xwhgO6a0oTrG8MnxbAfRKxzyv7XjcCb0VX
qISkGy1CxA6hK+6MMxYLz70YLppColvcw1dvYLJE5VnnmJAOFdaV5hLQTbb1sLi0
UnccYMFSqffXqZNa6AQUKjsFGdWNO2LIXhirOJt9PfNp/nWoU9rVScEN9UxwkUwm
5sx3WYuZrX5MIIk69pi7JsPp5KqyoRpdmQpiOvuurKhaJzWTZx0e9ye+tqzujVJA
cVTOWqQG4pPLzFbetaF/K1tJAxqNRaWlURjj7SVDVaLeAGWGfFVODnQBFby3FdYI
le/kV63A+4QcPyM+BhCXP3jmVVgv61hmCRMyLQoqUjMWeYa3vCexLmcxmDK5HIQJ
hXDHbdTiJAdMfr3WpHk81okyO3a+AamD4ywpoWWxd5ZG9+M0JTN4fAbrkZr20ahy
qoDeMg0HVJDlJ7+EvTzPS7cLHuPPIsBNJFn8vc4P2XO2zcHlMb8H5A+SP6cYQiPb
1nHArqAY0PuCVi4ULkoaU/ldOd+0Y1c3XD4k8QeceqcYeRGVi3pLUvRzGFgi/TBD
0bFSNtX/0SkF0+ApK20nsV4Po/wdPhnjIdkeq5OluUEFGdMdlVQf5EIxkiUYkPyC
O6sS6s1hHnd5CDH18jqwnZSAp7D3zlD5B13gHoQScAaDvtvgwkaJOKvJC4wy0ANB
sKT9BA9G8MB5G664u/q7jHgVtPvtu4SPXItKYJG7ArAeWErBILU6QmOxeEn8EZR8
apiDm+n5f+MD/E1grAS7Sd7t9f8W9n00dZ0qG4jpuSv/JLFNSToMbs8XUtzfu6lO
QbdAKOGewJxuFXKcCT8i/IBA8ICEe2sxxKh52myZ4/VNhE6CmZUFK+9azBWbeG8z
8JaEo6QQ+TumbThcpkMAiqOV6sN+7ltitt6mrKkKeAjtVgY5KdYSFWKj9FkugeED
shEyKD2fLIoHFFJmdHsa9Zyc11DBu22qsRvkK/nc77dhSa0QgKJSR47r5y65zmIX
TIwvv0+bmUsTkZylT1xI7pz6YaQQXMIAeYRCqQRTO5k7RxTQnlSK1vdbJaM5qIPO
gCQFZn7HxUiNHBi2M+EUoRClkFFfhc2RBTzAvLAilodahtZ6FWpbZTqSocN8YuQQ
gSJ01E5MoFVf+4JOIljAtMXP5gTCnrEbrKWW9ZQY4jSmyGtJ8avAzfQGh3N9C42p
0+E7KmxDX3FQufMW9GxsNWEdvpUaoJUrl9HPYcpufjZI8UpXj7fZoGc72KUCC5zh
4AXSdkO1w8RisodBOXmRQFtggMVGG8XDoPf/w+NK5gQITpeb7vSGXxS8Kwl2utKR
5exlHZyaq845Kc0E77QZ/DxLPEDeQbvLSX3NAnM64jPfyVKjEy9D5DtKZRzIJL9Q
T3PIEBk8wdIZwyOk9eg/L2lRNOnvz40TpitCPbQQ4fejrVIYhUYWiXzW30RWfQ0E
mL6ckQHH5THXzFpNi95txJHPybz8GxP/nbdVCa9dBVMcjPII1HWjdV0UlTLVgPdm
awegVDAJqnXvVIEr8ksKteOLP9JDpM2y+5fBwupbur+UZ0mdsMRJgyk3RmNcUklt
0fgSnC0WcuQc+w/HMS3dhyR1J0Sf9Xdpe6WoHQcJaVzl1sePZn28ec5TqVJ6oF9L
stPfxJUYbh+HEf+2PV6tJ/JD24F99JSp5uVZqYNUWCLMCwrIQMkIV1kpDkPlnN9y
zDxR2rjh3dardYJK56NLaZ+4JYO31QqZNLjFaQVHVD7ALbcmRG+g4duMVbP6RAeL
fIm5U13o/XgOF4RlcnU/w0stg4GJEFPor4jLTVtahAvvHJbu3eFqoAclPjDDL0MH
Jsu+922gi2y8TuVmpmLOcBQoQIGndqkoUAasH4bkJ0mFz910Y0ouRRTLhuiHxfXs
9oUDRhACYhN+9wwW9GFOAv403VoVU5Ag2YzQni6/GxV5wgNEfxE7YlK1IpKVmqi5
/ECSONgSw9X0IYJwrK4HGl1CoNgBrIJ1AaS2maatZ7jS9IRIoA7Rt3Vn84HG5CaD
ngaW3u4RcOr2lCKXDEGuzeZ/b/NEsCdP66Wjclbwdl9ABXHooDYxAK+CPwb3byP8
XwndqZM8TmTmT69FFKwYUAqGLTTdTCxbnZwS5/sdimfxTn72d1OCe0CHBM4DS9ln
6b860/GNxTUGoh3VFRjNM3mQhZb8AlTReGvpuNr6EMtVqvjnENgRRJZoisyLeCXE
wQjRAT1TKaMAatZ9LVXmlM22YLJ6Ockh5YBxinqtNHKCrgI9VpQSMzkZySjK8YvU
7LUqArHJVs9LmVBQLYuD/uYo74qOqCBz8bI5VPwj18VLeGmXw+QpKQtsfvzofS/b
9qUVWRitZWXkHrb1nszLjJs+qpTa4HQ2zCpIjkG0FVckC31gbztnfXcaGucZDXHA
2aNHA/fF3hufJ3//qz5J9JZJSOCDFGoprp9QG7mzTx/RC59xwucDh06TM9ANSiDx
O6n+frgh9rWCbo6J3RPPSVMwAiClXhFtEZxtaupMLBLLpLqcpcY2h7RFrkZtM6WH
QGd5+/cnzmALAdRqQPDyTGh1Aoxku2CBSd+40IyXu94/V7y54H5gpUf5Z3pBMAB5
Gg168Dym/q5Z9qL/Aoa0aNvvAgVJsQXOiwHJXFk65C86w5efPatd+uYrFnuDlORI
PoeN6RL6zxB1seKAgwkxnr09cUz+nUveNnvGOw33gcAgQ/oMCiCJN/uC4AbD/0Bg
hb6JtsD8VGB1684YNGGoDq2tFvysbyvj//viXqjrkRVP20yRuu0dONErM7vUxUBX
42+1V625tU643GZ1sAwcgDEWPLzMN+DzNjS0FZf6g7DoSd9BfpBmQbXd+zSzOZAg
AMUbS92ft36XM6o2bU/wYCBDwX4k4VbpVbst3nS/jfCPZ5EQ3IV73Ug7r3pLkPrE
DHgWrHB+ZJj/VgAo1ey88s9coqzKs5C18P8rVH/NZWHZks00bjWbNhJ3XGm0buEt
1KirDfbiESi0J8W1z0NKk0BHpAwFY/L5E/AB61cN62aU2xBlbZduKCtqYN9AyFnq
F/wpNQs9XaRd1h5ziyB937EXvu9SGN3UGE4O8rU90A/VIZmvvYI57JA2MBgAQmOs
gbmHAj5ssiEDIQFcvfgRZ7wF1Fvz8QIo6q8OOU+d9hsUJWGVE9KH+Zfx33NarjTd
hSNoVdJ/m6VPmxiByHqqPfwxlLQ15FqLjoQ2fQCWyUDKdF4MIYUt3sufz8Bql8aR
TZje6c1dO0MvHQVH58j+87x0Wau3myZVTSSXxQAmvrWjuBJ7pO1pWYa6LstM3l7h
yG90zYh2EbVBwYN9Gp7FnvpdifvLIh3F6tjnZZ3T8uXxAYxEHWBYOPBFtiGMR1us
8gskChT0vSFfsVz+s5+pQQz8MDZLFLkOvq8b2Al44GnG19QIBMjzedjha5vUGxji
jzIGlBJ9Mq7kWW7UVC4RLrQFlbkLQtlKHaof8aHebQHacjR7XX4a+4nZEi1pctue
g1c/eV7t7TiAfHxLHTg6VXxa9nOeYLHzwuvPxk6k/ckqJcbSuC5/5oP9D38jbeJK
wt6t63+0TWOsscjLP4aV5sg8uSnCHkTW28FHCJ+1gCANVxyFfKtdxki3n135lv9P
kwp3DzOHvIW6ebaikCSCu1o0vRYYRgZb0TzBXzBT9XGd24rIgjnrjJoGWQhqYW8/
Kb+G+oAMHeM1SrR4QXpNXHPhv3FH+daH37IsFmx+044rGpkFujkfWeHvj+Az4Rf9
xr1iPFcdHwHlUr5kQLGtEarapZDnT+O0DjUGZNVSQOnC5WNAopP4cPhdoOQpZMFS
mDYfm7wJyKXTOPkkMDPIYeai72DgU7KRHKOqf8hghF2AcbVrf80h0b6xFLERRU5/
BZDmgtaO5HecLME7lRwaaltpgyPQ8kDZHWNjQQXboVuURVlXYQXdZaDPEMekZgaz
tpiJB5PFv/AUAKBQku8GBaz22kLx0BTflxasXsEVaq+AaYvz16jrF7XNIl5OPLx1
T4LPBFOcdwnHR3Xzioiif1CqBGabD42GXqyaGSOfkK9jV98R5IIJ7MYk9lt5jjRX
K8riU9H1gUbTk/OdsppyD6CTtoFtk1CbRi4kyntR0u+vPacALtH71QT8iJzXizGu
yEzt1T+NVOSBbTbqUlhw2j7n8a6sRJmt0XXbkGZyboaDQzTOjysFQlkWYVQXWnWA
G1RWObVYalXAS4V5w7Dyc/72ZENjOAfy5o1eAFhtRm1gytj4Rh4mPo6sVu0iZT3N
/je5g3vpYgpKopCUklM2tqGwWMdxkv+tSuSnFEq2DCO4zw6cAgAP3yGWlqqj25zU
eGuZhfoNyNGOptaxLmHyAtUHl0jTLOg3hkhwZ1Q73mRUViBtF1j9wEAHj9jm2cUS
6T3pzqEahSpYDNcq3AyVLqrp98kItmF+16C4SEB+0OsO6TQVcjusTQM1E2XALTfz
ucvN4hnDyEZySWyv6pNgqYtTeQ/o1RLfZLEciX/hzu9vgHuheTbk2ny3VNo4ftdB
ilHegM26Em2sH+lNNVTOHYntPS/2xk7duP5YszkRSyzXxlE4l8oohFDuYvb2Bis9
9hYdg2D0xYUHERFyApQKVFKZKrbjQXX0Eh46poi+wOtm3moGSxaWf5Gg3eWXZt82
kiQVW4qiY8TdR33WrZAngxN6B7784A1EcDvQnxM2seWZEAuCeBVdanKJeP/9aFjk
tdIq32gs2WN7Z6lHCIvmTZ5ylNfWTjAgmkNAmiGZCtbJSvLR89FxsmR1CSudH/Cd
0fM8b+Hm4uVzCV6gXjOpdp7NtEX0rZJ2R4yVD0zT+PE7s0KpvnTH96zSHpl7Xy+K
5jmvC7fkscNAqkqanEhPkq5JBef89EqNTcXeoS6uJcw4JSV+NOf+TcEHvcjAnjN4
uBZJazVIi5dqxY7pL16iiBapaCdZhj8CkWvP0PlHQxcUHXf4vfjLcDptaycNYR+p
yfFpvLfyjJ8kK+7V9MLU0dWr3sKTBzPEwAj21Kagc/QpSnj/ZkGe2NIQial7RaSn
qYf//QQlfNxy/+WlM5p06AKueyTon0EN+ezVmpoFef4BGpN2QUI2yigF0vqwFaNB
lBCRhrIqEIkzm6E9kMSM3t6ytTOH517Mcp1Hq13WAzaTD2lv77tHO4TN9o515W/B
kICubOKGBmj4ZXTuOllO6EkHhp+GQOtZWNjHuMSGYUsrUdndXCDgLAXJVTE9OMbW
xz4UAaz+b5CTu8Re27Isut5UmL9PZSX/8gVLxJlCYKEBo4oW6QLWt9ZaFaf2cdVQ
zA6sgapNMDanUSc9FggQxYuW/e8HEGhA2C8bV5PwCgQmgpUaAWpEBmp6dy2pImOT
9VKHh40nysIItdU4E/tYEfoPrsJqrlZi4E8wuqP1oxWNd5PTCdIok+KmuqiGjxG3
GdJy//hMZbA1N0ZqYGkyqyamp/+zxxdqaF+RGQ2rjYpMgKLBjIUZ14WMVNRcCZYR
8oWg7+XH2rRLqqpgmjqqAAM0+3O3k70OAzSvCK+VquW95CAAVSncS3ziVxi15u8M
uK6g3HDdGIhJ3FZh35MzdyvR2RW495shgjbQVQ48K6iWDsLYhj6UJVr1LViKz1m8
dTqCiZyEvfHgm+dgm5zHXtaxdzYqP4Oyq9t3vPtKcyju0dJzx6aEJHj0bkGlEI3v
FppAGrEzyb/A65ltW/lH0yqsyAxotBsUHNGUMLvN66L+1cWwIHrhFhLjrassQnzA
QtWaYUYwZaEGwsZwCBq42DN/rwZd360svhC1jLDg55J6x7za9QUkl3PMAeOEiU6V
85untJQVqcRea3FJXsQcJ5ofBXmVQUBNRHqa0JeOYVWN7U7uqjJ0WM8YSLVCqZcw
Msw5TC87HsNzYzJffS/OdwF9R6WsQuZbtKqwdb8d0c3g7pirbfp5yF2H2nXdRSm3
E1yUEdCu5co/Vk6JtRYQFKKiBEb1oigQ9An+NvcBKR0h2TX6EVkL2oS+9i8yZyT+
C6auKeL7i4ZyZ9HXAGUCqmK2Ul9g6EgOBTvd6+Vie9mARtrNv47JdviIRNPTwirb
ZcIkb1I3sv8VmUFx7+9vGUQbaI5tcU/0ohiLg+aorObvFhWgXk6UjrzL0dtAlNuw
TC82gVkMOQYMArU+eXAgqA7Lvmn2bIKAZvPR6r/exEavk5MmQ7MWfvlyvvj9RC7h
szwkRgbsxVrYMzr3VSYy6qyGThMYW6CNorK6WFALctzdAuaLKRtAGO3biyJ9ttuy
Xk1pnFfjSO0eJ1jWECzXWxxdeTR1XJ+nZuWf4K5kmB2N4rxIPJodZCMvVGZPilMQ
1hSOBFkOvrPkgfrZqXRX5yIGQAv6ny8e5EcEUU5koSOoRtucZ/xpfJitKo1b9B/f
aw/FAq6amJO4AZCPBNYeAwSxYi6lSs9WCbLXuIQnt1lFM+AaFPfHSFCq+b2GnTeV
Mh1+GFk0GLjOQf550wLrtq+yTfGbzJSkUFuHzVUJy3SpqU2tCHTPJ85/UGS4H69b
4ar4BfogjjylXBV/L/hLrsJ1QlR9UFSprhyecdchJGg9LqNxXwm7nTjBw3Up9EcK
8RsEPYvIzkpupfY+p8soRo6nKJ4r06ILsk7PzLj0bCYsvjsiE15AUKiEpmbty+ta
DHtwVT2Y9bs9k4MdTa7EMEYgY6QkdqsyyLY5+t0+pFPXoz+xnLqOeV1L/zVUnf7t
hyMTV9ItMlb0FyvDNCuhN9P18n3pCOr99EhT28DlREA9kE0TD/RqQagWKh59ifNU
6/vdWXpBePB0qNx3XxljTuV85U54JNXGh+AKuhxXSFw21CIjky8Dms0Ar7vTs1BU
AEWfoFbLG1ZrmFgOzGjH3DblMi86mHCpfseYsVWHInElEYjfyw4Tgu3vPn0IqcnL
tE9MgzwgV6Yj0SWaWzczDmtYFDnsEBJZGftQkNd/Gv55XKdNd1HtMF7n0oIuv264
DWe+byZ4lvINFizxvxFva4XRSdzEZma8G9nr1Mq7bedigienSUvpYtLCaLRO2WeW
GsvqLDFlq3k8runNn1XMdNQOvoj4bUSCLLj//9XGna7cOPuyK462lAIpND4Bl8Lw
OSkKN9NzQyh4Ds4+KSTzlkQ3saG/r1M+zKI7MGaB6/ufPoZgJ0ktY71m+rbh+XfU
PcOPVc8uKihJlBLZ2IsdRShqvQRpdL/Gw/gPlQol3mLb8Vpo/3iMvicNFEPQ04TH
E8vmf/PQaVGPsa9C1thzuaauYqZmWtliXgtMnFx/7zzJxkfYi6jDGJF+WGOfP5zR
yBOL3vbtSeNHiz1i6AOmJZ6JQiPwTc6qjDXj6/bm5xUQR4YJh+zrgi1AB230hRXG
3j+HqIaEAWAAemDdieIG9vHvndlo0309UUG6VKz6mvHmS/OPDyzGVhnfeP/lycUR
4sPhmviv4aPN5pYs05qVfEG3xQ4q9SeEytiPu1gRkCp7v6U5PiXGbTTTfOqeadDO
29OPNAFw1c5+JeWeomtAjTFH9MIODG11lSbs1ZxgKFN8AL1TaDzhKg19+/+xkdLt
At3a4AuWe4YumA695SK1ScbdK6pPM3uiMZCjtuZmy6QPb9j+JxhJZUp0cqoj5kXE
Rylt4/D2ReRd4PLzHE1kQScUSO+2yFS5Mn/DGMBu3bDGNqL3i6Fj7VXV81qrDNeS
Ll/dB55cRClcNZoaC4huShBdLCF38+8ECHQqzSLduPH8RLMZqYsXZR96qM6zYoiG
2pj6YL3KS7L+823LJlFG767OTYMwSfm8GSE/bUoHCq7kzkILRJPwMv3rhjTMfjAQ
cX2TDYZFWPoPbpz4nr0bMnwUJo51Smt0DBTqEZAkIXuF6df7/2g6TUnDNOreaGfO
5vQU/VsfMN0+2kMGp5DeheJ1rcN8GYcqpTvybGSnwYdWH2WtzN4017DZ1RGf+jpw
+I/1+QDH2xZNW5DlTFZEEE9pzJ2gCYDWjne9ohTvogUG/xdSjQfbRInrZVLwTZb9
XNVqETrdf0zY8xvV9SXQcYhIzU119X5w8L8TRyT3ZWDj8owwccKaEtDn5ieQ4qwq
J82lCKeLanWN3VsjkRceurYoT6buHAxUACiexqOiTbpj5TRhz7Kmg7ePBtqb15Uz
vLBJoSAFK4YJPVs3Q6xYrKnR+3svwrrscxy8tx0I9jcdFWDSvZsR+gA5Izc5EHF3
Auj4TMTQ1D9gsMI2qw1N4MfGC7Aa5K2Hor8B3Pd/lVeBiYCt9NZO6irCyslzwef4
IoktZlVWiEkj6lx40az75oV+KDo7mvB2HrWsWDbs8N/+xZAPNJJmV42oDcmrNlSa
JxLw+8QR49nLwh1AKhPmV8Xe3Zv9nMobC0+wjau4cLZVY6JtAL0p9+Eo+EUVSAlg
JoFtz3wThlUyyzqFj47dzWKfHizVtIWum2ldqBP8WIGmGCI/Cwp6E4jWinG9WokV
viUiRia5kR9WUvQj95MTYqKF+M3tCqjNIK6ZUapytFXQ4db0feow1pZgHU2CbT0V
2lRtITfB605anfMTs2/RvrARtqKkJSrfdWQLV5H+aDdBV7/ks9siw+vySMzwMDtj
idWGk5soXwH4NEYrowlHnbXq47Wu5/t9dDnZUyRfeWF3pCNwCrDdTfGaxRF9CRBV
6cGd6ujznFwptDeFZLdLdLYnNY+I803TAW9wWHgC4SFBXPM56RQUPjtjlhtgtf+u
IBdHsttna5kwfyjStGiH2W9W9Fb5runRT7GPoRgnDrC/ES5sfvIqITNd0cWwM8Pf
Tfw/qV0H1Idmqv/Ome4UfS05GVRdYcwjrw+DMLIaLg00mkBLgDMmGmM6CsQYzG4N
u8TvCx4HsS19k62XmjhOO4EFkNZUjNk41EWVrHJzjuVX8+7ZNfuIH0q25Q/JGSTv
AWTQim6jDdhx123nH79VK10KRseAf0sUqupVfo3DYbeytG+4/9Iw+yjFXqfUtS3O
kYg+iWhDxzsY2EZASwJISmkWb1X/yOg8PGyrvmWET6efz8ctyYK/WVLNRItQTGsU
Tfm8DFg926fvUgAjtg8oNKKeHHh2K4zOGk8USfopUOdNGP+hu/smL4abdQXyXJHV
w9E/eMluzkpbMABuOlYPnxf2cLXi9o2cnV77JY3vnCJuevnxp3lsQi1LR3GXPEaw
yKoAVGFhFWiqxcqBX6G0SXAgTRaeXKUy6l/2DzLNAaXkLmKAxETLkPwxdYfdDr1b
bLBWiiPBRABOeIfXCQyPNSw0uMoPDTIU+qOLnZP6iBQ=
`pragma protect end_protected
