`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dhCV9MCmqMhE/FhBFV4PiXPTySdRanCfFMhhTua6OAeVpQlFodt6xwruzBi90MAb
6ItiZm8pN9TwRvanNAuefEZ0ZZ4BB59WhEK0i2LKcOG0fj+xfVQlsgSQXuFKez3d
zi60KnzCFQAA4S56szQ4+L/wp/X46HDisRTsfB2/HTE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3792)
B17uX3dNua15aYtKpzDkkZNUyDP+v/zabXs8qOg3zNIz1+yV+VdKU3mJ5LkBDJZ1
wMT7a7e55antb3ahEWt8pWAIT7xEid/r0o1YFKrN16jp/6G26rIFxhmOXkPFpOi3
REVgokNoiyr0IoZ828l3ZtHgyKq4UI7wpWEc9KkmlrhUloYwQuBsrIkOzsrByw0F
1s1tF8lQcAV22glN52czmawsNmlwjPY8s/9NW1y3uwRc/zH2vpgfcZlAuDczGjrR
mrJ8b5K5AXfHrYD/fRtSVnykGYguI6clSmGVxXqNZQ+07nU1IFk5N8FsNFsaOoGG
Yo/lF836cXrxSnJEhC92i95gPWuEc4AkgnVAUdB33SnSkfeiQ4hykCtuKedS7fMT
VGE/J/TbiMBA6rdCzrMz/15xURT9H/CSTc2HitexOTnjLKanENfISfP/zZCpokkH
VqFKsKaSSsMuhq2YTvfUT1U7947P+ZHYa5hI6ziKJv78SrqThk+8UOyXGBqqCG7/
NSBJWmrNn/2yp1fmvdXhJKs8plWDO4oLrRM0YdOLb6GN1AXe7ukPrZV9SzOm3KvR
owmOmSyrMXfNi3TUkr73AsIcdpe5gdAO3Oo4BwEYTOsskHlcSw1Mgk4vzEzlQVUG
LtVE8zzp2syDQjySyAklUTQKn+fAysD+OD7xZljLgwIkiyNXQTXl9SUNghfPlXjV
qjYrwMnYhgvResSuurDv7l9H/A6nxsFZTFwAWxhior4005gSDa8r/TElAcCl2GjA
YcLsVwzGmcw8wOX6cfxSz8F67O9YApXAcz+UV0LU8af9VR1KkJ4cP/BchQu5IkxT
nndMDqxCmQk4wknLDkItauLNa/odBNFDd9AnhzheBiKnoUv/Gqz+dvoC8s4B8l5h
LgbYJOD9fD215FTbL1wo9aUrI7PUGiTrZ99BsYH/6DieZJ8qZFOswIZxeUb/MeB6
tjUZdEW77tiHa+6Kmxih52KuHYahgBsMYXBt4no6Es0HSGaGwHFwRrje9xjPfMFw
TFq0AXxT18fFo8QXys4BUiZXsKLlQrr8ReAoTqoenIhtACYYYmM/VNn3b/jxK9SU
9tO5Eh52gzGFNNPIXWglxWYJUg56CPUb96PAKIeBSAZ5dr5G4La4qsZOHivjqzON
3Q8qIvHnUBIh1PYFxLv1BiqOvV4OypcjeYRpUcflhn8I4+7aUXs0dmWFiarHQGUC
5mD/gCUqU8UqAyjHvimWziNXNadWbNUrMBssJcWv21SGziqm03diDA3+HI48tl+1
OfyRUcrBEGF/A02RKa+QTISyCiuR70EyYcwwPcJ/ZNM4vsrcNdNj1phabT9dghTl
EAIHGJsf40Sj/z0IwEHtZ2UDZukngPfmJe+ElkrnzYPkAU92QVONq/KE5nEDmSld
QM9YiMHqdA86yPCYos7+AKjN7tHHysGiNNYiWpzmBea0l8NhKXzKTZ9dSb26L110
HCsNlg7beinDMCLdCk9qhAnSz/BBu6YFBjwyjYDhbyjbQODKXk5JRXgz//kS5pA8
Q4Y5m3XvUo6ounyh/4XK6tC5HMDXdnJ3CvgqQQP4VoOMK7Wc2yYmVBR2+HmbxT/u
hKyeBsihRRVX89dW3qR/HjfGv8LsEVl4FnfSQhokMozTrOvJHgQd6S62QNswW8NN
Nouy/FxBToyIsrjgPmmb+8pyi6oIYappouALWAccEHEpXfSt0m9lRxiFC5RbbRUV
3gIgaGiECkdYlUcxYTaBygF06mIyZfGpVkOYb6pfTz3KlEbYls1S+WSCR/u54EGO
PdlkCCr6xMIlv8aMVwcjKZXFvCd0ExMC8sVktlIvV3SmlnjjWDdcU5jidjiz6wMU
LaPy+/IiAXhx58EvhA0vi9Mc1RmiOi9S7sTjoug/SZCt0jTK5raFYdda2OYKu/IE
5JxpGZgWc3CKkppG9NWVY7Yc4PSHefbbMI5QrnQmNG4Fy9QPQNREH/0yGC0dJBKD
yRqb2B/938qKnjRuU399i+Wma/rkVijHxI/f7mbhy9bnbHmboMNvRChpuypQ9oM1
bHi9h6230yNNk8r7t8pLCB956Z8XoLZ7H/hb/IlU4QJvrZBeFSg/MTkPBDytyR4f
OL4RimSSLuxGszI2Do8NaugGzIFIHXvCuObbfegaG/QuopWUos4V2dQnhqFc466h
B8dypoUlgdJU0qPwbqaz/Se6YtAaU7lvyfMAXA+ochNScSQOJ5LfNQlrEH9qrgJd
UZCViX7RKx0u8+W91PMlsTOu/XynfmHnFjifZazdhrp9+FYLvsYdeCEtnEn1joof
78oVDn4rdxzKB57fY+irM9MEepoZ0sz+UEjaZd8hTgwqHMyt3bDrXeE/4KXF44fF
KIvWARhQm71YE0a6UZS8FWNhnfrP3UKD6p8swzmaHxASvKk4+/6XBwUl+DYUEG1T
K3rgWKh/taZVxheVoX0IerPCNdWUXFhQ2kEC0QmXX/zW2F13BACRW0TDaBdPkFTZ
jcWZCGB9LGtv/9uIsvwqfzHpGQvqlFAEItJe6dFCIpRipYXhLdiqirD6pHuWL2B7
tS9oNZTrWf3dJE8sas3EWfx9N2N/3YDBvZz61YaisyPgsm+8H3Zx7yguLlKXTJiY
sA1mpiicubMBmw2bTWdoJvobwe6TtgYOhatihTq7/Lvgkfay73dve0KAvzq7xajq
Btb8OP4wSY+LXFHd2P4pWKMTr0QSS5Vl2SU262HGvTFgrsLcu7ZanmbcUUPy+b6T
4ApVPldNcAKAAB2+ZK4SbrMZJozY1BKW4rESkfyMwYCSfRfDrgJHBSzpAczROCkK
mYw7ZDY8kfVTZX+vXHqkbvgiwx8ZQgjObtxcaFtZ1LgTWJkQ8iMvHcwGARZUWUZr
t5tHm35TypNMT6nIQlG9bM94kApjg/EpYfukzwzl9VnqJd5uP8k0GtNCSQUnszHF
N7qYZgFgoMpmj6h1W/YkbAsdhmYP0rAOT/RTRisWrm+uJebHXAvn3YUtAkjmsf65
oHoEYelLfaSdjvVQ1tXVcBm49pjB5/HnsZnz3juHLOd+FnLZ2G8CKqgbrwYqjazp
YMRFLYPPsq64MQFRl3uYTfClLfk1TfYnjQYJ+U5qxavJ4JV6RgbEbDdAqv4hO28H
Qyq1t+WfQYiLl4b8nwPacUP/FZgp+IzmWBuGAJGVvUmOoyAFaZ8wJBoPTbHlzAei
Ck4giEyWmb+5GWGXtvKwpV5cRvZL+YDA3BkL8XFmQqse9VUfKfg0bpL24YVgFvJP
bIixzTLKH3BlpNi2vkyvrZhQwMRUvUcdw7UlZei/jr+TvFZcgTahcPsilJo3CFLU
vwnb78XnSEL0pab2QieF+PMjta4E/hN943xKfoAvXrCumG8fft8S0ZUffrOMrDNY
Y3fLAsTxzKTSX51fCmjfNZbRi0hFcFUJQhtrRHW7Uf2MbsVMLiCljULzYoVYOcrB
myhyLpi5jkhtJaDL3YCg1UvVv8n7YS+ZUCGe0zWg/mURa+Xod5Jkeb+SkXF/wgy1
BaUnSA+Vuus951BddT2WsyajHvoDHvb0UMybTC692lCcLBsW5k5ge4Fr+vscZmfi
dYeedQ6/JTmY6fwFXtkCdC0pP0Zn9u/EaRW1H9zbWpJpy66zrsKcROGNEFILLwVU
btGUssVI6mVRVKER22uYqLxs8iX88H5R0rxJEnU4G1q1i9BBTFTcZWX2vHczXl+8
rVC0GrhPfc5VRCmzBAC6A54Obx9Ig2NEIwb46b8TrGuhkBvRqc8D+sFeYZshl91R
WYQF7+n4JdKG/73PD/dFE4j8AiGtTSHDDYGP/N/lRXV7nkpxmtbQZyJWHbhEzbvC
06+I0DI+0EW0vQrFT/wDB4IwTl4aCejHH2+58OG+tlA2aEEOuJmuGd+3SXVeRS7d
UA/LUOGnDgcGvfyHfSSWHQuyX5sJzp/sZ2yJ+GqMEIRRZ2XPiaArqb+1M2h1xs7J
l81YzABOP365cD/A+LeT5i63+foy5NswlcwuQCwwlvyXfliOQgOW9GdgA7MKgxHB
54pBzgDDF37LWSaR8FD22wWtAy/ieT7xs51MC0hjlpOhWyH7WwGrA51//JbCAw17
FxtvpVdEAC6RuxOGBo0KuiVmZ2nbZAakxala1d+pqPTwwr+UbIHQJ/uoW9kd4gnn
azsREteH5WyybSVRkbjn7qrd+AMX08Yg0Yrli5KwvaSfP46IEE/MlfZwACapgcDn
p6hw7JfIAGKVt+SyBcTNQNBABdmc/UgDqa8puKEbb2SyGXFa8GSBPnOfaZ8xrk+j
TIzhPFlYtOcYuA+bzhM9Diz1NR35Kl08p4D0DfHknUEIMscCovhur7nhCfJa2zMC
wcNkADj7Z1q2c/WOjcroK8dPUD3G90MW4gxspYim/zKSasy9FSPSu4oDNwe35cKX
uqo8+o8K2d7k4E7tOnDuobMNU8KAfcRRAB63ox27pM6k3TU8nKCnpHPPAMAEGxNn
dpHidAzmFaszj88EbkQNfxyCCGT2unL/u5plnhY803SemKo1kICY9IvdFYU+6bsF
y0cuURGuTh8uX2HjQC22g3k4JuY3cZEoMjw3rTnR7cmbImkm5yNeZ9COdEvpeA4P
eKgfko6uShYuPTi6LmnfH9hlohP2uWJa8GW2LXFXC3vfAUEfNtuIpKqc3kRgmKgW
6BqxVWa9CdgyeMxog0EIGz7gUqHLyIz47LbTXA4uMT9Ks4NT40kytbvqMeQOnHAD
NZvDR3oqXVjSNJrhroE/S8Ip2gMLmLCH/bQpgdEIMZ7kVpYBIpJjlKeIq4DpMGe0
YLpeeQ0q9EkLobV1kORuRhshW84UPHJ5rixSryQQmrJ4YDYuGjCfDbIWG2C66XkM
slsY/DejMEHJtJ8U18i4AMwsP4X46Wu8aDl3x9JX12hr3Epr6/TQqqMoIP7dw0tH
fpJ0NVfYYVuqybRy8Ar4w5oVV8R+b/adNzG7pwWviW0y7i4GBoEQpnS8eBE4r4Y4
I4FaG1HQJaQ9YV6v1hVZnNpW6PWXq+O9SPZ3RT+vS4HsIY4SjMnR1nYEN5kyr7VC
`pragma protect end_protected
