`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kFYQGwceTlbq0fnahQYDUHOKSv0H0zSqZzgyBLWDJFMMVUByIOO6OcmX9zo9hZZm
tIdyAgbY3GaV3j1f3ayfGxW6OfBnMMG+Tv7cSbCTB5CV7G0gAvFntnpFdTVeKcga
uwGVFFiByeQ5VvWJOfOPWL0skynqyGm67APd30wlNfA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5344)
ylfOPKcHlPqiSxm/D3X5UIF0C2H1JnCjvvdgpUEzKVrzTj46BqGMJHtPNSWCOp/1
HCLuorJ19VvuhmksJw9xt6/YLtNiV59AIObRAQ8XhzEIq7XVlhELI/swnxqUA5zb
pvL9xXl6J5+CxSHf3oR/KDIwwMAKsZR0iNUrt7bF9mEnh61MjsZtwmELgEL5BpQX
9zTeH4gn77/Byj/L8jMqtcJnPHFkunu9GoEUBnVnYj8SH/iD5wRWZMkq3Yf5BQbv
DSy/BLf3c1OTWvDxVmJWVc8gojls9ll9g8rhZ+cyBZZq1Eku4Cf35UEzU1HAT/Nn
NFFtv0B0/1qxEa4nW22EPvQfzoSUPAs3uurZcvQMjUTx9wrKuzRZZPY4eKhOvb3N
QcYzz+607NpkViQVwm+6DDbGQT5Ls0DQ4rdBYbH3qzNVeEKaEptS5OL6u01h0aNs
5tEkwp2zTkjHIr0kb0n0lxKprAqotqSi0ZGxS8TZSco7iVN/jY0IjFByCG018Ogj
fhEQEQUSksIxDqVWkFrJKhwTjYNAyDE2uHpV8QN6NmWZ+06wW+8Lg9t54U0t+Uba
KEYRFX4rHsCjRqZH8JgaPti5qpasa+Mhez8XJQNkS/EqkI8sKyfByXD0k6tRJqPW
c/dCEABLDSsnVIOivCmwIDiV3fDbJlFPfF9AXOlrAsI9IB8B1ZKX8guG39mvDZaX
LHsxEcvgaRKnXy6XhcfythQTQ49r8lpsepmGtdzKaedVQZTlvbPax0vGj4P44rit
uwjiinGvNzRgM/yHZHGYPP0Q3dlwzqln8/HZZIhAUfFV15cxXNImBYkSZO6fUeyk
UgnzaXDXQaCnYXdU7xixyBNs937ZtFporQ3cVpW14PQibsw4XxQ5rIE+xjATU48J
wt1EWadJSMWbCto0Rt+PvuL2GQkiTafClUHIEgohefk6X1x8tFzQ+fGYnwpyNjrh
7a6fadCOPiQ4evwcnB5xWZxSpntEgEtGApVIdi8Xq5cOXg+c3p9ebPV3HTzYHBbk
QSnJ0918mwwrzYKeSoP2BFCHIg1tyXMgO3l5IZnDw4zh3zPpkv7jK+lQSKFSUmmQ
cvoGn5l+2FUimrbZnHLnJyqMeFqQ01RSnOWFc6t96GMMabRhUZHoIAYdDGUS81AL
AAn4SA4/9ffGny72WRMp5v+5rrl1wCXg9mdJ+JYcWw7AFoz8driA1omtaPzVR3UT
YiDK5AOGov6EdGUkNpjcJozdSThw0h/NCzR6F9w/og9rIVAbGvwOHVCIqxoWIxq1
YJOFRua30P2KEXtY0K5D/y0DavnSv8CPH70FPE6pxiVysUTGtMx56XRspU+cPpwd
1oOxwfTYybxoccBPV08bCo3e6IWbf6Of2TAR265Z2Y+lUmhn+7D1MUNTdmFTxUmP
rVWseBujxOiPuUhLJ4DRNmtgIVtjgF8RcpImDYSoYPfMqrLvOhqtMaxi/bBJFTVI
0UfcRdX5H0RUYWtPYqHCNL9R604hrgYYKbnS9tyInnrnr79Q3fuSuybK+EjpNBXb
mHEzOgm0RHwDoR4Xj8S32zdb2POSATfJfbu5JxsYhDoWHAdsNegA/ipV5oT2feiB
dp2m5XQDmBcwtiIFracoVSSFLbgh2TIMh0VU8VDaTQwuS09zwFSs/O/4nEGFRYc+
mfIDTOilDN+bQzLSLDw16srkb3eJKZ+j+47l9WyAsMzsjzd9tpF9eU3yUpsh5J+k
+wOsPwYg/ksfPAeDOw5N6iaQn2FNykVa9e0DO9SHLp02Z3mglnRQfAnnpgz/IA00
mE3DlainT4rXTWg375mEeW0eC9qQVy8Cnqv2Yt79q7m3CvYuOny2YwjK2S12iexN
ufd1MZgqWi5SKU3SjQRUURX3dI6KQrPOufqFN+h8pJr9DLl1Lk5IKaB0/uJD29rx
ldPUIoeRq3qbyLwoMaG39eifpY2vwzyK1StSFEpVBNGs/lynhJi1PNRww9SsmtG9
83Pec4VIGIxgoinJbyy/PGU+BbZT/N5rNxKVme2NIcHEKEz4YJM4vE7oIKtVy/xs
PKPp18QACDVYmG/eIsRzNDFMxDxGY6ZiyBrr4NfzC/ZysHF+RN0rl0JS2lOKJulB
RmnmTpsxtEEhzyZ3Y00iSVl7pwa2VxCWhyNR14RxEx5fl2G5S+0r/+YVXI3CNCsG
5iqTQz57CQq5PgftPBU8YFUnsKswtTfCNwgQcBUbrj6KnjNjC7MtY2rJI0nPwxGr
kIUh/ATmZdiwiWAUJh/kXSGuC8+svzdek50MeqUpG3oGDJ7SWlYoa+9dnTFbXKiL
kkCLPDuPBpLSqwUYXGEFw3v/TxFOsDDdNgjk5XXmljuQQN+g17pJ//Qm3G/8Hfdk
vsSDS96IR3T2KoG63ZQvAFqRGy6wpNEXW6kkKVjiEzYBrpSFJLSxAushxWr7ANH/
Oq0NNxxjOCRLgAV9Lx8zo2f4SoT7Kl6bTAFpMtYiXC+dXvJwLt8D0al/Dn5Y0b3M
2eJFEgSpWM6S/g+iSG6Jzp/Oo0AXbIcD4X+DtbyayMUs5FKoIN5qC+W/1hxXuwHa
BpEX1ZnygFQkV8SgMrMhH6GI2F39Cd0FBINec1ZEOC6n3xGqeC4d9w9Tbw575mop
Q2cY+k/i+OnRAEFIeT0dW5mzN3CoMWtU4ir3q2+07DJsB5lxCIXG7uRpTzJIZYT4
WS1B4a4UMkTl9oap/T/7QQ+5weAuXRs6Y1ugK6wkpCI1AJNXw86IQIYXEV1B1keD
L+g32Yym6NVZ2MUbTa04IxmyMpQpM0C5+aEHILNJJdQDgLiWaePdakgJuNtY8QJd
DQ2dXEXhE6vATTKjMboPTVHQe3Xy6NzxIlVxp4/3iTrEa08/wmlQlOXD6B9A92hn
Dq8Mfo55yT45plK5OQeY0kd40dxTz4p81bf4cJJK15BuaH/E3gUS3KZSuRUtoJL8
qRLwuCjR5foEbDJt/N8pcT8gP6XyB9uQD/k6JXxqjPhura36hJ9vsrojNE7F2xHZ
ROlJmleF1k+WgdmAEVgHzHyUxvmq5XHFbnhdKjX6l6EFrAmN/LuqSfNwS393tomc
S4xwfPopcyavFVFAswu3DH/Q6ite397Tkf9UtF7cYiNCTJKb3AUm4lZH7h5POB6N
6LK3v7JcOVkhFHjfjBnlDHBSGn486GmqSfoGzamQisrs3sTuASZ0RcJb0rPExF3m
yX+9NftLceHdDgXIp94MUC/jwHALYu6p7JzHxmwuRT42m1Pxdh6V6f6oVuriLYta
50UlZjp3F7l2mVQcSZUHyQrL76bSCCXj2dyxNUCoqsfYYG+fuCqynXZQBDUKmAJj
iIQThmVV2IwPnDf2t5T/nUoL1TevBkrCso4dfp3Uwy2nxDvto5o2MTM7ayzUdczk
PnFZg+VRcnqt/+EzlH3aB/e8I8H8JQl1/DSXlEGjY646B7tW23uVYD9cyTUkzAu2
cQLzwWdpMe8fjqD2mGGSQ09VgMHra+2syY2v0FS+MCj37mRUnQ+GyO6L8a3/5R//
4FbnvgxMYCtzcDxM1ma6fqb2BbP+CC1mxdQ6+SZoDq1m3jLlrROH4xLftHbaZyWk
jvUIvIm2/MszJB8NVMgA4PEH3Z+SNSGX+tc8tsN888sxR/nfgkuDbPSgMbKxomV/
yA4sl4mAFNP4eHX347wLUEDm/SlIIhpu84w+99xJUwWIBUTZ8Ovs2PW22Sp0l5oZ
cH2s5PUUprcqc+tZjWvdr9NC4dFeQrIhnGKSHEngqDv4zbDuv1NGpyBo1wJJUCw8
BDdmBrh7T4aNC30dxCJlWMM8nGL1rztJQgQu8CyeRrzUBijKWOIYRbAODZD5+g64
M72u4z+nU6+Sz2ktMa0p+aoP8/GyeV0tcNACpQ6OW7i7s2KI7WOT7dAebIwfziut
E5GFHnnL+6PP/rGm2rfvXEOd7d3ctgviywNy6FF2ZfIP5Wi5COEWITJRj4zFQYa8
OpL/RMnRqhgGDWZDCdTjNznsOGAdzrbn1CNEj54Y9nW8Fs2iTu9ZpukGxe4BGeDe
0VvXJJgZwod1nVOXxS24HfM+1P1WX177kEjD+iLYolARp/omjgtBBJBm8QooAvww
3lCye5spDnup79ySUvSaYbILL2Hi9JDXzAu1sCCgPGMPJpb0tsmOiB7F52spMFQi
gsZDW3+KuZOn1QvgqK82c34MZ7GiuJwhqqct5K3A+F8Fsyf88ElO0aq5Q4QHRPO+
zUNrVuNe1ntorVfBoBH7WhBpFSMmfP3P3DA1AVi3AO91hvn/6oAml9j6RTqWPY6M
9mx/V/fISxd8TuOIfANLbI49h3z2TFNkD1uIePxF5aDfldn+eGguJHxT62fU5Wnj
rWx/N3P74LKYpudRm/a97e9b8hHw9ymUw/jqe0Uc3ioDNN0S6mPawtH5qZkmIgq6
vTSJ+so1Eb5HJ41dJeDV/hD3fNQ09tuda4UIpG7n0wHAZwfQAKwW8MKs6516OLlo
YEkaaHYB+cSMLygia0eraci/VFoKMkZqlSY+f+AFAuPQJtT6Rm7VreVZyrS/5QCP
SK2F6/xZLJ/hGOx8AkRRprrDrfHE+RcnTOob1EhjMoMewI9llBHkAYflvwO2HsiQ
RRwvBqUHZE+Ek7/PiIcKnHNV/KGEJBM/nlHV6i/Kcz/e7d2+D8HBOW5ig8WFMxxQ
cQzMN3vFff0DhAl8j4/P8e5yKj4ZZSjNk7tGFEcDBCRZyQ4LR6+QAJmcoSnv0LjX
0X537DL3/RrAhsYkp1Hu1j75o6MHjK1DHr4Rbvp8wrbH8zCwtrY2utOL37cetftX
CCElAybKR2f92/ZHRR6T+E94wV+Uj/1BE27QEHCs82PO6B27+z9jOD0GdBiIIXtP
UwcELdVgB9TsKJJ0QmcgyZ35sSFKFpPiFNCwBtY5A7cUkLyyGRNlf094q+OdMakw
U9sBfxkbmVmgHlDN7deFLkuEkQgXAMdYJct6nXsh44vyjlYNxE4+hri774xro14l
caBXMBYdC9QjTL2/7R53KJbL9AW/3agPRcVFhBc+lcOk5bh2yUEpL4SByvub+cms
xxyH840ahBDI91Pj7/fj2zCYTaHucY7tLCbjeSt4UOYBFKkJFuB0TG6LYQm2qJ6b
6/0kYD3YkJwPDBsS0GQ85KxTrfSuwvywbWc59CcPHCCRRB+I/FsUDagz5MaJGeIj
jlnHTnaf/6Y4r3dY8pniirppOrJcwO91/RTg4nhzq74QlZzN9dNf76nCkaXFTR5u
wHD4gF8hv07nwFaDK5OWrjCy7cwbbPwTcc1YGU/tDk4rRKI+RF6pY9mq4h400xH1
ZQ62H8ivARWa1B37b4InuzWZY4nuO4roWDn6KFYTs871WYsL/bm9p55iPWaZgln2
uwFZYzHAu0WEPJ/wkKuipn0RPZaeTWHKvGYI7MtuhaBNNsL31O3PrC3N0v5sUZ9e
Fn8i1kGbaJ4kQK9kgNdhH8/pKnBnqEKkbShUEiHD2bQcYFt7bBo9nC+QHZdCxRDS
XCHN4AM+x7aobp8qq10Qaij4teQUm0VZB8Ku0myEMRUOnlvQ3qLszAdkfLGNQQzS
d1KQ9vN8Fhl5YhT4OqrRjHnWGEYfvXa4sJS0z/aQQcqNJiqVtGPeeaJKMthJA4AM
GLNAXr4cN3/UNl0kvHnEkxgHNTaA8SxptXVs46KA5TCltunVKXTAfSKQUwJPk6Qj
Nk9l6cHESa5xk33QhhTA3O7yUQQQy8XhFWzH1w3xSibPN06FKSpIeNexHWuvgOq3
XSLVF9sBgMBe9U3TD386zKIoNc/H4jgd8Mg+BIP0UrzSibeFr3BNsHorO1fQ2a1i
Ff8nZPUsaUVWPysh+2FMEA0yRQAgAJkFnm9dCjN2sC4o50bLrV5bXRQY1AbV6WGR
UjJpvrNyR39Z2C7C8fWLHgDFf8bjzo5g1FMrMkXSs1LUttWQvtTn/4DoFdYDDFiY
RX0uixTZI9hXEIaBSclm/5sjiNupjEuCZ9/E+4b8EypXQ7kk7uajW5V+MAbf+dEM
2JWcQSBrDOzgnxFaj/gvW446QpfDpBMuL5GCpmABj0czBjjd2qEYadTBw6orSI72
kFepYhTDCtZ2MZPfSskFSH2/CsSSeFhV+O/nXOrAmblWxtNUk/0MVgkH0CSDroSd
IGgEGKDlIQ7fhzpagXCCeMz9o/SRBfiqGlSZKTLt5I1JCcKnX/B7bpdoZLS8c5Di
tZTiZHMcaCwEqk/zIJlG1Tr4xR8776u8Iawb4UGu9uqfVDxPh5cO+e93MkGbaENQ
CVga0zqsoQ7MnroVpoa4tiIgraqSpV8OXmmbXQvp8NDq9jNA3XVWU7d+DusN7Qyu
Ju8B80HUaTEfu+tUkW+2Fi57jsWRV1Ywkvi20e47sFgZLzgnM6oZw0c0up/BNU6M
0RkxiEP3l6/V57HJLgO6hfsYg2xpW5diOPlyPaiD369HWHNqrgngzIX6F7q4aEos
cM/mRSZHsZMroldZmKd9CLPvAL3TISQqpRSXIUiBgpBoxotkDVsAWjDJUH3cOYdq
5QyCDDPy2V/z4cnix0lgdpz7RgbePSB8XLjLSQKGdVj9NBN3R1YxK2l8Ugrt4C+1
+FyVAG9V/EAaY/0vcbsBwOc5i1mkmeRiTplOWjYa1K63a9zMt4bE7v82XN0Yt4A5
DC7Mgqr6ADesOsKsNpFndBvvjZaB67GuM8N5/IbiBNMyiOjaowBcjiLnVVQtATQa
L7PSZ2R+7fv0mCmsK+Yxg4MgKNe8xaYunmWDJpjo6dBWk5mbXAsYvF12Av0hnNOJ
k05M+5B7rRoKeXBRmESM18/Bm0xP1kRxo98EwVAxypCoifd/KN5L92iOWB2KUKuA
spZOKit/LpbB0SDKH3iWhY2qas29oBnOWhBdPOlBrqqjtJG22cqP1/R8AC7ZWi8Z
BkT7UrPmYJgvj9YZQKef2lTMnBwMqbdQHye9RjnvYEow3rc+tsG3JYYcmI7Irjc3
ZiJQVyZJ+h90ECJqXUAR+SNLnxDN3lUAaN7JapgsyElcY1rmNZMclSFiGbw3z47/
rLnA187LroA4NI2iS0D33QjNPJzS5YETwUvhNsULIrHkWgeNVpeyhrUci/xBanVm
ne7qESjLjhvENU48awnuug==
`pragma protect end_protected
