`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rZg3N78bFLbNTLb32LJztCBBmYyeuTczhcvUeeuhIRTkUYEWu+rjbshSD1JbRK57
J1wg8sqyb21WiYhVffVfU3BhVDLleLqoWpH2trUHZgsVvhVC2tH2Q32xS/JYIsOa
5wmO2V7u5MpWJcUj1QB+accadrbJDh9qVQqomXhfI3k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24512)
dFm4EgTbNQo5RuJYfgVdjKwzks2AhtP0gedEFsagg7/BxQeZE1/xFbexBOa8g4hk
AUiGDjLn46kMZsZaGyHoqXlCJT53bCsdbnlUro3a+Ikte30UwKtN4Htj/vneCAn6
CwfNtsSaPMrItk7C7cO2bHT1g0Le9V3qVsqfrDU8E5QAVZlp64aL6oIksLTqnjAz
Cmhk4sZepnUiqV+gnPnPst77avBZ+vbR7NvGXGm+uUuJFgjLHS8MTBbgxndG2ukE
85rDI+V45CuPXKJuRrva58udOE8yZFoxCqXQ8RmvXwdVDchACjfj6RDwZnDDpx2D
K76tu5ubfpDv8io3JzUUE1hIn1rVU+JwLCnwMhLkBHM+WyMK9IlFQtSMDVfXI+0z
pPAq7x6qmEbhCisu926EAaENfBPGC9KtzVaF02+1EVdvT0FS/uieReBtw5m4WiCN
15R05LwHOw3dXqQ3rSYCeroGmvu9HR6y7dARKIlPQ7najg7Dqk+86iy08uhwIp6i
v2ElIbaFi5krYbwTtWHVkwKk2A7y5/DvrqkJIC5jvVdVwBW4MK1Mjg6ibeD4aIfF
biVLhLLwAxVkgXsQeSvTIa+X0TPTKICawMcgfKVqEmVXiAAagNVCnAl2FRy1aN2I
nX6SbZNyxQgs56rFWw9Dhe8mIPkIukAD99l6e3sJWym9kWnjmMnEd4IAPy3oYVEO
OiDu35814302wbJAUhJRY8GJ+rV5iCo2jexskcOMm1U23WyPbyXaTp6JFWASOfuI
n9q5F3G0dC1q2RFikdyyX+puJeIW075aksK684iAPY4CNqf97rneVNNGhGVLQ5AS
JZgzKXHu2/HRMbwmi0JyPR8zN2PtO5wR/t4ZqyGCC0vu75jzeEjGQfMhUuc2Lavx
sTw5bSsNhJLHY/7jLYKsUHvE8Ac1r7uWiGpMJJQnQDyEixjHM5Ce2CqgwUdLTplP
ylShxsQXlZNizMxTQ0tlLaLvgD5CcEtf4iTlwKgAiVjxtWmUm97PXfoHBhCqtyII
CVKIpVykQhtMgvTFSypBUF/b4t76XEEglgr6x7BfT29hayDxzIv4zwnZjJ6X3CFg
q7KIHxYwR0yxbYomrTLgypL84Omz7b7aRctSmc8HNBwALk1k9S9PGas0aLrodoFn
PzyLkNgwQohF/mOBnbnrP668byps/Xab1a4KHIgorGsIW4aQP7M9OdAYGxbH28jd
ZvPbXRm1wgA1qWlPd8l1RiqcjFio853HV1mS+zZjqrsHGTQU+HZ21UVlON/hnAkb
FdXsxoqdi8HYukxegVlBGun5X2TCSg82XUQd0zq4JtDPP2Nb33F5ojnzqKXAs/1Y
i56myiFmjian+32WrcWCILQLawLnmzFj+TebzyxJ8ijKsak8rGyFKX/xBCkjb0a7
82LSCva8gXStRTCjGs5fhMgbyG5zXo0EzXvuinxZU+xTw2MT8JlQ7jZid9QAcyLW
JGhc1I2UMOd4Ny6jYmSobp29k2locErUyO6JDi6q+iXFYVKKNF5qJOqFeGcpaMKq
2+6KnUELNgAFdz79/+Uq+dLCMknMlIUSEvtILrVxr2zDZwOEIpzYSf6diMq/ewTt
wC3d3wx7MJIBnboeWTyXWiROzVO0IXC8jsC13CxoFfCJZFUTlIlkzHFIGEfUtY2R
/CaVKc2Rh0e4dqd4qRSGM2zhY8Z+yEczl8VaP/PEUv0lEhUIL+MjvCfi4HSDmPef
HlwvmTS53EBysLgvC5zZpIkp8gyl85vp7Z6QmSF4BlZ9sdTTYJF/mRUIBoEa9qhu
FHc6F8AtsEvWhY/0bQTsqS9Ps2YcM1NASQ26eIiXNce3s/F7nrIQzRHQA150DTkc
Nk0uRl4o7O+tcuNjlDq2efpTfaNp4i0wkKDMB10XPR5OIr5+5zwrWHByfMZc0KCU
LcLkZMlf1fO5oWJNlBVMYO+4GQ83Oe2SrJzAo7lDDp27DyOVtdOOXhhKEntBMnxY
c6ROik/rhrN93rPCOUyEb4a0WyYPqqSdt7t7C03s5vjDkIWtEwTXCpcV9xkHKqLa
NSTTxs2YG8B/pXn04KTIrbBKOjK595X3/PDcWcDJv/zPzSDnpltEaxSabZ1ttaIN
mLFWRSe3J9c2AIFKMMVyrbeXaI99segYYh2q8G1Hm+LdurzzTSIcSXvxJLnI8boT
I0kFCdX60/QwVJGz7mqe2ZH1f3dH3YKHNZo/jwfeCgSQpRq1IOIWQ3bF+JgVufYV
6Q/jD/fXcr2t+6X+wohb0+P9LlFEztoHyserCAZc/TlAneQ1L/9Dfkf/h/aC9Xlp
SVkObkOiYY2TyLuhHwIgyqYQnqWtK8WNVlx2Chg4PZmbqrYsHPbgUpfDEBts41Bu
dLl/cCx4uNJW85+8OuH1K46dTceZInd0SgrqxIFdl+9uvgB+/SRHpf7R45BIcaky
jxqDD2G2vOsebPRplPtS7VyR295YDnQWz3lTX6EMcW6qlb8OM04wDy5WpAwBw5aW
wKxKzalQbu1BUbN3aRhU+wZQdpiW8Z/eg2Wny+9lF8yly4F0Xt2cCLocael5O3pl
wGKci/4P/ZnJatFClr+/FglmQzr77qLaucV07+lksIPwquQg/UU2uC2Q78hcSqjA
dBJF7W08m78WPUnIL4r423jneNOglEwr46vD3UdVpEcVQQAA3N9dpngYUxZYA4ii
UBZUZ43iPSRso477uKcwxhuxLEoDamGTMgHdEBuYE7bK5KAv7bke1ZK2cTZeMSNw
ftXsET2srni3sOThevX5xOQzVEllUxWM/ae6f9s6mB86xqxqQngAeryCEZbB/86I
fuhH/N5zFYWjt3MHe5UbLakPgiXs49grnzze1Y/iN8KDH4jjLGKvbpNDLRxn0ifz
d255d+dc5bBhuWmh/X72drPBX8uXByp38RIBuUbI55apUf8F1Z0Ztnz1rCPkrbjs
tUXfFnkn+YZuS9jRbhUGOGdU/oxZIOWvYlMnONDA8QpdK5w2RH+EctrIXnUqFj93
XYmLAZME2brE7VIiqB0SNA94KS9IfZhazz9XKL+GzDW5P4GuveostXaqs+Mmuh6+
UYqfSkTDQHYv6ZtBhsiskUeJe8WVnCIQ781T+ts0ScCU4w+AttVn8OmTMInspPU/
uhyZ3W2xJcXUf3WUHjGMa1xFGyimCji8N1YqQaMoTnzWuCs17rTZX7DILexqogcY
kYl92yK4xAjRBquwiVyTnHozKe7wfrN9JL+NAmIDjdFiI7BcMgitlEpnOhJOcyr1
gCL0ztbW8wH5Ew1SiAA1P9EQjFFPPOIMU6JeIOIDhWy00zYNx5/Q6bpRqom25ZEY
BkWbqNmX9ez8KchvYiwXGArRphZum8+ZPZYRhJvRK7tX90HE2I0WTD9EtI+FducP
SnBmivUvjgS9yloHyLdb3Y9fz15C2FqJ0QDe4Lix0OiIRyjG+1ugJUa0v7B809lD
Qf4n1S1pZXp6QFCRkk7yUw0yH0Zu+4/5vqYCvh54KP3jbQGiAs7Rr5okDqrf/qbM
zrj45T88fER3f253tJmt74nrip4CohuaDSbDMhzZiiTSPAX35o11fgU8JM4DtOzA
177ckS/iDh7I/4HyU7ovYBeYjh0oM1R7QkOMLJIZyLqLS1sMvfUvKR+5H6ge3ePD
mHV7E00afgsNZl8D8PfOw6Tvk38NYnEKEBoZssQ37Gyoz0VAT40XIEaORKvfi/Pn
MRC5DmQmicnkEaAHhkIyYxyzG0Q4JAwRbsaJTnKRxJeMYdP3surTnDCeKZMp2ikd
fxvVsYb4I7bh1kY4eXxcY6jhGpkzz2XsntrkjJWQVFXu3iiud1brGXMjhzs4g78Q
Y75D2apsItc7T7qj3FsKYIjHF5muyWvQkhsMv+OE4A2kiQeXA2IAj+0v4fY9miDI
jmUIkvJSm1GpLGDJqLQU3/NvqHolzKNQhhyXMdAOHhvcgbxOccBoamYRk9WPjcD7
yB7Q2fdYj+OrR8DuFbK4bqwhX86N1SnChUvEm6LDH++TER12UbErDLDuimQfJexS
aRi7+VujEP0b95c+F5MxwDH0w1/OLhSkXitNioZKa1IfRSh5bg2v9PhHS5kZYAek
8Iz7bopSGixQPIWcTyEx/SimNvlcSTOxmU1RLaH5gogxNyTi+mle50TPM5rerFuA
eYAEl3vEOx/lMEn7qkpAytIzx+dvZolUGyOldnNwAqWIgY3gW6Ue/2Uq0+irGcJw
qw5enmBY8QGIsuTDHS4lKWrUX7272lTABNtvnhe4OMLk9A/vDMJmYLT3U/UKZ4+J
9BtDUuouCkKBnt5Vjl1L6TB+OWVk4Aj5n+0oWYyUuEQnqgzmJIKQpZE5aMrxF+HU
GIR2LoUTCMOLseydYC9QpQEuA+Za/0nigjzFFmcgLhJwagaCnDhla5jrlqPhMyKs
739BKxmgqMVm7Q6+LTGhv2OKtB1L3nqUP+xwJOVohvjAnKTtMHNV5W9wUhA7uw5S
bd1COxNeuAS8doVKe8jvlv8Q5jln/S99nywishutuSAG3VshisDpzsw8RdNEkP70
U4vt6/tZgOvhxlv1LKCzTqF0M0tZZzoZ0ZiCQsZRw7hv34Glv/C9N3hwp8bWb8Pd
YDojgupD04yknNWuqwfXTJLPTDXz3tJMDpbNdqarJekY9ucDMR9IiqQbj6+BkPso
nYm2UcFseMakJz4dFmsh/UDQfvrfimKAVnkXef5Po4HUptu2iX0RMpqLmJE5GC6p
hbTcnXGsjrKHa4jgbnE8USAbWVeLAbWrAdG0ExOLKVyLSvlaNlgZcickiAnzPjz4
x5CiUAs3/En8NsawzeM3weoe4VH519BSjB91BlDKQWB4obO9NUEImDzNzl4pAItw
kFq5tmpLcSaERiidB0lFeEIipd6Ci7Q8fCT0crOlapjzFcURAizeUcgWfnCkob8N
Zi4y4UaVn59LXd1Ro2lQHhVtFnhPwSG/LWLFwna3QVQXk/Kv9O0lwqrS9P81Us6d
OSkiAUjwRgXX5a86KVr17csiQQYjm83XSp0ASWezvzoa8EYAfn6jvbb++R2DTdyQ
Esnlu3BJnuA4OaXMibKcFj2t2czt1E+gDcP7+iscSWjkAE5i7k/5nKpy7qWD8moB
9jxgchZ7ndPUeNZDAvB2wWQrPUAgffS+ea3glEg492WqKQRvj4A4VfD2+iliKQpb
FYllwfrLB/sOqG6t079WDiKGM2Iq/R9AJrjzfhNweJtVIQAEWc1Z31KA0wT5Xx9A
aPdcBKTtrv8c5gDCQW07SfOoamsHZg0murqYj72yeXBwsK3HyOaLf3XPv7oomWN6
f6IR7nqqOp3uIxkSIe470frH6q2Z0smrEnwLkQZOs0dVAHo4D4DYO1sJG2RbyRl/
edmNEanq426kWbg0x8IKtj//lK7eHBS6sVi3eRbN0gtHVSS5rFsPQ/WUQdvkUjHe
vfdkCQdnQ9vxPKywMDCQQkDYALAG+kr2MYPhFcTaX6ujtl3drKWL5GYXou5EzYOJ
eq3N2HUb41W4E88wl4eltMMDZW2ZDVKu9qDQY/z6zlxFEOoDc4JeJ1JDjUx1m8n8
1xaqYENAaSVWEiHmxWB5AFYKk2/rhbCwQJhymCZkYFlFY1zg0B2R+hXSQLl+/zWy
fpg54N/a81jRlzVCZiUa4A7kvYidXvPqcCWM8ck2zqe30Idqf/3NG1AIeUv9ffiq
gtkvbYDs/ZJi8MPqq+tUNvtWyKqdrFZzUjq0f9GC4m/whbZmwWBgYP+TKyYFDOgt
jimv8of3StXEY4l4vsFW7cjJ/TFVKHvsylAR+Ae7mjaJtp28E3eP2P2M56t2E41v
mCz+j1GtzbZSRJhU25XDi0VJiPqgxRNRrj4KHE3fLya4637he8iFWeaCuIPJRsm6
1NxcUCxLjKH4gofut7A21nS2inPFdvy2Jcg8MkOgEkLWoYpIKN/wsCKxGnLWthrr
pLPQ5VqFo1Mg/dQ4EUYIhrzlVUnWZ54d7HYEo/E9+7F7/TxDAX/vg2UE91gT/6io
LTMwLblBHWIwGC3InuDr3QCcTYVgdSr9S1YGCJAg7n85ZWZMjQVV72CknqFcJCYY
4h72i9vx4MZOTQD8ZYFPHqi4xwoJIim7CEOQdKKn+mB85vcxa7u/Ks9SReqVzlDT
s5VNq+cVUm+A11eDXI+dY4RQvq5HwzKolinQZl6DWpSddwhGlxiTOJfNi2uWm3jL
jNsQsToHcVRUaRzcFKj+ZKHpzLTnZE/xtHEAo2i+0JeEshY3q5vDsstnr0w9lQ2D
DfJIP0w5AOJws7Rioth9vWROL64L58oPcz+rf4uoVRVlI59dnYQd867pTrLsuWUh
BtvgMTnYeNdn6ZblWjwC88dimGPNBB2n4D08OVEQDhL5yjEXKAb68iBY9iNgWy+K
8MBGko9+oQz+zG4xkjaBjWrKr238i53AWO1SMRzXmsH/W18KaDZLimfGijQBwnGP
YQdlFtX08C7xhjE7SkOjTTLMYsAWd0cQu6QQ2vfjCti8JKthv2+vJE6aL9/WrUxq
pCaUgGAcyQ/c2Z1xqZol+N68JxwOOQ1x9hd+qF6dDq3W/P5JuSvZDWVNWB6GyIy3
sdPU6eKbPIZsOKAna0OPwASuGhiKZj0a2AJ7zp1ywy3YgW/AC0us6OQI4l7SlI9l
QpCgN8kU1N1KOKQ+NfQ+T7rk7mg9mo0w4Eh6bb6x5RgBk760EPNpQr2CF7hhFJFV
WNWsDba+eNEG3Pa4q0WXgAaP8c6qDdb4qKkhkSlWZn64FQGcuLLsfrmpHuwDVkSO
q1rLD+guJ1p/MMX5HME46brGsWFqsCIgJPPMpkpRofnWn0XSOas9qHrips/x7CCE
/k9uY6Gc4DoDZSUl9Pm2kGUQFUETXQR6DMYdbdByolsXkc+ihlfkH6OAcPmTGqsC
+fe7v8w1qeCKmhg9txfAAU86noMwFL2WF5an7y7OxKWI0v8/CSuV5mLREdl8rLto
uNZKgff8ag9L0IsQlay7ZUV0FeBP7Q6ENLq7e62+azjgLdIsldk0yBVr6cnbGMLI
WgVfo/aFfPGby3orG/yWf8rwBldZyvRUTfrrjnBjywDMzG5RnkRWHRTToKOSd8nh
zE50bj2qH/3MXk18jzeNGq4OBQWFWkc2qah8lAWWIvk+pxESVUkFYxFg6FwKJZ67
vRWri9bAnW5P6TIbX6kghTQBaZ8m1Kx/qv02XgGoUEzci9qCoD9i61uOjHWoV+FY
9WE3dgn+YO2Bt0x1gJOrhmkSrurKeDehZY4R5qm3iPw0ZoSB3qxbFrATV8zBVy40
7BUrizPcFNIRSZwkTt7JVs14WhtmpWrq+CzqabLmRpuyR00ic2/GvmwbtmUkxI+C
Yldtzvo3tjet4e3RteZHmoaD+aHqBomCuwkq5YBbBp5a6J7E5NxA5zb0bmGH50j3
r0uNtm5JAUn9OdGEfNRvW3jX8Ws8Wm7qXQwSr6aDf37qFaWZTLmawqa4C6Fwy8Sk
zO/sW9RQiBvAqX+PwG4jjoReEkyguEQ1hA2+IL7SHK8X0rBf5Gkz5ai8Y77NPYXU
9EVqnsKkwKkHP7YrUyeoBm/3jelH1j35cTP74ONp4jSuWfXsv9hdDtjZOpbzrNeY
TkCUX7Uj5WMsbFqUUGreqQxVQLYskL6hpagX5/27gjOwXVBfQX8Iy1m6/cUowfZ3
UoqpeyfOpufQLa1kZMrwCGAV0ALo9kcO+g8fWMKeUN6h8aJW1DfAt6A+NbQKGH4J
MHqXydeiGvnOuy5vHWBLLnCKXu4eCmsZ8uSjeQoC9sLpuoEbPI+CHnU1cYCu1iVl
HihEx1VgN8hynFv974vFvsGm2UZ41vfvJJAAAlfAcPm/r12DwY/YWK0wP0sCHxte
Vb9YQgpcg/COtlQjk1mGkoGAO/63guFENQ2tg6+9VGiAYweMfk3pSIRspVLRyHaP
ecOhkuZhIVatmbuhGOu0aVxmFe3dBFdq9742MKHz4el8C4FUCLvy6yT5ahpC1b3V
+TM6hiKCjMz9TzIScWs+RAJAGR6A2Gm8SYFklTX9cq4znliFMLG3utqIX34kXYdv
Ki0VrsaVG4e411E3OINylNbLxypjvj9ePKi/KBLAk7t/BC93xllMW0h9xb/BypdD
O9i2ynXQZo/rkfwwzorBUACmsxHADkxXKNSSx/KoM4rkwOb+A/6SEkGlPzDoVSpg
/ibsLszxLOOsuah+SfZHVW3lJdoZF34NXPKIaPMtnYc4lnwSTNTYHSWsNhBeb/w+
04xFbNewQh3VhntYB4QVs/EKi/cTYBz/SpTQyh5ar1KbSSb5/V+WrlvR7OsUqi5G
ESh5y7fHmEh3HAqIEZgGrDnqh6Ze1uh7D8Y1t0PGmAoN/R/ORWBrhDAxWLyGmEt3
RCAnRetemMcgP1uuqmWCuSUKQu1Fa1+zGY5SAgIsLeLf76rOVesjooK+2gi1xtin
6blKtaiJdPWPQF0xZM0GWtXzGsH+lgQrVfIRqRedlEE6g7Ev83WJqvsgn7htXFzl
fhMD6ixQlm8ZbvPup1AyUy3wq0thNx2pBrdqjMj7dmIXZF8Ir3RJc5Tnz9QG0Kst
8jKrTFdlpdhsJ09Lc86pjwvswdg2pYomCWQYUAUxhWRIkVNASGEb4serTD9cZtn1
lJ193k5rkbG9BF0W11CA5B9aw+Gs/c3XXyUArQg+PjIx1p+aB2A7sFD3wElNq+1v
nt4o1BYNIYBmwNY+aJBqzrTmW4ov5KTctMXMeII0G7E/tCvfkO7QRbjj+2SvJWi/
U5xope1MatqEzEkjjSD6t+T3pY2LhdTkq6XNz0a4y/CknsJJEnnPLFqtGruztOFh
fvQXwPu/25Fz1Pnlz7wYhv+26gVNcNjZimGYpCmtuAXLp8S9soG9PAYCRkKekqdc
Z1cjBg/m9WeGM1+KTgL8oOFq5OmeRnaqZnkVQRgt/ta6mIZ7hG4H84GzvvdnDo0G
YRhhY2vX14jTlF3BGzG5R2+TkneVjYGEV5hlqTZMadH6dOScYn7QBmikvt0RdVgy
nYtNdzaHcQYV9Q8VeCAu+cPEv534CRvZ/yJ/7HO+wm3HXPJFAL/VEMDXnVAKlFW5
XQtOtIYfgUZ3WfvSVKEyA1zkGyfpdj3bAfJNKWXYaScsQy5VqmbsJX/rVpKrJzAp
f0jSXQVHyXx7zpDNeG9HDeAwE0aT6mqlMft8LyHF0A403I/5kuejx16uVklKMy23
SMJUiBqRPHX6lZ3+DglA5AqTdiigPjiiyaN8Oh10TJLKpK69jWrcSpBKwf8kk7Ou
ilkCtOCEUj8QAEQ6sRw6XFcHnBLiLOPorYu0gbohwvEJQXvaJmU80a3NROuaoFE/
jpFXyfICOUA6zkbxkdqWyKdVgKXFgRltq9ZDcHqtldY8L6tWIfoxm3wO7jb60U/W
9oYHceAdowTtNBNPQb/+uevoR1Xykfou4uMLd9jxqpTYghJtyoofMuDad9a679wA
xpKyoIWsQ/47soYd21xaa+Tr9SjRQ2ewzyO444ZnwxVG8LuOVi7f5+2yhH9e5lFv
3kL6p0AZmGh7G9E6KW4jYkIhOZa27TbP1ySUSdD9Ej5SM5BjIQ2laCyH3rHebzW9
psbhLIuqZsxn773lyUAN2b+VVL8+JQp8DwePRWtJVMk4slR8FVqYR/Snc/Kjwgml
Wl6nRjd3bxzwSjcF1bfmQXkQYh5a8u7nGy/UQrPV3C/PnbYvUV/jAOBZlpYg0hWg
VdNusKymWrjypxglwCZ9VVMUrqJOUhPJqItcyHn1uHqeOMjt2e7nBnVSVsfr2Cx8
RQMM1KCnqGdEutyfctU3GB8LW9UdMry2HeFa/TbqogcgeY10ANpXpapKwDde9J3l
KtbpXPjyHX4YrvB3skaWKu7nUBJVWtAMLSOu/qcwQquo6kpnAE/NnYT3oAkfKF0Q
QpK0dDOuzSJDUqJ9Zig5jqXJJkEzHsmP9juf9c6VMfoy9SAe3nmkAFllqcByPkrs
3UCeMCWwaPpNBcN8ODVWziKorF1HahOdW/y6jfVBHHAxRUYdq7Ep+ALzLUY9e403
6MgVqRz50w4poVlBsASoN0Z+8j/fRF0fOeyKZdd/5E+f53v2bvE+EK2xZj978bgG
f5eVftaE5FoLOsqbEwmrfTIVkZ7YtVl0b6GQLXpZ6SM9x8bZRFJg7hllZD5ilwyX
HEO0QSa3tPeZnwHb/eITa07QjhKAKsf+kAeNOjdD8UBf/jWTCAIzgPx+JRV4vD89
7hxqcJ4GK/nNH3FVldXlFtNPrfveC/DBMSJP5mkLJz+t7OfrKjEVp2xgifLEs0zX
gd2VqdId1RpcMVzWgImcGEb/9Pz8pDmTaAbxzv7pG1uOWmaHOw0f+E59P/RwK/Mw
ifyAiJmZEQP5kr6QPzKuulXum8X3xPFutgT0JRZRPw9WgV2Awo5b6AxLs758118w
C8ygZ3FlUq4dj0j2nFfvOtNQUwo65ti6hRjaD1EO0GJRnCD0XNcalqmAbTP8xApL
aqOZbzo1FMGDSYaaYg4tljIvGciCgUKfBlK3accySpfdOvElJ27p3rpNYQz1BHmq
chAGTDE9jbjB6aDTalW/5Ko6cXpBd9h3by0QcMSDxQ7EMCNlc8pA1y6MbvKfwUTE
ip54OxvUo0D8FJndSEZ1/eNX7f4lXrHSw0iA1Mi5SGo+gk0H1hQA81bsjdOEy3u0
rqodJEjXOKGppnofBY4sZVC+pbunZeYfOV+5Q30iDF7d8BfffkulqLvxXtz282Ve
b8xQIJki5dvbGOYQCYK7/oKSt2i9YgVhtnfvXmC8QsACDAKUYxrvVPcE+oIrB6Zh
X6qTEIYQgZqQsiUq29f7GHsAiuiuXvr4gPDcKaETCYwEd2GMtf2CN+SFsVn5eJY5
lXGKs6FGDfE5KuW9IjbxMUpYuiezFisfjb25GqCMZ4YUzCk0AmPDBfOQbeS1gqjS
jc1o23JMEJxyFx50fZhRvfqST4MrId64zQOqv0NWTAJFp/xqslfEAFQ6xSYuKcRI
Yp8Xq1LqIRcd2ZImpjXnwblsBrfneRTuP7sElXSMbko1fJabPed4XYCQpfhR68E2
GrgYz74eqMLJKM8jL7qt6LhsSMvHtju3KaqxrZvF9FCcws+DMwfr9UkbktYcutYe
kTqZ+RpT5ek3LcaOyNZdpGW2FV08ND/TwrevKJg/y1crFZ87oVd5ajli3/oNt4m+
ardKWpo/hRRzV0T+p228cK71fVK5cvzh8oCwXNSPOyQp4NsCK0BV6/EeKbmwBEqd
D/gaUAF/mzFVZm9uGIutvva2LNvI/2q7poh6PBPRkL76xJzaKejxi1USHHxZcB4+
i11hFkhwQHKQu8gFo16Y7/GnHtJIVh2apZHSAH4avNIA4RzO5VW0xnEcD+7KSrfV
Xg+IjdUYjt463SmEk4ArTYdk5aW6JcrrsWQj6go9xVRNwU9giEbzT/tU8ba1XLlq
mBCUOPhHeGLINn2ihUw3CUPALdu97hqzd4oncxMIsbIkUp8UAE4hAwy+nEZvISM/
cvUF/khSQs+UTcjl6x6/Ck77jyBiFx/aZcC1vugOXuugkAy1IX+DIL9VTjpMeMI/
wm2bxzcglTJUdYTFE00QVWSRTr8WDMBba7cGpOdqoiZ0I/Xj7u2GN2of4VnaHVOf
3Em0bjcNLkBbkYXLcD1Cq3xV/fKy4NhXhrDvrt49IbzDjWBvIkCU5k5antTtcYep
BEY7+Luv4eLHTvGRvhF016Tk0zxg/nudfdBA0fNs9JButwWFkwwdJpMv+3ikxgsF
QW0lhAOVU1U+Ul8kd0FAu6jmUlfnu2edhzOZqY4+POim3FkmpGy+QaN/ALmIRU/i
lyniXu8WoAneWVQ6Zs4ScIfpL9z6KF11dGZaecBHH7d/fQBkGN245dTAH735Wpc8
8XCm3G3a+o4xAMXkCKZuTb81TQPrxLjMaNC4Dj77pvIGjmlJnscKVIw3w3pPhC23
trOi665cU3CuLnpFf207TsAlSwipTGzDKJthUBUt55TOti3bXRErYsWtlXqxitHX
tJsPBky6EmTeYRr1zMOvGfIy4C4PPZNRhanWAW5RYNWWkzy69LKQ8lJa4rt91eh5
cWCHE3BDJMH8MjGg4lH5QKZYMts8/eURtBWzW0kLOlyjWNk3+c2kWZ6LZwzwdAws
VVsjGTkniwWzu8na205jAJYgOr+YWq2uTiZnK3gmhOHJT06seIgHGg+KqUf0Kr6h
qCN0vKBv8Z7W1aP/1aTEzScLOkQWvzLkzG/vF05WxIKGkm3flcgz6Wif17HjI1vw
rXAQvyTfyVMhfsArUTifHGtbAT9S+t24rZ2kfYvAeov7uD+BB81qc5jqEYSDyk3r
SQgdht1GqOU75sqo0zRDPBu2cjHd7zLGEEDtD/tHBVlzaBh0mqjCEApfF0eWBByo
9wnu3U0DTMECWze0hR0kzPokAyEQuis4CevSMUuTjTxcvy3isrYer8VzixxC9Syd
EF6c9nAWNjmX9oynJVvC37nyqZPbNWYvYMdk3IfBVzdt6aF5nNVjJ65TGM61HdD3
Pzw3oNeyJNGVJkAfwMXfD5dpGWvtCvh8ECK4gIvmeFADmtzlT1mSYSN1nSbJTmxR
vEEVTaxn2p5lo8NEIYyv3QtIBZutCpxeHrRoRTOI/IywytSyWnuLlBwzkg11Ne/K
eNI5VvTzH2OUEPGGNJ2s6epyZ2IQ96yKmvn7ixIcgnHkDOlH87Yi8CWebnlZkeOB
lNuplyXr05KQmVm5U64I78bCeb7N+xhlwgIfqv+yg64cELGmOMi3vg5Upau29qQd
wLQrmf87Lye60DiPqNdlNzcOsh+QDqIMfNrsH8JiOOFZa8o8PKJMiTWjAh39NG6R
cwibXdHNslnBASEFr7IH77Otld9BodYIuAfL571af8Blsfod0878NL/cGblH6KwP
MZGTj2Pa8ET4ebr06e/s5q1IFuRvQYddrcWHDuHAjJV6ZuTRv2dxIJns27GuiOZQ
BxhIxFapfTyWQWbiUUVAxAbRgFVz8XR3WGezd49H/XcMo/yto/xQ9wWkBySiUkwa
Y3b885g+pZF+S9bxOWw9zUykfKzktmhHdKm58E0sBVgX/VEVUGhRznmPlnvYAPW6
09nrrfoWKLDc+pibxvLgBWS5/VxdOI0V405/hJqnE6P5RTx8wzsf8jgdFMUL8IiE
XN6qZfb3g35UvNbc5UDsAlQeq7GQEo723GkhCUQ/PJqXPSULAr+v3+Zl3rNouW+p
NTUXvehPjJ6iwumfiiDQGfwCY43L0lnPfBVZojryIlafK9kreLakl4MQw9TbIA/K
9MyQncR+cVFM1p56W1wCfSCUoGkohPkDbv3xOtJzqTph9iGzPZaeGtCXimpbngk1
uuyfz6LuQR6Q/lI1xrsv1k9sJo7o2XtDCmNOeNy9z6oL+cNvIfyMBZ8Hga5dDZ1a
LytnADLniWKjfCjijQGS9CdpPTl6DxXkqz+DTAkaLVQHDT0OeZ7HYuC9Ukex+x3F
AbSZbP4BvRutszf67ELCYI1VZ7wN+9yRdlUPg8gxEZdayXxc6RqBPdj9D7OA5ccX
khBY1IeQlpODwfXCmorRyM/k+NPbfCgZrPX5UwbAoA7F4rL6fEj68U1apjLLwZnH
Z1kC4DQ0X/zcjV9Jvb2UVHof1Yg9xxcXOfCcxU1bYoV039EmjohlIQsYgVzwo/0I
fy/kqsutxftjVun8+VhrgI875vazBPX+xVKZ5K3w0d5cVtafFa/+hJUt5iD6r9g7
HtThSVm6TMVltzLcKWVOeA2SyLGHMe9mBmHTL2zD8bF066oUtMzmvcYWKUJjXX2p
PPN7q1mtQyeQctGDePT6oIQjqm/Iq3sKNDOEDDj8xYyU/WPnwYvMPOo+6PvDkQtX
2UlO6liJr55bqtbHke7lEGXSGIm4DXymK1Fzqq8CalJTfn0IpuUFtP2WHvRT10vX
7z1eXReLVb2j7cQP3y035zWKpvQNJmY1/JxoMylY8e8WNnvJVJQ2bv/7m/b8Qfe0
fBW+7286LeoKS6AKb4dnSRjfRKgJ8DwOqOAjFDIn656oW5LtKXoLNXDtUAlMb3XA
Mo0PAah23Jz0pTnRv8x7GtrwuWQmOh49KK8c0Rc/Z5d5ZKvV+HYiaMbX8lyvskVu
g0dkwF9KFm4SSfApy2vbOB+8ZmybCNJJrixg+tJ1mXf2+FPYfIm+mOB5yQijuoHM
9yWbJ/cHLNfru3joakT3vDqEJDlozSZW1Zqd8yvPjsX+Boi5omwVtOuQFRuVeVsU
2nhB2lU2ls0o57Zma+s/aGCZbiVzuNUrp1ztL2R8DuudSD2nZgEH7AmYWSgN2JvU
sQTHapq1BBinA5bvzt1dHB26q8LGMFlq30wHzOkLi3mkjSy5DuCG/ZRd6MykV56b
odBe5FFCxI6Vl0S321MeeyZpuA6iEX1WNNs2IhZGV3qO+zznCygpLzOEBYd/+ySN
2oNOa941fWKCRymjTFi/wO3KzIja45ACeUrlauLuYLWcUMO/oK5bi/FJwnLxlfLo
nSgJCWt5sjfQENI5/32wT90Qbbj+vNgD4Yx+gsQV9EpmAjmL3n5RaSVJ6ZDzcZac
1Uc/mZsnEeMIboTYNqAjKs+9QPrRm5Hvz6o19wGrv+T5jB0cilgOPbjc+4QAPDZH
58vDSWcnscMcLRSTFNmjfMWruL/oR3iTLnNBRw7XQFNZg1OOQsYKsDOjbj/FptEl
eFiC2pn2IGJXlnXE9sCo00Rs5BKWxi0vQWS3rMVsC1nPqt2nwZKY8+BdvsP7RehT
yBOt/qRyeJOlQL1BpVlM5xQu+1AiT5p2ZVcMzCXgfB6CMCzwyAH087dAcAu020Ox
bKQJGfyHq0E5bklyzCeECuvoYSDODQWWPhFZTKJqfKYUFiRpcv1Q29QtMv8GTjlO
Bt/UPomX4snGckApRD6pDn+Tt3y1q48vdjeyQChrbHerQf1JIPXIFntXqlWSxsdJ
C9RAr19tctBdY+Ns1jssKtZRkrH/+bpvuDQXm2lRzTb/tA1cEMH2Byux6YrztLqB
Ce5n2G2l458QmF6fgZI2tUehB/3Vmwtzopn6UjmZyj2zqWQXqHj675hTk9AjeWQZ
4sW1lgIi9V7Mh+ppJE/o8cWDoN0SpcislSjDmc1sBl5xbkrdeyFR3mgyvzUMdclT
IkxXY4fwCteuAAykWiZLfr9oo6w84W2S5RiHWNy+kpGy2Emodv96yzzSlQvTl3BH
YLzOhd6ZudfPF33xzMl3bSUOjFGHgPRPCjF2x7/mAty70T7VI7LNaH5QEjvIbQaB
WLCaLFA908S3OKgxaHiuvOb2INhA6xxVO/AE/sTa/xTt/8/gtKKkoJcgwxg6lcpN
/+kilw0m6jiSdicxLvTcWTuwph+bZX55/UIZXeggv2wh6o+SVwyJZdZvOPMxt0MA
oWh3DTPPNoGEQwGKX3ensycQUK9jZFXwletC0T/nR1P9pG6Tc8xgnlPbi/EyRzqq
43MS2faWc4mB+d6ORAkxUAJvPGjjzjhZKO8nnDCOp4vlfHVcuiRXftTR1F8yDCrW
O/Lvqwa2i7Xa5OBpJ6nGSO+JVWGV2+Sa0Mnmp0z6iFvN7RVuyPy7877U8r6y6REj
H8ElELdTz2WKjou0WAp95p7gxfEncRXPQuyuY0btvOvLhupf81dk1A3Ok204JIda
eOaOlDqHz1gL7tJ3ynwhy2g//2YYwIBEyfrKayTa+e3tStIvkxYiZmeceuJByYQJ
vu7mp69SrGOlfUcsCfbofINBI7hecxvQ7hD74LZ6GpBh/hxr3FsIoPxXKZ0Smfn2
Y+RQJSKtnyBrSMOaQ6wvKLNVuuoDB5ZeCtEYowd8AIQyL1auaVYHfLt0R2/z9Knh
w7MwhtcZfhXo+LHezjHFWQNLymw34GVlnkDAsEGBCz7S4qmaVUJoznSbmZnMqhH6
pLhSp0MW4Sc7fHxkJuYsaiWvuKgV8/bMPj8gG1SlhgeczdGFKwClt+yg0789wcNO
fu90OC0DGVRrjBlKX7QEvKL8jQG1QYaBgVraSyrlR4fwPkqkrMziAcjyyZ56svC3
jFhHNjDJyWW37HmeMchyUhEexn2BWC+9SksUAaNtoVrSfbRTgG5oHeIROgSeAR2b
2y9cGLwwAjT+yLghSe5QEl2w8f61J6a/6zLMce5w1R+VjKNNOPzcqd+BfGqk+hR9
pluj9dZ2FRMjGFVPO1MnalOgq7nOvT13vz/SMh2RZzxwySiZkyCWmdLxySRXO56z
WkAguETYy6ZowywMhqcbTxRCyisXAfeTDN6kN1GbwC2rIwmQbEfbpKfJmO9IrTQg
/3uJVGtOmthEqzY+MBUBE0EkprD5o7i5vN4YiyrYnKVsZ2kc/CluAWhh0jRNO/Nv
9B/Sv3nuu44FKlwwIKE52aB8O7C4hc8vQslZpkw+15VxfpciXqyCHo/0rX8HAJHI
7Ra3ukwBya9v0XN6mv0QrTC0kLBDGzhPU0UefLjfDVF4XMP0zA0zapoZXbR4DIFf
K04JtK5mhHYbFEpvZAZbY8J26LW3+lWXOWT+jMKWs0RKOuhDyPZB5qWcaXcFoQk3
+8lb5doDia/2/aEbshipZio1N2VdHpKiJuHCAnCthOd4IVBeCUD+QfjPFtWpJKtG
epedZoi1F7GzTAC0zXa/VgOH+YdVnUyB/Hu9PbmDZyb+B4dAKVhqoJAJf/lUuto0
l8KLcmq2ofy8AO0lqxdhpT4yLfvRqgbZ9fnyIO659owufyZmgXnF26t2DSab9Wbf
F7BbgSUcl8k12UihSicWwrfxv153fqVh42eU5mVb+12eTIMFuZgwv12PbPy6LplP
mLPDMGHFx0COidr+fBC4Fs72ZYzUId0sTOaMxxBkA/Dlb/O2BeosLjLZeYhNWzxq
awnWK9AKdwY0wL7Qirf/IqDF52lF3zcLqj5sAEcLBvQz2ymS3pp3dbtGUx616yMZ
5YPGU6p4mCoWY5ecbb1MwuE4pfT+ManBIFb9kQnqcx/SgMs9knax+dgiJGpH3jm5
pzF6xhNYFXLcD0qpZwNdKjGT5tiGAo/OwzAj9Ir+EFDLL87g9hTQgS0XSbnFExEo
1qtG/d9AvX77Lc5/u+k65+ULKI/GHQmf/OPQ6xjTjecZOa4aiGtA4xis8oZjLwAD
BPyDfQFsmLABdm6ADes01cWZJKflqA8ug+oJsv89FQfkjDnDqf8gKigqsn8pxggr
rldRzuUhmkm9gpNjNHieIISsYZdR4j1K4z2zob/CYNjhJfDIw/izR5Ob2l34u+vc
Xzz4k5+TKzVhD8oZR9rSpw94LpyX05C4h8H6FGmG+FQLvres0KSOkrrqMNhRKHRX
GvOTfoABF4Yvd4t+HqKVRRtrchf0qw5gQTGhSHjgJyxoaOJRGZ8mfxCB782tsSSe
IjTxD3a+JW7ZO6QOIXEigFYSaOboRL6NPZLfG055ZbKrYcTApPHJS0g2WPOCtusj
wDETehHCfJylxjPucq1Trd/5UwXT/Y4OZ1VP8HuaI50qlUtfKAfrVocJ7i4w6+uW
L8L9AeiTzMw9/ruHcuAdoodH3Y5cJAiBEwU1kOs+lZM320QSPf8/qhlwe5/770ne
b+QicVjlyw0featuT41rN63oXSKnNDEySRrkYkj54Y9zH/mO/Y7rOD56ePTV+zNC
mHd3n835Eu7mmjVY5HNNXLIMFvnzwShhVOV0bSbM3V8o+Ro9Lt12Vv0Mvka/EpQn
qih0DJR6FlGpx50fxtbffChvugRmYZUoXndgrvfAXv8j4i44oX2KO4Yg3A2xjaCy
FPoDsL8oPOIF+2t0K7iFRqDQ7boiCbilT+EeSFFTiTTZeglU+zy/j2DnIke7f1BD
rIkjzy2dCEWNjlzMhE5oU/gWFsSfQFlAV4j6gZru9QhIDpxiOpQfltxtXmxYLjxh
KtHpJTG/5vg9ECtu9EH2sr41g6pF9Dl9OaMDvGGpwly/j4tcmp0/BiDGbyrbpwba
CtaKz2gdhGsO7Kc9OPsjF2JJMEgqcE06PNJozymInq67jsfsvtrnuBu/KVy/w9Nk
jTJ4REOY9fbV1oxfRfg0r3uvqcu+fHFhIq4SrNfKEjRSFOU1GVvApM/Zom35/NfC
OZv9sxfmbDzRVWtFCtOcA7c/RpVQUTm7k3+Oz6c+ONgWiqkEWf0r+AAiLg4jTp9e
17vFk5H9JGW08p6Rq2OFZ7ApeRkG2+0QTP7nCYk4a0wRflubmU/6txVMkQ4KXjrj
/poTUiUaozVv+hocM660C9CPMP7GwZOgXqfMEWvSiqbX6uGKh8zlfO4ojCFkL2K9
xni6ZsbMmwmzhxB5IF6Slj5f8/tzS4n35qKBmocG7KmyF7verDN0KJ2JVZ8MVWrB
XA04bB1rOlJEC2i73kDfRdVw3M51VmOC1QFuMVxpYAwRwQsmvV+YfcSHsy8dQTd1
qVeTYwedmU7GLukTVPFwZ4eDvl13dJQuV3lUKf94z6X6afWhT3wGLoCWCHBBSZgj
zNPNjG5YvEN1SgjyGq+t9Ygk37xoWPb2PjQ1baL3wSTcu6Ws96PlanJxgMHzH+Li
H6MIJ4t+1dVs4Db1gLnqoX/AtFpLeCkCd7sQAvwSuWXkMLovsaJ5jyJnAPUnnb7p
Oov8GGZccR9d8Av+bTgeg6fanCHB8aEObzwYdfkZquImrSW1ywLuQYXyqJw9uHhs
J8xqy9LS/+OOuGehuaY8IkY1354RCBIPHG2OB7I/cvEaxgwZfYj4UuJdqnlkcAFn
7NHld7bmmvBLdYu43XfJyodz9690HPw8g8f3F/eE4CywNCD3ChmTC79/SVksglfl
oQ2yFmT01y9XP1UPZsct0AVZT7ly3dwVy1x7xTFv2nZYG+z4ruZMl1hOzEUvZvMZ
T/jt192d2oyYzNDx++2F1nmn1lV+acIFzGq5kLj87OLHp8CWNWRpNOVVAtoB+mlz
koVO0ppk64UT8VfBjIpk2JT9J9WaHRyUGDowJIJU4szisrPTyv3rpUSBCBfLe5yK
GtIO7yRv76qz3ypfl81CuKEp2BSbfvK2edfWdhaXsCkf3gwSFLoHAAV+eS/Kbf9G
Eu0+aNZoA5fvpZZ+iMUVmVCKFEBj71i+PwRkUzm78/FvI1jKiLu0L6j49t6Op0hJ
C4cBkoyC+ZTMsuwZYiMH8s+fVmlHtXnrpZV6TqeuPLFWIh+uDO7TjkFaU3KSmjCn
BRF2dMg5VL/0CR7VxLMRGDyZbzENEOW4FSWenCyRx5YI6LutKznuqCZjhCjPJC3O
WBleS8oPVsGHUSOSgXhQciAMezM6z5r4zqo32J+zIL2zmOThAyilDS8CKaGjD7L7
SOIey+iERsG1XceDh80c47B7R0Lx8oX6kV8DZVRONnnDgVtLBTVegi9WTPjRpIKT
WMVOc+9Fa/sCyqPzDPBiIrp3M3fluFjQiZCHp0s7gadOb3wcjC4VPXDfdgvKC7NH
l77wLAfpdq59zFli2jjCdf8ogpQna5OxzOUqvs9wSmtQuxnaJdfBTK1FTKw3CuXB
V34FlfLGIgsVBq0zNNExdHKP8S1C2SoguuccPWRhTIETs4Ycmrq9NGmTFbvjppG4
JviIH9l2wWoh/FoF1Mci24YQJgNx7fkPaiJAo8y+Cc3XaB74DRSko55y3G+as1RX
goQk5NYBHRgoqrN5UhrUEZL3zHu8JHUUYYDw+J/T4JStrdbbR2r4zkvykEAuvvcK
kQ59WKOmQhaG6i8gM1ztfiouc49VlZ9ErzlVLaC0JPit7QzFvnpJ7+0KlqiiqGgh
5hAY8W1yWghII9ckw7XdlmSDehf2JARJSAb0Ybi9/47a0jV6Nszp0ZhTl+pDJhTt
bAkA2zX3sjDcSgIXcvgeBZIHFtM2HRC3S6t7I13nHWA6UTX42M80KjM2TFXd5BPq
mUTK50V8PS3n36Ls1h/mVD2adPtlL/RFwAjkM+iAFVF2MOjW3nlwpduMl1c463Lf
7pEHmVW8+9CghhiZtsbEl9jC1qHvBkvLemkIBDHIIyNTutmAgA3fkosl0Bv8uBDx
ugPwTHPNa13ZFzRUUnktvNqWscBuPI/l776VnPZTxxBWYQXJARUEdSMrEsAl3G7e
e+ipi4RF8sQM3ob2QtW+4hCibCcs8ZeD4CCYib46x08X4Lr6YuiMzXm1p9e9py3p
QIS0E5YXxzhF3S/K7YHJ/0VpIymQJuanFnmNZrmff16GSFCrN6MHdvZNNb4QTlh4
kLjO6A/q6xltZ9Ma4ui0WE59f0bY0wo0jVgHGIICDcgZm/akCgIjuh0tyLqaeCeu
VkKCVsadGMbTZE+ruhJtJAXhGZ4Ph5K1IlxICsEELSZWmiy6I7I3UL0v5ZwbMTdo
EHOlT7xu+wBDoQy373ZyyQfTIMpI2JOwLFchq3g88fH5HZKQy/Ti6vTAX02gUt0w
YvRLzXBNNOyI7TH4zBqQ1nMdvcYYtTO+OwG5eZSNNtEHkmbIFbu1y1DPVXruPlno
IaoHLfGJl1fwqkdXZUjim7j0pxI2miXLCEl/jfzMN9UHNp/pwo8emImsVPox0WKz
VEIjEQaoqYt0SjKkNf0jDww52MLijUVE3F0eoOW8MuC4SgoH/gXi2osAV7vMLemO
NBAV1g5/0g1LIxfSjkeDDZFE2gKs/TZ6Ip4NBNDaiI4SUX1ONs0P5AM9+1FwLNrl
Re+lXVm00SXUxWUz3kD3YTPQ0A7I/Fe0n6mvYFwnArsBdAUTeMvnaMfvqLKagR5q
icExM4zWDHap9hSM0cObLt66ANmPZFEIQJYD9/SqTwUsr8iqdSqyaSgN8FgyUy/p
92hQgQZW4rYLjscK6p9c1x/iAWG6PdGtp20y6FafVl1u5Rn8KRcjrfGKZUlmFBxC
I2yA2fGoFAd3uXSpokFio1UjSsQtLe/1gHLuvLH9P9aKoPEV+l6+6xob9Sbq5TR8
8+hFVYPZ8Hp85VEtGldVKG4FcQP+uQB5yRahE0co2tkXPZIjBoxXAWKJAvpg6JLe
rik7Q61MMhJ9Tzg/tPunwFqQA4d6EGNzuttraa348vJxSvh3jEKUoG5v4E1xUJd1
hTCY98vdoO6DAxkFxT5e65WfX+KGMHBE20awN/j1JSqX28eT11jsGCYRzAdLJIQD
FeQqtz11Xl1XWcDipt/BpCygfSj+lnEi+N/qqZQ77kDL6rfZQk0ht9dz+BO96qLX
801c50LBMjotFnfPBIFW7N0+c6I6XYT/ThCkDRuJZyufBF5D6zZydiAwzjmFG5v7
8+uSOd7V5u4kXTIfxgOAWqRi1lvjnE9kQZZ++6iHUjMxMciTaTT98bhOI6mMRVuQ
RkMOa8m0GFzUNFcB1Xy1rpEC7GJt6zOYD1ume3zI3J9PcqmMc+iH3Q28nZTiZH/Z
JmV5LL6u1Om0yP4xt5GNzMqIcdPIsgjfLq9jcTRBxNjibd3emED+ElJsoQWugsds
PGvYYYI0ZT58ExF9iZlKJIJjIAFUGB3TNo+sF4ZxAsMCURmdCzMoXS7gzrMCkfxQ
CDnicqQt4Lm1HmsozKWwH/PcASmFo+1eABvVs2YWayMTRVN7fOGWVkkdOzc68ZV9
c1vQGfXI1/w3ID7gGB97bAbpQT6NvZvUVBudktaes7LalNkThIrYmOyBIJHq79nX
jzM9S9xrFH1aqn1sP6aQHPbcBiZN8vcSODviEeM4tOGSs6r00R3Zh1j/umiMWjDN
bo4itAhAG42FLi9Epg721VGasAotu7pbt1DpkUxU/slSWaNdfzZYnpBpe7D5YxJi
bAub2oJ7NMBazt5fX0K3t4N7lTsucqMxnkp2Z/94ckor72MEaUzMdm+W/mpXUeC3
ELz+2t5PpySXB/PSvy8jOgfTk96wKg7V8k5pdHP8MshUKyFthht/ZGaWUFq/mBgd
TtSxuAI4jT84a91f0LzXUW2hxQgcjprtk7GBAynouviswQLFNGBqOi42xJ8tycBe
lwnr+fa6LOamKf3XBby32ec2Y5rzrX/qVLj7LEoOjPWoK7z8DuCFwJlglaUVhYT6
hOdkFKjEiok/nyWsuDG/Da3JFMclxenXrUBy2G5s5b+fMrBnNYkm7NdNtmMzwX7q
czrrkL6Yshz1/rVUUJpmVQ4mXdnuXqa+gJLnNH7Uuwm0m9F6t3QuzK9m7GFL0tqP
1xygXX0oLBWAM52ozuTw/0b8FGWmtIrIEpw4qM9P3RLCxeRHQKBjTaEkEByUt3ih
7HDLkzjh167ezpSmw8iN6tOJTUjNbCtmE7gwpegdiQD3UODhdCKZmi6CFy5kmu86
Imu3thHQCm8KqyNPU4h/iLeWkwNwwwLE3MsFJs5By51tT/AyWnhKhvhH9OhcUrVV
aYt/LTwFWG7zmtbtYHmOtx2V7ahYgrFWGxy/6JDIgtU8C7SKuk/G06yPaDo83Qak
wiltG8PqSWZXFIXVb5JD96f95jh3Za1dWqZX9VqBXiBnl5v5OtvyF9RitazH8P7X
QL4AdRUJ333jJNZUNtOgxWJR6kwHWni/3Y99aiQeGPWogTRdoD80jeUvjSj8rq16
AfOJWLkq62k0QmUpoQZUdakjHGzWVVYSS5RyU23Ux3RJg2OOHs4TW9S2tsjTgzPm
eDS/Pzr4Kbqi4Dnc5fbNoTX6asENyGRE+JwnTVL8lpCkMt84Y1vy8TVGz3EtRfLe
srY13WUs7cuApDtYRSlAtPgEmcERTP9LKLR/HtujNwaNiA68I4DrJoUYlPJyQwoS
iOxuz5nMHA/F1zySfKP5oZ6Enq95g1iNET1LrPqyJuF6IsywectWi8LzJT6pwkm5
aCZHOVg19AbNJt5a51tzw+YgIFaZgqmSURpVWij1cckzKwU4sjtv4TaLyPjPcfAt
ECiuacsr4zLS9qEETonCNZiYphlTJGW97X8P/LZs/EGbTiSQYG055cmHM1WS27ve
QfTzs+7q4S/zRWYX8SAdTjVFjrIvFoE6AhQbZelq4Mx0G9nrP/FalOr9dyI/7mQy
1y26Mfrwd9kaSV4vdg+9JkBQb6q75/erCPW9zwxXIhi/bWY4h7if/Gvh2ku9jTyK
NJprLZG9Db0RAbyW07GcDLPImmU0AeWGRyRC6cCK48QndJJJU/ifmdu4WnzsipxR
hSQpQzkAMuP12ba4Jkv2Jsbe9KLe+sjbxCEQZ5T4WRfYPEXkZYbt5VRX4RBvflhF
HmmqhwhQAZRq/t0QUrvjWgYx/G+9hb6pMrhMCvgStY4WrdUAwJ7Upk6FgGlwoepy
Qicvvd+oWEdZxYVOSkUUl3+yIRirS6nyghtD8Hm5bZnFFh+UqGVaYixEqIJ67v5H
NoWwy3gAQ+daT/94gP1wk6F9c5EMkNq0XI1Ge+Jf50UBvpjF2bcX2i97iIB1EJ8j
Y4+nR0KAqCHqrnmyzGn9g9KoyKMcJ+3qwvluc6CC5tQ1q8Y4lmYVx0Qk2huenoh6
S8L4EEI84F9or+rUNoMHCVcapWfurFyWqkcQtVkzCnWXhicqiMPKIjcZoB8S19wa
9E8RFtyi2NDGpC9mIV9Rk2yam+RkB0Ekrg2G4I2D1xEdmK1OtTcXvVU8xeqxmV3r
ZAhctktBMY5Yxw25zSGC0EbxIdAGp8lWX/CGlmasnNkDF7eiGQK5Vxlp0PVzwhgW
SngeDITcUrBKp7yZKFoasBtEh7zquL2ZhooirNuVLxyeHvc8jBNwZk5+IpLc1IS3
c9ZrWYPTwVd5wHpSpvmGpC6PqQtKpNX4ickv4KlzwqMNIOY1tcfOuv75baRrYODg
V/8rpjff6b3gK5GnAOegJ3NAgRZHkI3n5bSLpoGp7WTudtMYs8NcRKO4/neHijMj
R1T6rol+5Q4UuyrdE8CJ7pasxn26TOCOz4sQ4vvqNx2LNIuYqQlb7oTwYLZ9Nbbv
aIds21JXsfhMJixgpfGAVIwt6Ch4NWK9xWh00RDNR38TyS+AuMzm2kZcW+uEB1Dd
tJeyxG35enrwLGfFk5Fm9D+7/TlqmmuDwQnNBcAczLH/odKlYmuDZ5scqpzJAzik
qgpgQXfObl8f46ttwP+ri7tUbNNmGpCSknEblkmkhlt+/qkVDRgz1XurcYinxQBp
y4DMMc/Lgnxd2i7Umj6PcKtuyTRsAfODg//Ob6kBoxwUa0uQlqrIM5GW8ZRUP5+i
tziRcEluRKrQ9WudE5Azv6Ybl/zYatkbN3WZvkrFNU8NRNTc7RXXm9NOvC73kr0X
pEWMsFDdTPMT+QCEaCMOXDtY745y/rFmXdDmlLRKEQAA41IvzTT0BT22a9AG0vaT
Zzxc4UjHK9xXrVBhSu1fiYHJ9AhHx3Mo23J+fbPzsqaR7N/yqF94ku5hm22YGEfh
fL1C5snI3IeTo4d2UW7SVoBzsJBu6Biix+fnkmTFq7xIz4hGw9wuXO2aJRUg4XVI
CeYcQx55nMymxbXWsPsn1hg65aQj5ewTYef1k2bZJqXBUDV4S6I9Hng7V4kHEu8s
lTB7P99DebBqgQND2tjmhFP6vSTInBA/BQ6uALZyosaqGv459GO0ZwrS+34D5e4a
LAk56uGQ0cTcLxdZHmr+EQy35jVRP1OuTNModrjd33q1UGJlcLnR0c2AbfqDcQEf
1N6ztKg3vehVDJcwyk3j4LzmI+8G/PhEvedI3zspjNG5EU2qZAK7CNE6PpKdIzK/
cI3tlFky3CPsfueNBJp3ELmDna9L3pVJDIOPfPyV2PfX/HTodowdm0ElSS/axTJX
yNL8eDePfqb6e4GiG0TsSeDNNQmFICAfQkabzErG7ru4ibECa60cNuvsKAjP3/aU
l9vC/L/t5L2/7Bv+cPxXCsXAScqsHbrg/v0luVtMqnlykWKqpXRgJg2G0MACsF06
6Rc9gPN6/wJTL/LLmltqXWfCvToQ4f24/Noqw7nt3PBB8tFlzyAIcp2poKuX2vNa
Vk3375ukhF5zjajFak+3nKeF33mW7vxZntH3b3YSrPdeGc1Ml8gUqZ0MuTZw8Qv+
q2Pgoe0jNQvwUITHlR1YmpkCL6HI2g0lKz+dnI9L2vQT74jgetue1nTirQi5yYcn
8UewrhCzQOcH09ISCBue6XtTl25pNRfLANQXrLREy8X2sUa6nbVFIpcq+sIGcA7G
isBsYSUBmYjYCvzY/JoTHYWuB5ImWYXhvybkARtE3AeGT2GbgMl5iQiFhKYvaVqO
Aip+U0+/5TANT+d+mi/4H59Or4aSVyp8R1VmwX8x+lb+vmeIVAIgSAr1O7kjjE30
WQ6mO2xS7aDOTVgAiUkTJVF5YxBvJmN0oebJh44ngQ7b6exrfDFLLgZKiqT646fz
rBBJyGBlSBqlc2jSqaJggnzzY66kLis9McDrkOg1wauySd9prPUJNErI2i1/woXZ
l3euSmXj9lRAZLqszlh/8uFkfqTyQRfH0m0U/z/BTGer0qx311t1pn4zV98em9vj
jkIWdA3md+l3THWCI14AZ+SkjKPA21cKELFvB8TcPe/1cK4qsbqTNRFsf4tHwQZh
HBMNipwWitXEj2y0zOq46BLvH5em4cYTIcG8Bfsgt17swD0dc9OFRk6033pgYTJn
3SQgTb8uNbU3aQxidyOjJYnxkHva+nDnTnkU5riObiXgSZ1VP4dXXOd6BZsgbPWa
fO2ReGlm8H0S9WPspZjtkLVZSB2kTpkurrGhXrVXeTVOxS+Y3M3jQQWE7OHGl1f5
bCwUuCSvpzpqKiCo2WgxtBFjkLkuOCs5YyJJnY3sdGL/I4ceGy08D5fEun83qLVu
wmop/nX4pnvmfYwUFi8PVAo9ddv7wJHcndKw1+R2ZrfQs28uDhKqId6sy/EoXqEy
nUW7mlX9eGqsqyaI/w6pQ4/tFnTySB8b1uL0gCoWsiOfUH3JOGpITm1FTYy32IeO
rAkE/oUYBYK4CAeoq/ubF3twJxJG7O5XfvBxGe+HItRTorxdSTam3FHPTjK8fCk1
lcGttbw090tdPMAtYFDNVkgkWcWI1G7Em0pZo2ky13NqKEGricq7zI9yKzE4177C
ScBnuAoKd4HSvzf7UWWTxQeZfeZNFvN7VObZ34DL63WcF9/sr9U53ZDCKP9TcBEH
+CN3ybameblWByl5YWsfmvnkPBkNfbWILRp3JfG2NDnt5iAhxjpxmNryM34QhP1B
nYUjTJr9s1U7w3tbu1cG9FTPbXxl2F6IdJut6OtQC5r8xBvw0QW3H+aTztJYTlIy
MqcJSrwHZ8+Pcd9JjrjSBac42n0a/9br6rSDqUqHW0xbCf0rGVF6toA7UhDUh/Oo
F0mJ5H9YfM6TweZVqhfBI11maNMSrF54Zk8RRr5Qcby19mpMUlU47GMYcfMFN/a1
awb2h79rjS2Nx2SvypBe6S+ffTQQbXws5c+QoPV2ReydsZy8LR0jL2NpSm11Nn39
gYAx2pP1w0GW1jL5ayNZe8uAp9yE2558zirOI/p767gk5om8TWSyaFoWi34nJpwm
Ivc4lIam+bYTakO6a2uwlh0MviXha29UahftuRPR7Uvx9uGIh5KgdaNC9GqTAUuw
9cjsTpSjSMIUKC4ZE3dv+G0scpDeIPr0x0PA1wzJGvSFrga3iwOVP2wFaGO3mTuS
pO2M+TQIkgxUPOdh/5KvJ+P9U1o3pcCW8FC8enAfqmNR5iBXwh77sCvCNSJDxOjt
b/0Px3yYzvlBdu6nDrEXQwdywLs907bpHhzEY62a2oxWYo+pnmdJCXCjUnKFt1up
KKTL6C3Lmvw8u1V22LlpnxgqWSnd53iWusS6i6j5vnmz8bO4TtZ39KEi2EvITIVU
qoi7sUJBLy0+OtfRyLEJPLIi+RGf3jSSJnFllVZDrIOTPhxqRYWJTPA5uhS6R/jX
1uinuY9ssryU/8gVAl57KHPV8BhU1VmR1szr4jOshyxacEk6wsRIY8WK274zApVb
E2xT/2yrwOpH74oGxwFrRJ8UctUy8YKK2dgRxleTfX4d0pnxKps/4ApAqNkTIlo/
40wORC+gBIrcgYvz2crjJVM8XV4MTCHhv4XVv3w+HoVkZVtOpdNJ2nv66aD7kWIl
UnlNpn47vwLyhfIwNeUYR1XSa7c34qQE6sE0OMmUTJMJDXqBjv21FRxv7ZJ33M50
MJboF/TYKeYLg/KIa6jX2t5IdVfRperlUBjc9cNuv3DGrXh7VKV8p0I+sjP1gjyu
QMQrmMcojuj0j5ZZzoKbKHM94GC/NYQrbp8sMOsKWs+Cf2dz/YlhOz7SgxtlyJvv
AQZvw702tPJ07YRFKdaCwjIbG2KjuR+txfy1RvN/t/tp4qdIel/AJrKYh4htc96N
V1C9/HggIwpFuIfh8LQLj4QdAUQRjWin3UYBWh1tWS5/WiY6+/l0mwBIleqtB9TN
+uZ9r5AV4rZqAIoYj6q2OyGf2qpFyD9ffe2pxoUmzA3d1uJgSKtop8D2ETbe+f2c
IHUWHsCZAXeMSNcatFwqENJNpK31KRgfJhKcQERuYBCWO+BemPLTZiXgI3XxM/Rh
hs3b9ELD1LKK7pg/rwFgabgom11AMX6BT3L6zkeIKzZ++F4x3vqOoOdf4anYP8hQ
RjWEVarwcR6zyKFkSEKPT+pyo1npOicpKCu7Ynmz9thpMOILuNaLjFXqE1Ay8AYm
58t+qPngmp92xJ4eJ+QXuE3IXTSJc4TesGvJnwugVZz6LH829Xh586Ks4oUTqr/t
g5VhigwMgJDICaBut9vQ1cLkwFQWr6EswER4SQJCPNsdepQDQM/tlXtg6Wk4kMfF
Spk0SEnBhVvBjFgpQaFzBaZATkjitLRt85DUp7b3pWr5yAYWpGpzN1ST0OmZIrGN
6unO5xr9YJWunMAwpy64ddXafy36FhPNytHnbfZuI/uRZX2tv+7/2QZ1DQeRi9mv
UfF15sujcQPwduGmnsHTI4xDHrDXCw7F4vakd63pxCX8Zy1UNy7ojoJbt2s453V9
wqKMx6/YNOYlnfnkz4vYU1jIPaWdJ03eeBzTQeQ43PnDEC0SkUfSWrQdWfFCbNP8
abw0GpDRe0zCDSdIYwjYUxG2Uyd5+HRSFzNS0j7XaxloQ+Eu1AMIy8H4dXI7Z3sa
HXiut2JxjyhWOtfzfH7c9hfty6bgrrm/C1Wgsqzyob+z8thNlH0QEy8f2mH3i8Pg
wfzIKSdMAB+m/nZLHpG5HPlLR1HNWsNPTTwzgByhfVjhF+ETCbd+yMAEOni+b0Is
I6IN6IxBcuPTZ0C1f4sjQuaJ3GvqWmsvGDDEEiEiJbldKygyUJHNSg0uuXl8wRir
PDShmBHwxT2SfAZ+jtVhD+XkTh9LuLsCAioVvxdgw3tL/w+aUHUsfJ/DoH5IWfxn
fTZUYEIpxQs3F1rLDm0eYGb1P5x5BWWa4TU+i4jz+1mYOPNlpkBua/YZzbbnC9or
zrLVlKW+MZ4b7/oNk2VrKehwZEEN3e0wucVsA6VsjESKkElZKIjr8ocZGnKTqUQr
sRCkHSdPfN96Q7MsjunaeYs54EAYuOakbBr5n0sn+pN4MSk6DeSS0j4i8xyJSEGI
xp8to0UQ9Xvirqi5k8nTcEdGbEyYr6G0ZhL60OuhRn2XlV8odthA+BB7Q84mhbKV
9ax9HyEMT+rAZcS54sR4BW5vXkyAaS/B3HZT6F9UIRXTuBGUOJ/gA15amZ8+kter
xsOX7QcOYtK5jLeF3G5LxQYbfNr3beQle2oIQPY64JLtlInC+7pmdOZH3Cqwy0Na
+LS2HOIfctaZckLkBkFBSbK6s5lBqZFgDAiijADseJEMKBAbR6ezAXPzsPDrWvj8
LvkeNPwEY3ICW2bGm5w6f2lNufdLGEFSv+JLwSvp9nrT76Zyzs67QWg9qVVuJnUm
lPHAlqw0HMO2St5okJetdo7E9zdGOgrrMOC4K+gCmX9Gb6FMuAXqzxi1M6irIcQT
BxX54jnYiM9vbYLfmLvUtpZHXakdF2iI6GhN6VHgjt0qTCLBzWmqOxS+SognxpFG
TvAYi7BhdYEE/ecYeepKsCX4sxGJ6K6AZvPF5x1UAnRQBciKt/MMTqt8+Rb87GN1
vzjBynFz3JZFE44FyZy5ga+BB2D0fkkV27rDE3d7tUeU5hn/M/JgpucTYEUBoeC3
R15sC8qfe8RBoyewy7ZVe6ioyyGAd8DKcn/FW8jLmSjg8S5ogUiwyU6+CqxZVe6Q
tyODi+9wfXw4fFdV2oR9SmVPpmMcHXy08w4364nrzqf6zIigq+kkUklrmUaEGFrV
RW8ZMx0tFA57sMZ3u72p7TZTsaayBYUiEX54qinQQ9iHN94n1ZmSQQ1eR6jEbsOg
Yz8UmvcMiQzYJghM/pwjbZfEtpyaPkDTMFDrp+1V8C8Z1Fz7ghLD83J4xW5prZDa
sb14ukB4AeWSGRzyLd/EA75uT20+XKsl5WpQQe7M9ouB0DWgQ0ET6b3JOYMsfMBJ
xSAAQ3Mz5FOCNGV1QI/v2DVrtH2uToH12jgZO+w4mGSOB3hY1qCFBZJsiSaPMry4
dvZTTSHLvHCu4KIlwlapph9TqwvQGk9yqNnW4GLel51cL0ZErAlwcVwNQ1jP+4L7
cA/MxEIZBoAwguIUeNNunq+Hxikqj8o+24zJy4gcRazC0LWPAOvGhyvhZpeLdxGr
VBC8KBymBo2AIkbAwjjhI8K1KKw3EohXq5SnETaO14hrmdoFhxQ16ZXMo1kEigeS
6XR8q+iuV23mIO8FqMfNp9qasXQOIWhiYIbISpf8Kr7tiI2WZ5H/Af3/jiaPRu/H
KwuTS90IMb1r7yPViCx4nkHMRR0flxIWSMrRNSk5n4eLWlXK9VtCT11XX9t0BXtz
FrtpGu3k40NS9Nfh2YGLywZHaRXiT8CKtablXqOOEgKttqoQKrIbgoE+uNPS57Kg
9kBWlM5wsqQgEUOlR5JQ057jo5pDFqw+cAcc/juNHMLVhK69zoLmT3vshji6CwIu
UtpqCPfL/pAQjTfPZKMjWTOaIFTyEos9pu2Vtl6IzoPoSc1K0x3eJ9dDfWk79uQu
o56iBaIAEQS1IMAJ7Xde/LnXwp4kdS5SbfJmcXIYx7/pnglOa0jDDr4lS3v/od7F
THDT3MfoQWKmzgQcCTitX9ivlXlKxuNutz4a+NuXcc9q/jimeFDTH6m9mwR0RdXV
isOkuQtgT7+VK/GipNUZ8DUyZv+dZJaGaVCjyMDMZMe+wVgbflu3bKF8CaHmYOmz
GrprqRKahinJwgA1gxGXvzEr7yftD8hUcPFVIxW+I6AvE3ilwYzkYiTv8YwDoBMt
XY6uX6Nt3Qoqm7rquOoBO7h437pUz4fIFQFve4hPFdyyjApqWD24lI+Yt2O60m8c
gijUH1ardWVa9f5IduJKDUFWNuw/8m6r41g4R0AQTW++Jt5O55FXwoG5WPA3Sxu0
2pbheHtqm7XI326hNmLVd80niDJHd9xxfrwod3EppdzgawNL/6fXdGcfm2kezbm+
qfJIKKsg7L2UbqbZ4pLGMhHkX8DkuzPRahiyyRhxVuH7b083EpmIz+yPhE9bPGeD
/TMQ+hq+3LTD7muB1EBEwNeXOuC3ujpYTmB0wQ2PQkw39iy+Tc+1J54r0X0ozokK
1Mc7u5I5/BiBbG+cFignlglpRjowg/k2NH7pvEI8OjkF7qSYvBE38EX2Z6Gq06gd
SqKYL8e8zTVFG0n422XnjzuTnO7sVYiHRJpA46OpZYR1DV6SP0nRXv04gXBx9Qgr
sK5cSfXHESuY/E7iPh6ZZ+kXAOJ0lrWmAfSOFbm0AyO0NZnbtxyH8pbXh3pu1RZt
lGkl46dqF8KClZV62QajtdlLvL/OqlDmyKCdapdlhEaOH+izsUVmlW3WzyIS+b8N
sdo316FGtgNswLwdb4YDSczFmCNX2v+acPWeFbMLpxXjUxn/INwhJ682n2kRd9Z+
s/kPFc4R7B6MOIz2lbO3EOwl/9fgVLc8BOfi9+Y9OwRVkfYDkr3Dg+cFX0Mw2NYS
54SynJ926GoUaZfcakHdKKoapsAur+iLrsKUH4RtBnlzEe0xqB96yS12n66juIgJ
dVWO7CjA88FIQLejaHTsGwVp/FFF62qv//szl3H8HQhzjX3f2RVedzp+5G7JYd6O
rxXHdAEhJq4o+sEscMHH0XpqXxEY9Wj+Qf22oXsNqX0w1XdSFpsnfTe1gcjKz/AX
J1N6F/l1fdU2DI6V5njykLd+QC9Il5YHZvre7qc+y675qub3uYKaTm6gmseDfeDx
qMsJqc+D4bsVEBvsaVjsStks8NCLhI+UdzOknrOUaXYu7GRInAhc1PC3fC3LHz33
RyqswjIFVAFXMs7GZ9qbfvn1WH8sDrevTSfdRG7AmRRsSe4vVfWGIqLaqMBjLzLX
IBUyWRQuZHu4eg5NH0FKugdA7FIJaSv2vPqYjr1Tzi5xie/+QBHFZHrOMaAlIZ6+
M60JVRn6zjsAVENuklLY9E94leYl0h8yoC509kC5xt41M7vb18gsLG0zK5vEmjlw
a1Y3RlHL/0Z+n13jGM4jI0M3kMKBpRVbHR74NrQmhxcX78im59lmazpKDxCNnitX
l71bF55Qz+bvSuoFsXPiewV2mRjv1T26ylIynR+TpuWPtnJpTlxonMH/1usX4UuI
e05QwqdX2NZPTsnbK5bqM07i2ilna3PXWomoTmQEKNQ18EALU/wH+sHJitC0hq+g
FQgQUhsktL06MzplI5im3uVc+cL45dyQKB3unjvNguYqhEBLDJp7xCK4N/ZYvRWl
IYOGc75yISX5JuBM8qZzw3m2SgUMKOjjJOWOfHt0ZCDquQjAhPCIWfOxsSKkn129
6vm8235kszSeEn/5Jrd8Qppzwu+U+9mZ1aOMzDIOfzZXJUliaclJx4osX4epJNZI
51Y2fndNcGLHrblR/BepAhipY5zXly58DibFSIe4SL0mTg8zQBjZ5xCPgzifbe7Y
V+0I47PKFZ7v8gIBVQScLztLguaoRvdYXfkN17fXtgUroArp4ub2vn3D5Q3z9P7i
ZL6BXrkZ1LdBhCxNuBI4M48FF0auTdGPN2aot3vAGu7ZSPWLdxwz/i9LB/ZfcTBs
VZuWzLc4g2dpe8Aey4oSFCmsBcNzf5BoipqMqziEiUF/jXKENCYQbmVISTbyUtXg
LMtYZ9bXjsQiD9iTRYsJs2W/munPmMU8RlJr1tZYO1KWqsiR3o2c4T743P6i8/0A
5qlyMNfMsBdtmLE+xr//erGpowgiQkQ/If3evhoKCnGG9RTicRn90+N1K7JKtYrX
02ChV2EMJbNsQS0ZRbFmyvOEHRh3g90xndJLuiefIvmqvlOTQqmyqF3W5ukc7Zpt
AuGVXKWxiq+nPPKtdOEeUCXPD19st8G01lcWWWwoI5L0XnaL9xMuLjxCWN3lSLS5
4N8UX4WFmVb+zgsKHxyxH6hyFFmParWLgY/OUPEm/ovRpxiZ7KNlSJWgZ/p4/0b9
Jb3x5TmKWt6yH4wyY6icjSsOwZqXHzm7Z4uySRS72Ov7NsQATwZwItkt8s6vPNha
eh2As6AEwApC7RxGhjmWtU1F6ScqyehakzFaLrXFpD9L3+q3aNjPUa8YEIMhVo1O
rOD+c3CtQt4BrJb9kUpmjW0ku1XChG285FeXy2ljZ0ibWak6FCJhwkmrNl+z+ExR
L9aU+kgLhuLDqfri2pIB6SyTwQRCre6Xy6r92RbjG6apbO4sm8Go0QpKs5Ub+zvO
Q4CE6s4/Wa8645yHTlqFuRwL/Tu6aTmr9I8P/TOgbnw=
`pragma protect end_protected
