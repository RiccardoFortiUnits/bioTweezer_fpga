`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j6oUHk1kDSSYm9ZkIr+LbrPY11d02gzSuj+/Smd1YK9e5pXPC9QCuM1igJFlTMKm
jPTlDzqjUxdFYIwjJnhqM7HgsmNKEExakmrs3EDMsje+LstjeAM7vIL8hnvhYrep
2tQPwNmQwu4ab2eBThWwJxKywhSePjHGrlGd/Z1mqPc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17280)
LjbHKu45cj1BRVsIl1P0ydK4gFWv56PpICDCugwxV20b2x+9K/VRzGPOY1uFDNC1
tJedCWIG6qtXRicj/auo8T6u8xkWnQppqdJO9Fp5URKQPfPJmi+bHox4S0iZ3HEn
5TqFimo2/WKbSH/bxAkoygopZeExKh8n48XepNHQs7qvmTVX8QLfr5fWoLEOCj+N
HCPjtwGCTFpcQsiZPNoLslwLyGxNJpEp1LXgb5+Ckbp5SAbX6P8HRw8XRhwfKcSV
HW6HLMMoyDBb5bspDmOKMHYXmgmhGYj2UlQG3+X8LhtrGnG4A70JUxHitGR+DzQG
WaGEtjgr68f6UZo0rEniw/MdrRsW0bJxCFBtQ8qgqee5pXtfHq6py0ehcuMnEmfl
rlNGCDjmpkqS5xde/CwLfqPCO/1noia+knvgAdcx8WIChjdRJGpDssyb7iQzDvZ0
Qv3aE32DXx3V11/cXHf8X9EOUiktxwQTxHxcV+2vWGsLwoe4e9gPXS9M0Oh+rqRR
lWnWMycI/fFIbD8FYuPld5q+QwuJtQS0tO6KQupH7quqNv6KuulsoINWaLUIpsAM
H8EurybA2LQu391zHLCxztXFg5274rGqoIQC57ZI2MXzucdKU6XMsjSQRi8CXTPC
rq4t2FU1LBjAZJoysowo4N+axi3ncyxNqgX9g9Xli93hGbwP5xRK4IUVFVKlhGpF
Z4DxgEDFXSak5PfJM6Bd5m7VBTyU7Hrk1zWL0nDAfL9D7UIeo2OoinHKnuEZjb+L
mOACS48xvUAgrcZPwbRMV6V8oxE/o4wMZqf0ZmJ8mzDo0SZFkLA8hYmTEDG4DFRa
Vhh1AxiuOa7cT/tY4rrE4sjdoGgcOGidX1MMVgy3pfNe0uRssAomB+7F6H3u7R1D
kexWevtjlNm1jG3hccYBlGluDk6IRq7Lpz6VrJpwnJjF5J/broUD8KkGS7hfd9fX
KIe3yfKMscRbw//Z2+iZgY72cCXCnl2FcEjlK7PvwqFGqp8rghSfDwWSzc5/jpNT
sa1kycZlqAfUGB0u5WwpIsCHgK5E4pLbudYpvcLrqIaAWMtFWQRiN6357YdoWbP7
sfbmma0mDljSe4uCoTPozAKwYhGLcYFJoXgKlMq7GCyu4LSNNYct8N+Qdlkt50aN
64EfMtBtE6/6gC2tltrxcZvxS/UX0ak+4p2bJTGqxv+6HIB+V0n+mJptfianxVBA
jf8SAFDVQGYVY/c6ow5VOYfyybVsgO+OeE+38atvWgc/fRQ04oYGNQh8XNJGa5/m
SeOJdzjXun+uDxRZU8lw+PVZciWmqm/zljkBcHYRncn+XLlEU3KqiuD49nhtgMbw
WeTomjRHaHkDXK+3ptzaxiDDrhI4txYM9AT7qXg+1mDXegEXqPgO1YnO2kg8pY8w
zX6ghvx1SodiFNFsjP2Zd2nBD8qBIY+0UZhrgq4XC/uQAE9o2QzN9XzLJwIPm2H8
Fku7ySV+8evD7AICMQU4kPyeXAo3R2XsWwB+C9RNS3qmJi32kEsoA+71ix4D9t8l
iS8H1nClyQFnhj5YSzBnKmLHDRy3mwq92m3jx1tWZHdr2MY9PBXBa6ltrtzbypQl
9psVZOPS90C0DwS0ry2mtqfx0yfbknOy7nQS2gR3N0N4/VOJF4Vxc9O/YgZAzOVa
n6I4uchWTxoBNNIDdnx4kXbyxlXUctAV4AKMrFDBj6y99QyF6KzzqRgrTfMItw1x
e1JYniQU29FmGvEVA7ZXhzvgWwsvdiXQPXim22j8Wu/t/LApO9/dOBIjvIHxvFmj
VBl8kyKi1nvs1F08anZQKkcie4wgue1vLGyZgFN2OcxSr+1exMqAed8hlaebAWlr
W1xnzf5Ee37aahtqUF+jX+SAd+8wXCJRoOGt25hPHasQa/p3XRqvfG2qxr/Laqe0
TUwE/zZn3KxVAET/lGEUdXdvzkTtjogGjmoyncKe/hI5fVVFbSL3KWISUXDjnhLP
gLNkec3BH118N/8iyoc3tEJ0wnBssMi/y2NloiQ/BQBxkoqe7oU6iElR0BW184QQ
OJtqWSMcupPfx9kXmq0XeygUhWyVSvXdmLKv4ecBct161q0Jbjk0CI09pwvNJE4q
9kas2gkPHbpW2VunI5gmtc0mA5ogOWIXl/MEEb8gkXYv8juUfrA7tkWAZCGW9MPp
rPNWj+R7x1p1i/HuKrCS7ffEA5OH1ASZcyOPyFd7XxzJWbHVvs00dOYaHpSctV/K
GEBPPazhwYDzmGOFZHUMu3t35YfVG7f13TSOcJKiHWExNYwlBHxkmyqk1a1RZYi5
ds7N1O1EwK1+ZpWIme2C1qMMKSJXgnEfuewLC99RGRTSF7gznCjMekpegFd+i2Ug
2YIAMcuQ7DO+UA+UU3WKYOYReof6jUt0DG9yydeP5ekKODk6BYcA+qSl6UhxogbW
Izuz+sXEuCrLZanKNA1pOyUfEBwQRXF/9187yMqWL2vZFg6uoFXBOSTEI6g7Ukp7
GPar7XvTxjPvVv1BS6/quqMJHWx7u3du2bcxD/FvxPZ45zZjHjew9lBr6WMn0DFv
Gy2RACvnzLXEIKZqyYR3e/RMPTeiRDjUzv4zeZX2GEf2xB+dfyyXDj19ciS//bF6
j5GmmqDbO2h4vmm8ePTuepyf4NLHW6exvpyrft0Y0v9PvBD6G4oglxSQtyMbgPzO
C59JNu90PJ39wrZI3b6KK9NUaWlPxXOXkCXA9ugknlwTp67gGwHQZAqVeBQh9arC
xLTy5Eu+yDrrWlXY5dXMgTiMLrOkV3rzoQTxaJoE1KSM/gkn55Ar7vkggR7oSOfo
G9olSjt/JifD/b7gSviBy3eWmFU/JBxTOh2T7WUE3DVVvDMXiEjOcYcYehIszzB0
oD3s3Gqwb3XFokEVeQsJGN1RBfRAaQ9apIEe5BBYLhgce1GS7by3sm6LtEFA5uz/
dr/j6LwitRuBS0ODEGcnkBremeQhSTH8teVWjYoyXIhfao35qdqiThcfC5/k3BGF
V2lB3cYYOJPU/LB21kVZ+IM/uOw0pYMpTl5tQdtdoYPGxVB36enk/oijFPR2JON1
6GswFLjMZ3WM9WuRvQiqu98KNQTxUVK9Ncc/yE3lv+r5INIq8h/PdoN2xZsRZe9J
PsJIQiPBbzNTaqRJoouAnvuA9M5t6LgVSHhMyQ7AFsE7vI95xR+SX0tewWesQf8U
dMSJbgwtUUw7Su2/VSrNAW6oE/3P9IESa6QAA5ywxThVugVg6NqU2OeYrB09RJuB
9QX4XanHF6Fn6KgrwrHjFFEzHaO4V1hZSH1K9/NC9mlkSYsVQfA9hco+PdnxjBql
QJUnmIMcufha/7rB1el3C3k2j4XwvrPdpWs2UaSMQIybRmGu+0zp2P2QJeuWp46z
SFUUqRvSBVLdgJYOyy0c7jmzVYYq+B4+wPl+92W/ZWfdHcGJg+ONhjbRxuTrMrDc
C6xWqnn5bFzDkvXQHzwc2Z/RN6HqftRgKyj9gNJE+m6sJ5dvr8/4y2r5OseESBFG
PdigeuIx5bWi1SAdzfp6x1CKDp5laij4pk5MXOiHgJtLjOYe4qV/oF29YAnUTrvq
NlZTvyDer6E7WY6+z0jHe4LPnCGjqj2sxdktW/mZ2VzL2NdS3d9AU9jwYW/KVoyn
+DpeowcGYOBU9j8cM/o8N+/ZROwVV3wwwkduG+11VHtufWjIbxpqedTWLjs5GIkJ
qA7DzF1iQjCHxXGib/El72Q71bthgmUnCzNuozRmgRMfN53VTkRt7UJP4n7scUcG
NDNDgB22+Fx5GfWMRubmUqgM3IRtphEgYbIiu+PYIuS9fXUsuX+seJRIQ5bFVypU
vF8OgGzj9pTlTyAXmE9KdxQICZznGPBpBea2I4Z67Srd2D/N2zdQ99R6Ykf3j/bY
wuH6424QrQO8G0tD8Al4UV4DkuNq1dTsOta5s+ZzRfzYgAS4WMHzljEaVZN9krDg
LceHPpxffc4i6nqpN8OqJzW+v0P7z1adF9dU10MX2RfMPFVnVk+m3FP86Jafx8U2
jESdzWFufxiB1u5QTR0A+CA5tgz4KK0oilmfTH7HkSziJq9bkZTTbLfpT7p4GiuT
iYk0yf8m8UH7v2JkImKHmkLXZ4nyCpVroPYZuwMWWDUNsKkiQDM5A+R0Pm/1gRDu
1eSkCSlKHZZu1Xe/eVisJ1zMsL3PyzHJgkKhpfByVBoHTtENdMIhVuBcPnPP1B+3
b4gpAxf02xavR0pwLBAaVwlN4IoMUWu5ORznBVzomkKxOpQYfVUE/56BBAY/naul
ZKc86hjTiTWY3xK1jyT++ZFLudWYNeR8x8hdE/7oAWb2nnpagMAwUrLDc05nXIVs
dZKW1U/jp/gG7paL6TmuwgpZjYtuI97uMSMg9uPCUlDPCPLk2kIm85R9ZfqVM98L
5I//5zcqwsGntLTJI0R1suCus3GmRBjq6z5ODu8wOp34ftYDXX1GhZWRjVENgPxG
kRvLb2G1eRbm2lG2YQMQurD/Bv0rTbT5AA/HVnV/1mGGU1iXnkWQWkchIa7tDCOe
//6bvFpBvwvE+jcEbtsOyONL/vX8hZl8z2mkbwGRESpqc2eU4Big2bE4k+9rJ18e
Db6jWyKBBnxGylTsBPBrbIP7EcIfOt/hvvc+s+O7+MTlD122+EIOUGd/b821AgNN
v9zc15CNn3UMdbp3Ht3kN/AgZjC/DWoZskCtw2ha2ANguvNhwDrKUbVnxPGAf332
Bg84fpJlStEstEIHCMRJI+6QuEO2KHjORy+PFpoRMoFD2KnJub5trrCkkr2rbjIr
mCcSCGq1XwTdjfKECoP1O8VA9//XR9Ln4QUHKfhF6bX3Z+5D4Y5YQpb4daTMFhqm
Twdgefgzd+IkYnHTZ0k+5Qac5cePBRMmjxWNaZG+ikh8KF+VbF6PVrI8fr5d5fMP
AUFArjc1URZrPeKym9q/ohpCw51IBnS47zg5Z5bK1vWHe+epz8d1tm0ZZYy+ZNKh
EgIbpsVhqkZOy02nteFLdWPm8FDNycwE+ACKN1cKTXlikpi0uiZCU/WKjoqyJHG8
2ZM6gEztPMP5ey2Q5sZODT8G+QtWXf8Xp8/28xsDg+/9ri/07YUypPfw/ypyMTe0
rtAQ22JnNTaW1lvZ6tZ5JBcZJSd48K4/1RAjZXnjz5GR9joDTCL+1l9BCxIitQ2N
ntTco/kzjYHnkFvFTfhwojgNZiItGcw2/RAjHlh0UfRTNmYQ3n7mDG9xjULKBDMk
osAckeBcM7Vg4Lg6xpxbtqQpBmrt+xeRpbt+GSK7xS+WSi9GLgm90si9nubJAtMS
LQUSLK6KgdzC0/v8hNmEHwRNAfTATuZY16UsR5gEN1RtoMf6EuQG761O8U7z8Kb5
aLDv0QqREePF0si4MwToxy53dvEkIrBIJ91qj+UoyNX0X704tC6XGl7Oey0x48Gk
xXe4Tyfwba5DsAHFwonNN2Zd9AegoNcNVLdMNBsGhJAgFvXLdZkOeVWNFam0iYjT
iZAJiS+WsFWom9KGBsH0bSw5CV1QS6jw7+WgCmG4NktVLpPITZxpCCiRRxWWS3rv
XxJzUDwtW4o5cMVoiJAr0/m8rYIfG3XzgIxrir9jQULx8KOS2AcgDYh5eEVEqdGm
tt13WxUUNcPW0re1STgfGU0gvvpxxx/MNEoDJaMEgnf+wnJuINI8WXwFsuc/GC3l
+n2fKcTQin4DxRXNTLA8a/1ijHb3G3KTO6Dbuwg5f1Nub52+Ol6oFQssefzI5Khr
QkAogaS720TwTor1aj9L2saW2pbPuIgVldReYvDcYxh5trlfm2itmLnQPYAzG0PE
EikkpGU7iBIUDiR1iCIXQ8vYrP2UGDpa27uHxrwWxPXRrnPcJpkTiDvu2PF40ulH
PoKpvXoxH6V2oMAE5VWNwKs0+to4kjrqrGNivc5y+OaQ41fyAavqBuMJn/m10bO1
/xtwq60Nytspu9+WAME3X8hbkh6qck5lzCMQ7j2wOQnjZ3pMs1HLkGqoHVBRw8qn
m7GstXrpCENPhXT+I3d6hOOjlsDwcLuWThXTbjVXQuvGixuP5URCq+RjS0wF5/pu
eMpC57ozhxSiDeqXd0uVOORnhC4IAUjQgaOrAnfS27SUxOXkin/qnDfiq2zRqC5F
m9sfsLM8Fy7qQ9RFmHbQBtxUJtpHxtwGwb7nHPSTb67okcmIqgaWqBrNiTKQTjgj
l7vJqLHq9hrI3yJdNItUwfvXBzMYp+bbBIvQpFcpoxPlR2frwM/64+blmqiXJl0K
tWlbvyoVXWGLzZS43haLFyIEZhU1ln2MtklmcV56zx4+KocV4QlK6D7OyewKSmXO
rHMWvXaJxyTeIZlk6cwM4blp8/aKp0aNG1eEoDlqdMDp5FLlFYiHOk6mi5b/++ev
dbW4OY5bm8qblToJFHCjgdOS01cEXAAbvUmrVo6AYqHBMkfKuBDMbPDM+Mvgz8vg
T/WD5CqcaHmFJOH0OHzCXBo0/OS1n2ZgUi/bdI8WuJeD99q4fjFxOniXSFi+0/vc
Mgu0B3yTXJaPCvx6k2Ar7juCSshP8iU1xhCxR+mEb6/nTMn+7Qa1t4SHA/wTTNwK
7d18+nMEK8N4y0kwV+1EUHqyOL4QeKmAACAiHk3Ve0QbDnG/tcELpbJ2hBY/2Rnj
m+wRUKJ2esB2u7w1baBFi0uZmFp3clo05CJypx8CtAc2Af9y85b4bnwE4VqHLjn2
2ak9HWluvMuH42m1pr6YL3L9Y3xvpbGCtbjvyKYBF8lTJExwLnFAbAO3iErnPlwN
iSB1h+mvyXGG3qQX5Y3sU/2YOk3b+olHJwlPzBVHlJIXkr+mHGmcfS6J7HtPEh73
NkLf5Dq4X/X7aRjQw53AKzdVpTF9KMftNQ29/75ftq7eNAdIDKg4IXLAY1Eiq6Vx
NQ5MDFefjfTJdu472qdWwEjtRwtW7ugWofBu93gS7b1HjvrJDnCmIVO9YC4osG3M
u8nhM4PDGYzIM4NdmTOvAD9aIbHqeTXX5HsbVjPvOsGKJHVljfWqy4lEnx1VhngW
uiAF3J6eDpw5+AOjNujmaeTdZHNFrj2DI5FONkfNf22CyA0uGkvhifn5QItbe1bC
grPPhcAKAS2yMmnvLb76gOGUO+4jqwIkETp2Ga1R1XC3oHMzzVpDZzSpucIXcDF/
513adZ/4j9u9eGOfW9bozuGIvuqFIMdck5sWYAdzaUEVCQHgV6ngAl4/9sdA80kz
RseP4mpoBnjHbNqLEKXR49QlhEOhAfROnEDNLqW18r7tCrpVDmbd/4FTjGe+DIVF
JDauN22EvVH5T7etY+WAG9TjwDIjeT7rHsyRSnrXU/j+uFbnNgHEaGkkh60U42v6
x3XoSV4hWiBf5Jc51kVIw54AivYwIdR09/GSR5TdQUstMZnS/omOg19R0EfnLddL
gPWEoF4xMVPFOT8eV9/+KI36k+QOMIblvT0+1vnWiSvgV4ljZ2VUx7C63OZVb81o
5ylrQNvKIZ3IjluYtxillHx7p/CsEBOKIV+O5j8CdrlyNxPOrhP9ViXfic+wnGZL
5q2Dp35OvXwWEdO7kOnksjC/zppnFDYrIxtu1R7rd0rRT4V2NkiQWrAQF6KQClzv
wmymLbDUzhCIxikz5znCknXujnR8oL7BVVn9N8SkrcttNAgg6dOm5SarKT2NjOyE
/PLDCl2jg6bt+Qm+qlYwt6Zf6bDMX+IFk7kEvfJ3JAEg3k4DM4u8uRk+mVa9Ahat
8+WoRQf7/gfczTTx+Cxoqf7r/Mo6YeaDj4kSL85zVVKxH2VmO9k/6Oc2eb1jpNP1
CTAFKD/wW6WUGtdirE6egUhyeh+RbqJoCz8zo9rFraNXwv9I+daNCosuMhou/1mO
vUeRUXUfE4GtLXKmQh3koxEb9r1DPZyoL3Pa9AXvvdcbn9zM0KlT8anjliPPfbRJ
BOzSFg+G8E+D2ZQGjPSFidv8CZ9lvI2rfCZEKu4RYqnZ9ItCQVAv75uVb2FDezG8
zYGuJZ9YXSPiy6yNGZWamelJP2+KK26Rq9xd2b0aQqxq7SudeB/h1ACRwiPT71uu
NjaisS2CXvgqdhXxoliGWvy9suu+OKoFQe7uk1WFJvNFDuXbifP7llR5fOPUcdHW
DFjuvzXMWczImXgmvihGUete/e11YmN1A/hV2DLZdY/9aKbcg13kOpKH7Cpe4jDB
rqC0hFvYQ8lli17vBYr8VQfMeZ50HSH7Pu7p1xr1YgAfNm/LdMy3vAPEqGMSa2vj
TczI0tWl0nwV+mtYEEdRKEZwc2JhpJQVh6uZ9m7/IesDyGmzF6X8jLJQNo2A9CR7
7lZXizOJrbkqonu+ici7d8BIVZ66quE4Hjrxz9u/dqk9vyrZNF/BsUBo9zGlpGxr
aU2JT4nB+iHu3ptaGgQe639p4W1dtjnF2V5h1k5wjkM6ajfNL/wfTvhKM9jFL554
yGoQ+cDVwIqGmyNrFdjMgV7nyXnlE3ZUS9Ar6ViuOYs3XS5+n0KP4UC15SgCrG9h
etBwvusCLxN4+bjfvg+562mNauE7kG5PcwjAw8K+pswRaN2gVupeKEncoHCgdIDJ
E4TYf6gyoG0cA5IXn8gVsUW/bpB72dno6VptGJZtEs6xue7FRJ9H2ffAv9zZjTTZ
VXwx5TsBmTakIPRKpVjh09xJI4G2flrzqodTS0NunMS+4JPbDhLmtdR7S2m2cdsK
k3f13uVZIEeqZkOmIAkrGHMjmA5XALJlrms1qolNwtezUWnX4fcjyHai7H78v9wi
ppeUOO294eL55AaIZwGUD6zWJI2Rk9qTFEiGA7OahjnzOdEFSNGK27H9eOzdwjXJ
7275M/1Mw0tf5GgaxiIbgh0+JkaOoUFLrSLP2KR0hcmBv8k+XZh6TOGZMjpntq3n
cpswo8FwnX/+3DP7Tut/xVWDtxmqwhkRvdqglMx7BuPXcD8HxXfBfwrNQOObWVIG
EDinmkIsKHlsz4x3ezH/VINmPoM0m2B7MiA/u3V+kWs/hHfx3oN3YFES+gAewu7s
cX+B3j/yGsKLVKNXRHtonZDksqk5NgKysXVyH7EsQFGmnvGCctVblwpeNTTU/PFU
p55kyp9tvPEfHYQXFT4QBcdpeiagzI+wPN/egYreLoXv5nxNsSyta0fJy19mTeIB
jeNy37augnJLJ3DljfNojyz8G6wRpppyt5GLdZJezokkYTsJnbPo5+b2yq3TOQ3+
DUZC2fnGZICnG/L5XG9GFzmoCu5xfAUHGnsczvfTHx7V0P/jzIMRL90t4L64VPvf
WmxPq/D69X0NhPLYpCvQdscM91QtcYD/UBMeZK7Ux3A2ELdVq2BoGmtqs9X86890
rn806zXXTopyyrwUCXJ9J/XAagR3aSQp3FgbQTDlJwpaOHrtebhVZtwAmWTZKNts
H2PtPuQscFbYvp9/TIWfnGqnpsPtElRY5vj8BmFU7tCsHNv894Ihjh68CUC4MshZ
WqLe6tvSOFIW+5Ozorxf4I4n13AsrXCmrA5VPO14twNO+JXf7VI/iyoj0IfL5fDj
5s+X1VUtbQ6RrlruEIr6LDSxlE9wg5KKOlJ9BkVSMaaeERpnzyYxWhPpnv5wa277
InacCnmIgopVv6HIJtyCBJmSYGkJ0GSr7SyCSAUW2FKL3f1eMnBBwUu32LMpzj6U
FkPS2pzfTUADfgRycV4O2iTQazNGHrcD2/llDKRLwdQtquImFDJNEsnFuoC3EHau
xKn6EDs65bQSM7Ws7WewpOTReoBlCjC72pgdFnPGtSgv0GJkhcoNIkNLEIzicHDR
cWtxkiZoOCsJWX6zIQI1+skNxaSoAN63tomEDVuyqs8XGQay/YXfwXsrB+4ELyDn
d8Qbb8PQ3RtcLz9gJiXb8oliaQRA6gfBUye5D3jTC0lkhHTRxnpN43+ktGhBOKnB
zTZn412fsx0nnpK+Pff9R2kV61XkVsYVUO1Mikj6Ti5tM41+WTvkxoSuceLccbjV
SwN+7fhmPsx28scTIeNr0kIalAGWc4fEG8Gs/gglf0phTas5HnY6oRg5vF6Vj1GN
QY9K5fhhO3q9Rr40KtCYKg/NBkZwXLSWBaHAu0lMnnGFiGCpoo2h61H3atNSctra
YuMmUgLrMUQmDutPWjVyPhBZD+SdyU0fDTwd6hRilXargKOQiPUGqC56O0iOkKe4
9cGNM+QgCNONkEzlTmyNJ98yTG5gD2i17o1ug4ME4FjDVsLLWmM5eBaKIBs0y4R2
zY8rmni90YgNN7XSYtxSjVSJiWCxU+Qo10TNGgrwQzaayqtURmFrLwV2rVnOhLoS
s/x94pCY2tLb5LrSOZz0EysIle6uTeMtHMAhbXyVYTGUV69e/Yu2HIs2zXaed+Ag
1XxB329vTDVTgaBMDja3UoB5paPv/1y1TCy9mjn3lxDTs7koL4NsLBDxL+SF2PSX
IcEFFknvtliojoAQYtYhpRstNebcK75PIQ7/hHK5BIzijgKRh4+6nQ19hV5lSprT
cXK8KoZtx9lmGVZZilSp61CeSR2SJ/XpDArf3FnUnv9IcwGury90d4TJ1RTy88es
wfmklHMsxMN7g6nRKhynln0D9Z/o2wmz16LElSOuq0no8TzrlYJOTlwJWHVa0+u3
6W76NSqdRWrWhzeM1AeDnHcnK+7rl0waGL+vEXgWXGbP8n/Vqe3nG61mIaNXqL3I
XhPtoWXJeZtALxnql0F637YHGrMvMpyE/fGYlila6Do5C+AjkdLLaMf9lX1YGy0N
DRxZsqWueqm64Y4/xOFSoueCRWoWIpsJT6nC7/PjYpEMdDtuHs6mNBVbpdQgO5uh
LyTbdSEPEHv2pqj3kHSybAuDGAgvRd10mWt5doOa+C/Q369HOx9iQoNsOm3CTevf
w1UxomISlwtEmV49HClh6BZ4vsq/T6s/5gk85KMllqaYZDEgVmc+xcgHDT9IqNvL
T1Qd3HS2cnTw6TrTKtKwwlGUbFNz3+1G44vpAKAeYkSG6aSl+Or+eyS6ApyYzU36
3e3f08MaUiTuF6A4n/aFERypkTNl6iVrBuSN+CaEu4N7JOoDuYdKedyltRnDpIM8
ZnSOCKTGqDxfUqUW1c/jwrn55GnSWvQF7lbSn4uzk2e/JzwcnaocqJExUK7Sh9dG
Ph/yTjExPU4YhMYUy0Rfex5TWuZJEjwAQeTA7mn8wODdqjAsv8bt0coZxF4aKY92
y552bw260N/5YblZ/4oUFT0nibluk8dxIC4U6DvNicXch97ai9HOy+CzadecQkFq
yrP90EL8P0uT6RyxTdl1JQ9BCFYWKY0OA/3NlRnBxECxafLltaEp2OXtKKRR0eob
nIwr2ymBCJQyd6jAjzyyKjo/2VAHPs1Wizh6Q5t5kIXKTtRbd/2rbUN4Ssz6C4YU
3R3rkWPNEpeNAsgZj9QVdUBFNwQ8MK7iFFalN79IjMdGbJtkQRx/3Ko8ryPUqS3Q
eR0YjumO9mhDj+9je/pVNWsfnhjAuKtiAOC2Bg8BZZhnWBNbP1yPMRGzHOVSbpWL
jgmRVhSuZc2AoT2uwChYSK1BNgeCczaTxykArSKDWrNXfkjWI/eiyHdd4rofxRff
85cMsvhIWsD0LsiVBUeAUyxm3JYjsaI2lFqjSa+qkcB2lKrEOW4ygDudBiob27+9
dkZEasWNRpr25Vg0iels2+uWqMVLtqk5ml+mj/6Ydk1ZcGlnQtq6BoP4fcirpd1g
Xydzi4jxLaWIu9uNh/n7d6CRW+k/iS4WxHqFcBip1aTAzcwsv4CnkwivRI6k8HjH
lZUQRa4X9T47QqkZdH4dHux/S4PDEVPAXwVOzRPyiJCLYXn3IqoT5PFXom+QqZvd
R84qtPfvQY3Oh3fVJmlnUqpQXFJ4VJ72qSk44o/nWEdYVCx1YxCirUj/2K/kAcX0
VnRwR5PmMFMnVUY78JiiNj1dJW/uiiV9w49FaQdQNjBIQNwnm6zm29hsRCK0LUSE
SmvITqEHtwHj7ptEUNWlFJEvRiw2qfg+AxUoVGUgqm0Hm3ptzgsjYF7jlxQqLTGf
W1zJCo9DP/ToByUQ474ISXfkN3tmSj5DjqO9IIfRtXgo88PgRDeDHHzUnFbiUteY
5Uq02mG3PyNuU1n82w97viviOD9fgPDmp+xxHSsxG3oZ/klIhMIOj18y/wUKEplt
oEXbhq0A8uCe37woSYV/kN7l0yLGpO3Knd5mcgQeUZANzvmy5dDStrH5PH9nVaCk
n5e8D3BI6WxeLIb3HdNrBAwNo+RsrNx0LPx+1AFRdDdGPzAe9VZgOMQwh6VFM8uv
ngS2sTVa9gZESJANvH/fSKAkZ+GhJfXTi/sPbrDuuTAEVNzHsW2HFH7nlTed/iGQ
DXQTAde2y+LOr7TOO+ORq8EhjvdqZGF0PZW0TbC867iY3H+L43iYxfzSwUMSkK80
BDi3dkOagiA8JRgSYKzBPdnEiI9xbqMYvRTnHCVcLqw0BlpvwPtNQlE2A7ejlqJe
uZuxXqaoIZM4VEKVTMpi1aNP4xzmQVZ0wTw6dn0tv7CcDUJFbkpLkDjqgq6LrcPj
47BO1X8F7YvjIagwp91y8kGYjVzXRPmkTOJpctzFd4PFWvIX7fG31QNedHNL+rs6
bAEnEYzU2LwH+YUUhS286hyNV3NaeDMi6pPJ01wZmZVqaLC8FEN8pOxLVz0sLxze
B+N8zHVJ2HOut4p666EgVtnbkUFiWsx+dX607pFkZK+DYbsHA7Nhw4rwgfOJxuSl
vlICP2E0wzUnisfL5/gk+31oYMfs+6Fhum3jNVQmoBQ6J6w7CpBUHSalCba6dpl8
VNqOoajJbCFMoBUShU9fJvMzJ1MLfAgV9E4Ebfaf0m/WaPnzyW40MxWABBgEhLUt
vrq4SBhsd9P/CsFq3lhbJfbUKLyAcQdCY17RBT5G+7oRB+MVDTjsu+owl4AKyYzn
NaCFlrE79VMvPYKEtXdBP1ViWLr0Lz7t8sssfMnqDBp6Qm27CWmpZ4dTVAtRMLAK
7tzGhfDQ5o6P88Y6kvRqHCD118kLIMx58KdBaftk9wQfJ3DtOOqAqyNOy5biqIh0
6X4dxYQDr4Ck6fjgH4MXpZMZs/YRuhNCQKEfM8ihM8jlXJp/I903PwfyTba5Ay3y
ob7BY0x60qmNfsqVBFbLO0Fx+lSmYwi2cF4miXn8ZXvMhMX4EgVyQI35NdUXqn9O
0+wa74sVpl91iH1ESbV2hzuHvhPo/SeRl4ZcVpAgcvWXIHZtA9dzpcMrvsiDg1Zy
BYtKlIRqFkKKmmzyzTktykMjB0oNLOaIbatNltsJfAiPvzvOwQtZ5Po0JKO0qPSy
lTIoDZ3LZsGb7wjXug14RNhn1GCCK00ZHAjL1hPI64+Aua7DIq35zEeBgiKicrbk
cdrswqPv3k2F/4teiTusO+CMpjAoRhKjeVxgv+LaRrknFcEzO5r0VRj4r8zP+nqD
HixHeUg/mOZXi9n/8Rn1ayF8eIiJQZQiKdO5mnXGS5PnGfpy5s7Px1UIx1VsN3Lo
4a/dh3J/zjUVYt5x9hIoPREjw0ksSveiy2b9qSVaaBBv5jlJX0WFzWCiGYgWbSGV
9JjIiE99gzO9Nk1r0MU31aAGDGaLcG6ow9DHGUJ0Saeo/DydZZbnQ2kxXOUElFBn
tVPEEOT8kfMf5iIApRRnr9HrfiR1EEE483utyFiy6kf+vtPrNOOZFAmtp2I3F4lv
OXO7lmpQqsdN+VQXs/Xj7HiehVTSKZ/4HTStIoPeXOowpk9oj4N97XqnW61fYj6S
CuRkkvJuM0wbxxr67DC0r4ymCOahxbmXNjxX5/fmUnYrRUNvbgVLdVBB/UWNE/ni
wl0CC/e+5snLNPjgseIjgScNeuuoj2uHY1drm8ksO2Vi+W56v02EPnQS9NDDW/TL
9kJTB4/IUWQNKK4tEua+UCV30CbYQ/iAgNpXM7inWoD0ZUk0zi1E8OyxpajXgWrC
B1URnnIZyKjGqwuEDFFXptrQxpuu+Z0Ifdrk0qWBAaI0Zz5gJWFBvTywZMza60Qu
l3H9t2ZvJaUM5jVT2Kqt1jkHX14bTgoTz3kXKkWBrYHyF2RYqR0IDV0P9J2h5/bb
WWB2W0xm/RMRh6bB08nuyIWykHOj1SHYUF7mQhNTk2wLOQh8kKzes7b/jTDVl3nY
XqE6/MMKoLyZutTWG6JGZEAevQ2XTNHuyRXvP7hVXPn5Pho76zT1CroM0N2aGgQx
Wt1O3DPY4S/okkQnSxhmdkwabZY+zkhBOV7YFni1kG+MPdMpsqmLSY0uSm84N7Ot
Om8VAXMEM96QDQ74ZfEq1voKyWtIVo6+qfkl0t5CB5oiX7D8LZbycXnQ0pBU891k
s+TGOr0QjSaVbPEx8tLfOIIDBUGmYDDI59ywC6dvkA66uqBjE9oiSbaj80cWkAkM
ve719CyD4u6WYFxUh8NDDbWFkCWcYLocS4Mf7stWynvh1pEGZtz7/d5Ff3nLandH
kRmEoD+wW7rI4eckdnSUQgUMirRvl74pHzbeesF5tah26O+WAvvlVpiedLFbj3RC
rVGRlSpPyOFlLs2Dv3m5VfbVDc8BoDWLSsQ9Oa85mMThxjTFkOxTp97e6uhZXbrT
Deq7Z5ABYHHZLJgL3dHlnAPJjoK3At/UznIMa682NuRID6FOxzLch1bjTnm2/itC
emk50VL62dgAuu7E3YTbnpPui9+q7Ex2Hn9nnj4dQWqevJC5/pk+6SQyO0NgtEXf
wiQIgJmeUno2lFkuv2byF+ACkSdCWMe6u081eK8q5+4Y8tEv637gS7WaZxfNmJxI
rL/j6bR5/XZZCS1nfCcDOPu4fmqKDbOjGWTtJ5IsPLd/5/EAcDqkSO7h5oPIiTWJ
MTkypu5vRYtdCXCw6jiOG5/g7iQlQIfUwdzJcYJbMVk7N9vzHXHOcuDw9pUOgB6b
DAsIm1x5fAvV0tDF1BvOmnJDkMsIH4WQanapScKJ0IeBh2QRMyJgg/chOOtfNOaa
XswSC1iVC2M9sYipK9hXbWYfP5QNjso4RX/qkBx1LhAkFjiUhOAp1C+l0Gq0sORE
bjGAd6wAiT3ZUqYJE5ZUW+dAc8YIreeAvuzhzpP4tWYJyE4uZpXWxX+7hwIO++xx
51Uz9uQQzMETCGv3WuhFAYj9f/eaoKyyhu/h32z+v5KD3dLFyVxor6Ml2VBTBxsD
IPNcCKSSWLFZlQfXGJWCUegoE6qt+QYKQmZPnKuBRPZ3lQRYn8um+PX/ipTvRuHe
IDcikqQu4uPVZ7+7DR8zN13vhhyojDpM+UUSi97/tfVxXAGJoTxkoSaEXm5QSzO3
S1r5I9Ks5M83h6d5d6Yx+sno47rBF2LVK2dhKRgElzdIhRj4PR/bKeYIvGFI64uT
7kQyKDV/l/a6l9FpbejKDWlJoYDlwUh/BUwPYR5Rpq+UvKEroj/61t7eWOymSCA4
z4sgAzXY3UsZ8erykCi5N1F+S3s2Pg+/akjyqMdEc01xUsfsXq7t2rc3+UCS+bnl
AdTeGWpwTaC54WWfIgMMrtk1RCFg2d+bHB2M2ZwuqPhYvw0q4pNgeqiABH5PQIwX
KXXSTn5cj3khZb46hDD7s9SouqSIvPKD4dw3Ia1pTEzI8et8vJsVKZLetE5BIhwk
uT3LTP+SJaLMl3/InZ73SjvcEFLRjpQ7AmYCM1vu5UchxjLgu83SOl5j6EQ8Lbd6
FyBCyGbZKAvXkKBQyB0sFcvBh9JtLLzM3fG3Vw/PbDiV+QooZyzEs+9ScVuCqorv
qwRF709pyzaCUadYdPib7+6TfzxD5vfI2ecE+grGPWM6l/ODPbIC/HzkjYiE0Aur
fdKhSXsHaMwt8/t13EtZ7Q16f5gOBfx/2WQh28tmlPi7wHpH0mGN+6ZB6FQ5Sbx+
deL6+JTA0WRGQy372GMSaPtjbFxFzbzgq5oCvYQseniN0pPCA4aXQhb7YUrcoCNc
BPHWA6MKdLSmSgzeBO5DLnly9kHWUEDkzVcysWK7ZEbT+0kEZ49Lb/eo6FBeLqy1
DMTWhLf1o7RstvQvbtFPsKFFpfBwSeMQWwoaXX++gs6SgUxPQMkqoes+9tLu2+f/
Dqz7/eVy15XEOuoK6+00D267ruuRsMOKjnYcmjpdqGfVS3fOUxnwlQRSYgr5vAtf
dB6GZAcm8KyS6MIVgZJp3ns1rs3sJKvdVAd8F/F0OuhGhdPUtI1BosmkDSPocE2a
S66IX5fFmeuiwXJu0S3h24I3eqSn3ECwFQqinJ8s0yGSCjRQmIDN7gV5b8Tubv3X
zZ0kxOQnMVF52TXsebFvFu8EgDLEWX3AIoYat9R+tE6eOTirZUx9CNUX56v7VCtv
XQR6z80kMZ5Rjj9NUceC4CdjjeanE9NW36KkTECWXewB1gc2fLqRKPE35RWzEE3v
RXH5Vq+Xj+u7lj+Yxov5RwJsFV2N2hDPnFoPc4ffjp7fHDRESXyELeh0ek2c9OZp
dvEAzvmWuar6wm8Ol84jhdeLIw9mM9g8yZoCcoGBvOrRAY6iQHFToNQOwl9F42Ct
ghAgPbUioWq3uSz7WgKCnIXwGJJq7OVPEoPeUSofdbSNtJPqKRD2jXD2+rIpOdWh
0ZOG6v4/E9WoGyaNDMGGj6g1NNmoF2DnGLA4LuG0DBhZiAiKxNr7506NmttivEa7
AYrYv6aSfiHDDM15L/OFvuFPQwftetqbCwnmkpo9sxoZqbrNK7GMRlgOQRn7tXEv
ITW4LHRBVmVn9wH4MuqxftVJvDIBHWfJbs5GWgnT3M1YLJ+cYatmRaxYrurhvGms
OrZYoLJm/zir8X1FreP6Uikd+PPIJPYLOGx19xY+b5qr3yy/DE5r1O5MMlWIhpGs
hdI2NFUK37Z57FZq5l3BP9dBxGbqsyqUB+QWBMKb3yvYiJIh2bNaz3dXUy+/8bGy
TberQsMn9OTUXKEdQpxeRJJbFWCqwa3ZuHSAvOsVdsI67rucfdSNbfA1GCwEAUOy
5EJhnt7m63G6bx2+MGYifRvhVyEimP1V0No3ZL7Wtrlkd2MfShPK5AOYh6/36+Cz
6DMfY3Z+GAV3tdXPVP2zOYpd1IT3Jl87mrnQd/axX3P4du9kbESYphQjP75EKHxt
uCS85RpG/YVFVxoKx/HbTQcJ6pS1Otz9Nufe5CApI35MDUpJ+nDvpphXCK8mWRoh
KA7DiZ1EDpsqiAA/Usc3v2rIkKrdvLQi3bp1t4FbL/A13bn51k5ydnrShGn1ZQH0
U3vO5eaGGJphxR+JFxTIpCOUz0wD7qfdIw9MrNRCosSJnHgyxNHH9Nh39l4Oeow9
HIXlri90Loq+iERnoJ9C4fB3DgqmTgPAzdA250cyGj9Dz8FY4Xk+aDFYaHs4XNff
52PL0vART0wfmHX6E2F9V2j9AAqeNgF4JW2zjybPpbKX+fXpw6r8OwY609yE1D4m
RS9t3krjoAIH54/ExOiYCmGRmdDwH0UNkK91BsbG3Spe41CjOqD1vR5IrSaq60ml
IWJLH0aDPlcUftUrnlVxEEDSTOR261Fv5Y4R84wMlXPyQIjhAIGlqpwhNa0kQgmo
HEeQDaFK8/y+UQpd5SVmcl5QldEYVyT5v4CUVa0CgrnLtqgehLBA793eOQ4ZSg+7
MqGf3p6YRWfXe8U/s0iJIy+7w1aagkSrGRbUDypSivtUDN3EhCmemN95tuFTBDho
iryXDvlB8fz8O6X+XikiAG1vSKjPnlD29ib3gIRPEyHbN6d0mWVdokglr+RfWDZI
EhTcQiW+hxTLrS8/f/lPktFaZe0s7nAx0p+en3JsZdaU6UXRPBULvruwi6JXSFoi
3r/4dweH6yOnhe459Am3Ib1W/cENnXA3XP/mHAk5Dd245FdaDiPBeqBAPCTPWl8c
A5pkAL/v/oXoZTWQwzg6SIzncE5cJfdGmV+Dji1ynhBbPI6NccXI7IwBqhf/NaEk
KFPJtKrAzXze6dUmqyfs9iXF7W+mER0BKiIO+9wbPtGR8TVShkoGRjs3xhc8wb+F
Fei+jJX6FSX9m4sS3mUKvFwkBkxI8Uy7V8uPuKYr5kYXQQ9e4e43xt9qAb1S6aqa
Lbv+bumzjL3L8DlRsvJ8VN72sLwhKHru0yQVgrApbHtO6dtqFDPK2DSLlZnm44rY
9fquDOmhajwtt/H5uq0j0TBaihmkWhyg8pb7kGVQQ15YJHla22sn98q6yierkp5h
J+CBeRDqGnG45BipVyAVgKmmfYWTxG/V5fOrp2+a0bGgqwJrBuD/6GMVFIdhXfQ5
HB/ZoFyhtOP08vnxRvw3y2LjHh/YHdgPvrv3gbNb3vP/wszosi/wocF42u+kOBFm
2xovZa1iJ1Bpnj6elzGMBsWgnWq4J2hKQqDv0J4UweHHFt4Fdn52QwO02S1pSIT9
kR815xrhIVTwj5IcICTH63a4E4fM31t0pw/GwUUAnMZ+VjV242B/fm5GUHc4zXX1
FF7dK5RMvQzydgh40eN7qj6+di24sdkh6R2t6SA8+nFk2tQWoGPtU7+IoBEEKbEE
Addq/nSH9Egv8LsshWKIuJAdQ2f857+DlI4LE2dyTZYOMN4IRuGm8VUcZlbsech2
OCHfn+XTDH+1JxcsSll4LBxOTn5ELIqAdO5p2a5HtYednJmg7hMCH7B/HAtzy1yY
okg3jahD6B/PSB5/hLXZW/dB8wX7TkXaWBSuAXtt0S8kcvMKcPNTks5iEBZuiIl4
GybTISj899nymYO4idyL9outhS8kiZuctBQUzGie9hdMei/mjSgYa5DWIs+11Gvn
OWorc5zqKlqHr61v8mzgHerbSaB0EgvDK7gbdNEBtnsz8p0sFGOA/eQv8Z/uDMHl
x8T+chFP9UKeJsO4UMBwmfmU3niivD8ELyacMXfZm0sD2JuarxbpWP9v5K1flMUm
F//0IpbH0lpBxj5VQg+s3A/wAhQYa0V9hf8vNkZlEUZDkYHovW967pzCc2RJU+pD
S8WA6tPeemq28g8D2xo+KSKzil1IzZksvgPLs5rwCgReXms56WoV1fyeH223RoXy
Zi2u3wugM7A3TFswz1VUtw5IU3ZS019efqlgzIGScNOe3WwaO/XGab+4klh6dRHU
mS2JgQ2NeQL/tiXu5u0BLMwL45Ule87rt9EhxIs2IN+iIqAAE1rl/l0i/oumDmm3
SsA0ZoZVYRiteioR3QGx/FefEvsp766lX7nHr/UDsly9Xd3W6pY43mXsieNWPhPR
/wvvqN38GCkAaqqiyjH3mgxjtruGIu6gZzO+Ihgr4h22UGv3JgaKR76x3PyiM+7L
AmCjBlTiurvOkF8LmCbdf7MQfRZPr/psgx4ueyrW3RKCcD+WF+4/mbkEdT3I/uY+
535e3cNoFWHeejYULWyUMc+j+1gQSnZmYG3WyAEOrHUgH2sNStInkXVRjk5ukurP
bX/ATHuEH9hAibcTdjANlLis8AES2mPM7CtltkMBOHl3b+VeLyZii33BF4sBENHR
iX+mpeJWj6PGxNNukYvl/t2pWeA8N4YdaeKKIQizBwITcubaK5rq9zj6gDtXQogM
wAWKPFtsbGo/LpZmyw3diKSK999ExEKMaahMXrynM+jmgZa9c/uRn/Kz3iD4+7dn
zI8VilEW58yUAWlDrpY5BdDN1a9NyKPIcC8DC+mM15zodDENSzHK05lvUrgcCBT9
IQ0YE9b/rNIKDYYN/jFRuc9ktRjI2q6YMleD2A44MU7/okuA6rrWOapjqgxDwVaw
lq+0i7qSZAab5njPA0g0TMm8yAzGEb/vpJSMxJ+8UoBExvL6NtKsUZ7okqNFnGZA
e7PvwJ3OnNRGMHLLYC9HLs52v4EbA2ZqeOv6p4by/IUHSsvOYsssZdDtUXpoo6Vr
vFPjWPOmD6EI5+sybd9AdjqlEZXCAvHxJTVKdFArPL30q9fjrBwgFMWF5aAqrfwZ
a+CfEebqcji+rQ9BmxB4U21mpfeKoPYWaqTjcYb1G3WZQg5l+CHxK+h2lBJDlsus
ZGPxp700aT26fu17r7PdnWPxiw66vQkKRbihw8jDhm1fObkbRwua9zc5Z0Ff/o1U
ai7ri9xixgzXaNj0MviPPDMzBUykJCQNMRJ8WQn+bgE2F8I1HNwLzXreyWRvg9qJ
AB8kT1vOhocS3wgDMYMS/Hoa6KcggXTH0dkIgzDovJ5Ot8jmdJRIsoEP6j2pqufj
aS1pHuiuOx9Xfbh39qEmFcTqXWHc5sTRjTrC+NI0w5lfgcGDKa/RNEFz56qqzz1N
L6T0yXlxujNtnl7ZM64JdYO0SIsj98EfJE01ukhcR7VK77IM/2quJpK+PPOI3hMw
I9KWSdGzZHphE8rRKLSS+H0UphXw3jkaeHy1MZYPM1xu1zfWicjt7ZeStZCzujM6
qujCMi6m8geY20xz495B9bk/oJettxVs3Xcm6/NQ8cSdlUJExjzbFr2aAXmt5DBe
ecvmCTvmSAsCV+u6rdlxN2G/p0sOjwLjgjtRb0Pvr2k1P9mk86CQuAdL1OXNQNbz
O4IKuW/4HdsJ9DV8q7H/8webyqP9XQkUM3JXq9maJdaKHPNH7pr8GBsWckczF3yn
vn3fNOugNkG5pcVjOco6ITZJJmFeXkTNBG5IuSDeaVnEEwPtBc1iykkI000wn2/X
oD+pM8BvB7ZT0/hgaUUgWrrQI7Vcg3zX/NhE7cAIKkxaFeyc5fgP6rGcwp2Nm/hm
pM6lyY+zSfV+6bQo1TzBflazXtfENcVwhtsYnEXnHaT6ZnBlW055kaMzJ+srNZ/1
9cmyr0D6AM1YCFzOXA1gJ0ng/qXvyKCir++Mjc+WDuv7XboM5PHjjx4xdv7zngbv
gSHAKhs0e3slGT2vSOPJfxjx5lafVElfAWCYkiXq/uFWV817JthsMepFJYN8w5vt
EogFEZKLdVsdHsjT01c5qwbb13ItfdLDnimgMEW9Qrb7TLCiceJS3iK8fqNni/An
SujKNsKQ0YDOYfc0K+Dth2R04naCwASDEhFdY8lvsHY5hSIxR5kz4tmLwxAwKeNw
+UnsC+cCnX7mPZJSVQP8XRSSbHrcB1uaM6Nb3fRUmQLIsQHgoBqG9UgsklboUov3
hwyTCgZFTcKzogzhQ3X5NEo54pJT5l455uqOazGB5dRWOpZmVAATrGIlx3PpTmGy
E2ebeH+z1yjmVT4S+FEIz4t9DRWSNfzdy9RXzGaswyZH7yfCSmP7Obf599navd0P
aV7pnqZEhhuXuFleKHCeVDnYbnAQwfM9ZatEg9te0s6pEWZsAlHD/IiThnYCruzh
EZAPnkhi/Oxnhs6CKlhGM8g3I1M9u0zJj5U8NdjSgMWMeVnEFv8DjPs+XdPydkxG
msF973wI/Bbcf84kdmj9/TE3yEOyCefBzjbA5M7wUorVK7734LAnG4iB0D/o6gGL
mTuo8SU0BPc891EeXG7YK9+RM1OOXdfccgwh065lriCG3mjM64i5feMFF/ZSFZP5
rq/WOsovr/7sfgJM4HG9rZXblrsjRXul5Z4X1GTgZdYqaNBnNTh/2cNFwYCfOAC3
M07q9LmVYfZRKu7YYLfYAZin6AmPl30cmYKhi2C2Urh6A2LqLeM48eRsv2swj1Ku
1KQCaFO6qEPCM4zrL2eNAfDngk5Hy/CAwfVrnWzlqo89EPW78LFiNOjGZoJCP08E
lbS5jiWpuZnmFGXaV2qHS6UcbhBjIvfn495UYog56y9X+BmnshwwipwD0XHq2bUq
NQ6tC7P169EeG1rrGiyVs9bF5OlbuFlQ9BvEGjGppDV6227WwljF1AvRRa6tSXeq
lXvVsQvq9cPT8X0qG9WGVxn/q+DsC79j5s59L4hdMxBKt0KSVTrljI2WG3pTxM1V
RIwT1azyLK9riTgUGSNlCntUZRsISluLdOu9aWAPXPqYO0hZ89bEnvKso1f/5NUp
A8MIkKhnW5nLw0Ouqg7mpMw00B9u9nq0Am8k+gR7Hhsrw87Yc05bqAS/WPredHNL
vFedibRc9FTdgZf9XV/zYyQKX0G9gsrYRykIT/YeWFZcTmx6A/b+9VieI7DWesgt
bYRlTLsNxHDu5NdqneewTQRC0mVjEvdzrItBJEGtZO5riqCvreYPEmt1g2LvXMDW
5BrgoIZ6s0uLaOyy/s3g9ga3v/P8qksqtE0/QGmkzeG3CRi6aPwE8M8pu7NWBKH+
Gtlu4rKnahg1unX9uCAq2fs9T5oP6Sr3vVqNGVJMgvYfd0JzJyV9mPZLnt5qWU7h
iwPx2ncVwPsCLyh2w6vCd+KFp/JRk79vCFjCSsmiW9NJxZOI8tGssXHzw1zg1ySf
oWqL0xCKgTsPKNQIW2gKFOT8jqP7OnIPGu2jB0TYXG9TH/GQuuIm/QHYzhzO3egR
bXsa+ZHfG8SS55onWrZSRRI1/aU5dbcnvIkbzJ6acZj25Dx7tk0nCkAqD7/2AEZh
TqolCzytmWb2nM2zK+O6Tz6aIdaLt4lvz00BbRZZ7PNPuIdvxNJVGGbX0hvgPl7M
3J97+g2ZZJQbHzS750qxK1QW4m6A3zXrAyUvU7SHQBm3aUULOluZOdNSnmP8vCS8
KF5odzDXNyl+XKwTTaJHm0WVSvtX3m/bjOO85VONgh752G2CY6vgXmm97POMWLaO
B4B0qzAwA7gjqo9H9Ong3CCr1XfYlzud0ijpI0g4QvdoXgvYXv2CkIM9bOMSvM6P
KKEv70ih+PMJTv0x3A3/YHbTtWnI1XSEV9jL+mnYre4lWFAVjQwVNy7aVsaWS4DR
mIPwoa+PQR6DR6122EatWdrvyx7XO/gTLQaBA6Ws6xt2hRpDCIokha9qE/jBP/vh
Y+0+AunwkSQnERpdhqvmM8/sZiAO7Av0Lsp9e0Bop1ihRVc2d5+Ts548Xcedt5I4
nd1U3++QPsSWXNKPWah//GoUnNnT4Gns8+i/WqHoQ8gqOr0f3giVqOm+oSwcJsoE
jiaJmmmDjoznsiA1toud3jzCE82IPXbN4IeH4/D+vpXoHmphe41JWS/l+pm2LuXt
FXOuv11U8Y4geGlU1jOE3jEtvsb/7wsPvV+afbXk5WE/wUB8CwCH3xwWQNVQyxKF
`pragma protect end_protected
