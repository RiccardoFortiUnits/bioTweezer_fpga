`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p/URvnie6qBrtkLumAqpMIqy1AHIvmMUMU+H6nMRSlV4u7zG5xc2bbuDZC0PrV7c
fbh8hHSdfXQL+JFjFALrZ3gReYLVWMoTcJKJgBywVERM0DxGi+qQbKB+m9R80e3y
EXGPzStkN8pFzr9MRBmEkiSJTC60gP0GC5ubaCe9Eg8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
P8v8Q/ulLWxMtZ53WfdOecPH2p6ga4EfvC6k5lzGv/+SwxnU8gqnBlVRwa+RQD3U
5Q1eP4ew1D65zQ+mUpKAJ839U2JEwGVcKad6TlVS5dBs7Nd+uDjAkzfO5kUMPeyJ
SMCSJo5GF4+kRMTZuFc+PDeRNfTtUHM4sL05T5etWPgC5+D3Cq6jboSqp5qs1kR4
mqOizVVSjrm7Gk6LPy1fOgGC7gJLVduUNK3FAioCdN35b3sPXyCGtRLl1ivcXqdI
JTJ+mDFmIM7EmbnWOeRsr1uX1bIbC8iP1t7ou0ie2Otk8zSr5CZoCFGmm2Ecjsqa
O/AlSwbku/zjqG/Cfn/XT7ajXqzKmSNrSSHMKGvH1YVXX6UnK8tFQkjVHLrdSbKg
5qpIHL/RMW26FqOWvpwCTYYnj0cP42N52DDHa5KSgSfSCpSvnwSbxnkBFpX/45tz
33rDvKLpb2s2BZL1mRQRMFx9sHUV+1NEGoA3+TXk9MLHA2inN2KuV1ftfxg2PEO/
+VcL+qaBxp3ZaNjG21PV0UWMHE/mfasjc44jBj8eakY+UNLJmqDCL451ijtxK0v1
PvsWfaHChr+9yQphGc6L1oa3MNUJfGU7X8JAnMjRH/sDORDaXgXgiD91HdmroFKP
FcCLrDNeggE4uDPijsY+VNLiWHjtlP+mKPSW/E6IRHYC2HY2qG4JMPprTceJqgmD
EgDfk1sar0uq1dTe9Bkl5u7m5zK/TUS/nyAtSgFHLeJ+yHNFZymxK2yxLOnc3Wo9
FwYXr7ho0N8z4dEMXSquXS1SlGh1Outxfe+FpyCJDvZ/MD4Kdvj4p2pURZvH2/G3
AgrNoNZxgM8pT1Wt33feAt0KEN1W4JYqJREU/g5ogIhjg0XUCZ4ytg7s0hhfnJyB
MHjRVWJBjbjPDDp0F6fNZivX25pIF3Pbi0+nyHyS/D9Go3xjDbgWWONP6fEAQMHN
RRsuqzfJR7fFGPQbP8pJREL0LM56PPGVbEopwZxCtFs7p12NqSlbBm2gJYxmfnMU
Ibdia/qo40B9pO72LD/zEutpqfCgmwJ6rbbb1s8J7skWXDPLop6YmXszkwOynruj
58xuwWG++eonJ9F4DS2vVhwdI+k6IHRisS6madO8v40Aa90QR26/0WhQXLvzjAyV
H36qHN+/25P7iVy93xH1bWwj8amEJOpkIT3zbfd6LWVcFdCLK8vOko0P8aTg5V+r
H1Q5/Eh8cP3CrcMQFmeVJBf+3iCzp5TFuI1RKyb0U7hwgtIhXOJXLKw7a05EdELP
Hnm4ytoIRt29Gycw6A+G/64lpil69QGIMl8QzDlPJ4TgITDoa9tcE8GLk8ZMAJtT
LT+8S+uN38hej4olCyhh4I5rdC2/m0k4qAF8e1BS+i+w0Rc2328H7Fzr9XOC3XRs
DgT/jmkRxPlM7ha+G8t4MSKBU3gQksAra/tRwvUA9b38QFNECAbevpVGbirVfHfY
6grZJ4O+/Dzmo/XO1qZOSs3z1+Tso7qHO5QAACABhHdDnQL8qhvqJlQ3wX2GiwXo
tv3I7iru1BOsTuTXQxTHXCVo3rkUPyRDM0QYIxAQ3jYT8HVNEU8aIJqWJ2fh8KY6
XC2H0OIwyMJdcyzC4xCb65mxtKjUwsQjoenVTTCM7RAu79Yx2jMaB4yHEqBJtW3y
RMSQSOnsHbjbCHkffy84vX/LsHSKyrrfl6+FyHE/z2qq582Tj8IIaMmI/P8GyIVj
npJFb/fdLqOQgoVmT+raIt7r/kqGVM3EMHNv1zRRcemMgKvackgQXeh0d58Pw6oj
BUWSH+o+Mvj+OtFr2PhJkWw8W9naVeKq/wpKwMBOkZH5O0kEx1e44IRaHBefEOEZ
g8TfX5fqFxT65zBaXN0JoLyvBmDMBoPwTislNaxIcLXcIRs1p7fg10t/er4hiDLP
l/EDugewKS/zsa+ccPmRWq5qa0ylGxfdYrMItEaunOHFcRpap+ae/bgFzC3o9N68
BrWDPdtUT7gfn4i2eRjsllhutjEnFUXfI76lYWUWxa0OHvIEELPmuUgM3XQ/aRbU
ErDSu6A0P5E6C08UytSXn+1ypcMoO4krhWXPZTj8H1gpQrghJuypEAVS5tQXpVL5
Nm6jhMJtDPZGEi2ufNMNa27NYD5yjnGW8dbeSctqfANmoidLSJpeaeQpxGl9UbC8
LOFz1HlivYAG1SzaDiaQRboAir9XuRtWAsblQ6PF+oT2NnwIXquvcwcbMn8ZpfEt
3EJoaSoMgPm5kgZr65PlIg/hrNxF+9iIQ0y7I5D5fACD8n+p+cd66IZu0c0HrWp9
1n4IpNMF4/pZ0GrQfCrJj23yGOYOBg2gpICaS/MIPrrzG1rS5cq2/s/w2ObWrKWY
Y7X//SA7qoRoOwrlZpGX/+LWOX+UuVdxHNKdCt9be5qyU0APyhAoNpsNlxCSFoM9
1VgVWUegHA9i3Y7vTHDeYPdr/tYC8P4tSl5XZz8UJzII206+HmJiMMZ4qEJ+V39T
bl2CGRrrzdFRO/yfAG5+Za31Kl4DUM3ZmYfVu3gD9eoQEO/Z0eZmUciFhjfomZFY
+hAOAQTf7a2QUaSSizPVdhMmWxA7RC7v3t2rOcricp4wL1BDdNkv3Cbx+TG72mFK
jkyBm+/tnQPUrOJfP9932muLTYjCY2kmybAfIPuk/3nI+BRc6d4eOf37MQYqywOB
+46DSdBi5Zv+xYY5knZCsgWnpn8DEsoBrSWZmV3fdjUq+wYA8whWFN1adKHaeZ/d
8zxen4GMrBTCayLRjnvx7f0vDxUMmcWhntZigGQhri3bpkiow9y3caIetNnGhDg9
pUfmRQAoGhdi5fZytAW14bGwgANx/u32GHPeNeMPZa+uCVxq48RQftrKy3NdQh3m
1YJdGS9sHMCeSkxjx6hq2PQO2i5xVlkW6j8KA4CvAJlptiu2fWs0oXujaxopCph7
8iXpkv5jSinuW06RkdnC8vZjHEX6ApHirbC3lWX9RMNy/jf3nCIUt+h4mP/hzI/V
RSVEMLrsWB6ABr22hrszfHBkr8d8kjAhbRU9BzHH7Nr3yO5l98bOtnpOvLHFzB/1
U+DkpqiYrVOleMEeuueNfzTAu8L2wBW9c1htIjuvd1SpfKvcU8j3yKfbAva66ddU
`pragma protect end_protected
