`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dALjGhu29wRs1zA4Tn/Szuiu5uzbCV30Sl2pIES9QlFyJ/GP+UIu0UzpE14QIJgT
0nmxwyAkKtR4l+oCEMf/sxKAqUOY8FcHhuejBC3bwjj5we4FSPDY/EdbeMJYt12l
3jItQm0nHR4sP0Lfp4Et3J/Ugh9aBNCvOsSYVmWoouQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
bScqhNfoM2Wmzv3gMJ0dXb7CwkEHx0/OyKLF/qz3ptnBykHjjgQMV3pBjfZnA0Dx
gVVDwejRyVrxY8DIrN5mhK6RrxSMJnlUflBnHDa2JkG4mF+2n8iXPoFq3bLSDFhr
RyMSp63v1YsMCoAsGJyEbsnooH3T4rCRLCbWYNcFVzD3jJ+Roe2VVjlTDv0nF7f6
2t9y1Av5MhJIn9y6hFTxObC5LOF/WnANr6WsHmcC12aAQVUZR/kPIvrEURPFwpHr
aq7RANig8GUMZiOyDixklmN0ARTCwsAbrnfgbxNjb60CrIITZkocMAcGoeUOPIFM
89jCWHvYPxxxeUgMBD3OVPsrYAG3Obch9xvesyD8SGyK44MegEZy4DK6tWV2bhze
quyvESsmYJUPydUbAgDki+iFhsb3kCvZ6e9owypQrZdCr9FxVZesDnO0MxjGcUcN
fR7xC0BV/Q+Y7Od/HnJQRrPOOXoEOnzWghU29vF0AzLgs7SOj+8QQvN1YLuEzoH+
7dEPLaBqo9v7QGK06EEV2dOzsaTIeYcOEPze6c+b/77Zyov/Xp3xaksbCUUhsv/F
MZPNZ3liyKP5HM18RAkSfvkP1n0w0X2tJOa0dp+Ilh0MVzZIBFzvGBL2KYMIEvtQ
MDDZgmUNjOiIb6w5AcfUHfwO23WJzJQHGwX+9mx2xuS5wdzygw/q/V8o5jcd8U4h
3wV/8KApGyCR2FiTI4PefzC31slOoAoJ0Sfglc2vR2zX4RGubTrAR/U6X6Ka2GVy
A0TGIXVESejEwq+ZK6giqdybogWqdgcDPmNVXqVFWVgUWXMKv6T0FAB6qrF0YdmU
m9PwKFD1Aq512IbWb+PQotMuPdn+odIaKltXn+vY3Nx9BmTL8xpHBEwXv4ujX1b1
UgOdal/2apsRWjz4s4WnAXwGjshU2XoEPSIEw6e2to7PUQM/0a6IZDR1FwFN1Yie
B1kKgovg8GKe5xAyJE5Fn6++ZzJmi6J7MNwCKUaOJJve31UB8jq9wNBDZ+df1JtP
F208S2tNXNz9BurOv8cWjg/8DiuMT8sMA+1XQfGOp3VBCcmrgotOI2vELl1W9IEu
vfRF+iF1Y8/1XbOnnBEbBYt14kEJqzdpIltzKn4/KlCb9PoYqhdzLcYVhybr4Mhb
r0l/NZHO6I+J2aAgIicucZGSSD4Qes3us8fBEDqurJkmJDCN3n7d2uVwytBcGvgn
wLwqqOjbEKOSxWRpvKZfKu/5msQvaVcAJUXOYeBIXZe+Y/wHDYtR1/9TiwGz6SsS
EmV7EtJ/nr1WeQfGGDJXxZtbcDeMdg/M7rD9c7t5UZWEpYutUUoSJBRlJF3X9Mo+
BUuNej8ZLqf5meIe3fxMhzkI7nucwBgcV4h+b8jGX2vWEFObG5ZfoT0TUtnQ1Fsq
KWwvTdwS9xprRn9lBHmxjCuxhlBSbJwo6mSKvxED2Y5UaTo27yaUvxxiKZb8RK3O
8+T1KPQWdWGQjw/NzFFIL4n7VSiGhAi+ewVeMvkwL2+hg+wt+gbIn0VK/YodiRAA
KJSgK81UpZ2jqLXp2eBCrz+LHNGJ6Yz4p1WKWqVZcghz5kGR0VKH2KIj4WuPguWr
d4llOc5r8enJrE2ELkqmYTBtgj6FRnK0gof9uBksu88HqMrAO65/hmdcpS0N1l6v
E4OgqCls22Nqh0zbssFo+09zP/YicwZv/2JeItPvRA9jflAWE7O75LXHi86Xp/nP
O13aTpPh509BbL80QHoi3Byq6Hy75j8pWuaAv/cAqrKL3ep+JxnVBrpmY9hJ7oP+
w+HrQfqMTnd9juQ7KC+VCEYmr1VX1PRFE8dihzdG9civvORP9HMnGZup+BjK9UQ7
C/4YT/Y9o+oVF82RaYOioSqKOcLrsQNHC1z7oT4R9RIxv7lkHggOhlO2Rfgam/sB
pqHrzcmScR5OGYgAk/o0U7gi6ca7EvvA4mw6e+dpW+xbUHkaHCg/ovzDKAN07UeN
K6dojrLo/cMQ2X7TPj2jaUn7i7iXG8Lva+UwcW/09ZFmn1eUv8IJNz07MQHOoAY9
GERP0ueg3rwNF7Le415A+sR/cpVcwswswzYV2029oqW99eqpK60PSPhpzAR7beu7
zHpWeed1qJABu77L/igoqya4REUwKR01g2gtxWjOF7RDZDBBeEwk3jwTyxbPRDS5
OFGLbVxMI62/GHXdtZehtoOrqRSSpmpqTd9iNvco+KdbSCc++8azKDPGkLlcTGAn
swcJOHIByF1JDFFyHCw4DaQBcNHSU5yvtCfU58zhmyVKRbDuusWCB7mBi1k/mz4p
ef+4PgDzFsiAqyEg3T25QNY9Njxszlny4T3ouzN48NVT+2nRHJmuih2owndb5CeE
8ZY7MozgnHJJdS5SxjEpr+GoQv3PUmW1CPdBkiktxfkhT095xw3sksSF4+XKQvIu
JWmosyNojmcMpxnz/A19IQt+l828JQqz7WTXlOyvAYx2xAZTXvOqdy7sr5VKBFfE
gMulfTn5idluhS5Iz5diIYmL7+MSo9bqs/tY/E7jAZhtDTO+pYt1wxGrqSuy9EIG
/DJ6fO4KRmZ19hS1hqrGMUN6urkJfKLK2YvIiN/d3f7b4y1yd3JUX+kop/KhYAu1
AedrnwrCLoM8/Jaw+Y526WG29y8YDQKpxf3pbUH09+Akd84tFIq+UFyATv7+Hs4y
xUmTKUYFaI8CdAf3gJTpAb2LPha6RXn+TAS3Pc/4lfZ+YFr8b1ARBPdOYcsOJdI3
uJnk1uFmlrJKzWlXYAlbuyRb76iglJ8qsQrev1l76xA9P/wWyYzOQpd+WHkCZLai
MEOZHfbi+7xusr/KHRejMQ7fpjoZt2U9WmzghuzymnvhUUTlQ/UYXn10XZxKbSXO
H2bzbjSg4EZF1kSVysyDylTJMXKrIAKOylUzGwD76lsds+0EDc11/WkIOg1J5ae5
/2ljU5Ocqt3AYYfcuIAwAEBZxPrZzo7BEUzi7pnyfowMBPqBdxXVGHwruRcLCkOJ
QKq035k0XuxGgS0aZNwTqZaAF1IkXnaqg17pfBl6pI86N8n1CTtCHpxQZXmqwQ+C
8Ra5DF9Xw9yfkU2z/uruOiN5Las0Bo9sJhHx5m8U5UzGN5bFyO+UTVKcG375TY7H
M6srDMa0eSnftXGR7ON3Zn92gNzdupG9PyUCyHh8ExajVHC/m98w3VkwcJuZ37Z7
wHaHsrasrAMHsVxh05eEGm9iHMYqCyyLbfGpLdY93RlaKVpRAUCGYYHyGdWbFbdJ
A+xJrdlQCg7XDgWgIgqzGUkTE4TvRdYkIzVw8dct8vQSiPfHQrfQV/1thhNARgII
lacxf4jgbBsz6+G1VkqT5neg7Wr2vhsdF9ARaYMJIdWABJ8kNfaeopUuA8EB5FVB
vPRB6V2d4nnvjkbFgzS5ng1BBgb1koWKn8HTINLBQ6ybnEWkoYrNgzPyTXBnRT9O
dZ6Gj9I6m5rCdZinHwNNvGelt5eKQJnjHvyjtMI1WkW32Yoh5n7otZnuZgZVI8/n
ld+gzGfF/fTBsxjz4GMFoO1f6KyYuq1PtmNeaqn0dRIJKdPeVilEUtBT1rdCNj51
F9drfxXsMr9Pqd5e/USY2pln9U0zmROg2SybOL9Ctf13QVsYDkZ9EmQAlfOZFgZ0
o9pqbzX26ag+CvIwXvtz3NbA6/+JUkQtT4IyLt/GFkjaImu2gbtZo5tXV4/Md5SD
4txAifW9YTtgFI7PK+ibBo8/QHmEJKDiNhO4fnVmXUnKQyIOMEbjaXy8JL5oIBSB
VFkWO+zTHi5jJT4WV/N8U53RGB+NLQY1IARKUn+LqgIru+Bpjv1/pBlgpTkHcOIW
wk5dZ/Abs+OofrXbTRp5cJQmfOz1T+NYksCa+KZXdYzxQhLL5ONPAxeQgdfLLvBn
TRKek1QkOJEouZRWmS4aYQhYwNVg0Hv4yxL66++lXU7DLPuG7cpiWVFa/AU3VJ5O
H7+NnzGnBL1aKRv/wqxiYsN5LpFGSbSoqEzrZmpGEx7MK9CT3MxctiMsV7fZ4/GA
ylp9r+Ml/U0CKSBqiuQtQ8982iJzQFSQNI842SXkGzAhqVRigfwxE+lPWxjo71tn
5oi7GNDpT1RSGDpp1PfrQyTg8kSZ1y+scWtOFU4df1mgJLMXJZBOHm//BXrYPrFy
1KaU4zkN81bY1Jo+VMtdXDpSdIdXqPh5meK2MSDc1lHIeo5R3yHXwm7YA8uiNQKt
3KZ998mIxc4wozG2pf9Eaq6ErLBBcYPSOdi2oZdkhbNd8Dy9rVH23nX9gBmPLUWh
KO3Su0Cc8KM0HKIJOLC1K2jUnBNKQGLCE/979URMxvWMUoS3HJ5j8B5onAMdyTn/
yV4H8Ds+l8eZpxmnT9g0eTAlVSFec5ko2vJbsZdboyceqf9V2KZ/tzfd0Xv+fKK2
ih02vWOM51VpfxDdDMBucVNlEGc+CKvprBdyEPu/vn6B/Go02aY364mVP8JmJ2xE
EGSy35V9GIqDAtwybRgZ0dWFU3V8++M1BJIgnj2QhACEdeHIbXXFNxl9URj2f+KU
5r/SBYEhpB2Zg01VomfpTOA9KnANqnb6VH80Hc77Mw7cxgZGolf0bq048SVHGVnA
HIY3X2e8e0mah4NKiZTHoSci2jBK9PLP7bqfexFbnKdwzTJ141KF/CLKz8r4SeMc
5JOFWjiIk68K+NFCBtiaAj+JsmoLOhCGH5D//DQhFy9cZ8/UNlv6C6QcGJvphm/1
DgkO9J6Ewhg+9LQ25r4cRkNgZuq++NeXoxJ4MeZBBK15G9HZ+CD/XWCjInSggQk7
iLLn4mZEvWoPJyIzH4La9sl8z7DvFwYv5D1OIuhnY5K15u4RPsgX/1KKuhzoYbXm
8LK8JzcVqPqIFAjRJufANxif1IRRTeK+o9AoP7jKn55r4cj1tMJHLaiOXGLPp9di
uz5knwjVytxdRR9+k+qyXReiJOzfs2LvjptYYciegsGlswa2xB22Hz1OD/1/IdS2
5eWNnLxRpSEd64Exp/hk4uhYV3jOmz2Ug0JkKLDU/P2/SVuHBAhEdX5uG+/Fd8s5
IXCWIhnw8nUGkIuyj6ydHaPW5TuqH79GiSCL1VvkDIUYMC/dgwsWlepHJ7/FoRLT
Hrouzj0jsFZqLiGr5Uom9wJ6XOXECeEakTVjeV2GS4yy07f8DejCyBkofxXWsgwA
VC3fdz28e/H2k8zG54E/n1P7bbDgDBZarAb1sxAbTKixJ+fzAX2+BXsx4NVrOctF
GcN/2TnqR95c9mqkQ5Bbwj8MFezdRL4UZhR5yfguLIKAfrZfvNW1FhNjc2yNJQk4
WchdG+0tnTN5za1+IE6BNkajpvzA6vHbfaj3ODBW0ztTg2WLbzxWfpIi9rkM9G70
trtjlr3VLOYPhUDHdRfW8k0xvRRIKLknWN9mR5VTG764TzPlP8ETzmeitPw1PR1Z
900Ebwa+FxzRUflYawPDUGabLNJdE+RZyGIti4ACbgciLMDhNzrUv0ocSv5aY6ZD
jlKo7Ro8eNEEn4cN06pXRCvEjDV3sh9Z2jLWX4DwVkK94GllQd2OSj3rm0cixtK0
XzG1G3ewqlfsOHuoyoFl1WTqPlcgmR96QIpQyyqwRYY07Mk0DdWAYdnSRgaNq0a4
qztf/DWoQzsUSztlhggjwEt994QXUmV5ejIsjFKWZ1yNnRZohyYC8/fb9GuB1tZc
yYrweq26C4gyv6mu60i3gVS8Xeqchk8E0D2Ien7YfJNovgi9Ryqn0WLzUKrIM7Aq
W/NY2Um8dDEfehBIienZaQuyFCyw6Z8vfuGwUd4UZ78C5o0LUnmngtY/m5d6vzRK
iXXrOgqwDLVtsN+BOkR2qGRJM91cuIwptWFK9nvl3gPZJmk1HQPsRTbGX+viv+EV
FAKTyveeBNhholBp9U7sKaCcEwHD1Oi79dC2kxHcgrAtqDjY0Y8FIlQ25gvGulo/
6eO2sEm3xFnvfyX9AiCu8zafSXk1lzFxdPrZIqeUyIVe6s+fcAK1KLqjADjt1oMG
U0JbI/INhKMSEJF7dwMJwRVWufmn+NoJAwJ+/Ov70yDoWXqe7yaoSyK2ZSDDHmkZ
IejQm81t+BJ3RuaP7jWtTxMJTNRFeHn8PDCBU/XGbBhW3l8sunWiqOj15hF4ewyg
UIfAHn5inoYTVUKn6OUfTguPf1/7Ia1nQmRql06FzhpN/0EVk72ub411iZUD6qCk
2uSCcbG5Dei1upSS+zWGW1cpDbROgquTIjedGgy1LBzSd0uUHaQdI/4LgZKhDM/7
yvcPHcOW0Png2YNK1eajw7a8wKCSs74MsfIOJsgP+aKTq4tYJnu147XixX9PP0Pp
l3XCXgNl3iI55LQ7rhRaj67lYEgBfgPDUanG55R/aXn7LfGj6ehpWMTtAP2C2pxq
pwsWnQCg/cZhTo1yuXnfdhHFQKQCqh+URdS+x8L1NNDDopJ6CcDaBmTMOlQav1EZ
etc61FL07K2c7IXoKC9qzA+zNSkxUctcCYNQewIFA0jStJ/gPAc2Vm0VuAj1yh6w
yVHLkcT1gYoW8dksHsUg3C743NISwriR6/CCVcbX1g0f6NfNMA2i8SUQq0l3ZpTX
vfJIWTMc5bS0koBgP858/rkBfN78SizhRlP5114fkVMF3iQvyjAbMqea4sCTlm4H
TodQ/GLeLo3rkupXoWJCXavf7ON2Z+e2iChJ22lnWcJ9aAEL+xzcztBQztE0VPk8
sPtG+Y+KkDuMDvYdum0TXOT1xKpj4cWbxgbR1aBGBbvUL1LGw3L01KUSNSVHMNzF
ccJv2PUIjblrMOteojHR7PYJ8c48UN5zUYQxIp4CKW4euQI64SNOqWJF221azIuH
gcZ8Umy6160RJSWOMzGss0QWtD2F8akbfksVtzrsvYtieJkp2xieJ/gY9gsInkaC
iWs/kGeDSVTMHwmepTKe0L2axvKe3JOnQS8XGuRtcQCvaIWEM49upf5mUpIByBQb
9zRPzZezb2rkcFnlHztkwdj0gvZxesH+Ve6iB3gG/+rd3O1Kd/WTHxtVgDi1EMr8
BMv7JoSbgbtUHK1rw4axmSFf+llrdX92zw2l23t+Xtfia39YMWnWVgf3sJanrZ23
8yxjCD8gNrpRAxOSkHtbmwWdyrkkp4XXf6hpFcxGSsO5VDw2TsguCKKJ7ke5eo6L
K33ZIkp4faLjJDNPCY3Sgm5y6TC0ytSg+a94EX/mhUFULZ7wfCkMMzIIH3vXkU07
nChPpSgtiCO3L5CdQU0jPjyN3tXT/xK+Mn3O4pPeys63MWwXYkV6ERV6I1/9nBJs
tOdPHCBGcQJnTUuiVPqzjnBvIFPxEW8ICuD7Vd8pSHtLTXsiIz+Le4sVkgahM/+W
5XZ0KiJtJvimkUfwsZU1VJIgeGN6sRu12QAsIv0NeLFHlitcPmu7mh3aeoo3TOPb
LIaUUrZDW+v21UxJzKf9b9KhChAx8YCwc9mWwNbHasMJyAc+xuNL1/qBlzcewfY7
tgbnk/fdSPXg/vCmvMMNbW94ayIhOhTqwlHWkOjfcwvjBvTKwlJ1BLRMQifnAPQk
uRsKUNJBv9KRlf9c52jWVHUiCt+AJ0JjTKOr5JU/zg26n+/5ggmsZziw60Ly4SJr
YQzWtJJJt5XEWnYFe/gSQYSTR1wkBzk4LeSFEpIBD6NOORynT2ru+XasBL5ZGYNa
Mj8UQH5jj6KuHR7Tzya6LzT0k0O4Gk618kqpSFiJvN8=
`pragma protect end_protected
