`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qz1KvTd1an+l8UFXeJ/Q9sUIqquf95eB0bNhEaUCIRNe3m/U1QtarnsjZCv8SKr8
4rA+B7RZQY5ySHssc1g1naS1DwqVCwo0coJS9NXJo3cBKurJMZ+GaQCk82OQlFdz
3oOfI8LomfmdHil78Nj/rNh+vvF6/hR9YrZcEVov3ro=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3312)
5tElGT2F5uR+4jYZgEQ7quPRS0wdHmeiMaLIpwtqYdDJHs60wEHy943MGHJ5Pc79
44KOV/qCr77u0Un/H+vjKQyDa9JXhDJQcnoIlsl3uPUjztg4mnfbOWbIVfJaAAYu
dvM23h+Vb/ScaAbLRcZ9NiOmfOOHCuuGGk13TsswG+OwCmpu0h4E37YR+lxi2yUT
tbkQV28Yx1IQ22SmLen3lJMfniZD7+oXKBFwA4Uwqe8w0CvUaziwD7jbqO5JPZn8
OvBVTCOpLFK2lt2KYC6p2f2sp0yCgh4nM7sUsJLa/d017Zs9Dimv/Wa+SUoKMQBT
0tUPw00OyG7CPS0yO5bwWiQD9CBNFSIn8P62IaN5QcGGmt4WMqclhCbkuV2DuwZP
d3DNtqotuEETW97bMHbSW7H32N6saiZqTgOeo9Kq6GLr2xtOXHVoFaLEIAnSn13H
p94m/CXEKvCZoqWsxL6nSQyx2HDCGFlUOwsPTGfFEqFSExnxeuF+vFZiTA3sBUxl
qELaErc07EAbZhJpsbTS4m0un2SPjfiCjh75FtHizZvfD0fv7vsBaxKsK4H/gny4
5LWxYQLFCSTmmxKkWWrY/pcCbCzW22Tf7e3Awv//riM3HSJmsYlnVpJaQ+PMrJ7y
FXYRvhybbXVOq5I0xJi4GYNR84mvlq06a4Ko3EzEm9Wjh63Jr99NQF2BQALIbsBE
wYGJfW5bCNNE9Jw+4qMqry0br8Fig4D3km+5Xdvcc3BHqqKhimhWuaaylYMuNqtV
qIC25punxMcj/vecBuFER4A8edmZTpxIi9B5cQl4la8vYmhh4O+Bui3/E/SITiTy
4dtyKabCGKL28JXLNq6T8qDEyrFkiNHRVmXI+2PUHDlMYRd3EUZTtKGAbRQM99ay
8s2trFFvYMHGqeEOcjuIt59G4pK2oeGp+3bONsZ5TpcAvsURQ1EpbAV0cMNqIgR3
SW2b7XHAt3O2ZLGhYFPrKp7xY8yeCn9Bzyg7tsun+dsAhEbu7Ljaab6BkD9K2aIJ
pWS8+nw95ulque8PavVWZxNsLWOEcmKAyA8tozKmPHP38NGHLaPFZy3BcreHElTg
v7/0QwAexs8SQiBoYjp3XyCkECX8CioRhD32qyoNnpYGRDY/OADeOIgFsHolRFHL
eutT9k3+XuBHAdFxNn4VzeXwj4YwJvu/fOU2fSmDtrhdE/YbU1+x5nPExFAh7iSI
z3cwcZIN8JS8dagKpjam3SrqqJ11j2z8UA+L1FF7AZdFDqsa9QzprWjHxNMyNxtX
sj3WVtG15rrup9BgGsiaw374UbRTXY81wY9HW3TqmVA/CgrydCALecqiE5Fc30d7
TgCTr9cSgOmoIPkPrR6WF0rNEHFhVK87BDUi0JXQSC7v10FiCxQagM6CBPGFL8sc
KRAh4FCrB+bIET5edhodEjnmiJZKgFduqFJN1eRGSO+CUFVkgIhl/wg3eH55AvKe
V8O2EL561eXvWVPXsnjt6tTUCI/3dgECQCXR0Fc/6qHo0KYL/Ey9v3Mw5Mgm6M8p
BLxr9nl0RUkInbesYhXEXlgKMepFPYEppeS44w7VgnwAqf5pxHwzqp/FrZz4JIX0
nocJ0f/siCLjy70ZYfe2D7IpqPBITD575DZ++A3oQCdey1t79pOuAaPX0rmO9I1h
xgCnsSh7afiIqjmmGOkPd8rQMhRXmRJJ4GUBU1yIeQIHBMKMQa1XkICz+j/57kX+
4dRKf23gup9cDCITNcOnFvyZEWfRqqxaXGw6TxNgkprgoTXyjZ99poESbgcHbADC
aZXUBKHeMlHaO9V6j6OFQYmZWznRZxcenQe3xVZdYTpEZjLOfcScpQ532ubOVrx8
wwHESlIv8YiRO5nyvLoPBeIHe1o9O+btb0Z7rS1j4wpvyn9C3ZSHj5/LxJqQwYBf
OmLC4BoBO9tToI14i/Xrz1qwSN4p9FTZS64zEWiRpx0cLjkIcuAOTe7rUpCQ41m8
Ooi5AkrMrdkUV/9JR01LDI50Kys89uGqj0PsfeD5y6FMwORs+c4BlcRLYKsP2Z8F
x5bGa6aWsIExS447QJ81kk6S13Vk3GndARNo0E47JoFFppA0iIFu7zGcRy09ggee
AXpj2/UlXM+z2HiZuN5bUknUQmsCMPxnurfdCEaBazTcJnNwSHne0BAp1+8Pqgqf
JSodgy42GE9ZpuLTfoty1/cFSJsNJrUx7pla3Oydu7oQkYmmm9owKnQUWQQ5ydH8
vI5RilMhdugNVHCy5BO7/xbfARTZqPX53kU6b1OmsdoZ17lgwrLJhMab2Zgu+HQy
XHh+/OXrjtjAr/3qLPxwn+yRUGp9uhWeEy1vz28z4DklyCdUn11p18YLWxv7LkbS
gmTsYj/J2HoZ+vmd5SFVNN6EdW9DgncfVQtjBGFWoq5qi8GnORIBHJsqnFkkGRkX
q8O73w3qn5d/xighmsnV+n6VPv2dwe8uZiC5Q9GJ2qHcW96gCvinIVAJWnBfF0rc
AmyUpCPeWJXUaQ0+ZaXWlVok6bbgIPBGdZj6Oxqu48NwKfd4/bP/fcuynvDv+NZ4
g8WmDgVIJpYW6IZO24o00hm1/0zapw0coWM/PU9C0wXJJybvx6OVELgyU55Ulnu0
PMVejDvxRSiICSmt/BlEWhrd3YGsO5OkXm37ggclMTEPYJkZe1d5yee439IVruN/
aI02qLz2XPT/W3qOy/5VpkA/IfpV95LenWJ8P0WkkXKulfi0bwsdId2AwLsYAUj9
Jw5HvSXiFPYmSv53qeMynEs2SRqCmFyAb3K3GYEotFDk1i21zXBL43Dx8wqRZSp9
Mubz6R1+zWKKysNk7TTvNEUp5/JCPY1mkt+znrxHHFHDP6vcf21ZxLouDIQlPJ+x
ipJJ413lRa0U+ICB9T4pD9oeIpF/ijnQaeqtwvPL06d5H6eS1R0fQJJ4GHGYSfle
H30zpm3eXJ7hLgShpjXfWTLeXSlUO4Dv+fE2AlE2r+4gUVJQnz63cn0eZ9RrohdV
u6CThYg+R6j2Q2nZAxD3rv9kkzJF6Tvc2x8KwegRhYtJ8L3AQIipJ1wuANBDUWGs
T/pE/2PBSO6E85T5LgEW1M2IoLaMDofrcvYmOaAADCz9CRjWwyGby7f7fdd66CI4
hK8YARUp6ZJgMJiJZH2yJ7j42xb+aiV6MlqALQswh+005+FHj5m7p8mxQUU3m1Ap
PUuT5Bw4BmtT4apJfnhXeKUA4/1xg7/EthcnmcnFVb8/NjhKIjhoHVlZgGVMDRUK
FkiLphtmF7jaBMpbrwDvHAa3UOj52moNmEaCsPDwY1TtmUmc3beHyeQGQAo7SbZ7
aAPHb1XtkYTQ50qwTs8nfFFbYRp0ppMDDRZsI0iWSP77rymjtfnv0lezV0yz/Fm7
/YmMyvGQF6qw3iPU9EDWkN+8Yfjt5lB69agCjX+1PDuebwi/ATTlXOW5Zn6iNjd0
QqaMdqVuOFJwd1Rp3IkjN8Ve9DrVL3F8GwbehZ+a879W4YJk5pY60wrooAXQ8Q3T
lQF/d7SoEhPzDNVo1mOGdvpCq8jIhaZeOzNYFlWqzm4v86K6WfoFliEckh71K5IS
sa/Dj2Z6w6eGxtCfmZ8B6UJjqCteFwo/+yXCQ8rY0t5u5GT8OVDLvfgJhYymJWvQ
KZ+TRZhSbUpJq+9BrxrnzprSCnIEPndeYJUdZ+YuvoWxh2BRLNdsI7Kn3NhMItBf
5GhVUFDes5Jqtdbqb5TgacZ1sVQNfeQ/FprACblD9x/FsuD1jB/XCL3YSauDJVey
Ns1UNXqJlwN8XXwnhEzpL89z++NbLZJbH50GaSbhc1StzFpGN/eOPlP95+JKBp8t
mLN8j3JsIXEIR/t5bC+bfNty8xfiTrBsbTMWHWEa0E/A0qU0t5baByGkf6n+mvM9
xRpAQZV9OyfMEL+4Z5m4MnbhxOSUETlIHYiHUD4h3fFylxrkhVYBMvD96LCoTw9H
1/3xFRxV+5rJeANJ7xAJ5ZKn3CrBQe/4wHKajyIy0ovqHvkF5T8js4Swiec7tcQT
DFazBxEeoT0VkxDN5EXcIOvt7NxnPm7Nw/BYLJs6Y8KvKQnti7cWPtqmyS6DU9bU
GULpz+rIT05DLDxb5OTO01vaIqgYhgfL+GVXqoTPl7TgbQJsuM/p4FqMWTXjgU5z
fbLPq4H9s+8XfSeDclmErXuC/XKysxeihlio/t/ALTdIjKSBoqkdMLvHBe86MykI
m6kMOD/lEfcMDxV8fObyI1wF2jNYg5/4yhF4qxeRygpc/WAUoFYwaJw5iSlPeQI+
Lq+qw0z16gQGez/2tPnm69ZbE7W3DIhAL37n5Zczjeu29LqSsjpgdxq3SH9IRAwk
iBAl20dEAYDpu/sg1qWLy63/R0pVv1F6KMRcpw7MN4fvyQX1NMbLYd90WkeZfvXO
`pragma protect end_protected
