`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e4gIIccnFX1ZuUk3rRb+PuBRyrZp0GVr5naUmFsJd8/+2m22yvYJpUDri2R/GO3O
xp+Hu/Qq6Zy4xQe+Yp+bXNXr2Brhu+i8U4UUjo0z9mJRRDhCuOMBIw1y4kUrL6ZX
fRbK5vhc6T8wUV5eXSRuw7sUKC9IilVWqn490wQxVoA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28208)
UA30ShWZSTI8ndpCbgXSphVp7U6IN8mKFJiEbVUCgf8nqFlm1y6Q8eVKIvTRF7gY
XiziVSSX9YCbLHdIMnvkCCIZMaF5rEt3WV6r2qCRXeFltoGTQSlTTGYJOTekTtCb
8dXh4ft47oO6QmkS+fuvNZpAzaK27yPb7CwnaCa/tjnRAj933mG5UgVxGGC8GgP+
KcUKRQHilNQiBAVLKSBcpGw9Gc3+mZ6p/nxjCDNq/OkFHJBu5FGFiCXwZ2umHhkL
SQUhXiBMyklwtO5NVQm0XFwSrbHK/xDXIWKM2vGxvbOjx1eKaJLsR11xXtSeTj2p
U+RHvzcWcSFR7cruQfk7bwKo0b2MRSCgMOanodG1vzjjRBIUPNJRfDQ8naaHmhq9
dSP1GNMEOHcc1lM4K61UW6pfNgWH4J4xOnIxy2HSfPgl8xobVXMq1yFvzP89Pd24
8TEuHXTXDu/e42RZdCVdhDYDj2CXmc1y77EyZx3H0EcaCS1TEILBsCbNxqchcPmy
gTH7P0npCsTO0Ts6km3zWfC67bXjcu7Gwa1UQ4UxC3sVcmqbe90Dh8fUXZaOzawA
3hM9L+EcIc+pILFpr9ko3+7TBFgYRlA02+8+vK1u1V7DhX/c4/lCgC5WARpSAme7
9zflQSs1Lfh7A0Moq4siukiR8MEsBtrEYEQPOMaoBVeiI9BE8Ohi0BSi7A8endhV
kxbNw/pHVEpWsRYUEKMIQsfaOCRaFmMCPvI7WD/c78Z5Vggldy35Wvz03eNvabNN
95B4RRelxpf4N7Cb+RxUWtPhF0UEOHXY0E5ypUW0UjbHhH9U/b/lXFia/Xy+RjW3
b9FpILzOiXFmYU4iymm1PZOD3Iqw0Tw75a6UNLjCk8BdKumQR3E9ENo/Md1INpHU
cDITf2pboPDsliyfV0DetN454izj6jcyjaupForRk8pnkxNhr85Swv7phTCjPYM0
IhNj70rI/8/HLr/eyI2rVg8lxEpIRuoo5O1TaRkt0rdvNW7ZmWOgYfZjvTPuHbZP
RGuoTbfI3hKd0InLDUxxhG2icw4c2IiRrZ74BebWMiO1TsC4ULX6HfJE/c3/8bRa
wl20xbLk7rmZC4n9viJ2kpibWYM8J749fQFVnizF39TRe4CkgZkG82phuUkmbKDU
txqESYePh6cebCly6uEwK5gtwIpkrLyjsV1fFW8SJ4reSV826zhVQdwssrhiKzDD
OGqGsoSm7JeqAw9ASpMCCzeR0qgGpHyWpnpsPlPhCd3gcgGVudBBZ8RgvvpSSjRR
dBHWzTe9XsJSR0Jq0x4u2lR7Ch7UJSoAm5OyTrAykg0ANKTemusYvsRlSfkGB4ub
0R7IP9GAG9pMdV55e9JJU8nisbSREgDDL82kjA5JkmmLc5ibxTyoU7BBeJQYBXM3
ORC3eJ/faTd3z79b6S25Z1vIlmY60xzjr74W4fX5KfROLjxcZoqIMpPXRNcjPBDZ
eouBfJK470Xq1O+TwsDIAdhpeNDsD5r0AwMR+khMkgEZKWracbwMLNuNPOfkFcp9
wgmrVjK2KRVHEMiKtSW8/G12SPKrOGwG6YNdaeeNXnkYSe0hIM9qtdM+ZiL4iOeX
3nrtZB0XEJtIJtRPKbj4Ff1SRYNHndBAP4P528mAqqThkb/JDIS7ndra1vKGaVXb
AGax8dHKS0+72bwhcvETtstR77w8rk/7ZXcz6+OsLId48noWPlBBWvHlEvrPKgQH
EUHpgkGf0LlRows0LqNPTlUdMmhIN8cJlTWDS4gMr/trJVa9/q5PYvR2YTQ9Yw+0
bcMRrCI7i5ivEeMd6QQtbyWYErQSz3NpOqBIl2EwyUTop/hTyuE9MTBoRsZXh5gV
nwSWTeY2HC4Sos4qeLWbCMY98558eZJQf9/+Xq33d1sw7lR/jv47pNpQZbmb4miQ
N+HJ0Hp3eFFNttbLCZkPm0unb/Zj0iurFH5u0qIuT+2lYXTNA5jQsptz15mZPQL7
fbt8dWsx1iEJZzKh2Xd9cM9/lYRiL0wJRE6i/pYvabOFSIo7fO4JCKCcvkz4Jfgn
KGZwDtbdQxW8p3HqaSfxrckYkJw6q1ImH0IFsjhbGQ7ACk9141W7fioo4K/lDrYp
/TNMlThirSo3l9XRlHKQVuQX4i3wkZfywIVJHRX/Qed7U+Shz9cZEXy4q+DJ9xNE
gAKirAsU+N/4f7Us8htOQ4Smo5DG35DMEHlvOg51BOxaXW/I0OGHE+vER2HNaC61
64F97zAbOODhj9MFJ7jvjRx135Z7YH6xNIj1J7iy3SlITpkiTwlVUaw9MyriZ24X
CHaXLkvN+VW905DCce95H+EvWhLqPg9tft1ngSp7TD8uGX5ZtAqbMzaPtenjrnOH
Nv97KR82m4my0lN4lzuv3iYgbphUnKMBmfegfyGnQ0T/TDo87IluaNx3hGtF20g9
+TmHEik9WUl1g6oIaNxRFceSkpJPZHWeTOGsvMtQwK/AZoAoiFutjnBu1WgVKIT7
9sT/fB8RMnhKndE2AaGzEJZhc40AwDvg1m9UvkGZI2mvtWq+vPzet2BI1s94wWyH
RJ66XLsYzmfjXVf50dg3ZWfPeo5QvTYOkpRmY52JEpQjblBRYsfw2OHAUymEvHNq
+0TyWsvPirKn1jy57o78SXovYQhKW0DRayIkOJIEuXEOmjMiL0qnhJrk2MPr+zQ9
b2djsOp9IxOMR8FCMPxeRyzSFeionQHqon1/aVOAFgURE62Jxefoxmr3F+q29klP
z8T7yYCuCPsUTgwDukhBLpywz50lIUvUETiVmfY/THtoa4RzL53EExMyUPxpl8Nr
UZDpo1YIMYxW7B3gQOukfC/vy/pKabK+Wrj5btngP9gPNnr/z7X2rTbh/Zk+00uH
YgsfSHuJmn+z0A31QOBpg9YaCh63CnIEoo3mvAIAc2XNAoiXn85ffpQSI+BzgRhd
wgqtXHIqfCpneyGUgi3nwQ5VCAuRRGGbcBysB5axthur58Lno+PiksMEA6AXyeNC
2tSxyXDoTrUYnU5zeSafSIzgRUI/gZ8sU1viq3w5iG7dpbprcMDIjW+TmI/1XPU3
ZlBzrLIoIue4iwZII+DpzuuTOtejDm3nlNI6FrjnnJKjKMBZC++kg/a/7fSiskGp
Ji3FgStdBqVSPUGllShyE7BPIhJLmfZNLlQ42Kl5etxEuSJAYgx7lJ8l6eqqW+bo
BDb4CanRh8X57TcHKe/1k2S06a8Lbyij/PQ83GoruKUHgCTQUNtTzoQST3EIXZ2L
Od3h9OhBSmFRam2vEkV8B7+I8f1b+JqQ3qncsxIHhIrEdCXtnyU795jlhvX+bBIy
DPMqNpnFOgz8EMsxCFFchLo07s5R8VOiLlh2ZWL11JDRuV86Rh7eS4Bbd2QfI//9
BYxKIjI6N1+ayTtSwp1hLO9kJrvC1X3KQUV8kFZZvENckT3XV8Ue6qCuqmEAiu6c
3JXitz87C5AZNeIzKZa5Ih4QLEUaCpyUTcUAiPZXAVtvhnacaT0Q+clKgH6LMYeo
QK+q0mrywamjx3qOfDxEpb+G5kv9k0NCewFSCRQaXaGsqzZPzveck3hsUX26EgGl
Drp04g0kbROYUQlp/e7hEZu1mDDpXaotQAIvoPcBXBh7eF5blWd+Z7UeiJE9W6CP
SL1rWjRnmcEnV43gQ1LnhjOOYO0TzsHFibat/IN4r52orxtFCE2P/Zm/PD0s0bY6
HfXShCjnDq5vQCmNTwec+MmOuh9mp4iIAmKLbmQNCaBBYfDz6/GNjH1K+Ne8uMP3
TYQ8XjUsg5+O633zTnhO4Tm6pB+gBiC7yOMmmNZaYmvk9XSf4yo3gsKfOttRcd93
6aZMKAZN8Qb9dPnnVLUA7t5NvlnEdw/pGDkkswDyMbylz0slcd81ADELShKlm39U
InkPfX4i5SiHqYiTZWR154shN8XxbzQg4EfXynuVIPAnmuI2awYChpEMfZ2b2K/3
DrcubQfwO5GLa9aBIsQlIb7xdWv+7l977eGzpKWXadDjUjmIL1BrR2L5XMcoZptK
dNSdSjHnxnkG8qo3qBXg9V3CV6mxKBwhOZmA9NTtzJeu4hvi7vOitFkLz2Irtrso
NcF8HS9K+gO02Y750JVwQFOQPW01rBapx2v+VHVeYwEC6iIG7jM7XM5ZIfgz8nGT
MPg+N5TtnLdjaU693IuSq3ci453Ck6tIgEc8MFicB0TCgqe8kWO/+mZAr/sMiaW4
ZiQWT+jTS28mCF1/F0zBej4P88Ac26KodOaJgaOJDcskLe+gQK3Hj9GDKLyxdlDC
Hzo0NMcmVkV4iHtvkCbbosSskUqjxB0AmCeRDtsSSJA16Rg6fQ9GVkHcUF5QVXK9
oal51q98fJRDf4vQs4+dbwifJTT+WJZB5ZIJHKxCEWlgyuNfXmSkdY3c7sPGJj+m
nh5eThw4LbLL8Bg9gjbXo9xqJBZBZvobTVxbDpHfsE9kgNy9KCl4vDgTu5hzLQMt
nL/TzJLmqZX501bFYbSEkFEdD0kZFSZbYvDOaUBV4njtNwILeliEoIZOABkc2Aux
2AH+Y6dA14dSL9GXCuhV+djbhnddQWQHR+qXkMOzdr2jSTbRx79HcQDsAEgYDaom
jrU5JC8km3N8C46s9JCsIjmr+Gqr2BzNeN+ILvn0Hot0p52VHmsjLD2Ef3IbujI3
FBJCB5CzeUNsJJKN34cNE//xudSn1758gQJSaMMsaYvloDEWlCFhDDKJ09fgUog8
fJqYe1bWt9XBXTtLgRZjFXF+9xJNkYBSI/NqYhD3TDY1zGNu0xb/JeN8ypShdFYt
VH8y12X7VC0syAi0bK/AgRcW8C8/YFxntIm39kWvnOsGzXdcifdP8NitFw1meEMk
9ioXk6B8j87OsCIXSYuSs3GiSlikI2hHVhaYncXyAFuHFdB6sp+9BAEtoxpXrQqF
LKcklTG/S7EThDrRSW3hKlsQw2iFPAZngBAbWgar5VCEVs+7t80Lqwj2jFxq7lcP
gMnWacOIQR42uSGswe/Jh4bWJi8umZRDtcNtMseigAkvIIHda4aHuPa51BkHEOiv
uqoQcSxJe02LYCHu1FW8L1xHx++gDXqMLBVxvp3INqQL5T2/+eKhQ5LX4MPt2q+p
txF/r6OXrpd8n8lEAlroOg8Mm1M5xCSBQZNFRNk56lM/V87TRToopRUnZ8gMtQv+
uhbNWi/sQHc339wpNd+nqq0R1cMI6oSW3jodxfzxU8lhbiPZmNG3THU+tNU4SDUH
owVz6pmzW24gZ8kM1V62DPE3XK2hAZIn06DfcOmcnQoMtz1ZcUJeY6eSGSdDSSFd
V1MuSN9MwbkLdMafqRdlwf5xrE0lJMwwtbUQCG2Qvnxo6rmIla9gIMQaF/wXoa0F
qR+X62jI86tuFNYPFQGFfPb1oT/Gb3C8p6uQ1DNqpB88OIvHhLVdRxsT4ByN4f6W
57Nemqdib1/e3x99W8cfvt0Bsc7C7IfGsLzridVRXKOCLFDlO9C5gzI5WsN9+jZu
G+xIMAXiCcymnTxXbUXUFKlYreIzrmrW1IquWCWagsY8IAYWtsRySs2uYBkg7IIH
EPTQGqm27KT6yHJvxWm99L7e/oMkbLVp4+GTCiJ8RD825mEN6TEqxTpefnz4u/sm
Ij0jSqI5hIOwTMEN244TS/1n0UrZwC99VgjFaoen1XMVUwxHKypc+KFk7DFLzz5O
GmndOFqtzTeGcGv5I2WyYBhoXZ2+txnQ10YNuOeQj6C8CfMtts2nFZpWCNqX/GxZ
iLUXODL0bQ38e8rIAGBxU78EmWhdxSvATUwpTjP4DenbD2gmJoQaLVy+SeDAMN23
y/kPeXLH1GVRLcXAeDdONnp0xYfepdFrxH0btZA758tFBR9NUq+1lHwb5oC3XIij
QCfKwjerCBSHAwv3B85uS26K6UtUXYEETRZ7HcE54gZ2GrbGSSkAGk6no+ugzuW2
DqC/sKMmy6uhCf4ZtvO564UysuxOcl4GeVpOJbGyp6aEb8AGubCwj4p4su9ij0Wl
OvzgAiK1pCMnEy3dDBeaHdjS+WEJK9QBy2YbEL7FBECHBU5+8QCtX75TtX7b15zW
tGYLa5JcHlJe+0ju5TnM1pE/13p8AhtEVT1sLFKsZZhYPzNLFtCRgzuU+k+zjUmw
4kOdM0IiZQWUFaLRhz/Nf/s0WbzQMujpZzX+5SIbG7HEeY7VYI9kuXjXqhxMg+PB
GokPH+Ltz7e4PNR7u0LfZ4mkaum/P4+uqKyXbLHi1ixzx6yUtNuBAiz2SVaFZP5G
xT2TZI6MrzhwmAFQlZZVJnZynS8Nh1qPRb6ZM7Espy+pn1HdYyWkVROZ1LODzhMn
42u7lWgpVT09zx95ZgUgSiE2p/hOTENsG8PSefr3TjWoiBkJhCS0UVH1WbiKu32g
a3KHrj5AJNgsA0ldP7EaBbfrq7iEdKxyUMOSXE83CobW7NlzgcxnDXgKMYn+brMH
+O/jjfJLxiSygio/zCGU2EIS7ua6qKAVi6CNjB8IBpSDd1KFim1wP7fQ++lbBqUR
PpS9caLJpySQAZsU98SD7qFWOqOGuQbMAGBXmvDSG/THFcKg9Vlzn/c3b3JN59O/
U0K3bHP0r7vNGySSEYbsbpquvvPsmIl94Bh+LCT+fnrrcueeT7EUdN3ak9KS2ePC
Wp2ieJshnYGQGPcSVQ9zmXNEG5nO5uBsbeEKuykmogRs4TG7uTlVgBfWYGzRwDaB
Gchx7jGlD+XEyyFf6JpA7IwI7HQ2UMzK8d2dd1QRLYCnDyD/LTOwqoy64d5o2MUO
m/nkWD0vceJpxMIIyVL/Z9nEADNK1kXE6wZodO3btl+kwvIomJ7+i8IrDYsMOdWv
1lEILUGY3EZO6cREO3Eaog374TzfFlYKetxhuaHP3TQvqBr90+UawZqMFs6XVXDM
PgBLrdG/8OTf0A0adT17cIDy3yLhidBoeTch9o3revrYjMZKrMeAiesqxYCizf7A
TvFnlfV0VUx3chKT61mjF2RbSYsNTSMxCTIxeKOMO4PB77Iwdh3CN6zB76nG3CKZ
4YDM8ms/ZhRvkU3SgDNtbN5Z0hVv5PTwj47O5oOwfy/ZqV+HH7MZkF9pWFI+qlio
Kd0BqJe5Y/8maCoKvtrZTWJ+7SJcNNKPVYx97JU+ZPxKrIeDhir6aY5xSnH/BG/K
8Cx5aUQS+Nwibrhw2t8ab2VPMXo43kvYWTNrt1Vs9CRb8MgVv0Efz/AHhy69ZU5/
AUmqmQkRkvWvRgfjmf6GAFBNMs7yZj1/i6/sXs9H5Z5JUeNIX6JqDaNleuYNaa1z
6+TEaRMW8qoz3NcGh4B9+JsLQ3GUU1JTZZ1E7gBU630SpG6PHTLIjSIXT8ynC0EI
ISac/NMsCxcwV1dzba6LXeUdRMwv2t/fjhtr7ujKFC8iPLm/vSuU+ND28BeEn0Xy
ebhnTtloU2jHNd2Ll3ostXB8V7srC1X10W/4Y6KYgU5xI4bhlPznYM2hBh/N6pBM
JzohKJv7oGhBtPpnj+/SuJG0vWUCJstH4nEphsDyRH00bDfIIQ0sFTjG6/DmoJgM
o9sSk+UAMHRBzS3vDG2P1ZDlvtvjJYiL5qBUyb5kVOQ4Ew2pch+dZ2SjOC1agu97
JRdjwESDCHmWkRPZQ/MdsFGcXIQyhrAuxV9UownE/tiyAAWWYbVd9FVNpU3Xzlcg
MT8wMUAX0nSyUQ65f2JTr2/WhSvoLWEORtUd5EIncq/WLZjVH21vP8blp6Da2e2z
HbpYn8vCkp4b6JJrifROSw30m61Ns98YiyTCRO7iQJvpe1z+dU8+OeHZxEuc3CUm
3mO1i0THUczuGX79nY5/oJahVceSHox2CO/MGK1QC5yw8p0OSTO3Q/Gw+M5D9bDn
kwGXKUIsiEkvdc6r6tJL4y2RCK52LXiz7gt2kMUkjNuhIhqjyguTkLRExG9UUc8c
w9ASj9J/b1h0d1PmkYIUg022pA/3+DTAoL1mmpT48+0S6RAKcI80KBgBwLRMEOAr
PbUfuMfZcJTIHYOUxF2JH1k6ZkLZFKO3sXfmA+pJfplCg93K8drFlwIvWx9D0O2D
gvObZmnkkaLl09cVs5mfccG+P1DtXtCYFrqBpI/RO3r+22nZvnTTaG06/M7nUzdX
ykm5dlAB4oQ5a4AGq9GFGu6hLYMSRU9BGx2Dlw/WAGGz8aMUGTsES3sKz3fwRXa6
o4iRA20jBhbLoElp2eernqZuJryh/AKzDW6lA1Ru890MVT5eVY24gDNMXKZF1odM
lxTFjSsWJzNF5a+TJWLNsHiN4Bre6AzmpVmo1zlOzm7dro+hFaBW8tWnIghJQB/u
RdnfmHUEZVi4tFdJGnqTMQ3rF568knubCwXasXtD0Ogdo3ZC1PnzjGU6XzjCUyiT
aOuMUGl6Orfw+XrfRJSUfu2OOkFXY8xwUOZ22qN1v2Hab0EMTFxW3rB9yvQ3gd7T
gmhM7ZO7cC8IVgYgZm4g+QCsoXIrAYbUutTmFHHD+U8eGop8XZP0/AmExFXtIbVe
ai93DpSDVtN1Drke7tDVET+CizwGgjd6m3LPHnOv/Y4Snvkj1nGrbDESkIvOn973
hqSbsIAdt3AiiJWZICdlax4jc+ndu9XptxmoZVpeDHjXLv9PkAQSjp1lLwE504l0
yI/zR92pm/pVQgi8SuoCb0Iws7lGyBje8fAnuJB9x26z5ekbPBN8WBnKvpZlvXDm
yJuTxPRENpGZA1ZlTVN1lscahIlvsvdhjVp3W/HCN3+hHxqaVYFOVQKDvP1AgCuU
1mIcWOQGxt/IjzlIdALZuDqQ5DTJrGphOPaiP1yWAUzh+yx/b66TeI552SF+taCx
Qt+4CQpwiypAv6abFjcmGKh5Ch3MEetwUJLA0DzHMCGHsR9CO6XeGjoD8G4DzDg6
t3znGsWJzQ8KNRj58cquOnWpnhev53PouCqt/H9OmQJPccHLlO8qrLBnp5Ybas15
9zP4YaJ2Tv3TMDyO8sBkVPvxPXEnSdOGrG8wA3N7q/6AcFwuq26/08gek6WH0dfP
HnT96ftIzjUB3UVOurUyuulFPfAd7ByFeiWfZ0BSZkL785dtdil+Bc7rhnj19grW
KowR298d1daOtf2Ehfnz9To5KzvuMW+V4hHEX2pKEHBV4ImIAZy7gGJxw3ZVWuzt
zsZqWVmGEQJq76nb982Ro4NWeo/GKI/lcTqflDA+GDtCgN54Og/FMMFjltDEDB7r
XPx0Bjv32he6i4lvqx4rbCQqNM8kIskfYsdfuiWG1c2dvFk+ZPwX4L5T53ShpV24
6KPxm8wRB3S4IC++PyN7fUXpxVgFoIbZU9BFRadfkpROsx3OFVXts52nOKrqg+Df
TTKyUMwmcBMu5A8cEe4mCdaIqs4yxdv/VaWGKWinFxMOyV0uaQh5b8nVB89e189P
7Y8tcxhx4ZT9AhV1exE9kifFdmfoSmPCGgidtBf8ByUUMHYhZqHN1YOQTU1dZV7F
WxBoUrdxybmaglCdzRcoRzSrCEp5U0XUCM425c4nH512AviXwriLXROP8/0L70oZ
JsntsRuKCgTV/1AF6HBn3Zqazi4iMCA1xU9wm90WqEtewKZbwvD/WbvvIljUqRf/
OCUgv9ZQTNyq4vZ4JwWlfmeWJmFghCd855e7YD0oLNW3AaoAjlF7AbBukXHnGf4R
pE4wrkLq8IL7e7pPTFlw7aJqX5wtJpZvF7o0z7++sNmxB4X9lCRNLjI7wlsox5Vs
mDUg5uc9fUmDpAI2XKcwwbGw0KbamXZEwjUflsHUhra7Ym3pfTUxLWba93lRqEwa
GF7ysbnQ63KE4K9yzlYtT48HD7392ctWKyKiWNrwjmlUAFfFU/+B2UYrrKQxo252
pLAbVb19YQOua2J4SGpGeG4As++tZO3qXoUUZC5A+wQU/vHFz2pWINHdy6SLozNc
iHd6PsaPp2Vp6DiZPAd0MbmEQD6vC9Ef3nDHKhDhJbnKwt/8KpLIatZFbEGiLA86
tbTX6ObobwNjl1zU8lkkFfFwVKn4hYqZ/oaqFeY/72/F4W11MykOgOTzinqkMb2Q
FkVvtaro5itrOQojnAJg+AMoFBAfborQjTRlxXIgI6vi5spD13Jo/04X5J6NyO+u
tBhd/M53mwrjd7A4X+DQV9uXd7oQaJw/qdODwfPImDZNcqIqGys06oDAW2CDaUhJ
F682ub/leygNLAx/XkjqTO8vfTyJDVjfq0QOiTzqhg3tUrdNOI+VpZGOS+ldMeAc
WbMLngN/mCMy7nPc7kNa2qtwtS0nApqfijRhw35z6VhnjZ3kA5Sj2lghjBMshCxd
61HDQB3q4XGjrC/kE9jbkWa6UQTn4BbAn76rOKpEXRCEiqYpWGhetY3HbQMr+EY/
tdAiqhOKQBt+CM6RfF4qsKKPHAcOOLaukVTmxDu0wRciUg1TE58DDwE/9wrPd13z
ide+IKcMI4wQLF8+ABtXvylE07DTX52EgyAEpTl17N0F9Zhq8aawGduLSzAcUkDU
Ovf3khgYalXGjZSpCtV0NGDoAZ3V+jtl/YhO4OehbQcmgXZnxaPgzxIIK3tX926H
L0OTQ1qri1KpqNaCiifEWSmTgKJP4CsGOUOAO+7M90gVtidOo15vGCKgQQ/h2MoT
bvNtZuMudN5v3GdHjcvVOmURSN5wSJuo3aW5SyncCRdHd6skZEJgOWFfaQp/sAWr
sm3dYl+6nvpWfsjpsv83lPWFiILs0FDXwd1xIyh1dTvEJmjRNOrEu0x3bEx9BMsb
rTiTcl5T7uq6mFasmwKLTX/bRK/Jx252xFL5BqJ0YGBTP2YPHi/CzCEWGs7n+DDw
ls2xk9zL6iKOjMSBhZ68v4oj2ZkmwPgecMmYq955/ILYFqaZFfcbitCPWRyTonBT
r/CCG5TcPYsA8LGvdkzyf9xAYSVdSjBiVBYjRy54OnVkYNdOAJOeB5uHgWxpfdSI
BGA6yqCWmXcDGpb3N4xMJ4NOlrPozkCuaG+VTv/UpPHzXkusP/PN1vnoU+rBbdlp
nkLuWOdK2JCN3RTrptmbbxQdJyAeRJ3HOrvyQuSgCqERU8trcMSAUKQVev2e84BN
mpPbqMi9Zd/46hh4HBudXaPQVApza9mTl3scvgs8Dv8TFoTcXJJM1F7nGrgNFnWb
fqQxiXObuiZavLIwfHbTi3FvnvPMQNWCqqH3vqod6G8arQDHZNcLj77XKI1v/h8/
Q0VuFN+SlkxvUm/bbSUZUm7m2AFi1TJ3TdwMgyFnEHTNxhRNjyWPjbcTTeN30t5q
XOFQrPDTcB/B6zg7U3fq24qiECYX1PqIiN5HMHH5JqScb09A7CXbB+OfSLilE+++
u0bOGF4Me5+vf6ajtaCJeBmYM2l4X+5ACFoL9tOTNLt9nXIy4UA8vGg5bnkMkWm0
4l1tXXHair0wkzZejKENXxjtQgjV0+dpSCzJNs9XRS36dfm8zLnXn+RHvvV7z9yv
F4Fo/DQqOX7B2F8mA9Q4m7lKI8d2+LdPFC4HrdIlmR8BfMofFTZ2vo7GU+nvsyyl
fqdcJ45ZwvFgbLjLMsVVipxFDIDBGWeXBF5RDTeG2r9L2dhDjIFNrvQqZ36pvFXw
eU0vCYLUmPgr4sVsMsBd4Pyxk+kNx1SrUPsMLGnjxzHlFf7edOCGHBPmQqS3yotI
WqxScmLnDxKwIZQHMXaJhi3n7yrviCNwYbwOzcg07GFnRmyqx+x3XK/DS+HtM2WO
8NtUq33hpTERfbAOcYvgKRN8mOh7Tcd/xlmVYBRlsYbU22OBIufBISDFtuGp53Fn
EVby7oQm82o2aDK4NTITOODso2D0Xgl+5uaFK2NhGU7H8jUtWfv6oOn6rsP/4zzx
CyGEE+9rgmaMfa8PBwLLP2PK/k4AVLrkciIP6CRs0Dhc9x2h0WQrTV9vf6gSqhNN
ay3uxLLVZh4F3OjVWvnAvHrBoKJwnUbifi1t3+8pwL+bHZI6MJemnfuOpG5XFMLL
KyYqKJstKIq1TJRiNt8sb8LROkh/GAQej0IBSKWlDWMJyHB4llEc760in1bHxQbe
ElRI3TteC9YNqrGL1Mc12f4I3V2rLxQEOfCxVbH80AMUd8V6hPEdONIhZGG51k1S
Veh1x7HZYQQeZsrm4fnpEOOLotXKBu0Ob8AO/dDUkmfQe0+fZrPJCVmCG2EjMDxc
s2ShV5woUPW3FefA/2ZONvNrKhccKADCnIWJc4qHwRVgYnVUIDOEwnQ6+YjK+b2F
TUn0sXx2zHtJWT4+ZhBUG6B00j4M97Y6jl//N75GIOeS9vh4yT6CfULCEf4ycrRG
52yGVLkDb+n1Cmo2ozX1acaHVkfQRRfPik/pCqp5Ch1FVTLvp5U+YM8tQ22ENHWc
vvoeKH8BW8/XdFRQe9D6X1GFIQCohSfB3sPG8VxaDAyh17th39aLb53oXUzN0Koo
i7wr/eRzWclNq79QVEVyTbY1fAJF9l0sQKYM/lljcZmeQuDeR8IkhsiJHDD+IhnK
gHGlDSo/JFKMMd1JX4Cxtsl9gLWTAkCwFKbgJJvprWmoeCkYYPOqQrz550mORVQP
s3DfC2kaRKyPVGRVCsfAFK6vGNO2W2ax8IEn+cBojQJ7oztueZldU7G6t0munByH
aJM4oTpLtLRRWbCLL1htqBiybcBsjDyPK+kzIGhdc/8cae+aHB2qdy3S0IRoDPY7
eN0Q77aYVs5hpUCyQBWZMkMxDEnNu+THrqINzAv+RHunSPX5HujBDVMe19rOy4kT
JpqURwRbtvSVJp8/Upq7C9A61wv80EzG3UJJlfW8Kd0wTGYC8Ek6rmrTh0lZFDXU
oOyd8hx8716zgkstZcRxUjILKQiZKCu2/B4yXrzEqVDNqYUKSHhrncJRHVCcv07W
+Q0QKMn6AzUSogdCXZ85nEHUWrJZpn1F47FZmvZIvkUfMSRDVXvyM+RMFM6BEhiZ
2dgL9+4w0SV4WDyqHHd5yUZbzzkK43D0HP00VgOZdkm7svWxI+vmowdXnI0j/nbh
rnk2y6Dm0yOX3Rn/JqzkGGsGEfCQhnDmC8KuFOFkfTrEKvTsb61cJ3QS+ynx9p0j
VP1GJ0/nHUCrBEXys9QcSLB7d4pzPrQpVsFhKDg0uvEsjDz2DB3sVJg5LkdvTnWH
r3yGyOOhl3ApmLQyMFr540NyUNGgDSHxjrjsVJEYgWiqq2Op7vCErstpu8bOrTny
/u2zSHXbmkFNqIgkL51WHIph3GyfuU3s21PaAmg7tsxjUoEtoJpSEW4yXsWoQfJC
HltJ1Q44CvQT0irK5Vz9CvBQJN7EWJ9gVzE4JmuWVpEPkcyIuz67SDd0hQ50f6dT
chEcKdnY5BPQOCOs4GKmuzF1H++4mrsbrbvtSeOQOyctwIng8r94JKnZiH8SOszK
wDBsgD1PdgcpbbeFche7tIalZg7jcyvqcdRiREZHsNeaBz2YZWk7C8D1aFpGQhi0
C30f0FGQSxJ3CyP2/2+ofUGwImZhPMT1TNLOhN0B+uM0y00V98F5LwzW+GVD4Mgc
EpnjHNWfU5BhWxjYDGq1Kaz7YsL4xsgwqedzWvworft7Trkaj0gl819gbdrse417
MTD+FvDQmbWrqQ/BEGcBOFep8iDn5vg+tjpKKoY+iFUzyO4+qYTGpLzDb8yMhb2G
daCdPtbk5v0wlvwgQZYoOdlgqW80EtzTF+KMB7xlTSe7Kt24ZlMrGx6B/upvgcRY
gL6xYras/15DmoufcOdxtKlddZ9EB6Fi0O6gXLZ8e6265TIA55qsQURwvnf54tT2
epdugzEWPwsEGxTWyhvvmLI5ZM7hhE9kGyQIHEu/hyaMgvOKTE8L2ffdANn/I6ze
R+5E0iOS6lE81+FTLUVJn6zDHNC7Cul4pIV8/u1vxuStgMBabLc5CrJVTy9Jiv8e
sMez/ba9qYXS0hh73xBhayWltICvTLO6grvF/8BYbN5iH9Twq7wlRHiOorHS4oG9
fUD0BugVWylEKyRvDJoinLTVO0goqxJwSmTN5JXNJK4fLAxGkle4N+u8VDxhBdjv
7Tzuff19fgQpl92FW/XmY0fm8lj7hl0F5vb/uSX/+4EmRXXB/xc/OzlLlLQ6hDut
5W3XgH7r7KTHPhVa/65uwT8DTG0pdaF9/XcGiPVSLBxiSVDca7fGpd7DWg0s0mRn
TyT2A4mAVDclL4uQQuadnCjecp4IkqFpff9mdIul2hCA7+fGQJKWK2EPeCRcwAAG
BObpNo7vuFq0CwQFivSXfh0vW5bhU1NLTq5UlMrjU1Bjix7bhHvXUYV4t5KxUE1T
gkYmqzpxjm8TzTSxDurihQx7kxTKDHkDnpMXpugf5H2YIZI2oQd4oG6ciwOBFgZz
SLsViBz4RQSaH8cHV7KqtqxVhhaTn7m/TqoeKnYsMWg1bQCmeeyhtI5fRiPEXuuK
gGh/cYs+ecW6S9my7x+O8VGCHcbjE6mZ7uVyv4BOWzA+Dt8e3OHiidmJGW7HZetI
YvAgFxbpugxYAATO9v0v0GZoKFfpmr+doaAqnG4iew4TBzpzvvB+n6GdO6xccfSo
AbDtt7oT1WqawBTjOoBMwtdAJSu9Y4R7+OFtHTv/IjlLsjaogcOHFesAivcMRS5B
23EJB7VRhyGdhQIR64vuatRZdul1+ULSTguU5RPSwHRITnp30BhXC4JA+qtFplVu
NEeFtxQstlv2+oL8fP4vSBgzHRdqy59wipcl5CC0Po3yJhg6keqidyVa2GhD0kZA
C0dKA8YQYrfbVW6c0s3b+74FJozLjWOBNYrOOPeey0bp4E4RWsrfT/XSR1j2iy24
d+GBstDcngm1G0xiCKKpi5FkqQVb6BFvLN67s22mAzDGxXndV+CNICFWLPJ4G9v3
GU877SFIiVg91D/ItIQWIGTP1JPehGD5e+3MJZ/x96UufS6VwXE+lNQqKxFuokHq
u2lfFnNozF7CD2+MIMnJApEfWQEVEjOqvrdMWWZRlvtu4s9IlzuhCgES2OmuTEm4
LDcuhgLljdcykZgrYa5qdoMwwJVfJddlZJ9t3UkRke4Nwy4xZcwVdKuvBSoQdkTK
xNMvMCxLzxdIIUXQxXx2QAnTpSVdeyDnxrFndBkv3OPokS81CJirU4pTwemBf8je
sLEqZ52glSeLfnfjKmBFnw3/CRALdUu0aWkG2XwnPA+jfItL9VxLYTc3ljjJ0KtA
ZlA6AaKL1RqeQnHDjiOGOAJq0h3/n9ukNnDhGRMAK8vTGnneZ63z8x6YAF97FvJG
QLe+dpxy6yHRKhz696KpJbMawf1F4yvyCwR31zd94c34wjHTuVeBrZtvLNejBwtj
rNtn/tuNNjyo6b9JqQ2dk9Uv5d2KnnFvJ0b9GPUj6HvUjCcFBQIbYX9ShfrNUnnl
auDYTCt+WVk1aBKPReuPsDQGhRyx0G6TAjR8v+nFIo2T7cLCE4Bk7JD6ar1wS3I3
Zh9r1iiGeLY6oqs4O+yc3kbRuGsc2R3WimJTOsV6OhV6L/2D7HwG38FAA3GGhlq6
WUXmtawrZ92k6QfsGRQqhKopVoPMP1RqzZHKHahNKD94t7q+wJ7JXhTMGzLEpZI/
7szugnesuEw9KbKSbTSwRHd6k/eSAMuaifB4mzVG7f6yT6WXAwqCdMaREf/RAUzM
iFRtw83n3mckjRUDvu/tUmOk7DQK9Bq7LRg9IaVONGXN0MZtNVd++m28BB2N0pJF
wGtPPa5zaB9/FAw8nfzvqmUiVd8VaUdC/ATZ13vQzui+7SYsNtAEECkXR2qtvnwj
LQJBwoF20fmah3aM8hLWUoX24RIAUFVD9Z6FlKduL7IHa+4R4mS4KbvEmdm6qQXV
fVywNOmPYV8TeAYKrlsCFAAC1YRvQXO4kjThOjxDRRI8HOm3TQtQREGqzoqVQSdb
5CxxOGOqb0FQEI+9adG68g1Vy7o97WaSynwE1pbE9tdqOMlMp5IaS2GH5j89WVwo
5Vl4sr6y8LSc+9gle2At9NKm9KownjFK4fSO8NKAb3pgkVWTxJcpZBOCXaEob4Bp
2O7c8P6mNWRyvDH4KuLIInlCdvSpzdWEDTCD2Ho0HaxNrsQ4+W4VpyP150Im9OKY
5cCHivOyyx150gWhQvDnohtwwOZkaal41h9D9bJ5bzRcKpgUpEuUHQT14AtB1hMd
FqsqlaORShxMZ7xH+GGHhJilmDMp8rOriSipoPNg9Vazrn7fJPRVrkkySXw/e/Eh
Sr3fcSoGwDMqMtYCcl9VZuHvxnSvAkzKhYDUdZMEmAOqZahFa9YsSlsGsU3E/T06
h6K3gP3wWGcMs35sXFWSva/YPiQYPyPs4ISkoxMDz0fh82GiRsq3lPT9pj/ftQj5
0iel9KvR3Kbg80ZXrKuqBIoljJYdXEsbUE2IT2zuin7lsIbRFHxqQxGQNq9MTULR
Vp//v7K5wCcs0bpirANUQiIvxpVGkp+A2GDwVdjdIEhq9gaUsqyqy15O1zIgvyCp
yT2ZKN6wG5ncKQWVQlaVBPpxTWrGvK3b1mzJRDxnYNADYfngWZQ1lIfyxoF4x36g
L0NTyQzK4A+Xj8E7EiNhCl850cPg08OVb73mERFm3MKq+ANrjYdDjIpyLePGYhrf
xgTPYKkFC5cS8xH/BtKHNh+KzF1WdAgA3JxswkNELg+iCYS9MFGrwbHZQJQz867+
LJJxHZ+k9ass4B2tcZxuwMO/3zN/trSeVLDE3HNIb8873BJsW3SfitpVYU1LBS/R
oWvOGwkd3nbqGU3vDGCMcKcJo5D11Az8hM0p8VOLbtDbqGu2P7AxH9fSdmPXNLgs
mIeY5lJAZKkAKEN0kQnxygvwz9MrvgtpKIqDURqxIfLKJ77aPnleNgxPiWpjdHkH
+tHgTeO90qyJErO9UvIy2gVIodngi72rby3ZSwwqJdcv5slzJXQm6KvwbwvJmIcW
eyEqIUkiT0+MeXEV8LEPhzJxpH4PLJBCK0BeVqjUKo/4McK+XscfzdX8ayaPdLn1
Qa8Lvz7WmWh/RoaDpKbgfoOOu5xr9dp5HYPRlPJOrRXFEI1jtU+hLQvMU7EtnhD2
gASBwUnymoTMyZ/xbzNOpKNbjo7m4Q50rsO/bkNWi3EPRMS0zSyzPSQNUYX1FE4Y
+g6HRKE1B7vAzXRqNAd0IWVtQ8x74l07Kf8FjgkzrLLd/Yo15qk5MES2/yY+GgPg
FFtRSutX94XinQyNmKNsDr/iYLoD+sIO0Ogl9k9zYAPzSxRyxIgdCOTGImxU7bxr
5JJZDHqXKI2cXTjxIV/943yO8Dh5rgO8CKIw+4n8STSjuCWfDiO6cDYVGFOQWSP0
YH2zj02QVYazjWFFYNvUOF++Lg/zBllv+p+xu9gem9kTbtxILHUCdYFRKUEy+nuI
Ai4hHDPGO+a5l2e3i7W1/JoDJz84HMwl0PQWYMU5TNDdJJsvIEmT8a/iofcV6x3o
YMD1GXbUjPn+dNGu5QVvwkyEfLrfIRzSDCHHhqc17qs6G/DZwk+mZJ7ASXwqWAZ9
TWYpwAcTiw0rXS7P+JsGa4ebV2QViThog+r0D0npm1/2DQGrgTurn0uiBQpm3Ule
LmtOQIbr1Yy7VNdmhAmcyy9XsGx6OlgUWuQ8BjrzjIQzg97tE/skDh3cP3a8aBat
5GESh6CZCZW55F35ys3G9PmxFjlHikUknWVuUGgFk+Vs0nOXUe99rI/WEpo1jw0o
nUCqh4QwMZFo+J562oW0dCNi/Qkvx3ICU7B9KK2vOFRPkNAOkTgQxBehEPNuwPg+
eevkEemes16jDD2/V6hOXtVSBKMGlTeHELCcSkv0pP23SMfUadEc9/4zJOQIcAqN
fGnmzP6Y/KUzX3ob6ukaV87rvJ/DUGBGAtWEB8GApKtGo7ciwHgbCxqLZipiZ/yD
lmI3bKrnP61nB8TlrQfSQMXJ6S7pZ6WfroPROwFLAroU0JObzjGXfZ7UxozZFM/J
LfcMv0xxEwuxs0i5Ih57A1FgSlhcuNlSxhoH1rA4kpMvX2JuKqhdhAgINTpafsCU
IMDYQSBSj+TIUmQHuB7F9e5vK8ibiUu2ZizyUQVyGg1yj2tIKfef3jvQ4+fda1Kn
1VomjOpel3yQf5qvxtNYxQrQwCLW3k04PCeXVAvbr2sp3/2Zirwu2gESI9miEvIh
wDbjRE33dRx3hXfimLlF1MBPl63FhFLotXuiUxQdSZqOuSMzndaPiBZWAKqGGki+
oTdb8A/3gKoCg8V07JYIDWiwPEPLGas7BKbuIlGxU1xRJ2OAUJZBAlo35ZuGbx1u
oUR/8GRLeWALzXoSjOTlL5Lg0q3d4ANg7wfnikmTrNXyNCQpY4hhhiDeHvpppfXY
IFAnfdSF+pW7N0cJk/nTLSFZ3fAlerYguwv5R+GNeCOPDqbljXRxoM60eXvsf7h1
wjL9ce6R7xkTU8XwZNKsYs2U89h4pUHd1W4wgE1LmmRbfTHo6l8EPrCtwFHWugDD
nuL4StGaECRBGTw0tmT/zOGsOnZTbQPXlFpkbq3TORdkVqAvBZ7JpC8JDMTimi8r
re9Ts8qqiO/Yn1BDg7uCDvlcmCTXCHD7sRtgK4Af+szalFYk3DLyy7zGfL3W24ZZ
1HBrIZZN7wA+flpbz0Cu8wks/sLx5DxNDRyxCykr+Ir7DeIZm4f9mGbrYLUeKq3x
5IVPctmrtOCVrTvjPX59yXBjN0FmHaNWKjnWx61m2hHsif8ERI9aOBR0sncLKhT4
BL4mGfik0B/VLCNmie8aHij3rc9tZTdl3gySE8u19x+xrx8dDPb2S2yX+ffdA9L/
wpKdrQWMh1kImwc7+7HYcYoZWvILxjlj17OTfl3gzLbYJTezoDQzghajtKqkYR9f
i5DXA2IV2O7c1SKun0ncvqwyzumlWsyzLZc27El5UfxC4RTk78C54tb4JCk326tH
RGLALG6WlN7rQsaSUqvbVkT3TaCKRWIQ8A8ynOV2EYYFpFZvJdmHujCUMZF2bjiL
6E0wOQhBnGDX3eHJrZc6GtW1RHolb8TtOsRVjmZDM08ONpnpJVh6QjZXGP1xn1EC
xvJIRI9oscKKei89DsoHaDY2ydsqLjjzBJ/Ox6lf8j3n3Urb6J/pgFpmcRALkRml
BDWD+wBgx7qM/IcckfKlyVnf0g7SP4I2OFOoV8jHXXGsc0JazSmWMLOYE3y8kWjO
sy+fgEEtiPs+0zjOxfQ9gBTEZ122zqQggJF3GqDFyIy01dB9ssFBur2TrAIS6PTh
IvYGVgH9GCVNaM+/Hqfpl5KeRPNvKEfmBKr13WjmBwg2kTV1XcaJSqCHRIklyUun
Y0tTiY0aKcH8+/nOou1T4t3ESTZiMPDojhgPdjyeEVfFaHYlZTUjea1hgsZMMB09
/8T4UM65RBwsMP5anuHZHjMkCvOG2Nxllfp6hTI6HOzlML/bl4KZTH5X5EWvqmBM
PACyJrklFGFuABIiwWbfrsPxUkg1DJ2s49kT4kOZ/hX2q926AuIgjQNJ0jUi6xHD
stwgbGpAx6hhzPWfDj/jEENxbw1hejVdcMuCgYb0rrSGUH4KsXMr5mfpuVdC0+6J
JqJiVVtU/i1kYdJuAA/WKGFaR8MVp/cLwomdDBBZdb6494UNU5gqJNcpZx9S3TOD
1w2SAI2vxkyk69AnyrPEmmzVGIkoU5izDAsDJAK2+W011rZtAMLTqMRLhZl1eh6F
6I1n/exFo5pRm4gY2cI1D4sMx6X+oR+6uYt5OcqN1+qorZAyb/dX06wk50Kfvhe7
wT/jff4bAd7SHfU9eNMzasZlPp17JjJ/gt1RgyE9LT/HbLakrPvJ1c7o7OSqaibA
5WL+4u2uI7QrDp1hPyX00o/UbrAhVXcbW5DHLZCm3RlgaNJ2UyjHmo7ZQU63JSPo
1hsMqkOMkPIOZA8Wavyz1j7FSTb1eXiCq+ly5GkgVX3dE9UUkr6khdLZJsvW7cKX
zbPWydIbX6oWZAus9dULiRRrrhICsFjJKRT/PqxTCa318WS49qdSmCfL6Jl9HPsi
bFspPuwtvusPhSVRonrkQtSEauLUCYCJEXHIoB8wQCT70/ZcfrpLBI1dDkERhuiN
L8kRk9wI5ivthe1lFck/xG5CJSUW8mvVem/lrzGSoD9B+48lAhJN1+67bXiL+hWb
iKH0wzhD90qPeH3uTFLPdQqCRbx0hPvcLQ+fTG9vBQNRGfCFElo4COFd5libjl35
tAJsPacMVPx5TXuUZGfbl44GS2lDu/OX8euEuKK7gV8LpqAsYGRieZqtxMy9leCQ
tyB8uFEeZVh9zp4fLEyrlD6hvzavRMI2g7k1Rp3uE+aYxYT2e4VW8pkInU9uK+J3
b/KyUUk2xGWkxy1xCZBagTD+ajD/S0cm9xyQQWUJrtu+do+GNBgNFZExBGdN3vF8
f3gh07D1+MjX0lCioqCwacNk8IldbOFcpXk9j4XurRPZ6f01in4btfsrwRAApnzM
8XVMzgqVj5RrCYMq+Cc3yJTCsXSc0VdRiWTbSvJ6tneUf+YdZOdJpkEG//6XMiuG
LCk/UXPUQQXVO4HkQlKcM9R6KV6/OgaNSJeqaDdStTfbZHCWrxru+IqCFrGBAFX9
Dl5RSwDhNe6/PPoXjCPogb4Z5llTKR3cvAWbBDCCPCa9GEgd68uHn/6TmnTd5xCa
kg+rEGMfhET1qYgvkNVih0OOmLym/ylEWaNxsKklAlqrjoPTg2UsyJ0oy/ppktp5
9uQPEpyBf8q7vn29RBo4FOjOmg6jyo209e4ZA8Y3hMZq2HU6vSWyjhd4hO7g+pAG
fX1W5g11ZgF67vaxa5SPKuHQLLlVuSs3oJAENdYKRFVkgErHVy4iJlNfVRi8Kewd
vfUG88QR9ENhIBI62PUFVeigAvhtQuhUMAMkCUDU23oGBy757CH+9ylrI6MRe8wm
GWGdoQl0hmlrtY78BNT0M/sgMNr26Z5s/jnO8yPdfrtcuQuqyywdZRL7c55C8UhE
1X6Ma9fWosceHzeLxjXoLJHUoNRcd4TX8gNkoovo6nv7B5I+lKYq/wD8ykvx/k4Z
dOLGTuGcBdJfQLdekmJwaZ/O0MWJq1HXLBD5KlXZJAcEclE1fcIK6Nxl7wNUAV5u
tDObvFtUzC79rAFkVinoRhAdMKu8TygamiWvOhY2EilvuN3/tPZ8p0v87AQ6Z3wV
KkVgxpprq0qsnn7WcL/TFtDwCA5VtCofXFtrRroPrqE6vOmGhcoctxKKLcXNgiDO
6OubURHqrnopYjiIppiBn2qan2hCl63hSWfJDYBEXGgAgb5T0OlP1UwIGvEgbj3m
3SwQHGzEc9At9HCa/qqrA/ECGJnNqaZ7CF7jyZp2kL+rDXHbZSMCZYcZup+Wlvzr
lLza7OMDUFQC5oJ5d589zsL9WHAIVGt2ob+M1sIE6sRxMcQoi5+dq1zfpKbk4DSi
VCynAwSRol/4kdv48EiBWqaLT3Xqe+aNdmDt2cUgfzD2cy/YANrvtd2EyGMIOUIl
0QBZ+7CueIBo+vbPfvPc4nAuACxgNUT5fEw5Zex8tsvZ4a/S3eLwXQwqoUQQyAq1
D7+sFF0vqozpZgI9+JUWqfiqXx2o8Y8wrdDqyA11Q+bgXxm8wDZuvMhIH2eGH+sI
AboPq/7TC/iewoCY1zu0STEufP+lwyNhJTDK9hKMQAtY7iX2i/7OyHcWwwpKwJrS
5fYsN0avWp+2ewSpSIn2phJ6kK5RUMG4YxrTJArVpdzNuQguTGIPg6X10ImJyda5
pZVvDJ1+h5Ebn+7XXqmZa3WgLBParOfft9iCEMwxMsSzwLlB54cOzPDV03trgHk9
XaV6SED8znj8DpdCbmkwklbEWxiMSzrklHQKmMnvajhNN0WT9gfay0xrn5MkwTTB
2CkjxpQ2a01If9Jx8djKcCIsHYrl8zBlMwOf5zdupG6wc5RQQ9t636+k1ZNpT4QB
FjQWheL73wE6CLn+gs3f5zBDyBUtY/1ksnr1YrbMDQQbVsH2zZt6GqV8gKzM8Vgc
+ya9sjEAsSVZ9y1L3vfJsuTf8pDxgXukK5Wd9w7yvczLSAZpLlxfsII31k0+jF79
tbKUarWKMkN19KxbfZL0BKjwMWOgn8kKE3ulGntL2lr3qVguiOZltbY0n264mlRN
GcXw3yJgPektAwpHHG+UzCq5rX690kioZLW92y4HL+yy/uHlAjXVJgZNc/6aL1m9
KcSO8VeGLgkSYTFyWb7w2J17PP3oJ0fxDvHVBaAjId84e7HBY/b0kvILxnt43l4X
fjwQAicFT/BLEt9IJOaMTPYq/F6qfR/eDryn9khgIz95cmUnPZUKpvSF7VqhkNfE
cLXd4RL2cYjEpSDm5NOoiexLjPgcdvPdxkBfBcHGEP23BqkILzPia3MewoDc5bYV
blwJFmEE7waS+SzUCkjf3vijNY2VdcjiDilmbHQbVGD6V9Rej4xy9hjbHUUpVpMz
Edozma89dHa2sSGhzcqExBIfyzN3idRfAsjavQxtajoQf6A8WoKlM/kqBzHg6ulC
naq+GST00bLQJR1lDf4YHkvH/tiHKaGSJ48CT5HCaackLPvQHrY1tAacfN1eJmmW
iXI2wP+ld3vh9EvldJHqVfLbatr4UgpnJp4y4bMMJAKxPJoyWV0C1NDilz7Jf45u
zl5vICYW8NR+df8LrbZfQBk0+uZ6Wmn8I06xL7FxMer31rolnYMTh4iktfyjBu4v
bVGCMZTssrnZP5RXHBho8w4uF+6x3JXoCHhOSexPRwfsmdQq5QVNhMsayYGhnHJN
AbzjePSFxRE+cW2R1VWvtYHfHAelX8OWJdTwwO/VSlApwELoOVP3nsgvWbDXgq9s
ROMmZGdjSD1MJOmHfNjGO/o4iuYB7hPAQmYhYlpExpJ0efVsLf+fpoot1F6gJxZC
2Yc1NW4KVJx46KP7uo+nDZwug/foS1ICKuKqkdYbWYmr8iETozOyflq5bClkZVmo
LdZLJytxwbtpnw1mIhxJ86h19HgpcbgyYB26hbnovqmmD7H/PXyMJVRjE+/+M9Q1
mxvojJWF2db0qcfkuRJX3xu6MdOjyVptswucosecjguRBbVnCGrwMVlYcz2+hyUX
HclU5BKHOKoiOLaaCd7GcOlaF059urL98hTJlNDBgTt+V1BUWvBwjVq0fTc6VdVt
hNdtiODoMyzy0zsEgFneR+MDnWZdFXXA9dqcZIUnmHJ2fD3R1L5gNzuSucukQCbu
w8rGXFR06Nbo62qe0qajqjFlfTgwR3vkbqlG5YXLQGShxPMJEuI0rWFP+XFchC+y
Z9qbY3Rkni7OpVjcawUbuBR6pvg110KkGUpeg53Z/Am1/6Zq5iOZAnpoRwfRaZZ+
QkRognxTeCCho+J5yvs6l7NenV2onPhHe145QnHynY5o8Ir1EYaBw9rPHFCUBx1n
nVdFwdfHeAZN1h/WntPNdFcpJZJnmphlPDTYlKHJ1PdzXpqJ6vEn61bxzqQNHhp8
B7s3Soaltn4tMBax0ekKXFq/8AHCf1co4DYfXfDYMqOBOMr8jiNi8KuoxWX/7d1Y
wOWneAVLN2SZgVugbsG3ZyJxuq5ZbFFcs0JMohxmd9pp3OUaInsKkDlqLNp3+pom
NqpdQfkS9daGSp/7EUfVlCsDdVQ7A47fQZivFdFxtziIWM14lmutDrKnWVPW0Tl4
uFbyCOw05i5urUHk4iqxbftt9wMw+3KK+0fkupzIRJRBRnZ2gY3esotGz4S8eKd7
CNQhAGL9C0+th3jsDCISU2PA9++sQtKQ3Vjx9FJ22G/yvzIvSUta3eqEZ8JNZJUn
c8AzYGX/3LBqucszkRAxLOPVmAm8tiHbT1B+HgHp7CjAW6DXAYZVIOV49f4Wf5ot
a7VgIOZ0sP9Xp5+nztNnSXbxuMNg5LZYDGxRFhR3DFtXwrfF9Z6H8npvO0UwnGu4
fQpCIZk4FagEgL2Me/5juaQoYQJUMuj8iu3yQ95VAKRxdIvzg3ZeGAST6AYmkkcZ
Py1JY3WFSYSiqOnQlWxg3sMK3wbT2LqHBc8777L5XLT3NggzlzplVtsn/9X9wCO1
ky/g4xQtH/q2kRwsA2hBnuaj1Y/krMpi1++AdroSj40zRwUENpuNpKrjFnIfP6Yx
SLQe/n/zJpDph4VRDI/YK9lcYYa6BLCeip2BWz6m0Ue++WeDAVfSCqsCsu0rkUVZ
flhC/cZoBSMm9w54SzZ/IaZpWySPsDvRxR4kh4vy65iqzNMa1IQUcgclptqF/Kjl
jezMOV1iFUZbJ+xvekmafezj7VKUIg6HMs1dKDedyfTsCZTCNG2prUX9YDFtybFD
cDvyfLbebSRzcTDysnRqzLMXnVEgxH1wM0lSg+bpVzM6+R87+tFFrdKYR3to9PgT
4ej2RXdqMoSZ+c5ls95fP8fh4Bn0ZXpeKK+yTne4eUC3f5zS/ORBtJ+2lwcQ5pkW
LgBTK5B6+9uphTPzaDOp7dzPfH6V15JaYWlPUY7Vjya2yp3Khz/ZsQx0blLxQxTu
SxqSq6cQVBaTH8qBqfnUMw8DCC0cML5KxDBTtY2o7khNBjeWYiL08wFJ9Iyy0VSL
Y12GzvPlREXc4Uh1tj/VX4PeSkTgQIV8pBwFxRejv+DnLLNgS/9uZD0WCeIkPQSV
2FxGOzkSSj7uSTFLxodYjBeFJU+Dt3bNSE2VRep9c2iKOa9p7kwRKUggC4CVUCsa
jh+w6ShF2s88SNUetn7FXJod910KDNOgFaWJGUD70OC0Mm0T8zlwTiwAuwBv9FZx
pQqpVDCrzVeHqROjz8/353lWciIshAvQ3LRMXGwZRQ90qlczkShwArfNtgPd2JHh
fU8I+i/Nq+qh8CAC3/qj7xgn4XiJUVi6zo8cv/OI+RMhUdXEgsFRuohXpy7yUGyJ
vp1I54s9fsmNYYdACao8eMnIX5DLLCkIMBxGkquvTdanhqVwaoHNDYJxwh072wgu
ChVxjAPNuCqOlFKS+0DoEjlJ8/R1XZT3Y4ki93/mw51mSTaUHsHCzcsUO3HXQOuy
Ha1Ytnm1idAh4l/K4P8vl4cf79XSZIBHigCdn6l8YraZLZ1kXtY1izG2XDgtfjdQ
Jmaqox+GpIgDLndUeagWjS5Q20jasanF3YbqwFQBSJ4tDhTuZaI/eFTJeWyvwQAs
jhreFLBrBS6WXGbJ9pFekA8y0IB+F9t2dBWDHi8+rkZ6D9T1w8XkGzieh2TWHYf7
+QEePDBubyh3ZcqkYJqSfrsazoXNPIScEGPx5GAY7TS4rSSaPjaQiq70Njxuudnu
MUwV41LsZDhH5tly4Eej5jNt7trh3KAZlXGP815q6xLq9gMIxi5Yw/YpfKBtQSF5
LZ9G349NDlv07nTN7kf0k0hNvsibJVuZ34imlgvcOwq5oGDt96P9HC1H7KReMXE3
W3q6zrshyxRQ54c54C3EaT++Ay2hU+zHh0bMz0KymnqXydeKrSZcxTQoGpIeIly1
Vwstdnuy+gcW/yX7TK+XDS941y1VDlDckTr5PdZdyXzffOx8ZQEdMwWuazOEYjhD
FyFRICZqIsrAOAqCPwOLUItxDpynFseTYUS4OK7dqlJIcxu1HVb2MPAPigZ8nxi2
9Rb2j5Lr4U6fLtRakjN6NdzfOYnJZM5Z38xoxyQnQ03+bwYaPzrYLbw8llb46y3t
ogrB62mmeT9VXfTmtmoF4wZJobybULfsJAFhI2KBRvwcGN3Kuekvxv7YStPSl5eI
qoIrylNJH0N/eQDoGpNSW4YnLqpBmhMhUx4VitthgHjSWNwl23CHb+KGnoOoXQh9
nPd095jg4rcq0yVRa6HMY2rkHVe94xADdC0buZy+W364S3Afm1CxNUxmtyEWsdgq
Q4kLfi/o3KOMfrNbMJHIFIZxN2QmXvqcVOFTrJVkHwDeRwfhqgvzniC/qGs9TAxx
dYNlQ/xkZKSdDjrhDfp9zSmfuhJQ73WzpyKLufQwp9ON1rgCZPPinJefk8FGiMhO
YxSRImcSY49kIaNY5StPX7q5XYyCApvMo9lMa6Tv362Rz6jbbEYPi6XtxOHRL+sD
MCdewzn5Jpf8sPFZTh0n1EPOSEoLYlMKFrpCbhwZG/te+kJxI8FuMmjVjTNJVWRZ
2X97lT3kpqZrlwxF3q76BRvm1hbu/Kc8D6dfrCKiT2J7nrpBPiC7aiYJaIm1wSOo
MLEeKtIlQ+rB5cGKNX+sDx0ugFcfEgxclZSdjlI5Gy9M9OvSv5yzIfLJPPlKvJ2n
YJKFqrb88xhP7o9YGQlM+yBk7dE2DuelGxeDnTLAi4IHjkp91VUy/OVboiaAWxOc
IXOgpIJ5HjrI6LRNStiz3MNHHrIXYeGUH/uNz2a2ukJEMqh3Im8NX0Bsf/8letBS
KoZiwoN1Y+BdiSoX4XQmAXlICl3HYqil6pt3kbaCFRbrsbZ7bUbUv35HoT23qwRI
lZBtvjnancMWB0OzshjoXvQJMSLlfN959/lYnweTTBW2ZGC4fBQ9VH6tf4koLRVI
k+5qfmaIIYiXi/0BZh7d9krfD0IdM+rEtZ6YGzHqSZ5f0ukd9DMDmsWFmnJefjB/
qZ072Y1x7hT5BuhPjTUs9Um1anKccArqF+hsYmb9/3VGgtwvS3Jqd/5yS4y/rBz5
u0atmXf83xh3BNM+UT561BZtDCDjdgRCzkv4gVoR5Q0CkQLZjVeYkvAwTVwseYwX
tvruUiJ3FPEgqJfI0wqsuxSFnNC70cZ/te7oLBOihgB8FdBmU/0HvNc4joEIp48p
G+GLqUQQ1f/EprWwgl+nOOfnEJ7Qio3I5vjIqraW1v1Cbelz8fJn0qo7qxfSHbpH
eo7V6PhNSc8aEyB6Vi4/NQb9AnJf4sSLyOCFbR2Pju0MQxnBGAIMJRP8hg2hO2O/
EmcEd97xhJ/L1ZK5BgwuFI3g1s2tM25lx/aNa9dA1zrTa/8KifDCSpZCUe8LMXf5
XPzJTT2ftOyKPsLS+32u1wxIsLsG/Fo0yotIplqJAWjRO/ZS97MH4Rl7SJrZObu+
TuY8BCxfvf2SVNf5tHEAh2mLk+Gv2t4ZUp+66Uj2sQHLNAOy+t7xxB8M4Y/bS5z8
aaKDxhYOJnyiSx1Iw897MuYw4mzzUQNHad0TGn5I39nQQ0brwf9iUYaQbDNyBk12
4PDhz7PWsgtGSmlc5TIXFVJgh+5seI2+aDesD4uIlMrgT1VjpZMzdJOxa4HcAP7J
FE0WmApvY4HVeYIzs9PLJp0464Ff5DYJ6EZdUkByrBvbwAelBle0l0CybxtGNA4j
cVw48IqA1CZk/xonqM0HflCaR/q3MztLr6SsG6Tox/c0G6Oqm/7XLJvk07EW8+eb
ZRzY7OnPMN0TftEl4uY/85ES6xAj5/znreSrc9lsp2Zufwnxlrprw0itN8iH2jvW
pNzOcuSdg2rx1/5FtfBBVdVZ+0ENFn454/awB1yHLo+2zCR9o3Cp6PyVN9bTNR/V
1f2N3VfSrNheY2C/y3awgwcqqvnY8V7R3eouLa+teNz/4HAozJFkJ3pQ0wYqXPVD
BM92u7sglmozqb93f/QEs8ePeY6iopHWgC+YN/OvJ0uPFTohm4rG6AVAAF6r7RY2
wiPJOZb8CqpujLFvBCGtuoVZcdz32+7dOIml8nBD6ZxQ7C+SjPLSQfhQPdg8jvsT
jNFmdA9f0fwPXHX+kPcd8uyDIEpDZvs2ugkSYUF3+ALM12seeHJ4XrPbPH4JaKRq
57r+2EWHnOYhdOjTe8NeojeQb1xgF3vQzQxzmt1N1K/uZFZmfZ6z4/hSEwk8t5Ps
b8eIVrUntF/im2/YqGASRSrmkZ/e/RfBCtipQYSflqctZROSVybyeIx0Fx9Gobk3
kf0RJCI1jR1LhrmVv4mqIlq0AOMZFJNydYXfHchL/6J9zuB2utMDV6KSCajakoGC
nCX7NzJE4S32/VmJbJDY6HC4HdBkZuVKl51myxszu50IDDIHMnf00PnXESsJy27y
KncB3CYTsMwxoAQVz2haqB8j/f8wle9s93GiLeUylN61seonjZBKQEOJ3gVYaHvL
JNGT/Q7+AspLN8G/gmKzpjH3aMYboXDdtoi4QvdjBJlF+lxQsaX0WDYP/t3DBsKC
Vpt02A9v1S0v9cOAG1kWuRlyoUepvrBxhwN4P5G6MJWr1uVC0LedV57gODSzwWge
GHaiHXzh8M7goSRsyVt1tJG1qFdFJFu+Ov6Uz+fXOLpJJK5bW04/7/1xfts3Wnsu
nlzPCD/6Vqqmu83nJ4yoZl57xhgE3dFPvJ64hO34dlhFFDt0G3hriEsY8ODtxkOq
v+qvwMifcMwBanjqfhK8uc1UnOd34VkwjJ5suTWNNOEZy/gAyVAc7+q+/AWtdboq
/EJFfEdA+0AzIy3u8zQbgaHQ0PYhhEiJ8RR3NkJhCjsQDzsY/Xjg5AIbv9t+94ri
Wqob75HT2J3pkU6wjwnsBoF2m6XyVU0FAMRbf9rcUzG3lT3QfbhpWhEGl1/gnRQv
8OtbNIUYhmsP2gVOxR9StTcK+DXHjroYYUwTzIyKJE6UKB0OZj4OjA5gOyMaPgfl
dif6h2zK80ZJ3+F5ApmvJBz9uqpsNdOwo09cULQodHvwJxWyBCMwSSNBNA+gZizT
JCCE5KOTblUqERGnnWKTxTjautZ4rE1XevrHF07VHBf4OZQXR3g3zrmMmjEfo46B
/u1wS4MeChnU+C2asFc0W3SDsPIsjfxWlC82288u737vgpxf8XmVHr612ys2BA9g
/b8jRazPyAx24VOB17Iaqc6UhszmiMMewXJVQF17w29a90yHCMFBHZ449ZYPf4gt
rm2Et6EFQvtdy4CGrdzq17+z9Dz8m2uSPCKTu21fYMQZmmFwx6qqQuAIbiV/9I2z
+XIKDLY/qhwgXMpZ5MrPpF14gbuH7JyfwMN+CaF7P1lStMuhAJV+Sg7UNmTCTgsZ
PM0vO6qdwHhomYqzkhmoBA6tpdzRbzuYbJveJogpOrzbb6CKplDe4sk8m9f9X8zq
pCFYSDd154SRhl9yAv7vi9a91r83WFDi/Umfp1UmZAZjftlzOjtzyPshleGTuNeF
+dMMSay2rmuCyciTrnSQVplrYTjbxRSxy7NzzvxDJ/e3VqLQJWgUj2K4hhBMiCGB
MtkGZSMpBBSnSY+bCaMHe/yFuiuTU16Dt/KG/21EXipWJXHFXoJi8jnRMR4QUs/J
86XmGvMteVR5ASHto3/vYiCzK0FqLAjCcY39o1qZgNk+h44MweYquXj81Rgv4Rgy
fL5id3reO8CRK7sS+KfjfbRG7bhqy4sQBw6IcBuFaLED0LEVvK1vvPFiXfVrToFr
LupTwdD2/Ji3NAtHR5jyLtYjfVbyNgQas5a4HTJfrX4cC6tcAlDBnnk4nHIgxF73
NiEJDFwfoonaLOL3n1MFUuDu15epLkV9+RHbwkWSFsoin6WCHCnDiFaR1U3S0q6W
ujit+Asxi04KaqNwmRxMzGqwbHVqOMI2KdSPWO0nKiQpeLJePsFLAcFiQ4hKYwp1
0PXWlveM1Ism2r+VVWbLwE59AqFOLYs4aXqNxP0Vifgyk1dTihSpcGlrVK9WrbX8
yUHLOmHzHlb96mEgTwi0SNDkT7Ki4pkrCtvuwOCWZTMH9nK654Mk6G1QDtjcXgbz
tFHWu3LNUPdfSGXpf1oeSm7S4vL787snp3dcHOD927AfuAvGmD1aLclQ7Py6Rryl
On5mQ72fuJrEenQP+82dyIHwmh6Ncgpo8QYNDKc+Qus/nQ6gMMwCX5bFPrBqtRA9
yBRhCuOmXgyH6iZkuTchwZaDCnHo5BTqCjdjgoLVHfYTl3I36XFyiG7rauf1B+vH
AweoBHCwh+BqqLfKGw9WREK+5Y4bfLrov67oG5XCKWM26B6b3sHZVsDQObu23rHm
Uc8sndyjPIYr1/chEslVktP4czZK/qns2Nj2u3zdz8luLvIeIi2kNDS4t8HKXAWo
VD6lj4LnBlwlPzsSkydWA9IbxKHHPutWMAPFLlRc+0sPKMsr1+AyGQG0Z8JobC61
5kUlxAfTqpsX49EB8BYxIc5aZ5HDh/1PNvHTvzCJe8umEdy2HZJR8Vxe9AweJAxl
BJpeMY7RW/nM9B8wzxQQM16xvSudTwULugszyiycv6j+67O7Qz/kHNbSUU+cE2gd
e3ElnFsk9XTvQcrTIjHFgalSkbiDFAk957WcTt7lvOA+K3qC73CaDZW6MMrBIWQE
fUqX64TjlonBeKVF5mCv59qPj3py9M6tGgU6nlYSnHhll5iki7oBQOAoHh7iIBvC
v1wrNClfvN9l4uGXaXEycuLee6EqrjX6XP8Ks81QAauw1r4Vw9ZT7pabIdcfnDUq
rInLkB649PBXaMOP9vzR2A0Ld5x989ZAAD0wOqWBuEQFaoHqpXaLOQXYaWQMsRuW
RAZ3KjgC20EuBwZeial7MivGwciRyNc3OtMcJRWFccr9I3rw5NvBayoVq2WmNHWA
89gh7irvesdrlprTF6p9jqOSLcu46nQj9un4jvwr0P76nstqWDCtqOknxjsohOwN
tP2x1mvx1z9L3Y4czpAK5oyXEKk6bx4RWuya1qNvbKFbFVCIuOdkJ8/mK7OljQAX
Z7BqP9SgdWEs9FQLaQdjm2MfV1cWTQ94IEzy356ox2LIIPwe0D5P9wW8dTG4KJOh
Gt4hUehSLsovrPdhB/IykL8dC8lw3W7ozXocQTk0YlR274Ivh4btc/yXWhkOSknK
T7/GZ8a4NxXL+J2Q2HOmv6fIxgmjZInANwp65pb5oKQpv19C84QS2uMC15a99im3
hLexS7YrB5od7NOYeqhVjCr91BI+OQgV/plrCkVRVUjL35tNgbtH640j4n1GK9dj
pU8Eigdlz66DnnuMW21tc6uU/7GkYnJR49d9T4+ubpLRVb9y2l9/dqADbwDwiBZy
01GYRwrhR9M/B0V2Iu316vE/srXOar2MnrodVVXMY3/+IBmt3CCbMbwVP7yBqljX
tNZiHe3DH0Tn7uBN8j+uId3tmEpMYpBu2g1436dR0XnA2yEEIZczZcfwf65MbSaz
/FH+NKIc/1OKqO611HKENDI7i6o3OUNfREr1G/XZs7CNKsQY3oI4ywIEDTuLUawO
BFwncZf/+rNeR7xFivh5MyK2G64g1chWMKpB4qwnvwTqTRbsxICmw7vmX6MsqDBs
XHr2oAftOaS6GXtOlCGmeJRw6LioUXrbV70+ObahfCyuJw67W8agnAa5DW0hVunZ
RPNqoR5kkhxEt2r0gKKqKXie7o7gD8Ai9RRTT01wX6m9V4WJjCa/DrBttFb5SQz3
JUPv4GJ5HFuBbyflIBuZpvhHBwXGEHVaxx5SLbe1sSCp68pgAOPhDv4Of0lMxjo9
2wI8NuSC6uSg3aoKVpodokjWtzCzCRygvUAxNeHlSBDWEI92lhF7DRW3GvCNg6vc
pCo2KOTguKzCNyoOoJtY7BPYJ0spX/gzJgD9nBiOZ82bBrhnhyFpPaNlQZ0koX67
Kl1x9FU60jIjHWCOm+c39ADoq/78Ft95y2QDvYEazY4duncdohZAs/0pahxGAFxE
ih1AXJ9TWn/GwiFjZQqqs13cECPghPbxsP4R9M7RVlCWqB+4+LmnbpJOO8S866EZ
NASmGZkz/XiieKHH8Dw4CA/yBF7an6TT57GjDD6hLlTbSloqSZbcASmoODwzhF/P
ENKxUoVVl2IViQff4a4r396aZ8zHpCSZBb4LN2w75k0M1dnz7hUt65IZqil+uCf1
AmfGlmtjBJSsm+RDbbxEEYVW2Em7RzL4JCBMQUImEw0UDe6py4wabV/OuP2at7ip
F+nuGYK/sKUozzeDnUo8p/vlIacHtdje0t+f2otMbLSJgzQsTk48rMF6B0VfxcaR
A44imGDY5yo78exktYGkc3swHIFV5ory52iJYBzKR2udzgrhkaphLYb6vpl2hRqx
dOV0MEjn9O/1qkJhpSqF6ljCKQdJbYv0hxmFs590b4CuB/hgjrcFq1+oL8eGDHt6
JhtHhbsGvH7qxOuwx4RWinm5xvo8SHSI396iS8z0YxK9mfHHBBoQiZZ/gxg673TY
5kE3y8CKNXb1p3nPaJo1Nikp3F1+aMKoHzqedQH2SDcbDoXg1uvrDirN+rJbNByp
8mdHz3Uh2lrDp0jetM6jWQ0UP48arw6SKUJAh7sdeCuOeTbNFFLDE5nVCV/Qpqxd
AKZ2hchYTXDVTVNMNSzBEvxYKqGtrpnAnKbyOunFoI6zCpYdxlXMZo+h1fgMxACG
c5IXZDddK8sGvGz7TKSgysQwoOlDupHGq/+libcW54Q5qRQD87BdhsWXCxYvNMap
OFceJKEuqcGxfTtGG6XIMV5DUC+S4WKIdPDIkwLeRpjCFEDeYkSPZAvafIgDetXy
O/gMZE2mQ0lj9Rsj7i/msb2NB2+aZXQLJrT3UnhbZyjXhV9Rwjy1WycJQ/XF3/37
P8VczmLQavUvKv6T2H/Zew5wFRAUP6+4a+NA6arOa0WMj0WLL9d07zmKGAUrAAkN
RnkCsbodfgtPcF2Uwd7yhAhIhDCLfIGRzLnELo0XBUo+36Wj+J1GAll72UQZVlX0
RH67QFZ+ayTWiPGuG2FMYruAWAXVUZFlrJaW7jVU7hKheZbYkRz166yXN+S0F5Dq
2yvxa/CQ+ItO1POdxQUR5MZVNwD3wFOIfXwWW4o7lg94GoDN74h2JpEaHaLSy3y1
t3fzQnZeDLtLjZSfiHLbvnWbWCB5qguK/U0wGzJ5dGB6/6GRbSlyN0lYNPq3ftb2
PMVW82YZDd2khEqbh8nFLyAU3kcP2tID6VhRXAGkw7i50ML5wOe9tSwbcKJjP/+C
ZBeehytgRv6LC0R8yzJfDfsyZJsr/Y6XSBqd3OUf4q5wNjQg/FOdHAzXCV6WOgMD
Sv4o2v8LYI5iLiabriI1bSC9NO6raT2m9qxIXiBj7X+BizZquWkNMGbCJC+s93Zq
5fzWM0tdSPBCw+viUvQxf3zcI0BPbxzUSbCcCHF1z5MKdObXHNEGeO1Ktb6eBgFb
addQjh0NBOHCucadrc8AXSkpkvOJC+PsbpdZtKsC0m0W2/eUYOUBHDd1+3PH2SBw
bwHgUieXsVtELIw6yoT1gLwCvmAYDPoBGhtd3OiiPqq61wict50GmM4iTDWtRCxi
TQCrCKeH0milZ0SdSlAYLFy0yST7YZkUaGr6rSx6onOFTmAS3LZPVPOqxrg9daiN
6AvnCVQvKMUj8u7UYRJxh7i6Cp+53GnJEOxbavNH7z9Sw6nzkImhMjb1T8KX3r1h
9E0GTZaEnLPy6SAWMPo/Xsn49lUpeb6z2eCuNg5srl7E9xAkjK48uW0cjI42oOr2
MjbikwmkWVQ77s6+KtHK9rWtigOj69NL1scZKAH8CI/uiLlsXfZf4F5ynQk+J6K9
FYnd0otPFRivYVmT/dN/iXbvRMmI0pGhqhx8McEjSSNlp2jHAumF+u3BuROFmKi9
lFMukspBBkKnjC1/6pLqBgpqMdWzRsFa30I00vI2el4AWWyf6RfqNCG9YOYsGU/s
piMpZofSSLwA4tm2/jTklwWamOLmdi9ICbQjLUqm/jkqJCsr4fHwQJMtir0H9mtj
mJwrQfq4WTLgO5BYpcLXYefgTn0OW2APqkO5xinVhnt8sEcDUwq7gYHIqgLOkR5w
mm57CA2c8UA//+f2jERSp+ee1PLSDxe2hqnIMH7q4WsidgyAH918p4Xv23zkd1ff
Q7ebDXzfmxjqqcN0U2AiGF96vbOFEL1IdreSJZeQfgb1Xqa0haPN1BCjeYDIvxjM
3UgOjcPctcwMFGAcCD/DfvrAgoyDiB6TDX6vuggluQVXrW4PmXMj5EcCIWkJVg0i
YMBm9zROhUxhQQZTvvxqlIRzYPqFPJWAlEXu2U0OBDwrtrA+k96qUmjUDDoL8Oye
U/bmN9Ro4GkaMV+Hwz+fafyTY/aQJ4qqUsrCfiqDT27laibk9/EaQw2nXMBUU0dm
e7kWOgEmpJnB+ayaAS0yCE3K7wu/yA6ZGEIXFKPwgaiq/zcqVVtWrMsxQVJQG96L
7igcLPNFOijBxwrOtrSQpNwQbZ1Y4LchKsn08jJ+D7COmpoiAVtg/mm2HA/1smYE
J5tfxwVZyW5CacU0BK5MBPjuOdzlBzQA653JpxtZXFgTucnLDe4on4lhDiTyXLOl
/LkmYmtiUU0XUp6zmdapptW+IXgXfMPibyHdSYa5BrC+8oa67dvogobkqX1N9zWk
KbKUCbqPhZyHJ5jkPRgN/F+TZAsipAGaTlELmmW/i+yQZ8DfarSJzViqOKtM2/xM
pf67EhP4Qo5oizPrzvIiXVkbL0fIgarS3HbQGBtyfcu3NwnVtI7u6dhzP0vy9OUa
FIFPS8qWDCveL6tXVrj7szJdytoK0dWj8xhMw/SXGykhL61f5Gb4XIfziwWF+Gou
VPGuBCag1g8x3YdcvOIWvGh4nSa8JRaogyrqfEo4fOmNnSZ5h8U3pYhX9XCMWXz1
qpJ/6tqNVSLCa2wW08Kxx+hxG9a1maskmQyU6IuFRlSX/ZbSfREzh2iW3QZMqFae
pbjaFgdY+MG5EIe/7nBaBZ+GNBXdaszg2Un2kXZHJsD8X/5gpJ8Q91xdp5D0dKao
TaCLph2VHEXH/PR/Eyqn7awlo5EvNemOfpkT9iEo96zBT86XrLby0qHUhMNb9zVn
sY/jgDI8BbFSlkoeZ1i3nCix3fOLq/TYkHBqyY9RXTAejcPeQR8jLWAIR3kKeEFj
/vwxbZW2jJx4QdNE5bladE+L90lZVF8h/ywRknsyt4yIFvWg/vUwyYukUYcbUiCW
s9rbAtWUVyuEqCbw8WDfsnRaocFhL+2iFppsyTVoQ24dhpM+VaTOeJPi1/gugNN4
rJaxzBSSJEh8hJGQ4ZUY98zPKHVzKqfMbFqG0A2LHlKD7IbM1Yw5jAKoAehKMUBr
+CQILBNPqPFha6bKsHWd562rVkJLCiIbN222sO96SGYWRGsFz4MiXEgcjohiuDTT
03qGZs+PTKHXp8Mw8Ce+lNNtxL5xnbgnB/H8p/MCPgmZoYVpCj6PiiveQKbRhhDn
c8fuLj/UtSPL1x8dGyriEzQm4GZhGrz0UbirZazDbCg9qD8aTl528TUxpbL8gqBe
1DFTZXKVHLSope4qF88WKkdRZxMqzjOgKNohRR/6LmsRHtuCYVzd0vjg49P3XVxe
mGmEMxxJZxL41De+K+rTwDE7H0NW3/YPYxPdSlTStKUmTU0pMSuLW+3IGoM0rQ3a
8Yz2shFwueSvbuWHpeRsxkSroE59KhCz1Q2DNSPwaegNuzhEdynxqgfStjrPThwm
K619jUdwAU2Qw9ksYj05+9aSEcjTyL07jQgwZRCll2CEA3YrMgWmNIujFonJSnTc
wzIx1zFi+KgRxYccs40s1PKKSroNcrkJn0pZNGtdMboN7u85I1ELfLhNp7s/PtVa
F2zfF7OVP9f/FGScSDrGDGckl3qH2HY815AckaKjStIEFLz2fc/ZVyqQHMaLgauS
ePvLprzJZ0PT0REfLlLMxdvfo28nAYC8NuvFGRmFvXoyEFovAqgpywhZHSatAED+
g4kDWI+ZbkDPyYXEzJ0V9QaINP/0MkvTMlrll6gEOljsvs/6CSt8C9HxZU4Y+gVX
xs4Brk+1FHSn4GkDVc02Ylu3v3Dz+mn/OAhmUyEPGdExeGM9q9HdPZjYBYN6YTqL
4HdfLMb/fMPLauWkkVg43rDHlqK1OWrQb1R/8UjqH4uYNapdZdXqCFj4LtMl4g4l
ooM7icmCpfKJCHHOr5fNJS/mjcq6eHt2Ua+y0Xsiy+q/xZv8JE+G+o1Cp4WqVM3+
HiNxRgBY0D7dVnWksUHPdxffXQ9ftjP7YN/izSJez9R0hPFLMFGAlJpdAXOPmTaO
xkuX01XIlJMZVBkmo2vyEUAHzDRhR1g0ym9GCUcmM8QIoqYV1QGHbSYDp6bnOssd
5uC+CCimDcSu/xMGqxC/PWWSG8mr7tbxudnJbGW2qBR5C9Rg14c7tgzFJJdqBpye
n/4chTBVsLXcsLkOOqUW9FYdQOKJiPZMwb2elqlnoZrTJ6FEzKTy2eEh9Htu0BL0
dnve7E2YLQmg9fBF/8uKdVcPzk49KY4593tM/Ovw8p1OmL5i9tlDyNLzGlMhG0/O
WCH92T1fngGB/TM2ERgA1KGg+mkmgO7rH3sZ9qwjzsdKX2nx8fLXbNzeDK4fELjJ
kTQmOzrzylXsTnyCVyBkcpftWGQSJEHGGrtlLrZqbttRMKeOEtZiDQ6xs41wnKvP
7QhQ4JUsrHpGk609zKFymEuKjzH2M7u7wLbRWExBguH/PdjdK/uYKp43f/zCXJFR
ekWUv49CiC/ivIKt3gXBY1yf3WA9xcN4Qu3O4TzNS4q3RZSI8N0dHR3Qjn8DUdQe
1W2lyehvid2sOVXfSLKgfg0aSUPBYLywTIc4i4+cbks2H9HWE8wGV8lFr24yyYQO
SJKuh5NXKhfGPDOciyV7rT252Zv+At4NGcOG+/p32dZsuHVaGSa9L0JVPUQD7F54
t0HJQEemNB8xGWpEke88K0AO9eiYXN+jQFB9Notq89M8zEs/v8BYAb3Is062VBQI
J2njXewZd4ZXR5D5q1H63ZUNVG1Pp1Xih0t/v+/r0t+QgPU1Hl3a4Yy6mSKU5BF4
/WRyFY2fiBn4XzSRJrEcUGe8PgK5HX5DeMPh5nMad3M0Ui4f2JCJFEVgWGQZBuLb
Kol3F2fWZhtXqZB5QYTDwr8UH0ZA4GMEt406k7RQqLYmsEYfbmSs0nlnajmdFeQS
zM2+tapGne66KHCVW3dejXsEBV6FGJdljbObzM1aeFoHBRn0V5GCOixC01aPLEu8
9RTzJX3qLgMfqzRIPdOxUzwb4+9scFW1TMx2LX1kw1cyvwO0XzFLG3ue3TUs0OHJ
vhIVteNrDvQ+KxlgYGNIDi9L6F2QeVrezoxHOT3C0UXyVoA1+MTByveOwcezH3Xx
kvmyBEA+WYdL+Qnmwoj9LvzOPfQwke5EZ+qxAizJ9CAia0lHciImoXwWg9Xyu6Xs
TxGGH0yc4pxh7qCZz5b9kwshZ4pA32TAMJOT7PH1eLmsnsVuKBKkJImXYAh2I4Iv
4IHxXTUtRBk7jXjA22FI29ejnX3qsTjsJZ4xnSJ8BtdTOie93b0AAAQdHp+DaJgL
NAmR02paJaLUQZqBSG59TuF6T+1TSQbjHhWMM9fIYPgWlvWPAcooOMpq2iuoqQ7K
O4VNOFueCnOOxTWRBK/lWDNjFk/IjBUZoQdh2v3Ups18DHzQOI4wMNq76PItMILj
9akr4cn1exnqyyy8oJOZSb46PqmXDFLe/1HT25ggKLxNI3a1a0uOZOaoUDEF3BUK
vvAIjFNQnepuTHR6zIjlSrYX6gYIlo/33JXrVUvKFdhj5iDOHqBVGI6GTcMnD6ME
EGckjD4hS557Qway++K+YOwznd0L3CL06MwvrwY7ZMkVxbwee9Gdmppxax+GznHQ
w6y6KC0PpsX5/7O2ASz+U/H4lsfRg6xEuRfaXs3Pp46+OMpfN71gwp02w+W/FVkp
qXmUFKI4ynOh+1+Vr+pB/tUVltG8H56Nnn74z4vFBPEWXXPdLpmJOxHtOj0feip6
Aqgr6F++r2rvwt4mdWykqC9m35fvLbpbsyKEvyIMvL4=
`pragma protect end_protected
