`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RsF6dNeGf7NB+AOD4l9+RZfBdp1wsqkwz6+V7hbpL3tmBRR3jXY52nu6tvw1ilXC
aSEO6vjJOvvvJG89OqiNXEh0a3UBKTLmfg9l2m0TLW36NF8rq5kfw0k+k438s6UZ
fMWwz6niz5uaUOspuWfjV/r2qrsyAJ6h89hRKmqyyTU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12432)
p8rWFwa22MNCocJrkke2mnxOMTpVerNfxPNuJFbhciPtwXhsrhHNRtzqsuo1FY6l
zSPq75gvdZAZ6n7/n4nHMXYgmqz6lZJe/pXRM0LVvTG5jRVSx0cCQkNlnMX6V+db
hMcFiKtj8vHK+idZG70wY5WSIBMkkBqcAsDzALMtA3nZQKQ8ZWzlmnPQiOfAlYwE
YWqX4/QIGQ9g/cnuUAKQlU6cZ2vEUQV8OmaoqE5GfyBR0qZMUhIEdFMPREprUQoo
M1bJaEdFJHEu83NNB58KogRIxGbwYBtYIDrtuf6OHSTXbXNjnW1BkMjLuOmAclRi
2Vl7I3vfGsYcNCQBQDkkWssIVC4xe4gaG/48bGN8wD41P8pVbwRCrUGBgT8Hmhyk
Y4utWV6n0YaG1P2sLdPoV5VYH5/a/NzF4uejo82Yb34uLBX+0no1Imy4cHV1Opsw
eo/OiSoM+0GAalc3AKMqZCeXR8H65o0rmchxDsJscfELqopwDk5n7UqZqmk4XJcj
zIPwpQy5Gd4b2Xc00AJsB4xdNgIhGF4ap1gWRcIRI2wQd1898wIZAmNJGp973S6R
JvLZxHBFiMWksAhMU/kW3p1oZqTQ4zuf2b0pf3T0wZ3iOHWJ5GpCZ4D/l7OdUrnX
STUNydvCrQTDoXpQHK0mLv/CcOiVbyFZYyki5wWpNpF9qcYJFlNaTnrLjHTPVALY
vSHR5exbPTpSFgpgKXyjsbqGHEKVGF0Qer/01rRQKwtnOeZOJStTXEOAydPCia+P
kovTLrlOrFQw6G/99szS3FRYK6qxaAjzpgL6fAGiW/KYafkfitGTnOJQeY7cSJUO
CkyIDaJqnsKnS43IFacIaSRqti677RIZziEWF3WsfCOgc6cDnH23aQlCEIc8mAWJ
cA0QC9ab0wk1XUdkUAUuSCp3+6XkFdIOrtzYc9daZfEBwvW9oIdGGRbMHZLZXaPV
/msomxB4tGLQa18xtGzsPEDu6QA+i2Cq5xOYqCxAXS3rZtEwuSTgIKOzvhtMrBVy
Ry4goWD1MpI5o70JLeJW0saIL38pF6mwg9dTIa79jpz/gfKFDvhGK02XX5ta0Qq0
R/8J921MsIhXctvie5mWNcOZoX8UtXFFSm5f5XKlScpgYIIPN3hijk9aYaM7QhCb
zLJOTQXLJ2EP9xHZPo7Ig4A922/somhzutb3QpHZCPGkxgrtZrLybW5kUV4KuJGp
H9RBwAcmlK4HLQbTqWpSdBuVc0zkV0sgILAnedAJ60CZif/PCi/ttU+I/X1RzpGt
VN2kTtoxonqdr2T46jOUHvoh+6+2P/pOQYyAEQMKQM2EjrYn/OSuQnBRQHOcBnEk
iN/WgPlF5ssERNAExtUkcj1qO6MI4lv3iF4yux7PJvo0noHgc3ZgBql/M7HTR74p
v7fz4ymgvexAuUJjrAKrER4QuoZW/nLvobxRwIxHHunamhlXFBOtUFqQLTd8ilmO
YXMFi1EwZOU15G7XSowwNxkgNRfJa2nuk+TP2XmMN2d/aeubVoicQ8bua3iWJjV8
vkPlSM8QCPuYflMuD0S7qqv0VXVRIJAQo5Ma2n0x5ttMiIP4nEGi+Ysin05ewCon
MOA8r9b/8PHNKo2EzuvR8KZIMqGMXBMnT4K6WLIGzKfTcfBjyQE04Xr/6RDzKp/D
jblk8OT3rjlccvoQTCJ2Inzygxj2Q1BHXgWAHqoegXkh/doRW0M7JUj00DKb5bQc
N+nuoVNd/1h2NFAy6NQ46fvtxtiVctREwsmphqLgeHOJZyrbp8vODc1YD7XsXuwG
IggU/WdIa+fwtWLzoXUVwWQ2LTzdFjwlLkOg+MGIPSsGhOpkkxiAJdMQZiTgaaEi
+UD2IZ35kz7BZlkRi86ibgSBmFFavuM18hceAaCFYKxvUQ908kKDkG6tb6V6OSRQ
9DWNac8f1zPdpn8BjDfFHiu4A5fnv82SBOClkg8m1McG+B5ukX7/8U0kC7YpZZdT
aiWwHb1Ew7D8BB35gDtvjDAcnpf3+cd3KD4jagxm66H7+1I/FRMZPUDxVJGG77nd
bZrKaW7zd/cII9qRZm7DQ6Ph6X8Pe+hxyGlbIkiLbeAOmyt4H8+pYAF5AzQb5Job
X/QZw5cilBamJ8VCGP9MDJ+/0w8Z3MElZBforJTRG3GPWdu1No6qhplJQB6XTb7y
SZnZkfy8naUMC2aBTj+8b4Qyvo0Q6LNViyD1mzQyvuQRPwIYiVvskWPDrPjAEZG8
31U4HLAY21wBk9yALklg8w7FXA6xUwDcHzqiwrWPiAOMGWeF6bcCZDereARxEFAk
VS/BMxO6yy1jSQGdEdtLEhyBT7EEaliT1hiPeVo1LGNTyTnyNxhoTYeTIjSnE1Ik
HBjxPjMsffTFkKOFmq/npvfNbmutbQYiCFdQxmNb1v/qA2iWkwqxfeBbvJ+bzPtA
LR9e8gRhjnjH0E8NQlKElwnnLkAhkmK6kYkKROT5BKR7EQ+wG2xM76/kI5NO7VDH
w5j0h5fvklG/ZaFJ0aZ00IHZevcfcoIjLMTIHThOWbYd3BFY0o8z8abUXfCYVyeF
imgY00+7mB/ZMXrdFnr2P5LXWLAM5E0DqPtcyvds/rVzHyI4ADxNyUqAyoTxTtXo
s6DwTjJ1PuAT8wkkvVD7O7BIvYz75crsjG2O675aYseYj7nsNAOcOnJkJkAIM6wx
iUT4C36KFxgzRuo7B4V6m/QMH6TvrX7RhLP9pd+BvKgLu3Wn38xFIQtLD6OxoC7r
akB9ON3ZPnpspRlnCAt9YBPbOSzufb9Ww/gCPnCqInYZXQtm7BmDSGXsR5zKOLv0
UIHM6DiDmXfUSxIOzIqB5mOBPZtb+bM+87lJ+/ER5kwj7gxTBYU1ZChNN0+5hXOo
BqD2ULbOg+JlgzJ2KfvVddeH4Fy4ehEzh2iT1BoEERsxqqHzYBGavq7xP6FLovwg
Vx/jHY5XbrARzybWQ6hLQer3HEgrGohzNkCEU4gyeYZFWlfwHgSTNvJPD8evThgV
vqGKVcjtVJmCSbkvoq7HN09CcQ1Jw5HLSIHOUWq2Ex+bnUiW3hvAbMhCku0bzB+G
jGe/gbjEz8sMlSBvV2CmH4D3YHeB90tzRONZ42qr7qv+jLWlmUOt9uRfSEGooZOO
5p1LvHXKhMFDlPBlI0YsHsPEHj053M2jT6F1VaOQD4VBrlDWDugXK7t58uBGCtIe
293qlnMOiS5D+qkLACo2VGNsFCV7EpDTVpW/lbLEp/JqV5L2T6giQLpVM/GXN8oO
pJmJqqAY6NhjYQMqsLi1Pl60aJNghtvkbVlF1NTy7O8S72wD0F/TAOwJn6ZkDN0L
e2HsxqPpBZ13PSNcEAm+NSQFNd6iQBhXdWQ0E6apo0MNi+7cTMNXabvfekN1DuQP
RRo8pRsT6al4lzyRgEZkmQIfM9NFVC2hiYfmlmJAgAqdQxMi7rctxQMfsqIlyFhi
jswgl7Jwbzy9+IBWnBr8HTnh/ItKSWfxdF6zZV5ViXB9zVCEEbhA7BzTqpMIerJ/
m8KMbUuLyXMiPGx5t+/j09n8Is6r8nqxd2MX6L7IXNQrYU4dsq0yXwzXero5sHWT
yYy6t3tTi/P2E3gSEd7GBOv6BnJLZ2ul4nLZtR1Vb7XEPgeoHS+3WN94cf8/fSlu
ycDNC52Zqep5235BHpHPmLaGOwQW+ZpuhmtiHOxoSTIFxpVbzCdzw7c+0r4Qk9tQ
omHWpg2kHT7KKDXKDpTLwKlq3HB40GoitBHe0XAKroRZbjwRLKt++h8HLxB0Vx0Z
hSxrzFfBf5/+kVy7zZnRU9v3krYLKKAGEyqVXjlrpDDh3FBG+zBDuRvTdQvxOp2B
gd8nmX3Jr4Jn9/dhttFzv5b8qM54yqvAmssNiJh665N7nIZ8J2eUcZdTnADcIEnm
n0quEJMWL+iPYuWsB0HbZ5uD7uKOyvGNwyLB9rp87DZEY0Qg2v5hWXaJqmQYpvRi
0A65CVIvC8yxGMnwMGRnbTABcjgH983ivKzAkz6602jzhknRg2I2VAnSJ269mbHD
aE/pswlc06rG5oa449wibwIdx9UapKzLztQcxlBVyfjZ/152Y6+YXyIy1mjUdDDj
0mRS+ZOleNpfVtN2bXxPVZv+UmVXTfNYODmwb+S7vVOW+3FpzrdbrRt6wFm+mT6r
lqzrV8vtqT38ApRC82jyacKspCIe/fxIBPTYRtsOvY6sBB4Nmmesr8Nr0w0+QyrN
3jTBi+gPWfd2oggJb5KP9ni+2fJlgqNQl1Uird4jZMhxAI/Oh6/6roT4FhSLRmlS
3FQr6TlEtns7o5RekXUZDD8AkEd6Fv8Lk0fwfLYyAU8wieBflfncd8slekR8wAsQ
htWspicyjxLN387qUbNLr45I8UcUsqw/z5bk5n07KXtSU4PD00ZizfZiVJC9MN3h
4apMaKjBzUw1RbDdRidPvDj5RTSNefyQbI42TD3rXayRw0FmsRwxlwa3fiyUZ5+y
qneWAfAq08IyORny7KFKc9WmpbKdd+fjDASEl/r1b4tyEj/od/K/NuE1F07S3b23
vmgee/dyVBJpA4KJip95S9yMVRZ5q8vEZun5mm40ky5hgLvT4v7hEnvYP+g24LEg
v0dd51RlhWf09udUnx5/Rs4oS4A3jQ32TjQnFkOlSGjg89vrRbxH4kS3Fegc5NAr
ylqqo91BRJw+cu9SrKL+et3h7SFZMfhfPysOu2eLRyNtfmEOmWR6BgYSgKjzs2k5
lX0j5QATFLhNhkTQ7VEXRoSie4tseqHPIqIFjNZaQtgbksGT9f9wZDORWV72LwOK
MDPYC0I5Zk8vpbJEkdYp850bit2sOscf9UNbJe3NC5FNsKgHcdL+6YhzIf+P/7Kj
zlGNEWx+Xi22rjvkrv2mNG5SsDDdPzCDrTN692DV0KMMOJiqTX8KlsAAydjzJ9kw
Sb2kOxDEe3kp0Iz4PJB0Z+DOd9oOTGhJNSg84sGnRHPmGLbbp1oHjuDRLSM+Wj7I
BlS/COPE2hu2xl5kXdwoIaWh0cWO9EbanZYhbMYunehHI3CnHEc+AQ4nt0vWJR2K
HfecKixtCpqex+kD/I61rv38VO4ZUOV72L64CBjJviowao7Cs2CJNvbekweDV671
VnW2dO+ZSrANw/5rvAxtLkNqxu/y7IaGWGHtopoLK9C0sSziEg7bHN63G/gT7Zth
WArQKn9r22GOuZxhQolVO/AyCEuXc9uw926rzBm+erEb0nJbyxiQbBK0loU3NkHK
tqdOAlXv8OoQeGfbt7XqocmwAh+ER/qMwW2h6XM9KHtWSvfPO3c2IyXnZ2OIU3y7
8pyatuJMNf/KPsXABVhGQy6hV+MXL9g5qEEV6zYR6Fhw3rXqQgxCnOIPOEscSIVT
jPt6c6qFvVNF7BJTpuAqYbLfLomfWH3kaEd6K4jo1IxDdF6t93+zllK5sWr0KHCV
0XYOvjev4UQ93fWjBkil5lLJ9MTdlG/0j6neK/7xtnsWKXo7G+SJ5BpPw37Yrlyj
tWB8RSrON/T5uiJssEmf3oKA7VPOOCL/xuTcHMiXdLMg5wzmB07RbD6d1cqrYTSx
xwcyORxAbuZkGMMk6Lj+pmUUSKBGFC1C7Pv4fj6MJ6f8tgx0c6B4RbMelCtOUVkl
grq/99E1TZwKLLpMoH2f+vIiRzZtNioXaSaV2wt4uHlcLA9txudepABxiI92aACz
wd2FYR6nwKQ1+tIBYpuetNuJLML3JzEgGMkj+2tC+Sq5xEF40CgumRnVXLFXVO3l
p2+I0sEKdHT6IuGNCnpX4CwXUBm4xlUoXd3E3xWjFzOc9X6jK551fRE0TVAt72uh
dltz5AO20rPUQGQPQBr3okI0FkmN2cWvLxDaAMByoCY1E+BYs7SfeBjjatQ5xkmH
CH+9RGatVhzCGK384WxBstX+7svZLv27n5WtMZr2EglOXmmujBHsP1CUHXDySbOY
Kuw7ZOeR5RSLlu/lK8isEQqCdw4+aSI5Wlt7rZ+/VLhEOq8Xo/g3PUyHuwcGBpn+
XP6WjRsB/12RHaxcKXUKRyjq9LnA8AKrL5QTez3ibGQeQwnew+Rdo3G1hg9kb3UO
iIunBT5Sn71zkMjVCDFIEAnnr0hfVrN3JIM2gelT5koIGgpKcZPe+x2sPxVjbEJx
P8d+HF1XVtmrheRq6rDiBas/4eG4W0sNmYS/kUsmKzdKVFI8vDA1oez7xLWKSQS7
9Na8epVAmUfJad7QhmKjbeHPZajIU4vb8jKcZikiz2n2cJID7s/1qHWgG6Srh/Zw
ogJ7NWKeD4Muf6mQXuD0NDfQXL6zlCSn0Tr3M/1AQiAbUAWhCmGrla0A24o7ju6s
Gn2c84dmDi+WUsVnLjOHATYFqpZ9D8pV2fLmBk8JwXZ1+Jluk3PzyUTnzGX3vzim
Tfotxyd1EGn/7naz0St4JnVU8qxfkk8CQJokyMIa9CI860HxAl7c3N2YKFQXVhzv
v9UZ1YYSFnovm61VRibxK3X0EXHTYM7z7oSFCLUdGpQJakjMxjscZ4iMKp8PH77p
zbpBFl8FrhmNLnI1bNPn+zaRwbe22eF85LvlZnJwP38b+uuLjcekkLqdlb0V76AY
NfervWC4zuvk0O5H84xvC2NXbfcNhW8Ecn5HX51qEbJuqfTBRP0+cNRdO9NpVoWA
evykgZDyz2ayc5A83opAwEwou2z6StGtayrCewf9eH/VCZOv0P5NJKFHpNDmn9HP
hYLWMDnzyC55UUY1URX7cnnpXG8xtgD1tbwcs8xOEH62EFaKCIyt47g715/TsDOS
cey4rMH0OUXbQG39ldGh9vSYRGTDegQICxSdUz+8PO6sLBrg900CSYY7dVM8kYpz
iGRmEroTNg8/lBfwDZoNo2BuNE64p2IHLGqgxYxKpIZ+eNNAsWx3TGeZDt2DUcT1
Wfd+w+9aLH7Y1Vscyo2RmMF+bHCmflpQWpoc44SO/YGz+cEvGgAl1KKh9aFg/5NH
9XbfgHlnjJfIu2w1J9OHOBWS6Qc+we8m/6+R3LWW42JgquST/6sd8wcoYcTnQAKf
r5q5phDnKTKY2X6cW8wJHVBoC9wZoTO98cVStbJsVlbOxYgwcqzetdXCf1XSFCy1
WSM0X2DzKEwxtkiqxAbgcXtuYz+He5mIFwMigkHll3GFjEFZlTNHdZ//Mfq3BuHr
jrHJbxefA0gSLdycmuTGYEBYZQlQ0VK5hPYAVKw51Fi9DkGz5P9ou1slcbbLKCtm
2VLXmKa8iPF+A3bVdFBdKoZSXq2jwZNxVxZ+vj5dR3M/ZkJwPcPjW8crBxthDY92
iyZ792g256FtKv39aIEEZHAsKusoDgpmj1dEVGLJnuMCvl85YO8LeaMXu5FwXmT6
WMy9jHbLoHKHd051YOAdj1Uc473qau8yagtfcCpX2h26CpbUjLh/U/zoVpAUBsug
G1V1xuqlrMZVgXVaO7Zm09sYK48B4zcwny+lf8Yc1C2XmH+rfJOWmOcoFdSdjMJq
3Z+1d/r+U0fBRZyrRtGUw2D8KDAMmdwBhiXHSW3PngyBIc3uJuc+T2UWNME8pCKU
EG3mPO3TCcF9fnFPEIFR/hRdfqe6M2z+lX8ic53EBHdvYM0E7oL6e1j1hjC8VC8Z
RD1c6AZoVb+veVya0zXq9nXx691SvMQ5MgUjFc/o4M+V342jwHBo81Fli31jxPt9
264ZHEQxJxWHZ+l/+TOdKoedTg/4nPOVVjrutfDaCN8chEx7Gh7HsKKs5rYm47qq
o5IoSq9ybkUFoXotakBk3+xxRD82V9ZI3QhB2vMPP2FIXtjp+E/N/z+bC7BnBq9p
CJSuyXvyNOimP3JaetYZmyAFQGbkJ3k4/nApZhLkh+bdKgg1QdGRnp3HcgpiWpUD
Pd7v2eHsWqLbnSicsXo8Be8/zOwqqYatfl5We0PopSk6spihuWeU4a0utro9ck3a
gDH5eaEn96VMWgSq7T10T1wOjWgTqnfHlJLu/AFaHYlJwtW8epC3JVb6pD6hu5H/
PXnPoa15OThzNZFbsdQ8XmKrZjfQnpvZix5QT2jvSPupknAcMMwI15R68X8S8mga
C6hVUnt5Px3FyuOxvolzLPhZ3eXblr+4f5qvCZ/1il6WMTEuF9tQt5z6aVXCURU9
eruQ8LtIDm8AQG+lgtYrWVVF8gFB/cf5AhrDdqwofzkhmPfZRB+8ExGlUOmo4HrV
An07rB41HZmXciyaJjGpJm0vJW7+u/apJKDGzTwa0FVHm7J0NGhgPV2mFY2I8Mlj
HgniqzUITVchkm5gczO5KqgJbb20Rt3AruMXRPDizSyPE456iv+FggJl3orJb8ue
Dc7Xr5SWhJskYgolCHqV75/mcp71BbY05ozBoTOXQzp6MxO5sMHOSV/qW/b6og59
1Zz9KRDXep/V+VY3H/fgTrHd2AX22GXgbubPbEle9SfkNKRyWNKwiUqycu9l19Wf
k97q6a0O7MlRI+CQR0r2rdKazOHTPHg1dR67tN/DT0x1Xr+uC8mR3Ryk8AQCDwTO
44eWNkHFClE5DrpI8Ey53N+1ur7cwLBqF5IWupeMV5cQghOHzhhQ7Ep62GrAfWml
C+amq0YdrOoMTT+1jxS9v/kaLSHbSyUDrIxOvfE8F8pHumAIxWuBeOUktrhmM0/o
lBLsijD+VyMiEYqbW/PV+BSv3pQgiTNSVhpV27VO2SMvfHQ6Bs6WtbfBawlnbn0X
b6O02J5ZsAjLmctCb9UktERC04xNb4lPfWezOseTbLVmNbYaFYemd7dpRHc6GjFQ
5rBP8ABIfbBbtgI4DShDZuAfbs4tagd+wMeIn6pxDPvY4EsZqLd5Yffznt+3GD2p
heU85S7G38QzTSiVbr0Z0MEwcmqHXJNjJwYjJi96tu+bzvpRcdTcDAXbbdR3c7lI
bwDHkTO0TK1DBRh61W3gcQN0wf+tCu4QTW8a3cN4c8Za7NRONKskaI8TdO497erZ
yC9ga7z7u2RFawF3zAUps7HDVUdBwqmp31E8heqBWFfGNR5ajKDeiAofE4JgOepD
GkWFmEZEB01+mch4sMXNnVoIe3eWkIHpsyBp61sz1cBGQ42r2SROdadbhD7GWkYH
C6XHjav3pVfZmAtI8xocoCf4IdcYnS/xr/rIyuE8H++SmGfbLQSTEZ7At1c0HCkR
59NKSopNCVbVQQq27OopRR5tqWNjaLPWWprUZjMjZknaTbc+YwyAV4DWRsXvp7F3
gmewhwWNUCbh8rVpq5tRECdRdlykCq1No4uD9ejdeg1Intv8EinoaJdDf8PTgL1S
YXhFl8efSsfJZAXdb4VKjWIhnhiWGJbfVAevIZICESul7FsTEZWdBwazpq3juWSg
w9+h9JPZWBa+NbaUI8WwBwAggbEFIxOeyvu5PB3JjftM4rZubyP1XHxy2ebDnBRN
48D5HvOJiU2GI8bQun0RUTlrD331bAbtyiOC1jPZjaOuH3O8IuGtqasTo/NrPprX
aagy6kbzcqgclqIFXXUU1i3bNcVTHqMrMmIZICc+4Z8sr0A6tvipzI190EsYaHCi
TcODCA1nwNo7VQvVlaWiEM6TUILjtd8oRgPuXXLPPhM5ZXk2mZeDk6pqAJRI2eRE
r95NUq0XbO8l9/ec7V+k+EJGzRY/8sZbL0lHLla3jCLdm/iQ5HG25U+MXd8fNUXP
iy+L2Uu+K0gRQa3F3PcnyItgsftO7ucyAUt42Bn52S3aEUx4cxQWALLsAfV5wvG0
5mKmSB0xFbxhNm0nDF4JkIgv6L0U65z5R0/sz0vrRK5nsAred5kG1FeRDBrRcSb9
ZdtUSRHX5z6YREmPhKATkW95LylFXQ8NGyqullrug2IwcpNmsYbzM4G6/SR2rFR5
tHFp0PWSLVXAlONL46kK7RVtWDz3EAlHq0zR3g0hyEJqXg+1gUZlhwwB3AlVsUZY
qABrU1IoJgn1Vy1k30w7ZM7+9cX8eA8oJEbQRcD58TplZuP4y64gPo7MDXuQlxFk
CKw09pFOqT88vu0ci+Zpq79n399rfARe3cZodmt7c9fEb8l5AiLvdzVjfO+hfFbV
rQc7UcAakACYlldg5NGGJGWayki604BvsFVTZMl3Eg8++0/A/kXThHL+rGe1n/Nr
K1HGIML7Gqa7+/rrirLy1BXZmQFkXX1LWCHuPDWas/M4AJaCKDwQCw2kEh9Is7Ox
Y+fPS2ZcapxSoOTouR2HaZOQYMULbQy3id8lF8D2S/nmAeZMwBkAD1fvt2uxxwqb
J2fRk7dCDVzDZb2XYsv8tLLjGMT745BBpYEI9u4x9kg2L1Hk93vGk3X8MXFdoJ3p
TQrKC+G+qD+CWh6oe7OtIYCd2F9U75NMDPxA9gGAnzUeids+YHZ8KjmA+4NdUuqC
fkZbXwyqj+qy6+xmptutLOeEMawolkWK6ZWxZJJWtrxY+1Y8uqFjaNxe4jumVpAv
7ZXFt2+PRuMdcC7QlInEdI/CcNIbXf5+AWmsXbOk4w7huf3GfykUpeDs9sikyCQo
PO17pRKGrvzAHTTgV4UugKy+IYNhREZEdTdNPBvMh630xQiZPiJiJboI/4gWbygw
z+0ERcR/5lrWP7GiSbcWE1qlJLIzkpNu98DKS7qTtuGoWYd2gHohmQBu/0G8qqJ0
OF7aOX40RlGwH35oEQkUmQs14CmUbqBim1ZZ36vVi9Tf1AVOb7IcO/ibPl8h7wTS
+fWBM0AIquuR3L8WVVwFyLW/9Jmoi77RA73u4wzevpnJH6OTyGL+rqjUV+HJNyg3
QjzCfNP3reGNuzKojXhP2kYLee1ef+G6QN8HmvSOM+4c3e7T7rnfzzpPW0HZiMrZ
O87po76mXo2jmfRzWw8wr8bQ5jrZcfMiXyNkBeuTHqA7XZ+pSlOQkwSXPxlMRdu/
lVtA9jwrZYiFYKvV1HdHqtncc/1rro1Z8KtIpddTc7eDnuSC6lZrBPiU01NWYqjs
91n1z3H2bxTSmo+S0yEW9bDxSBh2RtEI6+93Js+zKKvCGlNSo8jcZuwNdakV295f
hB9Iz61MI91+YMA27LkaeErwak5zEUgOH9L1AwTbocd3H/so/gl7EJ+WrlNfTfEX
nLoHbIFFqGtcR2Sys6DHFuvzVpLaW3P1MJpAhL+TbEvfM0F3dRmjgKzaPOPvxUZw
Ekjstmh0w7bQD/MPa7TGIndv+fXlqCv6+7VdvvESSIzUV7qilomfayf5G/7GAXVO
nuAWswBpjhwECVc8mV6HSTj0zrZsY8GLMmIuZL5PJdq13DFZKKG4coCm5WaKCa4Z
C4gy6/aoOaLlzu3lyBfL5M+AnxsXmxX6ZvDdoBpkv7k2t/rvqhcRAFvqsfNjLfDV
T7iysLq3m9YYHk1jjPlyOPU/LFl7LKAN/DvK+NmHbdokNJgl7bYNogRmc9l5XRhA
gyreOXLlwXscyMzbyWnq5hxp0wutw6KA+IhM+hn/kHliBnifwG5LfvH8pOEJQETg
3DoQI1xhX6qAQ5939i3EAirL/ILduVMrENV24x/OfsezD5hW6XzCEce8Jf4JgKbm
LgERpyHS2p1H5MYSzk7HsTkc4rP/ZCJM/IBwugDaGicPWwCUuNYVjFOnIvXaR90b
0j+vX5YPmDdqbLbxZl8OMj5RlpAyS9Or2O6/sYJDTo9GC15kn+9iuSzk4pA9atG3
rAzSqgJgOAUP8QxPYWKx3Htmdp/ejph0zWAociUoNb3b7GD4jt3P986iA+eCRcEg
PnEr6DVYl0WiXS1709d0lYJAI580mWAFoaL6FCWdCzIaS14P++TEj2C7HQD+WJcc
hnNBTFgpyDHS1NumhdhNVIS6fmkc7qJlud86b18Kywy86PO9Amm6nbvaN8ZQU0po
Sp7l3gVo6xWwTMPUOgptvPiLvLefwpFQ3YG2BeBzOBfji8YdyOs+DQlmjWhm+MVx
JplOJU6yHCPSXipuCIoGrcBBb7pbrDCNou1kyJ0lXGQB/aNaihWEk849ZC0dU8wV
AeA1K7YPSaV+vvzGZsmZVpBZYmDbitSvcbEcza45RALMPrjZ4Vfizp9y3iNBToNI
2XYE47u0Z2Mv5jpWkuC3XQSu43fwJA378kzOR03zvRPUDDPJRpkQBYdU0N7jHHoB
0sytRm3DGZVBMexBODFM/9yMPqIbwRF7TOfSJsRc5r5ZWSZ8rZOz2BEp7j/3UADP
NmzXooR6EsDXKfKJGziMsJQ3AqBpsBFWLq573qFnaUwpoD8KCg5CJaohj7yo339C
erhibkmLJLAxzzZzJtUREo/JnTV+3xpubBcJdDFyXByjWp0LVyyZkt75QCthCQQ4
8g/DfqatbK9yC09nbFmT7uOio5M38OVu/7NZwFVw4LxhNI5UkJOoaULK0OTUQhZl
U9arkxQGUEvczvdDNPVuIzPe6fdGIc53bmWQv2Y6RU5m7rBHLtZZs4EulAkDmIJ0
kZ0mA/IHKIX12IhTv1BjEXkDeXED3EdPlM8sRQTG/8qNO8ZMk5D5lH7dqXEMmZ4a
Kunj8BFA8hQFqYAKlnymvdesDbZQJSF89UBkOJ540SFl4Psq2vd02CNph7vSA1k4
esX9+W1DUqwUDVT+rvBKs92w1IIeTEiCjZawa/V97eYCSTcqyqq0Z0SHOje59IX+
ycR/UbIRF0J0P2RwDFKNLmww8r5t5sIWtG/pYaxI6dPs1AYy/18MUKaIrY3RVnGL
gYG/oM4ajVMQVRlX+dKUxAndsb0h7p/7igHsFr5YlGQavGiFLGv6gDzyIzAZXaJv
QOH6z/ixrU7K6OgtQ51PbkPWLQbdaruqODXf0Kwyu4BSYGE3bnK3z4mX1Kx+2xAm
wF3+B8hDSEurNJtfnrCKN/mu72v0yHTAVKYzi11UaSmzS1lMAUvpo/pLUxKUOdla
t4VhOVmecGkKQnHh+kpSH7UU7/q8Ow5hUodbwKMz70vEOy2/kQF8ophBpM8W4SQk
ddAf1hQaIXb8OmNdYKmUzxjatrk57m4IZOqXXbkIt7Ru1UE7pAFhkcfGs0P4RsXT
beCzK/9PCkN7GTwZQ0fNv0j5B0RP+g3dytUWlnRGnThMVFFfrNUt0UihIEGaCNPc
q18ZCTnU4IZitcAdTLnQuP9B8KvPyHdZUUG4ECCM3OZH4UtOYed1Btr9vwlffVvm
bMO2fPgiu3x/vgu+GEvjucayB5kwMmQlSZRyHnqEWrR7xuCuOyVPfWbSfh4HWtbr
7ykJd5YgIy9s3ZxQZ8cHPFdUGdM4kAG2lDo/LV63CzBCkqe9toznpAVYq3ecB0Sz
6K8EGBAOJP6/Y7HKK2167jw5tBCIyr7EQkBJgFrIuTg0dol7fGALbWxMXcMfCS5q
mOCWlXfB0Dfi+QB3M2sERqBRWVZmk0KljnRe9HpDL8pmHvchQS1OO37IX9RwoQqe
SVX5cZLbnm3oh1ZPbEnSOMZNSE8OKuTWkKZi6SrNTs0yt7k+NXyWvado6ZE9snGF
wtG6mPktpzwWrYvhi0dcU9Nt2erdrubkxH22WeYSzcsLwe/wvTk6TR26W9KJwL5w
BbPdxdyp7Ds6n9243/ivXWtIgnu4TAe/+OmgZRqyF/6WrxZDUdjFTembYrAaX7mp
UFQQ8SVcAMGejmKzr8bvb2YOrHVMBZYSSxkdY6q8b27pdaqdGeRRaYETDt+qtjiE
FXt7oq6vmPMEslswh80oleyMUwU+kMS1SMswi2+OrhQQrBhCiDiAtX3s8WpIyFby
CGEKZiOIFg64xsyQYr4/m1k0/NaQEsDKNO3nJzX2l9kOJKSXKywIRjtj6Dd8Xx+J
Zs62+6Bi4x6kOWH5NZLDOGvTYZNuYW486vqKDVLumh55hQ52L6fcfJGA4VrDUvpj
GOjaxQgCmtJwsxFLupUvwNFTgXEzW/FTIX6qql4De8K0S2h7m18cRzR9VgU89Yp4
P6UPAYt6yozlInNZhJ+WfBIWqKhge7ceNswoG9vRoOf1JlVfB6UEPt6DhFaVsHDl
68HgCyuK6EkZNhCM8gUDz/EsWab55mJZ8F/XoZLLd9f0zthaLXHPI9ynLQtdVUiK
J5XwppxV0sb6uzjfC1JkxaXqScLl+oOg88fdBDA5oF0OZ7tmu+7j+rFaSOqvqOkS
RjHLrluCuug2Yxj+tstMXl6q5piWdXHZG55Fb3ZOvQ1ajz479YxvpxfSX3juU3Q+
VZM3S8neaABFsK/CfpkwAHeGYBw8WGTnd8QNvgyxfnJ61v0yKfoGKEFCcpNcXaxq
I2oRdwY6w6gCIWqXfGYki1SdsETGRaFzSUVbYHdNtqAYunpm7lA4Q2lSFBsDqJ4v
wWqpQTZS4b5IvjKmAnj5dZ2b0y2ZgfhUdeZLZLcJpajXdgIl8vNhbk6+ZImen6Tz
bjKk2v9cGh08//IOGASozLsA08hLafkzMq6zR1IR8B6kr1UkfIuXp/wyFfhn7t6u
A71sFSgWqClL4EIUUSfFFNFM91l9//2nuDSFy4cTFBe03Tqyl50baBGoy5fMzUwA
Kipj+Y/9icJsknFztD3gmsaAjl6mqdHbBpfpil05iFAtJRuMLNL9cp/JiBSZKnUS
erlngpCWTt2KHnhSAtA7jveX6yYGxwPsp5TcJ05OtPA2pLWV02g8cheNaXhm8xKn
knzNO3IHvyWHEbJf5LoWgPxn0DKap+DzY1hQoSMqGRs+xDnP8cA5SCXqhA/TwhGq
CUk72umlhKhwT5xcBLoBrRpH8l9Alayonqc6jFJ/Uu22iKRAXCYpmU0hQp6AdgeG
Wz+9DG3gVZA5JYXnqH7Tz2XcbxedbbzdMXFZlDdCKcMZLrjXk8xElf0BxQW/LmYa
elYnlaWyQZdn9knOHSXTdtT3GlcEj1eiQdTZ/4CNdzBWR9pxKt376GFltI2UH2tW
k5pl2W78NnYtJntKV8Dbb1+883h+9vxFF0hJQcuKBR3JCmbn/KDp35+aEDDpLRwA
TARkjb0T6Hfqf4ZnrPL4TuCLfNODymYgli8Nov+y+yQLiD7zqDNWVMsI4In4lV/T
i5WRK1m92RuLkUtQfGVeTPvVqwhf05I0/RJ4DZqQv4cUwPzbHlVOtGUr363wjb9R
iSRNmTwoKuzZwfP946eRfZrvJymo5GP7ql41ma5Adnd3AJNMZnhbHYFoVZNy3zNw
92eoMMCygw2YkC4f3ntgI97bOG9rQgpoqwJUu20+SnaifynQt1uMsAjdfIPdkFek
m5ZHyXtA4dZby7CFnmGuXTlhFhj49dFd5xhoLIEI4HDw6mkcyLFXvZ9VZCcdBlGO
Zm8w1ET+p+UiIONKeiiqtYrppEPqQG+iCL/IvahhENqNN7aoyfpZ1IRQF/ZwcaTV
uAz3JVoGELrN64mrRvOBAGB+qLnqzSovxyTimuFTwvEiXQfE/y2SyD9OOhp84EYX
L0FsdNk4lbfko88SZoXALV59YEhKdECxDBZO/lj3eLG3GXRCpNzNTwebYR/0r17T
Zb6mcTcDMIaPLQx3lCaOQJA/1UG4PkSgxPwfX8LtMEtWphUixXigqME01Cvsj1rA
CTlW1cY5FiMynv5E0IaIgSP1ZyqLAuTgXPCNNoUVWdM6r9BouO4zgvEGnbhohany
N3gWsc45jjt9QazoRZo8OV5oTtuRrdLDLxqbdxxiqe50VtRrRWhUS+fB8nQoqzSZ
8xMZtiVz20IbvHZbEM43tYsurX7F/v9GEeQo/jl5oO93ds3rUbUlfrg5Z0upsh7q
HFVQoBwZXExJ0q5gSNtLGXroW0CTg6pxySTl4bPTom6ZOCCSbTMIbi1NJq+KZxUN
JVx+OhFid6x34XyW2VohDbLRO1NOHX2gtGcXUjhm4Yv2WAeUNrwFDeiO3+DhLr3U
e3otJykoQiUbDW31pRCaHb3kyyCANga0VtQS3ef2IL+jJZgxtqSENGFlKFX3atAQ
3SbUh0bJGcpPj9BSQxiduQnb92CNvTe5tC4rlxjD6XF3hFRFn7E1fVJa0D/eqhHK
SW8MDrqEYHLU/R4IkQOHFy2ewAITljweeNLFTTSWVmdMzfzFCAESpjB8R8EaTYqU
1ZzMT/4yIZXN42aU/0oOQW/zVh2z7g83rBAxCRu85meXUTh2h7T34Wk1zZOsxIcp
dnn4O0hSsKrtfeXJaxRmDERe6wSyM9TkxbPviRgG1hJRbfA6atX8ZzY4i/2zlexn
c0QKDVXGOi73y6KHAGwvTEHuaL6rffKV6J9fHNLWGfdCWs2BlbY4H5nDVAPqKvN2
6npnoTd/8fKN4w64jx49sVou4ti8Qm0uBk+cedjvzhJ3BwkD7rHcvXShxCodOkeZ
rsSsyQ+Dg0eOtY8v4yjBZ7RrlkuKzrBv8zFoiylOiABNDhAB/+dXAIU4i+i+1gJY
jsN0ZyfsMO4aPt5OBNWgo/TawtMlZrz9G+tQvRiPMys2WqxtzS6K59k1hPoaTgDQ
LKap8tpaL6lngEy1VzqucQ6hnGDmTN0DQJW6l9slktypJkbEX/jBa16HAxunk3ju
tI2n1XDhZsKpdf3rstubxgNvJ2SDx1nAOGdHGwIKgeHpu/UT3Tvw7RO99pHnqgqZ
OJ5SxT1EsDO0Msuwt0WpcqWnhYEBt6i1coKlXknXG57sCrl+GsFkyIeUHE9gYN2p
`pragma protect end_protected
