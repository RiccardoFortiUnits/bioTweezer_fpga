`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j+Agey96UawMlYQKQOqmpPXkZaB1z8Ew8cDhIjyXGV1jpuFvPEn2fb6Ku9hy12m8
Zp136XPG6J+LFx2OvtWPYbXdm5DWlvcuStVcYZ7KbPgH5hYH87QneXxGCin1vRRs
6eMunpDkH2IQt9UWriMyu7NFzG0wLKFWICC388OAe+w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8304)
WuSZUk4ri8RNY8OGovWod3YUhBPi73yfY7oeWPO3n8rhF63NAmNKTiS3RdTqHjEc
G4QLZPgnBcyIvjcawA8Ez5s4uQ84GTEeutke4ZjRF/hq7zLHwINE8M7RNQddl7Ws
dvm5PkmyhAkGxktevZj2mrFKbPA+TasFFc3F7esA45CIzv0KoCAfkn87pmz/2QUm
mx29Scu5zH3Hx9YAduPIO884n2a2Ac1DqrcpvfjhgWGoBFKCLy6/I0FKh3GrXH9w
zcQShbCrvKNVsmTUoSL/HyL8q+4tem4G2whxW1pV3M/CWU6Hk6OyRCridA02JTuG
Vl5wEblRuLDfU2+slIi4DpTU7WQo/hTEJmmhRHCi74ojiUS4VeKbZDxiYVteXqHI
IuFDAph+jarM9LyTlYN0Hj50Veu/lQUrFG+vjLk0+8TOAra1hmnF85CawxeUvbeo
dDQr7vEX1DbjujrEYLE8sAnWL9J3D6EpfltTAAqLHvCnbbd3P0zYbR4ClOmIzWDn
IAqP/MtuVd000ZG+2UJHRIUXy+hzW8N+BW2urO2cgtK+yWzOwAacTmHW1BKy2l7n
IDSV4/FUTVhR53MenaQ+IEE0X3NLp5Flc39LrHCZvN7WXE0DeA6hgQWf11KlGtMU
PEj8PqurIimv+L8exkbPfkKr/3uxKEVThlHXL8pEAbZSWkJWCxtlD0Fex4N+nWjD
7cDdbTIeVyHxx0tbgfyapDJqCRyTyppkrgpWr+u2xDpyOAyXglEOd7hlKDrWLf0H
gPN1UNPbEKugqbQ9IQ+W9Xfop5Vut8SO63ZPypp+t2kK708ZWz1qrZtmfx5uQFc2
chmqJiK7SgWfZERo0MVu4gVmNcDlun3n5CDXEvgcwrbEs4unGKcr7HTz45s1oBLh
qCcyuiPvN35S1jlrKU8QIVf53aEyZWL2l4NDrU9MIKg8ddkJSXZjZmXBdHaXeKVR
BDWY2jJPdHYea0CWrnWJu2p94Jq9xg0OipkfEMySLUVTY7Z6H6kN99cUit+PWo99
27yFxWDR2ltl1vaR2lfZ+Z6tWqLMvQdeFFCFtNgP7OfxVKfHVF3AyVWIWx5RQjyl
9jqycMJo2+3dJJN9XUXdnyfGHYmCmrBk+sfE3lyGENRoW5ZxV7Hm8Ees8rR6KXk+
Be/ZorxVrGENR2lh9jwdABlcGaJHpWrhR7YfbTbP0GhmuceazrkYPricRAdjHfoA
2NXo6u1IrYq6PjIpJH9xUg5bWgt2Ncchr/sDT1u692XSB4GvUxKTQb5VO+k6x7OF
mcvGEPsiKx5lqXakHW6s8trcxdI9Ef7ksp5mc9HEe5pKl4ONlkTC0tOHRhZlnNON
5TQryhJDItcwN5TsEpu43WYGdJh1hlyeTsrTrYfzHr4UUVPov75YHBvejJ/UqALH
hZtL5f1aRiOVx7YoO6plPZlvNC47I3JVHN23alqk0vZMAC89RWMU6Pt5wgqEgA9t
p45YWjG/1Avji/AFRlB6htNKlBCHJvOX8lU+yoTObtVWKqKKq576CsSlMwE0oOEf
javyymvy542a3XoFnCix4cAWilEOglSXj/6q2MrpHjSBJrwx9U+/FmFa5SCplcdD
L1J+YPtKDjFpJDmYbfsqJOJFO5I5iq2drPcupbAwWVLIDqGxtMIdr3tduXfR/fXJ
l/kEMoictUQ+tYtbvmFtqG0UBTNT6ELd/g74khktT/WrYQCVu6hx2wXz0tX5JIRE
aITl7B2c2ImyqqSRDUUh/0AOMmgGeDZrRYKRBy5h9U8XOAI7Eayies2LlOLDEIod
t4XmxODRxhIdFbTQFIHBOcUkp2M4doCNgWBYwF93c3z89+fBH2JGzvYKeS86XilW
gk+qNOEEZduatmIHBhLe85mBvXzLLI+pXa/CiIdrcrB5VeFqK90wi+vMRvHz6QR5
iPXPHJnsfxhNIp/9SwjQOUvajdHlpcwHuqy6UhSHxxsmCxaHM5iCYnmXDyyTgaH7
51d2Gtz5KzLUXmNM9mqfEiCTo0Tz9e0qkA2X4QTpv7WHmJ9/osSDJ+Z5I22pcIgL
RhS8AMMqtxwiXBepHjwIUVS7UA38sF9/nNh4iwGN4/Ux8L9JfP/11xYpz+T5lCdJ
V8a/BEabOuqeTmuRgY+FK414B35XyZOTm3nk8c0K6RNZa65YvYwIlkTKXb+HHDpd
0wht5GJ1k1vmQacJaY0WcaAhmIsZ0e7ohGcpKEDuK3PArGMLUpqZ1hbkzGHxy/Bo
1ma1Etgld2GnmMxpwh4BmkO5o6/qSvpOLqwi1NzKPKOq5YsiMRB9OXItOG6+IkIN
gF09ABWF9hjzPkneissHiJd5FQ1OnCqFbmERy3zv7KiWDLP5nq+wYMBgotnNUhHT
VLEsEfhFj8CjMXHOq+JN6Tvtr8iLRTIilC0ECuGwPj9YYjenESilgoW+qkR2gfb8
UhAxz+s4GXY2Jz+LoELyQRe5UztM2C1nzjc47cbuJz1GbmzULJAnm6bId3hNAezW
sLwmapeO5yieUKADOjm1qOAWXrimCSqKzXgc8j4NgXzH/UVk7c5DHSPKkpEkjsBG
ImMGESnBBOTEg674aiJjvgrnAf1Fyc/g3kvJXYkbBGCmqPzxU2gbmASeLZvR5BdG
Xky6gxTuhsr3lKzfRq3vWYiAtmNXF4OkuP89HKQYOeFjKieNEjg+PpstbH3jAhJ1
TxkdWKXYywgRzcs97DgeyVVpFveBtW4kxoAud1VcZAv26iAF03RNSkHtuUCi1osv
MmqSDtp/OGSDye5jvqgZZwvgXgl9Nko+xUkBnSyz9PVtWAylEABzyXqC5vrYb8Ww
7yag4de1Xc0QnNqUGc24Tbu85O+VLL3nNJKT1Ys8karm1AkhRWFtWg8agzsrinzG
20Ixiur9h7DYG2i94pRmxXmusQacfyPNInOgNyr3P3mdf8aA0p5DhWeQILMjdETQ
E0EJ0tsmCyR6pL4f0e+hEIEJNqZAFUOu8Trk+ZhfADx8Gkukm3ChADtQQU9bib0Y
fuNO4HV9rDf+CgHE6vH5lb+f3g2H43yj6UttLA3rYzW3nCC1Lc6m7yJb7IkBpGe9
LRc3ejPi8mz1iHfkFyio6pCmfrY33mRZorhwtCO5MSM29UChbjYa5vqO0LnW8sZ9
FsPq0mKsfu1avnW2qJTkbn5BPVXEXHCE26tkXtmYSe3O3ZDf34rEj0x08aEWpw7l
COczFCPzRgEGB+Mu7Q35Kghc8InONN0jM62Ks5AquF90pvimf7NVSqE7gbYJhZYa
wTjB2Nomqwma7dcnwdpZwyKHMLmCm48IhcbbQ3plRWnRF1CH1mDK7YhYD57+8l1k
SkIF3WRxyqiCf0sjeoRVFccumpaQ9yJh9/rOqXhSwdlGgb39sFMblY/50bVKXTzo
Lx6S5afXG64O5WQqmEkpmgLLdMzXUd1IGeN+m8Nmna/Z6TY8cXVudfjiX/J17XEI
Mgq0gcLpbQh6JO0SjuJ7QFmq1whAyt7elmwOU+pXkc8RofUeDmgM9bEkeysbBger
JK9xk1w++aqnjhPopIY6cXsd8AMhNMqTKGBShmpHcmT/4oWYH1+hor5tEjCIwmA9
v7k0yiFedCmFUkXWVnETXtNs4thV2KVGLf4GXt138Jdxpp3XdChc45LcVfsQ8gyb
CmXBaCkTfzc5G2Lym3zFCbc6T0KrH/5A/XqRXsBTQz12vtmgTQNpOwfXOinCh4Ob
qd8JKhgLQiGjOoH3u++YLG/LcRofZ7kN86HtpvC2c710I1ndCl7jOTqcViMXU2C8
tuTJYOcIu7I1aLaaIpgrraUrgeq8M3UOCe7wwebFx6qIjsxrbuE6FkyonSS8Ytzs
tXPE4Xr699aBnRvDbe3oc1vw5M3GknlnvrnG3VtvLUizo+qZIhvC+Sq0yaDomVel
AwFzD2LAcEUNgaQ6k60Py2VAJA+7edz52rKH9ej3aAmBuOHolzTYHTEBIyi8tlmn
nKFt0Q3VRcoobgBgJA8Wr716ejWGoLqpnshkZPBPUwvmupct9WG5H6xXaCfoTIgb
9FK68f8sk/27IdVYry6cZBmc01xeQkwqR6Y3qkG1VTW9f/KDpB37iONMsFlF3x8t
Z+HT45RIQShq0kh9OJT2T0yC0zb3QyOiV+6itJcWS8wgpHTUTQ3rv+8dEAS/9cXQ
PxYkEtMURk5hjHRvU0+dkQrULVO+RV79X8SPjX7/gywRpitFiNig66br0t1/herl
LQtcsncb53QdVqwIJy6KDIBtqag65uOKYnTN3u20JlSUvKi146GRureyH1SFdjqv
IqPaUVSA2Ko0czcdCyXp/Kr98XXuWPDuf2H5zCCyPJoG6kbBAFFCS8EpNsXMbd8n
EC2l+7IuGhxqVEgNDAzbcuLEaQxHCcdX1nRFMoNglW36sMQTvgi4SDDg+eVZ3nHW
vHRwdaw1N/DW2MHygmmbkr8IkKQQxLgV+YWta0mwz1LAubyaB1F/fTFSvCYma9Yw
f522w4Wsj+GpoFnwQ1GPaFiR73C6t9vD82mQSbXi81oYSp2TNlhb4YPQgxGsMjxN
TFL6mkNw13UjgnHcosibE/xR3rzQVJOVfPMOumr61PZjYZzotLaKadQJmxOYE2My
o0DCywQ5NrPRB0joLU+uK9NcyuWPXSSgzOeVpKFwlsSc6jARSZkeF/U8zXvFDQ+E
Yb4kCI6y6dcVh5Ze2OgZ10M0sDhgAisCxaaPI7NquqdNM2x/jINqPT2lYjlCm10G
WqKk+Xu6HQa0ypq8/IEoFanKOhNyM42DUdNviOytnb57z8f00DBxm6v2CoqyW99W
Z4jvcT8FJKJrcH0duMPrdymflaRukrfa3JMNg3PT/fcTtBg98rGSuFo2LSlOzhBE
KF6yLt9iEEiQmbZ41pLamSClEKnzx41FTwkFxIH9ZlxEjxGji82DQMpyepNKn3ps
5sUyeaQAoJguaLbkP3/u4uVM0OzEfDzaleQjKyeV9Cpr0zxPKQhdgtegKC+CiPk9
8pA2KA+4ixKDJ64eDQxrklxZiTRM5oDelgZAJiqL37sUc/qzBcFWaweE1EkaUewK
lA/ah7km/plbgHC3pCGvwFt+DwkSURKhr9DfrBkgZGWGEMHHmR1e6v7De6cZOUzw
MWwA3eGYm/sBgaFeaw5M05BT2WOLfYkOY4kre/YqOiJMOzllNUaOwkX/etyFwp5Q
VrforCO2PLFXIVN7VzjTi9NuqVBaWRBwlxABnJ+yk/xMhCqrR/ktZauunnv8dYtK
oPZHjCvbhlXf17Gqb6uH97Rf7J8WU8cPRLyj5quvwmLqprnf+kaBEjxtQ/gGysy7
ZjEd7mYzmpumzbID2CvLWjAH86qG5Pc+UYEiFjVOt3Zpy6U10XExHGY1xCy04RXT
1izwKHBTwZNwpHAmYVsgfdzN4z+jh1O6JSfqDHRB5hIUA0fBJIBWLepMcxXf/fMR
VdEvv1fUYhjKECmEmZouXnCyc9Id3IsMTwoGkP1inKpnGY7fdAxw36rvd/IIE/vb
VMEhGjgHG+ddEA5FTjXy4QU7wuXqo/pB+L00dKJJS6LegBwZ0b2EeM8MHZnBjBfr
3tM/yhKM5OCtL920aqE4clYbXmtDWXxybzatxJEkxePaZGwfqIa6hG0aMDu8cjwM
NgZ2+drmenuNE6oWlnH4UXsNtVju8Sh2xiLkcLsM5p5QjtAvFhr8d5BUPmYYF1pO
s1/n0XxSuRUVjOKp0UTArSTFaYMAsnH1kqldgdCtUrZkp3kpIBDZUKhVmVh9fIEg
/3VtwD7lXv+iWbHkcroZ3WyJl6WHrxoYMYSLkM9XWC2RW3u4WnoUp/Qbf7TTMDWL
eE9oJ2725HhhqlK1MAfzd2JCr/6wfqj0cQBWZu0jqU8zpfuG1b7+hrxec5IjkRcv
H5kLaX3UxyMcTj2YqhwisrWIiPXcmzFWEGilnKEhChiaBsHeq+Y2dihTjTcrGFxi
mGLxonD7ygv2/5icD71qny2FhS58aaqT2SqjAocoOc5rezPuJONafZlFbmsUXgpX
TVyi2qRphSRd53+Y5AKl/O8Ws5MLaCa6xS2tX5UeDdQyL0txskSool4hmfcarsR6
ySzo+OvL+0/1PI8mEzu1yIp2c1ZHxARY8BrR72LOrlHI60dfHm6MYfNkIdu/vGCx
c80NJF5iQO0QDgAB0oSa+RA+h6CXMDI8LB4gJ18N63dBk243w7EOgnW2fEsgrkc/
Pyo6mbCezipHCUUWgHELoBfsPKmRAZZnIaNzgvvIZYCsvpYR2Dvge6wwPV/neG7C
WGgQgkP0311gkPgNshvGWdvl/PxGEc+12SkUu2K7gZvORNlRv1RFG6/NuMtip7xH
J4eOqE9yAsVRh5rLZrWmj/Q1Z11DOZmCdLnZQH4PzzAO/MM2iyxytL5/EnpnzJ7l
bchKX//nRbde+DkTaqs2bdi4lTIYXJrjqltcC3X033NBBkCvUhNfuacjJZpDfq2e
qW09GwdCE6xJWgDCYhkirX3XMtVNV8kgu/zWWJ1jooC7BlyDhP6OriB0ZHzW7SKA
4S6A49zfRO2SfbeJArLmy96J/8IV6WOrGvLDYEwWjawEaTesmyyA+TrhCx99snc+
VUiMe/VKup5TV4zTVxxnYiIgm3LAifjI68lzeYGegUWTmSI3jaTcjT49kCwpfFSH
PE0JMnSl7nT40uGLtw3MlPwG5kHxvIDNIdv3CmPYq9fmuVLiVgNZLIhDSOb/xA1j
Y9k+0pyiylNd+RysTccCZ8nwfrQld9m4p0/KNSPtJUN/oxlsct5L5bq9YwWTVzux
6CQFw1xl0H9zZbP0Kx+e+n+hywMbMgtMWWThSqjjhXNcX/4pZLjRqE+f2EgDa4d6
g+Jpa1oXRVzZdLeRUstxRZT2iswaZRfftrpufZFH8jQyL9t+zefghOREXb1R+MxB
MDgLXAXnfman9cn0G6ECv57VibLGhiuy/LRQbYVa0b1lwRqlB4L6KXjYVQ5TvIG/
qGr5fredogA+uwEWvJAl9crWdk2OBPDoiq6C06V/n6j9rlJmjm42PErXbj2Cm1Gg
zTDpdkQNQYwvH9fiq2jviodaI7XOLUQ8Ryg7hALbAv7Ozb2WIcBQGiW3/jWtYXoG
NPV55EmDSzqL+qiiv0mk/TgJ2/sb30j4y3uXBcNvcEyNb00DeXWMPouaLf8Op138
hz9APba8tYY6nX0joNwz/dUPnbFb3rw015lJLYl1Fhk7bY/H3rbgCJJqvFU+g9fF
drEnbonl+qGlLJK5uULa4nsXm1mls7xbABbtvAXrC4d5u0QgfAJIuDha7TxwHr4s
EIyWhqJduz+53gc7/ZPtrmYb4XK3/tjtDMIdgYnIwXEFUKSIaF7vhDOlT2Rpq2t9
f/iGMeXOHDWUie4Q7vU/IrMK48wX9FQ5T5HxmnBs1W5tYiXfwuaP6E82bCgMDnIS
btDDLjMPvazriaZPh9qDp/BcgQzfxwaFRVi/olVIMkaJFsB+8S9L6eVyqBRwShBt
p8h74Crotr9WE4b20v5McmR1/uEdbS6ZLbQrp+s5bcFgHY8x0M9Cor9dyJyqBTu7
qgIOqr8vIxIb1lNcS9xUvKrH+xmz36fV8A4IYqOPNovvpOS2LOBamKlGpybkede7
776kuW2IchdmBHEVBLohXaPVvN+8Y/cFm3v2zsXnSOlaLqEpAO1+3Wxl3I2i1Btt
dTcUPDFAB5Eg2nQo0Q6jv7ZgXKcvaLDzZjQVPfuc8CZKGIRp3dDipYcc0v8aA0wg
QrSL7GcoPc0a44AKGC3f1aH4EuMtbqA2NfWCwGUkWamI/sgCmoESZX71TKtIuaV1
KYRrJmTt/7tHN/ryihYaA/S6ASPHWzMmbAAK+9eMVI3w/aCeTtIsZ+aDZpkI+Esr
psjYwjTWWjs1wlCyJqShVedbkjNu96axazYAyh52bCLgzl2eEXYsV5brzcBCgHDn
qLy999gCvaPHV2B6XDeCVR2KPWisIv1z0Inh/k7L5B9tS2tfeuj7SNfxgaNaZi5G
ETyg02jFZttW8vn7qGQNoQKzjOJu0kuezIgpIvbmNE4IJaBKEcNwKKJ2womKh98M
iGDaWpEJKiR7R4PzpSBMvB2Up8h/RhL14eL5eqxOSq6Mr6CaK/KijN9CnRg/VTWM
kE0pEqRJI4dgT08HOIXQ1Wo3iI9O2Pny+mdJ3YzkoP5EC22WqkuQJTP48PBuWuAR
mlEeHpd5gpSdre6zsDHLCXqJdgcGlDMjl7qeL/ELJkeRSPRZUv0MfRIuR5M5AX4T
zCi4grYzRBnZ5ecJ/0EtNIU4rhBkFByo+Vq+/MgCj4jf69/E9p//R4lvL7uKHjaG
rE7mSKUhtN6HEU8DuOx1X4OslWfQkq/rdZ8q7QgGfbM69iNnpovUrnIxMFO5A421
qepY5ueO3gqkW+9CoFjLf203skdmhLz+NrC64nZaz0rg8ua5LuNSDiyr3+FioE8d
kOhH5JwZ0cKLtwB3u/qKYPaauUtxF9aqQ7iheKMskyphnnq3RXc4fjnA/ZLOoXEj
Ay6OEhxGyqAss/b+q+3H0rfxzNuiYrbcXrAf3a564v5LlJA3DcU7doL1f13LvS92
MuThdHIrJt0SnxoWHhpoznUJ6Of0ljIiBd8X6hMvTieCBtNsgihsL18k0Co6TtIQ
0w+tsG7ERgv4lAIh2nksLJJSR4rT2KHNeTQ6AXYhIBUJ7panCQ3hdp6acmY4vu3t
9M8VpKqzPqtbUEBm4AaNbSoV9M5YB/bG13qSLO+o81eIz2WWotfdwqDn5Q9wO6ba
8+x9a8lh5VeAFkNU7n2VFpiXhzX3+AS2fFK0NnRBmqYZTN6Yq3/lhyfXTAEzoHZx
asLZ2hkZj4Vbrl6MmL2u/W9vDM7XDO2e9aQQBqDCCA6EMGGpgks5ETRxIi9aAwTH
7p/t/6Jfi/ZQnwHrzTa+v2agU4BZe57RzlROlVUmWWYAxBdKvxc+PXQGtFI+uqCL
VifQ/ctQc47pMU5s7EGTZZPKQprkprklEC/s4e/KqSRLeuyjTe/cDo73BW62YPie
gsnItuLi5BKj5MymuvaxNC7KeZdsLPXFQZuMH/ATVe3gaiAGgm3J6rOdfLuk8h93
Xs6+hlZrWsLcMB8Quc6u6bpHso+voOPOUgLQWDcUVKXoU57wpC0nonJtyybQUZEX
E2/+Rc7NR5eZuA7JQtDUu8T9qZEZQYl6qBe8YyF5Qo4ZtcFKVC5+kfuijFcJ4gEe
fftrqPrAz/ARucspwTi1Wes+zyZMR6oQbI41XsMNGJsBZWbxbj5CTfOeeA3ANicA
41YPydv893useVwn0kHCV/qfbgzwHWe6NalDshxTzGNM3fB2mjFpcRkJG6a3L0er
VqqADGAU+DtdHB1DRdclUArHCBtqO5S1/zb53dGJeTFb9B/F1EhxMi0Vz0UryyEP
fKXcuUVmXRnHmglZE90jK16qhi5j4/PvpoRV0+T0WuIJ/T5CYYgzsThlk8lN3rh8
lnAV/BYDhofagliDIX366FvryfcoAtcrGGz8YvHOY0a6+msSUbexs4DELPC3juM5
0rMVdeL8dKLENu1Gt/2VXO3a/On5om91cp9vl7k8bUcx6/RW892nxX3dnTYn273o
h1JTCsqNj8mXyWIOOdCzicSHN5tWs5tVWNV5e7a9DTZNKLgCBCsNPxCAkSeltmAz
C9j4PT7b1IebJ7s0moJFImKzGRt0HHR/1iIUm0FKBdYsZj/B29EqUhp/h0VDeA1L
iDZ2H8RPQrG9i1eubFpFEbyrlICXQMYaa/voWToQ6yEsl3fsI7O0k5Oh31g7j74b
UZy0G945zROYC8EPkDzGRpyKtjOZGjiA67xo+m7EQChotZHXpP33JDgmYPEHYchX
py1U7Q1/1hT6zGqi+vpzlL1WcvXsRdp7IvLFTWHlRrZYDIBL98T6HiEynMg0MpKp
4EHL0czAB86FLzgibcHUxWZHM1jVBDxt11uV0MfnLmnY5P9mO2B5QKN/nQ4LJaDF
jyi+bPx5ZQF7QBITssOA96BQqPxUo5Zcg7nPyPGJXK2EfvAlsa/paCetU5H0ZnBo
up0fwD1zoZFwaeQrcxVtl/tbD7P+DLvg6g8cEGCGHIcYK0SM349ZDYDbyZBEPRhI
IJ6bzRpSFh4Z7VgnO8VVIHCrIoKRJN+4M64WmMxgA2PLOu90P1IPeGonjhYVsoFE
C/In9Po0Yz4ifg1udtPuOCm7l/+2hgQ2thKqdNfnZRMPbjy7fCykf7FSov9QWtNt
ZtvqMyE8g9fbEtkPK7xgNd3hjCidCBBI1nI+fj8WRF0J2uMWsZoP7PVBs5pMM2FP
emTapU9a/VMEbYz1QZq57tBfQtKhofWgwXdBtP+6AMrItfwAXoWSm+GsmUDuf7rU
oi3/DaUUBksmdDnGDNgxDiTMpNwpDo0+cOZsglLnolnvzdxuAjkIQcKUYh4d0+sP
cvTm/gR5XE5nHRTHwowEKLEtkTd7d+lleIXEKTTNc3xXlcwFLLbExPb+d331lQA+
M9uxUJfJUybEHm6kv5TUtBcuLkyG+qm49M4auyywe4JonaMNUUTEiATRTSRqbGMq
kVE02fl2cschfSVMaD+165jD1TeAYHA+S/xzUWl6+g7YHJiRiOT1wVeaEmnOI2Pi
0GBZTLebNkysjxmDJ9epK0dzsiW4L6iGDp7QBhbPbIlht4VMx4PQ1xiBFVl0jD5a
N+tpeWxGBWENLuLc9G2EKeGbuGcdY+bG62inChJa+L1o9WgnR8hSzJFYSCHBaG9D
ymiysmgUenFHywthLJtU6/MwDzpjcVLE72edVMySMkn91dTsao3quopik+Xbhva1
eLYc6NT9xMD5uQXy+P0wVnbjxTEeh2E8XaGSWnRFPAMY7MNsM7xOJBGviWQ5JwYG
J0u08Vnn9EnHNQgCYQAvCH8QDJttOJhUrCJlPDZKk5WJ6dSIZJplGMxBvMDaYkuW
OeGPNZzVz46rsyMjea9l24E/Z64weNRyDTnwMiT6YdQGfD0sVq8VMlPhi8cgVot1
/sSPspiXbAx+cdcCYwM4V75htaD/Vq7L7vI2yvgDJXSsPP/b3NaXcscsqZAURvpX
`pragma protect end_protected
