`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hKYToNIY+ymKtYBq2WYpadHbCDScrSho4QX3HrbyKo7xLLFWxKGILVFE4f9W2qx7
7Y1trPLulQY0d2HDlyy0NMcgx64x6S/tedxa36WXfo5BLFWa4gC6CNKOSoVwFGc4
1wtWvMm6wcNoJr1uXwgp3xzNPlXJykCd/2kVeOIyltA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5552)
Epni3HgTaalABQ5xvyoduRdslnOh/tlsXwZNO36mgTOp6jb4i/75sqSx27LpZArL
3/iYn7ieluN2qPIbOCKeIeiJ9fxC+8GaoEL8rD8Vyj+1lUAZlBB2tbskCw6YvTGD
fJtFZAm8Um/g8uDqVwHBZaEdDqgrUiNlc7Qqrc+l5loJutf0OoexddEViPNZDBFd
Gg9lsBEfPmtzICgAbI6iKoHTXzdjzVWJrAddYer9+6xPeRxoHjUsLqIwHBWtcekQ
GLGR+AzdqPTs3TbTGo6oLjte+2Wtm6lbE/zyo1XPdJsPgQ+5+VtkZbmkF+FCVGzd
R0yTcF3JRfXYu8TQK1TMkMqTWg6VYfQcycKAjpmsVD09ilJc5fQ8VvL6xt3Wy+Cc
6w+BtcYbH7dCVnZo8HIOgNOzt2T2YH2yX4CQuFhnCMIIovhuj3j+aMrtuGH4uL4O
iiXgOdRmhC8601f8ajnt5c19FUxagpjf/nhiOk9IXdafgSYxbfHbiry/2fwIsYej
MSNcwtI3tOLuH4YNflMyRZL0et10nmWxygPKdruMzYpfGdSZrcSyhBKCiHw+SGYl
C0hJRZp6dohSaoeUiZiDtWtAUx9Dm/ylOP4DH1OqoNYUv1Iub4zljlTFegEsC0vG
V+Q3VUdDJvzZTQnuBf7lMBAkBaWUnwQKfZ5YzYi8sobwsdLRE/yfxnwhTc3YeM4O
Kz+EmTWjLziePqFhx2PwRoIbzGC+owahRR7Qs+2g9GqKpUaMzruB1Prh0JMF3Ibx
5/78MEpB7LjorPZERgiINUEfiYjnX7om6m22tROIMlSRO9sWi64dBm5iVQlpk5J3
UYhWsvAeiGRRRTdXCqAe/149VWid7p5AbGVQYNF1TJexZQXaT+/2npsql9t6uLlo
sy4xYCxN6TOoJbhXMWLArgPYa9gurHyqc8znqi5mOtQHAirKvT8GBHGUKclsaRx2
maVpnIMqWOpUri/XOqrUt/k7TtXutUCpJuxc9LY20SAJrVvBvyErXJO54e85snTc
2xEeKqNMX8s+Z9P6MSxeoiDAE6lPo5QgB/2bqdwZ4eJdu1sP96TfC3gW/IWtMjfJ
gsrIfLL4CYg+o1AsLxP83pMTOmtqaxUY1kYawt6532Q/T1ZtaWH3akb+dYkKe6BQ
frLnQ6uvzKaFxbfhS7fHfTWsZYLtG/SPqmRI9Y59/jRotJ34ZAZ2PgnlLyCaV6wZ
ZfvIxJAsW9KAsZqeN/nsI5sdN4OFcHkpZnUdfFYcsrTeWAc8hdIeSXAXV86fOtr4
6glg3nbyBSzjE+L9WxLihXE2EY8bGVmis8TquLKu0z9GCcC+ZGKg8DpPCzaO+Vjp
WPI0HFzknWwUM2GEDowc+32jLI8BJFdRj1S3ePO8d08RkMb3bxCqFgoT8RmSocY/
P2aAGIWYETWHlYBhUKYGB2RNrH1AIhjfzGY8NlcMLcpkPJQ6xPiNjXmLoKt/n/e/
XGZ/a8jlaFIwRcXO7wJtjKSGsr3GE/KzBqrTZ5VGP8MKBYIKHctJZsVNHwetvlJ+
t2Tt/pizkzGFO5E+Wak5RhIZ57vwLu0gE84/drLZYFSJNRTQRsCP9MKgJpIog43M
XyiSQYtSOM1njwnVQVABzRRH3izXi9GzaNiHDn05ucR1w7WQwSBgB1ItdeQT2xJG
p3+4y9NCOXVhXeW9v0fLHfV9xj1OmdXQXRwXBUalXCuxwZ9XWP3xI6PRRoUiMXgm
Ht93CKQI7ubSC7rFeEj1L0YVCGfbIUESR3qEO5BCKVVWwDfivuVvGrxT4rrLHbD0
HrMwnsWUShuGjFu1MrjqtHp+JVSV2gfn09ZswzaeB/087blIsEZi4rH0IesvMjK2
xDFPHAT+mVWBiw9nM9ZhQrtLEaJzWAEZn+pWX0RXK5CDbXp6OwnlGHbSoOnJvh9+
fd6udqpaxlWWDfSo7jZhyv+slPOb64Rf0b5pZ3jmjLcBEvddudr5/ZojG646zlAa
qXyMB47zRwgd192kH6XvEmMlPB5pu+MrHl05AJUgh5pcUn3zqVYi9rb3pr549GXG
kO1wVx6ebmsYLTcqwcAd4jiGGLIKUYSwgp2e+ZzMc7o2Dhzqv4mljHL2lRMGFqU1
Gff+2Ivi/GGLstj3ZvuWwkDKAwDqnYb5L/eFJUqyp8CSfmob5Rgix7Ra2/VV0SON
mjGuqVSv/5XqKjd1DP5P2K2B8qR+KzLBtT0Zmfye1/sMw7XJwYBfzMvsB6+agYxI
Eai52FkJhXg5T6XxQQ1gKMj4xtumaU3Uxrfr0UsivnDxJexlyLvbgxLdnBK2Lkab
atRNs5LyuEKtINtdwKkFqoJMQl+xoqAK3PwGfB7n315yXmPgy34hp2f88VrNgiPm
hhyxDNxQOVY+fevtyZqR7BnWX7NcXcZWMl+H1vUOqG/QaEw/fyHTaWl+dgMlA96h
Gm6ZxhJBOU9UxUdpgFSGcQVroY8t60f82ExrC5uwCGZygMLJYZHSIWCOodMgqHTM
wM9anNS+etBkL1C61V+F7nJCVenkpvjN99fx0/nl0lco0cuTW8jC+jjMTj2Bd9eF
OqFFHvdULK7VPvbuQIeD8SCDQ+c3vdHimUve8iELI5EnC0YhCk9RGAwjSfq7sCPI
3qOBy652emz8NSaGlcQpavytvVBNQBDjvMn1ElF176Emsya3MOUgJCX+xSv8nAkD
xLd6btyjBcoM1mThUqMnycYF608/F2doVA/gcuR+wM4pyxUslURJGmZx1fqB/NgV
ys3ySYC4LLn/e5xHAVlmytr1udrNMiWyB9+myYPJI7HsBx3jdYFffmP46vqC8FEK
szv4leg93XDYUi9n3xmaHkRaMmMXoVQunPkdlT58C2P9gI7POev6tQrFIheNMAj7
Wp7yiclV4+ISzuq0FgQG8Xj+EnUMguCdR9/kno2ddH6L6jC2+IJ1717maewfPk9O
QiyEnC8YeEiwO1jP0ZBY1yrBh+ZgAOvMsiVp0tTf8Av9QAkt6VVlnNK9HV+rYyeX
BLBsAcL5Gzmo+9Dxcu7SpiOXkhlX98hO7iDhPFBHE0jgaKZIocwTjCZZU4cVW1jq
MCaT3XjkeiOg1n62XXRNEyCQRClZ+FHfU7Ifv7nCQKsJ7Z9DC48G3NpjlQiUai0N
I6wvWsDnjKP7S/2LUaDTKcHDHskA+npXU9iCLcUAyD6V9oZ5+Vn8yfHQ5VT49XDl
+0OfDCHOSdTmvo6T2Ptbw3oY4wK+gVh7O9I2zhWaxAtky1IuDPj/wIE6h8ujwwdX
wRCQOsDKRWpzCn7BN1ehjdooRq1nofwu4xA0qE213aN2iLCSMx48rBQRQO4fbjWd
iok65+pCqrpTWuc/MAP4ll+mMjT9JOH1PxZHaZI+1Hq4dSQT/aubpxpg38sL9en+
glmBG/ieQDIzXJ5NLVNiDXZLDbc5EY0A7Q0kS3OxF8psOBHECKtxkefrypPXyupt
+9mMdFBwVpiiv3zEll89rl3mZRR98MxK9fsCEgkXlCnqmWOhjaGz4+H1Np5IK7CF
AE69II2y9+r9AyEWD7hElFDeJmW3jEP6+ljkq1prUjN6rEjPHeCP0yE4t9ybyAto
nBhBEFh6RCObpIv1f639HsUqnrfesURURx9gyqRKqtcf7g3Z/9kS/CIGv40VrWM6
TGlzymwpkxtsue8LtF56/cmetYqpOHMx8KIKoCRAeHsQe5o7Kh3ImCXbEDkzR0ZT
YV5IwCRY+T6Yso66NGhfJo5R2zNzo2z6EeBleFN0u33Y6z/Ijc2uyOLRIvmMe7Zf
6xA+LsbLcqkY4e3hKc9dllHzdcjnayxOk305sjAXgJbxq83OzJwAZ3SdBr2Xb9L6
gNkN5iX9KaZzEdQfGJ8BqHL+EUB8FrlZ9+ydYP4wVHb5oxtLE+iZ1dXbRz58CF1f
YOvoog2g0NHsDQ/cvxysSx+0r7yJJN8CvzJaieYJaR71YTV0OxfBThIM8E5itE99
w+UydCpM5zbqV9/dP7Cwijar0/XJVaM/tP+aWylfkRifWScEWCC6hVh0atXWMLy6
xeDDsVYfYGpoR8KsVv05mRIH7rrETz9ErYywhhrgRws5G075pZH9YcRImIcX51ZR
HqJz9yZzZNu2OCCSYAPAI4vfNWrNl4mOin+XsEuUP7d3BFP0OU0mlfm/FroPWjZC
tQRK2ueBOR2YW8eiQGC/krDbWFFUUG/o1IDOX4r3LnhiLpPgB7kqkHim6MW7oNjh
5lefogEX4mqTca7oVnY/Gu+UR8KoCs0axUGaIhd0zDPwIvmlBDqQuzup9bGr8K1N
Ae6osg5WK4bJr93VrQ5S1006f3f7itJqHgULF3V2RrIm0x2unRFgjNRU7TPEI/Zn
K6nlLVcWSD2tJjp1k58uzwPJgblbaaq6fW92pnuuu5OgyMy3HeIDaQx92I4pEtCG
QA3Nv284tHb5v8wSEUR7lsjno64bWmOZ62XwVfjtCi5/jTkH3jd+nXfkU3gdYLwn
Lnf1aJPKxel8hqi5jrn+NYXks8P/Lg0e2mLIH0RRjMTMmKQwz2E1rmR7ZYgBD6sc
5aWcdN1mfK6QSL8KNkT48uekEQD0SC85RVbVegqLNEBBMBJH3Ao/FWCLKvQNXqG/
MVA3N/2/pyxZ+5JgbCpugk5EQAT5uks+7aTtdxRChcTjCtM1jXhhoQSUNBab4pJz
sC+Wjx2VjV89SB7vLu18QKiVlLg2QM6ZKIPF/vNXiNG+uUPImCjsDgs4pXR43IJa
UZgiXnCrVCBuGh4s+p8k3gWGJy2Crwa49CSK+f7GAgwPsFFdHSTMIL+tpRpUFR8k
0nIbjy4GeXqVTJlXzTDonnpd0pTmQ9XeaMSwr6Pxl6fIhFf3aj6KPRSEwdouVzqK
WaHLO1JJZUXh4yFlzFSUIO8UKGpXVGBtnorGK1TpXnW7HmpiCiWOX8jKzGVGOnf6
hWkc+4Ni82FUCrWk1wZU3gYsECEejCHQ+2EQ6AEid3UoMqYoes85K0zxU9oSte7K
bXq0B3ke5XsW/koTSXpQNAwSIgeVuSwiU3hPqMQk+xeugzOz6WBGMy0BWwubtmmV
eLPPgPfZoDrsZ24OHkZG7plUeml1VhwCz9WXUo99p4QgAD60NwrPFd4RyOUAdlAd
1hMLQIJ+6/YrjSbdBOtS3NhUZLTbCN0ficti6QNggditEszk6itSO2kB+Xx9djBU
c4bCnO9dRtfP8w+an7Bo6fN6XfXeBtwILeaLr7f+MFFdNwaHlzlVtZZxTKnx7whi
ukoy99LdiEFsHJpqq0O0cPM4kiZS5vYFGjyefobXXrEI3K0lYQ/X4E6r+C+rpjEY
c0dqJovvaAPaPzOZZ0Oi58XN+AeWts05umCqBJZYkI9B3SHTsg1xvzLkzXaHSD6t
6W9ywtI9kbz/5OfOs70kH93OH/ejSs2Xv4BmfM3abXbUJ1gLs6gWx/+o7xSW36Zy
dXQp1HMFuDHT1QY7hz6Y6eNmoZgDSyGSn3nDYL2H4BemltF/KNWGzZx1X/hQgwdg
0b/KmBfM+pvDXc5weJ/IzOaQ/MliKYoa6pSMdQNpsAw5o8KgenFHKI8lCLjTc1ng
Qm/GhCQoNNitdnChUE35r6K251xx1wBXhcRTQfGabmD05n3OVNIkmtyWe3wKbzZZ
W9/tHnN8/xZ9gGP8aPgAl3tCANhdgs41UpIF0phQE0cbvRphxjb2kAqyiWzmm36x
gdZL5B2dxNIRwMfMRs4scqtO3aXSCq7toqvVmyp8y8tiBeVKDcE9V9X9j8s+9HkU
ERVFUPApzpQwyHDFfdSZWlMxlh61d0bMdBTgeI3AIEX95tG7CGXcJej6V8waXHJH
8ox+79c+iBLW5t+jxlwtSqBfOJZ52C1Jh+abhzIVMJTfbvKvBn+4tMM5YJM1i5hK
gv9AzZRJvEi8lIGH5DtFZSl6eERCNriTQ1AOINA6AR3EgDKkc/tn9bCWu5P6Z9s1
HOp5oA5rig7vIC6/5+AwsD0gW9tiucRHPHzKrobSekwtzv0jxdDPPLzH7flS4exs
vQvtEAxJSMMRyFIQa6iOAgDahOc8tGiCDxu7pP9MMhtfmKVER60m6qPDPu7Mibzt
DFdwdmG3fmoQyBz8y+YuQIbiO8hb3SF4OJdogY4XjRD6PQdfYdyHSZ2/6DZmpQ3m
Cy+GEQm8G0BmvC8sodFJDiErZqAi8Af8E4usKpg6zRA6lI1oVyaI/JH88OiGQVpG
J+X8Twgt3P/QL1BHdSbDHkTBvB7klr0vHsPxNWEeIOK8Sao1+mZGw9Ixu8sWZ8JH
T0WiSSPYMuSCHUMYybPJ3wtgBVT3BbMBV87lal9B5jGGNCeVVVLmN+sTVySjosgq
DzI6JeT54QivInVnhwp+cZ1OHBcyuwjdKH0acYQnhXUrwxdw3L0dXcTk0N4wcirZ
Cw3g9Ju3J8Y9O4rtCgrnY5B4mHyWaXLNGsiCv/KCZF0THz2iEzmh4DJaNPFbgHBV
6/syNn6GtMBX3bkkgTwj+YKfM7mvalhYRMkRVOk4nZPGg2mrWrxF40lnH8mPBsVc
Cp+fPBMq3q6jJ5wM1ABKgTks8H8GbwiNVcp+cvx2hVUFGw5d8OyOJ2NBfUEThiVH
eF+RubWfK4plnwgeuViMUkDl7BNAYvZXrNrEaEUm8Xyh6mJEAcTiED7PaG324zHs
eiwmXkeozLbrmFjIvVaByPaPGgsrKLxLqOqp/tS7yTlGIguLVtdhP/xRBlhmtNnk
HqMQvqGYsncxNLC3cXpr7DZR2UetlNjnrtT0sUKTIoDHRFAi2t9pPJPTvluXQmpv
flruVmY1pp70HgcrG9SpMZNiVduDJWZXHIaqxowF7cU62xlE75C3+R3Dvldq/I/5
xkClVE0to6DJFFs0He0vp/EmFVec0n52h6MoUgFibR2C+QWWsWY/UZcv+KO66A6M
lzpK2x3lQfABgiMP2nSVnWTWv3OfubxKn126/M2P809aCO/HFIJ4DVRA6b9sDXuT
I2q5FlE8i12GBfYYHLxeXlOj6GBcjI5vZtwYT3Fot8N52QwG7wpSek5cTIFJXE0T
o6bWPH566YS1z8SoeXwjyNrQEQiG7ksfso9osnHBshjT8K4feioYXCqQGjBIgYng
AkwJAx/ezvHA57xpY8pJ1J3rPIsan2uBP5Ycw9bxHg401ELZDsTeeCg6JewHT1wT
Tx+cYPiiitJAFJbFEdSSQSnjcS+SMBhNnhd24IYOqjMTxl8V0AONaqzYQR+kC7tT
j1eL52Q2QnqQwjzG65jIuW3JpLIMl95c6ht9A/cNsWPLXaWMsKmEE2AlW19KMQLZ
tg8mnIy65yMS3ZQmaDWuKtEtFjhsu9Y0q9edazx1i0LOnQwUYpiJze2aOldi08GD
3DfkVQ7m+ucRYGeQivvWjDKDWSupX/wpfRe6ZjIcmAs=
`pragma protect end_protected
