`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k94RlANjPtofrG6YacbxJKEyLRAraWBio9+RJICuck9DesnsjSVZxINl0ti4uo29
OyoZp/1nOMjoMcrStfcI59qe28R5O+ICA9I0eBOvfp16DpiH3o/oEFaLZrc6JxwH
MgpFz2KC1HWypZvXIixTSLfdh4KF++byd/53RAjKsWc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7696)
qStoW8IUl1ALaMEhMYhVOpO0rj53KQjzwJCJtbAt099FANh8PDBgnwDI730/zJ6F
LA8w6C7psBgKW8smcVB6CRP21teyJPuYtR3w3s71mgHmDgk0QoSNJSq5lO27DmNY
SEHxl8bNclaqOjQfid+1muB9y1JF/VsoL9O/8zNpet1tj7qDmZco+UtRUNfVs+1K
xHscJKWSjG9FCvlgkLui9L1DdJuSYLXPHIYSrHkcnW4pNNsKFcGhKV4UKSy0YlVh
lC2MmHuXEgqBsMrfEveksDa+fECZV0B6JpVvAcAPOAJIes2S/vY0jqcktroovPqh
jD+ws4tVnJRd7krVvWl9HvFX/K7jsVMtSK4qLw/SS5tf76/Zvc+jGJib/9w3SskM
iZqhvIHwJVErQhyHLjGLszwJYDTt16dfu67CKb+lFWmc5whVsZHD+9SOoY/4X8lZ
Nz0ze0cQ2vprIoK0mnogd1fYiFRJaEBcoQGi4ppsoCenMCqHkmDTKAXA1WZUtHtP
pqJVkZjoBIBhVoc+XCQpFesTJRbA8rL9utvzonDyZcHRrzbWdIdoRils4YKGrkAo
dt6ryyHZO3AAfkb/YxixeqcLvtrSahcwu3yCgZ/nRPfGi9jeNNUdFQLdtmoYg9hp
irbNref+tpA4utiQy4NfSKvKHyFDl37rDELr3tXq3n3nIBeee7FKo3FoAhgYn8US
orFvdNSedbndMxUtccXKMWbqepJ7pP4yyVtd7gUxk9OAA/JFY56LbeygNm5soF+H
PXtu9M8OgpWmZpCeefnxLK+cu8Z/BZZF8TifkkADaUmKt5glNJwHstKL8SEKIijM
CeiCyL5swc1XjqTD8DeN9RbDlnK0I6O5ITZ+zXI2Dos+kdzOCvCP42J7eE+90lQ0
J1662FMo3/kHSJwp3RfR+j8zfeSeRygkQ+gKGy1OPucLg7zr/FOxp5jFyjij4ngy
yhGi+e+ZifqwFHGnwf8tg7mLbQ7SOAkBvbfaXhqlDshqs2YeO8QlaAcF/dqKJuCs
5joLdl3Kk+vomSeSUeusp2HQPs3giBHee9nrrR/jUjfe6bg7nYqibOC5GNl91RfB
8M2rLJIjb5s6yQQ3r3uxjsIfowx0Dqtv647SAJBtmNI7pBSg8aMCqMraCOdhqHZI
Ez63Gm6B2py5jUsrR2rOcypQV1IRPs2Xs49hQ0/mkZenCs3yDhiBR01bbuPsUBHI
HXLjnXH6++j56b9m9HnZKrzxje474AjDekuqYqiamd2y8Bb1SiBrzxxeba0d/Cxu
hpDHNgtkmydvM57uaXrw6VDBCLq96annvjXdeMWi90d3bGG270qYitCLgkNF2bjn
0pbEgieftIPQYczI2yLI4m1j/3GTsMu5q4I371Mkv19yg/mVBw+fPAPM5DYDIXvj
mArvM/iSvhxfImIpakXOn0eyLCV6IvmIafnc9zLH9PNRJHpuQ8flW8rpm+4UOHh3
w/tbq7XKc1VfDyDM5xn7jMVn7AOEVE/uRmRbaf6LHLC2FhxQ+tdGVspBpIZFvTiD
t3bOZhfnHIb3gLBtgtCezfFgfCbxSObwZ3H0OGMBRWE199nFbUgWUWevyeVRCMT/
iizPBJhKoTGjj3n/hOf1UsV5WJTwOqA5M8Dtow+uypTCwk/FsTjLTvW8bJps2bsg
bnWLXEHTk25F3p1BAPt7T6IirJWqCD5XmmYNqIEa/9XAQtlcPT8E3Pb7Ao6KOdPP
2OdtVLp3CtTm+eYriILZIxU4ood8ykA9046Y+/8jJIuEkrBNrbYTxeS2leyS5+XI
hecnfjbYuPiWV2olQLCh4VgtrPKnKlCBzJR3cxzinIF55uioANIaUjdCTJ4AVVFP
AH97n0gHonG7u71QGrSGlMKyOTsrLhqKnSZyIuqXyjYn1FiwdqEXTu91dDbtVdqB
mdZTKk2XPRiKFJRf0qTyvKV4TyZgEcvnFqwWF21ijoSldrH1j7Mw0x4oCXYp/BD4
dT8QSaR8ZSzcZQ4RlUyMp8fY+S9YwfsNcIVw+ns0oIuiK9IR00t5Sjfe4uXQObPe
5u5ljomOeRNW6yQ3S44tI2VJ0oN6kem5BunBO4yp/ldfOMJFrCPtUj/Zv/90RCcN
WzRxF3JyuzNUZM0ZUzVvnN2MBS5VdmGP6/YTlsOIK4oROkRUcnEAqiLsAoKasWuy
821uconFZ3EweS5FUUIs+YrBP/yDy44sAIQ4HJqDzoJMgc8kQedw5j02ZacpeWXd
qxPIHjDbw0QNgaRXJyUB3zpfpevN83lHS/Bcq30ZvvTk/hIRvEi4n6rIME00Vy1k
f5BW+PtjrHObBBTkDxMaNusqWNxhVQlDrg5XFKLYGJx5zVG2pManxU0H5qQKFsfn
5pmaqc0pL57PUcmQg965hEIssWwUCDKtUXghALM8UwM7JXvRVjTFaaiIpKT+jOpP
Iib/YqhreQav5xwNFBWfKtvl2VvbYhUuchTnHeyVbF8KXXNXf3f9LRveUlyO8/qa
kscqcee8BFmZrTxyveafNj+GC+wipDVwwVMGj0/pHeBLo7ZkigzUUUwF18vdYY+1
mnTILiMiXPOBIVpp3UwQXPdsMJrlqErUiGYZjIaVErJWUqUaX0IwdCiXIlu0fmRV
xVlCmK8wa9mVLnjDHcYYAuWqH5rKErPqdEyvdA07/8oKZ5IrwerNRLbYaYr82xfs
hgRxzjv9tdXbrJDKDxVHnYEfKbvo36Tn1EB9TV8hz07xLEyNlW60YyyxceRdikW7
L23CqNyFxzntMZ0q0PRN27XAM85XSA61ceB1GWbqvQHS2qCG62b+ka8qJt+r4QaV
Ghg+uIyyDeTg1fM9w9XPbTMy45Mt+NEay5Aqfaeyd3GqHsA+4ZDZvyMa4RE3aKOW
TfJ3ZdM4tJ2qazsx28LIwlTElOViHtax92C4ZjQNZ13S+UHECmoT7sm0eYTlAlcA
i6SxxIwUgnTiq6zu3d+E0/p0kP/WnjuhwuzeZx06rf31RAGrC0D4MIOJBPZ1nCka
n2sBEDI69rRZfZqCe2sOVttnCL5vplV1FPeQAC9avubCETZG5EKVQZcr1bUISjMX
xrmNKYGPXcHOSapMX1uN1BTXad+DyeHflzQ20bDpf93nA9aLwv4SZc2dbTAXsGEc
mmu38KeiqQwlnMSIkl96tYSyMOHoR/sL9iFPi2QzThXWsh0yOW8IMsbzgHVRP2lA
dOBK/okNeGJj6XIRU5B8Oo7cJBj8lmIBgfs5QBDt4Hk7+/DOBkVexlHpQL6dJBmI
JBdYdrKwYXBs7qOqIxtYuMneEO+21hZPS+UFA91aXfB1nZ94z3sUmyc1/SAlVEiA
Xcp2BUpo8n4UyCDPCSwBVtjZuN3ONw/kd6oBm4Q2M1Z9Y+X5Ng2irwgbEqfBlwFV
Slnh5aSmHRrNI1Q2bcdxlikDWEKtf+0pFocOoUq1s7k/sdadwnKHSAOy8fABJpIG
h6OldYIKli93oVQIR+g8htkB6qVVjmQ9fT/edKIs7U7ek8M1Qf3YwBhK3sWneNwA
NvVZilz0M3NRHWBcV24+Ai4x5b7/cx4fE38/+GRCvv160oCCWVZuLA8vVJZ0o3cj
Auv3ZKFNjglo8NpbcraNqMDZz+OEP1pbcb2aO0fTNqWBDJu8e28DulCxguXK6YRI
fwa3X3SPntK2DWdVHav7a5djnAiq0CKyNp50ONvcrcjwuvbuwMfTWdPvQLq7O1m/
iFlPsNiuuWDkvxh/nwPQvbABuNMzO4P/nGrg2xVHNdKOGugaDRpGgSp6V6LxfQop
69bBZ49hgxmxsuI2Z3UAxyhv568Qf2VVfn3EMYgjZK/6SV3sIuylXX44ASmaU4pP
F6JIeXf2r+GPfkSFsjyhNvZODP5GXWCmHs2dvMME4rTiKUISoHUmh8/61kgU+9de
YOyAhGPauY2+D6TZXuCXPGM/pxC58oFiCvJ7RrBb0q5EDd5eHz2G0SYl68wG9T54
JzfuSc7F56Ms934C/KsAWbMtlllZLoncLEFWJyK3K4f7WE7CnfYFedjJ5elBWDOu
QM7rsHpl2ubCf60mvBXBJuOyEb9o0yG1UqzazOsopf2PmUUcq04/5R2sTNzHIHra
JjSHV+UD3z9hYTl8wQX1cZoFCXY/LWJLFjeSsv4zrgl7B5CF6SPDrWfcX5I7WDuM
CRqurtx6Dir5HnfPVxWJYbsERYEs6kBA+Dnn/rGkLHuR+Ej8yHzbmydSJ+gXIYal
ToRJDbAMBdGkt1Cpj18Vxb8x9eipEvtCerpieA1t4RpT+s/sjo0Mr1DOI6QLYp3C
sZwAOmHJ2Kb1IhXnlscl9Vlj2WCiBK0hDvEvk4Mk6ap3gZB+Y7FGd9OeEcr0QH/f
Z0maRhl7ordEGjryIGSvV/oB2mvxyqYKN9ZxzhgiDxIqgvW0tcj9d0P0mTltELvE
B/YQgY7xwNFGQ4MLoiP5wlY9vXPQ4dNuL4YUIAGttQulrHQgKosy/Le10x2xdJ0G
UfQB4j7mQRsKQdi5OZ/qTNuIZwMvg4RmdWfckAF0lZjPmJHJwN5F7Vjc2UZO3Ab3
gs/GntBbrY80Bmdf5zMdAqd+LXTNTDCzgwKdvND1Buw0OrnkHslCXy980TZHm8VM
yK7dOn/OzN7bfqJEiBir6iITr1ixU63q+ikvVhuiwUTkDhTDuHCc12ksIBW8VGnS
0gx7eRpY5wUH/Q/2hFgTckx3cWgKaDXRml4Fkv+Zl6CtnEWzunPWwMuDElIBz7ws
8ayzFH0MLzPDv6wiU3s/iKBHRBiNHqka6L25kzrTy8oJDANVrCpO+h4Cey6vJs8r
3Wiyu9O49pACS74AOXsJbN3+icyLS1eaHhxH1+qKt3JALobkmXKr4rN5h95PX44S
srkT7cvGFY/qJxhE2ga4UxR3OdXYdfHyq2XWkwP3GWIvUBLBg0vD9U28p1yiNzw3
AWQzBl+szeBWxrhGUKXaHewMP6nLM1Wq6giqokqf3aUTW2ZaM0dNX8j8UTBjhISu
ceyrU5FQk/1wIqO/54YC7dQeR9c83O0CR/vNh6Fn5hyJhkwkNduyoS2cP9HkPFKo
3uPCcEVY4hOZI7/x2KDw6jfPwFJcTs5ykIbeAcIfR3QcfNG3QSHnJsrOI9lD8FfD
1th2pHjyQCPZs0t9cPNzqPshoXBjhl0aZQ6sa0wGARRtWikLHWaw72Spv+1xNgSf
wnE1CYZUj4NSTx4SbIfSeALjdxE2vK0XfzfsMx9xucra8cjoufLZmPRmqUihzv6D
l3CvqU3J02ithgjwy20/7X7dnhT71qGlmERZxDhYQsVs9ej7HmVPMTXeJWoxs/cy
qGinN0lED5SzIyoyqaZ9hRrmIQo8Op+bdLTv1PF8eDIdTASggcm9GlSGc3QCeHsg
4MYtqddczmOItVQfS69osI+ctInsm+9QTtmVpBjPvaxd17nOtmwOYXjHR1HSNltq
uF0kMrW2blUkrL+V4FLeZjm5ySFhWfe0G/DfbWBRtRGSAmgV2lB7Qw6JNbpf1SXz
R+52GjII+mRhClLKXoytlM3se7BC/yNRmVlC1HCpFwN9Av1tng+mgHIGU4mW/6r0
gF9p9n04dw0jpl36nM7Vt1JKGNM1IhrYyTHZeWlO8D5yACYQRsyoavZdvC/2QJhu
gpUhB4EPGjJb+3GtALNupTacHQKZtHBid8SQB0D+62I8kVw4WixhlRFEdBuURbdU
hoS7yHy9yCa+U5ys1wV32aBvtFTd5jkLWLuO0phM/UApUZrijAB9o6ROi5AV6K9n
43cdx+IoGBDai/Pj00uBE5N2QNrO5ebg55YIcBIQSJVcQKF906zsUHQ6f8bS+z/o
ZmIZdledP6GdJF9ihs+meCcVFTX8tyjVf+CnA6DsRVxkVc7xxeuujyjpCyEAPDBq
hu8L+T0lFW9ABqsswTZIbMXmY2v9Fpqg87iNxVuWBGXkJEwehYGETCRE3dkc4Rqa
YlO8Gv8r4TR+Ju0UDyciHIJ2uWcjr2w59XBhOtw9vo6KIHxyVavSp2D0aaABwUCd
SrfUSBo4ug+XbRcrs3SqmpQMs6uoYJkfu628jR7qSDsTGB23UDVF2IEPMowRseaf
RbWCce4LK//WuLXfuLMsS2oSmsvt1jPI0FqnLBju6sIQSyIKOn4nnWgkZA1ywoxt
I2Z5gh9/7xhPOhbtaM7BrMtP7/nI50y/3oabT6XWiIC2IgJSO0NQg0xGhT1PnLz5
57JHyYldSGmDPJVaihnt3vNE5Pv6+JF7PEDwmtkKsYUnjD8LtoUQoKMPzbH/ZVsB
dy0lhP45+45A+OaGAmUrb0aUtGprFXUqGujheifw9LZppP/aG5fYs1dtRfhiixN1
qeIIbG2HTy7WtmXfqI0z1f+VzKJc1UAZVllN+2CqhNBlgo2nBsfxhbJUHoN6NQ7b
SLGAc4NQ1QPeZeO1IUtDfazz/AjuncwZmMYcVEmPFtRSPTleTz+vDkzr+C3hZjfs
upDUvTGyj1vtie1IRC+GkL/x80UvmwC8HxtqcRO6OpHPI5AIxyY9ccBFShxsXPwk
2mEZ/6BoB//eBBoI9/S12mBpXSNxe8HMxG3Ay/CKg+zoaNUnZFqWR5FNDdE5Vdfk
1VyIb7EdGm0T8eX4+RHn/YdMrXx0dDwTo6U7KhYBGeF3H4c+w92vbu++Oy9Kd8Jl
gNRfon9P0mzUzGyg3EHl+Ttv79pZA0wChGu0woiFUFAGBKv07mmhXDyvR4EOHONQ
WKy9t9b594lDxMjeXDii3hNjQ/luSr6I8VUEO3BhIFefEQGvIsyogGnn7symrhPs
fCNQqz3Vn2vtPgTzLEvUqYThblXitJSjq/52MExaUzDNTOzGIuMQY99COhRn3GsT
9O8wMiFFPNWEmX7kcYZTvDX32iWZAzkiQjDiyCUOPJxULbQoADouitejmrrE3Ful
VSXJ1IWCHAmZ0n8SyhAKVd4SKFCt8AeWerIdGzw9vPq67QpIl0GPPpaMsOGseKBo
tUgkK2immXl0OQMIvY1WjPadQ5E+vV01JnRbXF3TNlDUnHrnBXSrk1YLqdL7hFqT
jHBIs/REOWMKLjP/WxnepiVBARA+agP3Dnbw6hb9gcoNqEXwffW2z/X4T0QBpAfU
iIqvQCi/T0yTlvLkPMZvRwg4m6sSisfKDzN+T1A43PeKppN5/12/itSHpy9pH140
gvKiRrpBRZ1C9SJKiLSYnUKPI0AYEwcFw8izPIYiCctRqJeF2sS+ep2oA3R9uuM9
YZ+i43R2NwUqvgdG3Qu/m7fUkLTGv8aUb5seo9pKJpNkzUf70qBwf1X7dy8Hc5/u
S6VBBSqVtNwQX/Uy2X8inqjGW0vYrnooAwnM3abPE+ufbSKkiY7YBEHpv63qLzBY
IfhCXsnN9Yy5VgaSqbbAy/41NVa+Q0t6QNPNBM+NmGN/hU30PGTRATXeIbmG8K/K
lnpL0Dj11SzN8MBafdtpwa41Ag0FGjAXJxy3Im9hXxUpwmsAVVB+BrHB0M2RFp8F
kWZUxV8PWtoCOLwHenghfhMU3w2p/c0/hf8Ov3NjMES+EoGxrkG0yCCUvZViYzsz
MzOpjuzESW1dut2IyTUeIYSz4yj7ZQ+O1iHucUwSvCybI+dao6WpaacTRjEuDYlL
dePe6/Ubq1Ybk72E4zreZE9QIRTUXS404X3Dd4KmaQ/G5b33Bvhg8Dd6WYNPuzPm
qcCa0fuetPu2TwGU2fE8YWhtw59LFW+cU09RZ8Dau7N1HogLiWVDC/rcl0T8RwA1
Pl1dLMnmpjcg1U/D0XmoJJix6g4uYjBbLk2G/LpvwYeYENzk2Glgz8Hwduec7gce
YL1pEIFh/r7J80u3u8d+UbrQR/77dZaUJKDisGvITOZCXOo7KkkO2LYCAcNzTMSC
uOWaYdMHKiVhhIB47hHwZ9mfKr1cYiITAn23jCb37tB5UFA2xsHjnWlm5aa8KvTn
GLjNGBbf+Qf0KePtMS20sM8ak41OPT/Gn6PDfN5HZPRLFBs07wmU1+f5BAzgOfgg
eHQDePXI6FG/p1Gyw5ZjnYyU8oE7me2NxIIIx+dJ0fRBC2YD1RuVu0BCY33qQJuc
RGDHhdqtYH1BTHRrsIYkCNk6Hp8aAgLrSyaMHfGJGQmtKwDgoqGU0Nr3JbmBjxE8
+XTZWJBqu9KxhcO/0BMOYOqGS7GjoNrBUkCbVsIHaHMPrVMDu+xIZvLkN6KgMfx6
B9cL6UtwH9fHosxAfBYwb9jRk0jBTaJ6Z3wMKAyTwSghZAI3PU1aPS59QQUqSg+L
A/Q27CYmrd9eyJDzkykNtKROFZc3eZDEPEEvAsg7OZxeKyr+SlH24wel91Amn2ih
EjHfHEqYyTRlCtPOV3DrbgCglhZIvQVyZ4kRvaZUO77Jx3PBTPM2nRlv8jEo1rn7
x5UYiNIFzjGLkg4Jixzp2JikalYLSpHIsUL9kxL0ljK5lh4H1nKZB3zA4HVG94vO
HvMz6cKWs8mAnBu1nIOmc4b6qDl9VTBTP8H8P54bI5Ns9mnri/8THXtN3CE841Yl
rCuirxvjfKc97teH5m3MracjUIzPxLiptzOLytZqn7/xzvAzzgHMsqrOS/cGwekK
I8RsbmniuY6VTH0b2u//fQCY+UVtQZ8PoNlH+Nt82DpaTGvA0o9fd5zj6svV/m+e
VpQZPgmAY40+mGRVSTMGTwlQdwr9MA3d7y0VkW8S1uBR4QkEYtQh7fQkPsBDQVd8
14YZCNJ/40ne+0lwCgHBpaOIbcMGoCc0yVbXcXBPU7c+U5R0tKFDzradozEk/Rcz
6LOBa63/0/e0Nvv+UVcuwgSswlHVhLY+YAnq/HgeF1NWlCYkd6Cl0DElXOSVOz+b
IGe6jgpLPI4wbz1HVJUzX6lQhovfud6sJnpbyfV59YM1K/Mw4swQSzz3lbvcCAM+
i8V8vm7dudILgwhpuqol7BbFW/boatZ2oQEBfm75RLN7Xz+24N/bn4zzHO++tbkb
dslO4SVM4jmdYRRTjuosKotq4bNh7lmD39rFZHyCnwALiOlI4b/glnZ2mIK1qr7R
4yJhSTg3qMa+lwdquytkLO5Ax3EH0yC4jsO5utUQQRlf5fHZeiirpPtsS4Q+uIwO
EIdjv8jsXZQII/W9sIrMgcok6x61pit2PaAV+xMGPKhWasO+q29rqbijKMZY9n5h
HKR40r8CtBxRy/mJ0heyqcTJ/GgxoBE0MmyTJYJYX7WS07v9Cdi3jfq7CybbUGeb
WBu0quqM114yiby6WCB2oi6UpfjL78dbcksLosqMga1GwnR2xaBSWEe4J25Rr0ou
sdo1uBfdTA5xYYxAp6nlCYRZ8rIFInMIbGfNU27boehSfBb3546rFFhieyj7Kcsk
LGYUEYvq+nEN0VDP8/cSHB8JVBhTe0TwDyx7Qln5Xz6iX7/V0gcmnVzF1yilf3V0
NJqc+EaMIuHm9LA+nS/vw7qiYNY3wwtDH/hyYYzww4O4AHpRJJJBj3jCt2vq6jmb
E4HJGMwjntMJgd96SkrApO5as1jXx5VA7JAgDnvG72n4Pg8zukambghP9DAc1k2M
1m6eh8DPO2MEh1SoX9J5tGImsoIpZsPRrXAmYzgTQ8hDAdWLdbfBXa0KiqAXVd9D
6rHpKR26RIHh5Dy96Fs56iRUe7XNcGfcMrpDs14Uyh5jGYLTsr/f7Z403qDyyWTj
PwzawpuwPA4sK60oMjjTNtPCIs2g/yWVGFkUfb51SRwqOUjXMoamraFVmnXpoTxa
vnT9tFKcc4CccaYV/PN5WCzSa8w7LxQnoqL0hSYVgwb6eFYwYhNNeT+bgyxMntl/
xKLgNwY11kIGWf1eHC/8BYDwzg2HW3b5SDGH+pWv3bgvhLI+5BgODf2JYeR6Conr
I4RBx3CTaemRgGNKOpboAYULVhYfpeN12e2Q0CWKVJysu4Ch8Zm/J09dj0cFFTzV
c0FaNE4AQxr2Kw/rpNARpR4jwmKj7XpL3aLBoBAOaYOcVbSpzPVJ2H0BnqMZXL2R
l65mldvVzyukQ5PHuQUXxO66B2haNc2vPZPWyVHWrdBJ8PVuPlQPhF+l8tIOUjGW
snAKGHCuRT07Kv44xgrAeU1CiqSZo7xvRuly2vFY0Pw3HR3ABR/7gg/rI5/qQKG7
en/yAfoFHnzrQlP4oaikEF0zlYIyqHwHTGifSTj1mwFQOuPRPkP1luHuJLj1FMNc
6fkxicIq1QTYheM05RJbppgTXSxMHZskZY5fksYuibYAZMkhGCU4Pfu6QT2JO6NQ
FofU4RGNb3v7LuBE0raliQ==
`pragma protect end_protected
