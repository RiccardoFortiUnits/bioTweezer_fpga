��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��x���9eS� ]�_g�Xh3��1��63�A�1{Վ�eb��9��d8_��g�G�oWs$㩕�䫀�*Q���7е?-�@�Z��.޷�0�Ȭ�*
XL�1���-ec��D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2�}���i뉚��Tfp8;Շ�-{~aqag�ES�bl��뻠��,L�3�
q���/R:��M�Kܔ�[que����u��H~�6�,vS�a�#@e�BハQ��`�<f�
��Xt�ϵB��9�m�sϗom��4�3iY'�יŮ����1�F�%�~��Z�~��ҋF�g�nʭNW'��S_��ҶV |)	��';f������%��h�8��OqF6��h{},n8��ǝ�aB�S���̓�R�&\�O+		{�o'���~*zI0�ֶ�b�v�E����d{h�����s��'�!P+.��/����+��]s�nIHǕ��� !g�?�Pk%��^T�I��=���_�O���i����6��-���+P~��$���C���ƽ��Ӻ^�h�7�x4o���f��]�_�8�?��O�XVo ���mk�p5�?2����O�W���8��b���zF�$3�/՗�sKK�z�[0RKŪxʂ�v�3zx"�z���h�V2�j�v�3�9¦�����Z��M��2��5�;�Jj�crh�P}�̎@��G���fv�+b�J�'���<����O�G
v"w��<#狵뺸�����������O�E�_��5��XAok��N��Sc#Y�jgd�ȗ�I�������&ѕ;�
�ᴋ�T5�8�ՊfP�.�n���<�v�$+.������l �5��C��' ���Q���n!�2��! ���}�t��7t����5jP.�m3��ٍ���� �9� x���<O��~���1Z����~H�֚��ٜ�bTM1`�0���
�NzJ���'xA���u��g�E����>x��9w���B��b�kL���T��Z��BV�X_�u�4723v�I�>��}�O�<�=��Wf>����>p��Br�%�yA�������c��(�+�������8�"��D(0����|���|�ω�؜_	�gE�F�-��0�����hK?ȴ���z��<����pZd_��;�CP:X�jS�����gSԏ�j{�9�Z]�UL����h���Y��A����e��� '/L@��ɕ��)]J+V��҈S�P�z͈����I� �e�kg�U���z|k@��R���o��� �k����T�T"ܭ�@:��+�d>��H�'l�~ad��|ߚ��#�����	��)/R�DݩR�9�5����i� �x�+ �VJ�	��� �.a�ė��,��1�ս�_<�b�ٳ��Q�4
7���%w�z���R��sa*�K��/-C�4{>��pg���w=�7>���rr�Q!�u��g'y� 7���T��`�%�8iĮ���mQ�H���W�y�O}��O\QPd���ހUR�գ���k(	}q�ܥ���
?�P�E�1P}f�@<]a�+��c�ֹ���P1Q}e/Z�!�_��DǄ�{�'�i�/��*�s7��
�W~�	�M��4� �ˎ�e�߈?���ϯ���N4n<�,FUҗ�󪔏@cK�K�NB� }?���~ӺE���s����,��_UQj7��s�#Kc�6�v���d��{��֙��0��P�5��%�$$�k}�g��`��z����s�pn߼Z�fn���j'*���׮�F���!y..�d|�5
���O��s)��ԕu \�M��֛��n�`[�3���H�zo;Bo�S��ݤs��?��/�*��\�6	k���N|@ԉPbįި�]����!�v�}Z�f�����j�������zR�`�P��w�'\�8�S[h�	�nv�@�s�����s������.Aǻ>j-S�o�i�N�l�t����m���k�a�1��Z�]*y��AdY䏮Hz��v����)tR-��{D�$ٚ��a�Z��B�_T֜$j�h�V�L�v��=oI���l/��A�y�0t��ݥ�ל1ݧxꭵ܉�Ӆ�)���)
��53 x�ϴ̘�l�(k����Z��oT�O�!�kE��G�d�q|��~kw)D��hʥ��r�-q���ܺr��'Dvz�������z#�����;ۨ�qM!!�n�M�À��y�s6���KlZFR}���2�7����ՙ[8��6l�b`lzrO�ʍ+Nܡ�R�x�?�Gk����>.y�*a ����􏰃�/�9f`O2�<��mz3ϹN�����=m\X6U�}2tM����ǓR��Y&G����q����Í\������C��&B����ࠗ����s`g�c���8��%�d���'��ɮe���=��
-�\��1� ��!8��6~��ĸy�V�EgG�*�#�F�اA�RH�>�N�U�7��(��{%4k�U��o��Q���Y�A�6"���
ܞW �Z�05i2%o�����B3Ea	��.�x�X5m���z�B�r[]�;��{pL�y���������J�.Q�3.
ES��&\O,�>v,#���?S\�QύKT�/�7,@W���4���3��VH;o���GZ'�r�1�m�aҏ�-���I�f~�y��+��
��X|���b�!����y��(����~�I��7���g
o�V�2B\�W(ES$Lf�M�؏���a�d1{'tմ�\�~�C��w�0�j��=e;��M�9c�n����#�UxY�ң��v���� Q����FX��>��뼤�e!g])s�B�}7�
�d���s�(Z��0��a*�|a�V�-B�4:���ق�Yl@�oQ�uFU*�4J�MC��By�:U)�h�8L}�f�;��|��T���_^���f,��c�Z3�/��=��8%� �B���J_<U� ������#�q�c�p8kV����	v�r_8��Cm��L�
`�^�J������?"Ȉ��ev��>��4�|[�J���"%BY���Hr5�M�
�R�<.5���������pX���Y�L�� GK��6�gs�HkEt�W�zݺIAd(y�n�v�؋�qj�q�0�J�8\b������:	.��I��Л�̛��ϵ\gf�T)P���H=�=�����9�����?�5�Q(�g�KDN1'�z=ѕ�C�)�9�\"�؟=����8h�m��sTv|�&�\��ی�L[�*���?r�j�6((���h�xwF:���D"$�Y9I��(�D/��6NA�k{WB�ز���	�.R�
��uw�+�0���|O��/��I���A5x�}�1g�����l���;!�P7 #�Ғ����Ӗ�1�"w�m�I�K&�	̖r����F�@Ee��χO
����t��?Uz}L��--6��^8�+02΂x�m�C�%�EzM$�b[|���\)���a��D��~�k����y��+�i�d�i�il�����Z��w��{�ߡ� y��� �h�����$	��=���Mc�m���p\w1�A�Waa���l;����[�7x�s��C�ͽϵM�^]ߣ𔄅�e�V�A�Iz2��XQ��ѽ�[g�gu_d� �>��Q���4&��3���a��>U
q�)����)43=�ŭ�P���]

�Or��M;V,6���/�/��-_[	6<��tC�?��)u{wf�������(3+����åKOX�%aa��%�m@���BΝ�ӷ#DZ��eزÚABKv�������Y�t<!�m>i���&j��Y���� 6�N�J��dK:H�F�>u���Q_�'��J�k3|����BX�����A9��|�7�f��05Sen	�3��Z�&������Gjk7Y��綏��y>pz��0�`!#Kڢ��<��f�����W��eEڻ5o[P�ۄ�yfp�t8uV��v�2"�����i���!�v���^�3@��Ҡ8 ,���8�P혟H��:^�8
2O�#�E��Q�\���{Ԣ�wh��H	�~н��_+srm�^G;�K�_!bO��	څ�MK��T�Q���f�����q��D2��j	����1,������ F���1� ���-$@��F
C�H�ꇜR�Ӗ���klxYL�K7�����<t�re`[m����rC�(;���������r��,bPv�듥�N\�feF�E�c�4w���9�2�Vw��c?�%�KL��-�|>�pR�
��+��Bh%:�ۅw�n��������0ˈ�x���4�f,)&Ln'�F텙����k���T0H��uGa!4O@�&#�*�(��x�G
�&�D6sS72�J�ݺ+KAʍ���/\���>�B���l�g�p1H��{��j�o���P����]��.�А�n��h�<�r�������5��~S'����S��8��p)t?G�<Y��A�ETa�ύ�V���_�(�(=��Z�'2����]կ���B	;��NB�ژ,y��j� ���2���O�:6�H_D��ף�f�:��k
�$^����n-E�wr1����i{��ǂ�Dz���"Z��Y��-ò�X�U����I ��VԹ���.=V��g+�J&U�ȟ���|76�=�#iG)J��-,�Ӽ������
������"����K=W� ���쳄L�}���DUZ�u�����?������I]�K�Ȟ��GA�^`W?e�����F���g`�%;m��SU�3;sY�w�"f�H��0�VL����h�X�WL����&^ B"0
��cjE�UT��zY�����7�