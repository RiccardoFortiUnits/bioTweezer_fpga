`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iY42SLn75gYA1aEBGxafRnxZyX7w3J03RrWC4j74/qpNvf90c1V4B8tB1EB9NszE
awG1tm4KQjHtP7Y7zhMqB3THI3H0vKXzb/xk5J5fhT8ry4jMCExjrsb/xv5OteNv
IugKjQD/wnszAgTAIJFjcnKcyWJczO1pCvLbAk0jcFo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11040)
5wtfBVuciNFb31y+VrOsc1C8vb2D2oXv47TEbG92EgWKeM8RIFg0J6ROVIjqVqYc
sCMRVtA9wA4Jcy52/yfBY9G72KGG91ATWtfoornhZLF1MmaIeWxEE928aJ0y5H8k
mFRI7GEXZkAGiVApzOS/1lrHhl6fsYTUaOt5o0R37OC+PWQHa/wBqLCfxp4/N8sg
RHyOnUPZw00zS/JroQKowDx/cqkkXa1PLJH/iQ0iea4/4r+uF+ZBmHT5KxohP3Y4
CxzQkrkGIMc2OMVoT4Mnt5c8fDPwBx+/+/PGtvtG/ayMsmWwjH3Ye9SdF88GCgVU
bCA6HZPqmVNCsmP7gdBRhfHeMD8Zx9yUEB6tJNBkcdnUQelAVQXI8I7HvJxAWEPm
+u/wy5zccE8+xe0wZVl2vBS4Q5dkoZrRAYnnskk7QMscCd1FVS7+9G3k3Oo02xzE
6Xs+/AwFUszE8tgDOa8a64zsswaY6WDfYfYqOJqMtxW+WXaXKgS00gh2dyT6UoT1
8VEpmlRZUy8F9rTmzi2v+akxDmd/sVzRUJIL8zDWu9zA/paB3P/BnODVvZQhtNYc
zkCocsmN4XMUKUTXOreGGrIt9lPFcNiTL1qLU0iWnJLOpsjoXe6vr4rLyk94H650
GM0ccsBHkghn2oWX7ObXeQUhul4caGEEwHKuPcmGs70WxNmHuZxs/6s0DM1IF/dt
gBY9fU2s3SDX7+cKz/7lapd0vdejKuocQp4j/gY7s0uqZCQMRJtyZmH2RdWjTKjc
hRHNSe95HLiiuZNbmWzyuPOu3pStfutSiMn9SzsXpFNEaNCADt4CE/h7/pqH//CY
y2DAgFtzk4v9bEVucUW/ip2X6gvdhkXSjTgv5mmWXC80tHf4ZXeBnTmWlQUgNC3/
j0oQ12EFampTxZHe3hLPcFkWfTrJpSsVjgHu06/UewvhOx++zQlar0VRgENBWW9x
83X0sm6p1wuMPXSHQ98/38OBpRNoHx31ABxeM2rXZry87e0sYsURsEfQ7T6EGeJ2
oCk3xXX7QMZ0Ks9SDVB9qWXI5lT83i0d5cCNMcIlQaW0ieIRElcAIcuwUEVivKLc
BR0BxPllD8Ruj0kHdJ+OTtDwO6I8d8ZG4rbJe7XcwUTaMIzkB57Fk0g+aDMv+9tt
jVsAc7nmyMtaTSgLM73hzzP2jWyS0fMZ0nmoXpNMBevMpTIbJ3kY3+Kjl2YRWEqz
vn60PxjwUxgsWsXuohZjpO5uLCZLCcxg+gk3mrzuTNsZfGTUj466AEEcGHabrBKT
i+QmPgoao997xd64RD++17hhEVgjYCANrPCCZcd5PRFQ7+tZVsIDRWY8ceRyBzyl
JRXBU3KojmV5Z9y2IbSzD08ILf9K50rtv8cT2m9qd9b+00ZkKKZc2MUluy+nBdib
UCNCguqNkqzczIZS2bIuEu/MFNobz+YEamZdVVcphaximFQfIuhLynYMVkoLB5ar
h5AdpalkMnUvqFt535kVTX9MhH4OCx4AiWXc0ZhDCo+V+J/cW3xOmQC/vmgO67Pd
W8ASC9kuLnRfCtz94yC7GhuLXIg47+jIH0XRQulpHmYi/onkZPe3AkeyYyLus+hZ
ndY7fc0HhQsljEKv/R1vtve/uwaSoA0DwPE86tBWyM8GmMwbXm5WZPM7VebFAAIA
gcSDou2B1nBtVPtG5/E+rflp4hSDWazhHfXnM51OzXNtOPIhGMOSkP7E/NzVk5yj
Iq1l4jz0B7wKdu3ZjC+DsDckrLxzPxm8cT3EGrC85aDcyH1QLlRoRT5X5WqGHMFh
EUQIt4gEg7+xrAEt/lDZ/4rk+uU+0zosVjv73DIB5PzfYoBJLGpo1I1Ge0ienh6q
mzY3Tf+pCwhk6alPy7GH9H0klp+Fw8IDqx09Y1jup9PnqgUCIhBp5fv0Yihen8FQ
gZ7Xn2dK3mGoI7AevzD5fjUcl0ua6dubbQZb1c/GupEObcb1XRgAdye9mNARVlgw
gY/zXVjDwKgOUFQcDPgX5bGCjznfuI6hJjZ+BUnqYKjhB37tQjt4WnzPhXxONxFk
oCMt8ImmPh/WXSFNVD2sEob9PR0O8l3UqIFPXO1oVd/q9ZPcxpTEaGE6BldMypIa
rU/IZX9yjBONnEvVrDUmuhjiZV6wgGDwovGbJcNpYvno0mWFqBmSDpOxkciPRKiK
Ir63TSTvo39Euky59trV7uFsysvvRd8aqmWOxb1nBaOu9XKgYhMW01E7ep7aGStf
8+52Y2Gh7F/aJx8RPyH78RJf+P08BJsGgzz7devFZ+qofoA0WePykAhNzahCn2Nf
UX5JSugzXvBqRPGVTrEAJB/lWtOXdE373j0oRjv9uLqsivDvWk3FqeS3ybauri68
Ed5Dzu7v+z1s37b1CTVx83DW/hoOcwhvSdTKlR/oMCPUXUbpFEro7dEbiTypPOfI
D/Gxn8YcayTRrFgYssZ3Od1Z3V0xFiLPGFbaTXBWAcZaVNiE7icaEjVzatBSmrtj
t/ECq9NNdmgtCnVjdf2GYaunGUlUk50YeYveXKeDuRQ8jejTIDzJBpPdBPxAZHA4
F3c8wd2hxBPMZscpVtA7oqdg92n5IfO7oeXAwpHgv7733W1XTlrUgAo5ineEUiOl
L/C9TbTvl0ylSpH6Zx2yy8Ie6Z7QCLN/+zi6sg95f63o5oYaAhOSkREYP+PeNAzX
X3WQqF5L/EQxApm+OYmAq5KVFQWyXu7bkZrgqH0YfL/C+E3no0FlXUMKhy//B8cF
K+EtzjgvSpAvGat+CVa5JBWtVse2FGpHzGvOoZqwMKG8HHgLgBBX0ArfugXy50cC
WV1X+G5jDAd9ndRYnMOWsxG7z53Rvqw+FQZXvG7RDaJwBprU7lvz/PyiA5AocTbC
kSwss+8d5n9H+y1xR0gP3+nI9LYVNo/Nl47wOwvzVaIRgXXNR6zQakY82GnXo2Nb
qiCV73VRfUY4PAMjeZpxzgnxcwoHIHUuimcU38Hd/WeOhRw0u3HazSE5EYzZ1bZ/
UZV84ZbKOK0jHUAaN2hcZBhCZqkNAmLsOqSjtaPJmHfYtoQBsRQ2DcIU/siRFWva
LhnmJGtwrSxYtXhTVrK2hx0Io22Ow+21G1Rdt+oJkRF5C7HMztMYhfcezONE9aD1
lUBFLNFXtb/jFJA5kt8YEZEgYWJNTnJVqtaB8gpZ9ruJNbYrDlQ/0yqXfzEQa/rZ
Ju0ralr1UDLdf/tpFOyToHAPaobl3R1+354d8Y5XG/sh/g7vFQWBFVmPsOG5dxHQ
lzgFhnneBwzN7uXelZsw1VCdo/Zj3SW8dm9D6T14gLvZltqxMMr68cNDR+lkHqgL
iydhtDCyy0qSMfSJbpzwokjV9oXHl3MLnjIU7XApd3tte16D+tZxd45ZPZNY9qOS
2RkBQ11cP2BxxQngiVzU1sZxjRRznUTo8VO4/K14KocYLHEDQ27/PFbzBN5PmI61
6LuiYMI5cDZsrFom2BO7R+3qrkF1XZA3PkynFqearb8gaLmJi/2VwE5IvafaPY8l
sMQ9xJfIX6n/JzU3Pe7ULSKRdHtscLpnw9UQ06zqK+eo55yqPkPcRK8FtvRBtVQ7
1V4DBlJKZyLohFAQ5reskA/e0QecZgqwv5nrabXZBRbdjkonV8vs+OfMw3XDOjV3
0xhIC3eyBho81BZeJQ4dhZ2I89zEo8/zq0VcPY37kAs+szy9JrasM+kEu6maYbRr
M0v17Jz2fs2RhINN37l6ZtUhNDvY1oxKA353W69mbBwpGmmsB+QjL7cLWLGkoT2t
pHdhQVPmV0nPpI4MGECkkhMXENT53uk2CIx0cr+LO0xvJAUP/ygA4WmEzsQFXqUR
b9rVFjbHKhqLfuX8+ibYR3Zosbaf0ieopBWpVRzKNyPlqQm8jJdsiAfKj8O6/FyK
cqwjXJTHJsTE1Si65ysMWOJcZJ4Lguwo0qb1n/J7bz2toAiTyKitlt6AOCjzJ3Rs
3xjzCN00SWlTiFoEB8Vmy1VsL/uC7IZqQs20MlAXX0QGPN82ndyHjNUgVLg8f6t3
zeSRPGMkxkyfCeG8+omirPcTa4aH39Lib7wu+mEkI1KrnTOPvtNzDHI8WajpPPCH
fSACYyyQ2E2OviLTeMTwFSYULde7vkE3WNuPjQZ24I37WPYjlV6N7K4hoPhSSOKw
TU/lQASMKGMazkU4IPnFJwD43E4ItASzHW1CmbLiAt26EIQzwhAzjX/eiSnBvdVr
sRsOvsAj6g8OggMW3cKiGtvuVAtnX+A+kF+eD0fzdKsRBVYdEfwCSmRvIwNnVXgq
WDeQiTNk2rNw3gZ9/CZbDi+7iiM4R1UH1/UWCVe8ILMmY0A56eXwJy925MNo9CvT
+6CJaEonfI4IiUEbeFTBO9S4mGBOqAvgH4Nw7fdGm6R1ROX8NFxJLdsj1cI5Gy2P
lClNkT4vEY4gFAmdbmskEkUbk/sL5l2c/Cyhg4YMeJ1n+tTtV9JiKHx0Gsk2jPfP
IllzXKG905XuH2GSQKxVKpxbFZif/E4QdX79j+R/Y8Sx4tiHxjrtx9DcnHHPv3Qb
cgjYUFpVhiiy4evOBtgswaHH0mz6xRYFdwjMGYU72DbKHAll2NSaMY1oO8VNrkqX
h630pIMwijfJDfllWfiCy8r/F9AMhEPX9gEebviWxcJeQ4tGJ22cwTQv4/yuOjmf
wZJyZoY6fsOXRSX14VgvDhn3L0Bd0yrupROzFH8sh+k3zInyWQLqYEuchPiVZguP
MPmlE8QsKFjKtqthT7MtJiA8uKZrF6qsH9FQWPpTMOWu6gIQTwFjCTXTzz5w76lh
TBrNBQAiC/GI7vzUSUHuIiokRJjS2x8tiBN3wbD4qxVrbvpsaWrKWQVkUoNGGoYQ
V++kU4LtzOnkGdfDuVfyv2DiZNwV7y2eJHu4HuhwAqitfqJswfwONzyDudYW7To/
0WwQeZf6RMEEvRhW7RMg6mQlzVvoXJQJXhojRLujiSHbGIZQFSxr2MJYgjxTQyak
MxDwOTWSaH9N4M+/aTtbk2TegGnz5Yj428IkCv4waOdmg90y0FCCUOtrL2FJux5P
eYQKMPu9YtZ0PwL95ZQMADDhrNEI0zcrUa5ac6HVZ69tZnZ9I7IQ2nVv1V/pVPwr
SN93859xeqGM6QkoJn3fJYMh3lWwZkrU1c02o5ii3O5G2vcvr+Wyt2yYv3mtUrGT
XvMpDAMLfeKturrZ6OwVKzj497mf1OeW5r5byzXBWn6HNsh+ll963mOOzobHFJde
yuazdC4N4amhqx9uBgIrYp0BzQh0AP19flc/N1gew8lfz/3xOh2YKpoON9Ng25GM
VtD3MCc6J7A88jZFXq7oCxgp5R1SUPznkrCMx0AIxeCM6MBEQ4hNb22b9nqBw7LO
MaTr5su0/PQlMedVsjWT87YfrIb8NvKw2+/LehFPZbgqZWQlVsbPaHv3u27pt5e4
mPchrmAJqLGAKlVORwcnBK9TlJV/OY6X+crw0P1t3RM5pEcywf4pct5kQYN2yru7
x9G23NffFQhO+vX0VQ5J55C3KayS35VVkhKul96U64f2YN3eQD4R1DYg/VsRCvbK
HUm+t6Yc4jhL7+mR2VXAbjDUl9k9oMEw87C4J0uOhxAqxcIa+t+g6ux2KfkFlhCB
PrQ0QEEzI9JfUA+FXF+Jt81ZU75nNNhh1jHrqGJNj6A/HMXEZrz80XPIWOnJpOkR
W3lliTVkQlKiF3SMrwzX8puXglM0k5JawXlm+DDshJ6T5W8TqpoTcvYFRLXecL+v
TmDwdDmHCX9LAS3dz2LrDMVC7nGpO9vI3YgeJt5sP4u0+HqBSrBmeVatOXnLjBKZ
JOQrg+qnAOApzqmllMzitIoE7I/bjBvdsfikqBq597CvCx2E2U6JkrfmYSv0yGw6
Y+DUQQUN6s4/XDdX4U5pGBwjGSBzqY7tqT74DGHxH8BnRg0OyeZwhw35LnCt7p1i
kUg4pyTMDkk5yRl/PlHPIEfacvxxRHqnVUMlunYIOgnb9Z0vs7Kpz3vrAZSzKK/9
KtsrVvIQjPbFB0HG2s9iRdITO4KB7mrGfDBHBVfK8aRVfWIfw94Ko8EiUFP4Folc
QuSUrGmzQZnTLs++Thrh+kNVskaTb2T/niVR/SY2bkEGKi3ly4siuBVFko8ojr9K
EW9e0Bu4ITI2QQ98pfR0GBVDe1UGuD4z2ooOnD51AsD3SABkltR9zmF9PETsRUWS
fM5pXCJtpnNnT23T7Px0lMxwvTI1jhqkXhaPg4MHzA5XwZi4go9kZ/9SlyrQQGZM
929XbgldURj19dFo1FgS2s2mvrZ9mFg6kcs/HBRU58gujTl35daKIuKiuRrzFKPP
cKkiwFpvDuS/wBdf3JGl1DvSRE2hh3LPDQyz75YgpU3pW3cU54/np689Sk9Uqa+m
HlrS68QaX+6nfPcEngq2c4EUIHHn3deGvKTnWZRsMHObZA4lRWKXI81ffwYl1poV
+2CKeuLJMd7hKmgbzf2tRc+0etk3KxXv1gPVoBzmUNGDGV7ZwXZwIcKvw/rMwNhI
ebliaqiQ9dxtuktz82oiQbG1KNX6gt6CM99DNr957qAOc+E6To8mH0RY51hC9dyU
wCY5FcXH/s2ls0OzzQFAjydqB36Hse0dEhtCAt9p67FFXfzbO6q3BMCwyEitctSw
lNZGdslqcLqIzODKuC9L+mya7vQI4ZERTzCwtoFjDkFokjk+nP00NoWh2CQSPCc/
lXFyDkt679hVBz0fluGlxZp84rq/kGAamuCt/z/kAtMHLo9OFQI7HaLQs3D0N65I
mnkBbvwFk9g0I9p7TD6tfQWz+lxCgqaLQy/nnE0zgM35UT5EqUOmPJD74IaHtcSO
MzfGnCK2WKd9jJ3tnWUZMfWP3+4cfKuwJByBelwa3BNfJgVHfw9tm+xg0JYg0B/+
ZkNP20K/Pua6fhy8TW6mpUz3KT5/wn1P0U7JROUTpjVlw/Nt4egrz4tRLgu91vyq
FMG4fEciRA52R1w4+84tb5L54lA/tA3tLdozDtLb41jw+KqaI7RQMm/jLi60hXrr
uqHuU+gOiQzc9XIrYJoNq0Z+o6q0p2xXp10I+6MjHYGC4SW/rlL+8SrPWUppuDHT
AXuF/XcIGidepF+lCtQ8fdRBtzzl2fXAAFGr9lX8K2pehnZYjmWwl7y70pGKOhlA
vfqJu3qbLk5f6TjZgQc5D1GcektgReRKKZjbYcvPoUtpSYLCVRIiYE1StETdXvYF
rsmE5VqvaR8dOyLQFX6WoJ8dbYQDvqjTQu4yf451GK+w6418VW8QO8mTU2Yo535C
+6jMqJSZAx6yvvcMmC/BportlAQo4wZVGJnZ3MORz76EqfxCveUhWkMacPEw9Q+y
DQthcPfaLHaqNscJ33wcfjVn3exv53Y8+nDtmbgvJjQjFcexsSzUgrDLxyq9wzHR
mGsQ/bDxaM7rYv6PKg94q9lrkTvgmTXRZ9RRlkURU7+OlUhIK+JegC/erU0ZWDie
f9HGAq653QUHMXp93++LGi7xQqXBCUoi3P+HgnpX5g/gEBbCWLRjei94vEb+bJLP
Hy4Az/9+euRDr35UJagK/VrVHU36UUqbJ5orF+zF/nLWRmhfK7ki+T7CbGygmyAn
PvV5Oc7F/KK6rTOvbHYHX3MA4awdMmSfcLpj3rH7BXaSY64A1ywBPPnSGhV700Z9
VpLUlSnYVYp2ynG/DjdP4r00cABi8otzY2DBDs6Y5CCJQHHnu+IY4aaH7ZHHKVPc
NH9tUTkaG2wgdGw3DGPECBR7gUG4pr0lsMLr7296gZEGMbr2iPxdFl9XtLTslfEo
V+tmKRqkVDwhmjQ+McNsBUlWPq+6wb1OsczinREhOoeAy/wwYbF4X41CgO6UhUFh
Fgw110gzFKbNloXTmB4/IDIjR0VSR0YfVxQHZoL3zOntt1CUJ7lOQu6QNW5PJcVH
E7IfdmXwIK9yBeFfNAJZicDANre9lf9hirZEJV1ey6DmeKb8wZCm8pdn6Blbw2eB
k2uaIqWeb2SJwKQryxG3pHGU0hJoalyzHpnrPwDs8uDmfD06bbLvvliBxo4QdtAZ
JKSxJ4t3vxGnB95HccC5TopJh5psGVJTL9jrP61ke6OShVWqTvGM1RaFzgil/tR+
QrWOJCorHRRhXRL4vEkDPxmQQRB4nLh/k7yWP2fAMYtShPA0NQ3PTGdTlPgKKouF
iadVfCQdgah6/uVf99C4s2hc+KNkF1YAuxurhNpIBDPQpPiV4O33tcYeXTrQV7+s
MZuh1eR/IOGoqtl0GMKI1ivTVGYypo91bV+Ve6KSoTu3ZpSwHIAU8bRRw5XPBmJ0
wUD8tWD1AyIZx2yQyqgehVLBQ3Y4LExfvlW8jTN9p+BJN/3VXr2WsAXdWH5iLaGp
WTP+N56zQgEDB2lwWphXIovmdIMtJvs1ucgPx5u7S9lRWk2paTRgjvujMCaNB5nI
PuhyRf+UxyMwzzMvhCkpQUY0ctDAUHL5SBhvab7jAgdo6OE/xq0HqjdUtyEvpNYA
L6Xy65Qo1QCKUc/l36Zq9ap3DVSOdnPnFV3rxIG0WU3plbemznLBIK71ZXSFFHDC
OMDOHZBoOtAqbOEFcc6CHh8N+bFhz0bJhF+9UGlCj/o5PQkgy73diaWO5UuONDHf
X6uXPICHCRlUApZ2vr7Ws2/jdKdcWkShqlNG2QE6j9PXBFxcvNYrjdz5DQ0LT+Jl
covBBBFVzupwxhOmWwpXYkCxJxPTYLQ5S0hAzxj6IE1wh7xwjMe++aioSb4hb8CZ
UC1o8yA3Bdx5IYzevutN5Z2q4oF2s38J0QcKzcVEoZOqJEgPaEpcfHmv2jQZ4IpP
sUrR4T9XAFy4Z/safv+R6c7TBlkpm1caGwXapZLp9csYpKUcHaODblJiHW76f+s/
m3vwtY+Niab4RFbYX+VVGEreblnO1VGlRyKCZpIsBcyI5YTJGEnQr3lHWQKT6ZXo
5/mfKpGtoQYk6/Wh8ogOG+KfIY9NnwmazHgMhxcUp8Y+RI7i98pcqG7bEV/yVnCh
Ba4YQKdl8bLYi8HQ8d+AzQUGV8Nf9AMVOO+REpc6dIwg0HCWz1E9HG8Wr/l0naGH
CmZUbGN0Ddm/OW11CaOp8GKURaG4eP96tixQ24Et+4x2msGXjVjZarA+ihipTu0B
tqnx9wB3jKqo0w9Gz/5LQYeBFoyK+xa1UP0dFmrxl9SP7Ut2RTID8Nr1HTYh8E0W
La7ug/1Tm5wgaDPnlOyzhcmKkVNH3CrqIG0mD9cg+gE/qh2ykbbFALGEsnkpZmte
HRPECfI9oNqkAd5OLelehbf5PAn3FIxX/SkIumo4nV/ixo6Nx0AZOz9IQkLhF0bF
yprDKVuRaUgVUT0yU5uSBcOrUnmn57tSpzGoWvK37nIRR6EZzuXCpSv/giHniKWl
457rjQMNgNQcjnS0vJf/x22a6eMonoS77LgbrrQ5lxZly2xi9CmqCqklu0ktl9y8
jqyJlMG3NzbeBlgsEX1TJC6oxi7BovaLoG4/bTrlffe37gm29r5Qo2BUFgvu4sC6
K3m1+zKcldqPvtWoM6OR4Yhhd+SZGpBGtZ1/HCb+c8+cSHIIOOVZDhz4g72sk1Bu
wiqRlr+pa7k18nnfyqwuneuI7SIodeUIG8Dz7eD4h3DmtIlGDpMKDq/rY16uy3CM
fnkInp5EKrBuLp3gQi3tYW+49xXwYfDsmv+6cBdJdlT8lcCk2EISR74cOPDCHCWA
Dp+bl2PYpn5W3/cx31m82WGj8NjXzUkqMq1kGoHNH5MuGUrED/+NP6Mp/2/4KxMn
WgCAdAP+qdsnoa3SDvd+WgJTXQ3ZecoTIgBfBuN1JrZkI1QeveDO4bKL/HWuCW/Y
w1NPn3m6DGxEpB8tUrmQhDG0Jw2XHTlzejMoILUhzCY8Xx+DmutzisPLF+Ell9E2
w7cZCOJFu/Fpk2wJnMGgLP+GfmuF+FqFNoKIbVN0QbpFa/Pq0W7ns/hGMvTQv7mK
6TGEkJ3RR6Fgj5ZEoDxocXdwzoEoh3g88DFu04S3cQIWWtkUMyv/IvoSceHLENix
oFeRzrB5qz0wZUnD1tLgNq6zH2c5GbL1Easc4RYaq7h+rv15jvdXEZkqUcozCra+
/GyjvfiqdnPwFmrR8iRscKSqbS7RzBkuy5JEteR66hw74AkCI+fF+UfE/PnpG7nJ
AzU9iD07CmwLNyEXn3mXAgHkD3pAGrfjKKn6uVyIISQgJl4zOZZXR3GTL9QwF/n9
+8ZDoAR4EXfRik2pyjEGDHYSxpQzIc/DsnETRL7JR2Qd4nJE3OEF6PC35z9UQ+jv
1TF/qUewVQ25vlshmFTAM93XGTB2Xzc5CMd54lz2lJzhZCvlkx1cLEywBF9KvvJf
bI7y2/zR8LCPCTw1tllbph04Vcm+2e97yg8Gdv+NVBWXlseQ7uTudeEvERSvzv5K
VchEWkPs/GP1XeDUDNDed04YgZBbE29N3rAVSlaHX28p1ojqbtwt4vV+L+sBLWq0
3sKLA3Au7+9Bvye18WejXVJ4WuBywkIZWNM8Je9XAknRuRVrZROtJQ/rP8OW3ei1
nqQDLzDtZlxzNV8q0KClFSzYBcpSq6VXVTf4M9zZzm6AEDlX1/iSE8sOiQQ5jXDe
khIQQgznUHhjnBK9b9oEF+a0qMKu5usFWnSITkwbLx2bdwe5kf2Je9g0cFJ3peMl
DZ4NqrH9FuYta4KsYtvMbSURSAqKtO4S2gkMOEk+W3TwJCtcOmwM+gnPFEvOVw8f
ONh1YtzUwMfMNWA0QSKbB+r9hwIPHOdawzJQLEDCnJcbv8FKZwNv28syxQa1ad3i
v/puSYIeHsU32CmlsRuulZP1IzHRq4GE0e0q2C1OWQIT4V9MYLNxQ21rET8BgZUi
7uQD/IOiQDTd8BFbaIOD4da4nEZMmh2IjcnppHLILQFo6E3vCJQbHodO0MoQ9Crp
H6Q5UvR4XI1y7/NhwN2qhIq5PmWoI5ChsssOPC6IMJ2u7hS3Vn+SCajLvFsG3DMW
RWvLVRTc9RhGrkChN047EYm6fG5bku9UAdft8/z47LLEVa8L8N11HpUGrXn+UV5o
pg2XLKxxC98MnmYuiXADYBuoR2qEXhXLnJ6YxU5zKJyD5AcLxP+60krxQLmQqHew
xHyviXh11Yznm3b5TUE9FI59xY0vvQoSU4UXQsKw7Ft50ED2IylvnW5OGR9gnOIN
KRXqiW9ylvOfnhdjluhS4naOL6nX2ECf6FD2jOMmxf2pKRGlxAiLQmfmZkzKuFb3
WHHWI2dZBCZLYMnDwysjYq5PIdCifh2HrVr6ex/qN6BW35cNubF4nbE83tTgDfDy
+f3sF13GyxdrbPwBInlIEyPzftRXrKO/y7Q75fixWdUGit4yt/D2He9nOcnzLxWR
+ZL28IWZAsVtf8rOj7BCpsdaLpgYG69KCQwqEXn6GaaFxpWxfNOfu4cf/cLtupwt
ilCdeRHEXgdVQAXfIHsU55QTQQHYSfcvrXk7TD3156hO+rPgL2mDdNa99Pz4YXel
tjZoW53EK3w/NGgeN9G9LdtVXppeGoE5Iu+vFH1Ba93ORrVcuEC+UIMW2IRg5YXD
fEnyXMUbi+9OI0pE+H0FKCdh9Ciaz006E98dhco1XnmVyNPTE1kN98gvua7cmrmJ
Nfd8oQXLoBf5YPj+QRA4EfXcms82pOnHSFafrKC0UUK+ZbMxzgKWF82DEh/F3aoP
6t2HYl06RoeDoHEaEUXmNV4+coeMy40F/+NqjvZsO6mmt0cd76iWTevF5XWC4xhK
YzHGSUGViobAg7VmCFPAYkNqAC2t/o1U7CdvIu/nfLjbreS1NqJR1Kyj7wLWkbRR
1HEhMGJ3qV4fMjRMR6A5YsIl00jZ/0F1llqlVtwWzcoIF5bjFedpOh0nXJwbFdH9
BkQpSWFTVIyMvUzOYwMy4gmRyq9kwlK9wvdBVj7m5SvwUeD2/H6YW+Ra8Md4K4cJ
7rte3Of4FZOiIqONYtrRz9JcLM2KXYDeQ6xXrOMjaEwLPAePTasVHqtK2ZqTpmjn
NjnjewO9lqMf9u0YGZRV8KU7CEQt/CYovWCMr+vh9rdf3kxmn2s1LeM7IBSghGg2
BRrdAlfJy1USZvTMgQ7Z+a7Dh4RLkbE6lrP/btA5XWstmqDePwJCZkdkrXjPnF6d
SHSPTwSokGfP89nlOD11NxarVPLUkj5TEC6kTSGX5bvGOaiDnE8rzIeR03J30xGg
xuePlfnMROeCDqMmxE4NyMiKV+C0tTGDAe9N6iG4JSOsgP2601DtTQGTkvtKcdi4
9zRgwwOUVXhSRE7bDTFdXhuPW4vDYXYH9f0Q+D/GJ/294vqjshiwXQxaa/IKBgD6
5MRSKzyJsvZPLM55rQ3jLcXvFD+qofwpf+K4jgse6nbaQ4Sxry/hurJffsI+Xn87
JGqFV0P4LeWZgnr1OwoejYxCXWcnxvT8aS/VRpaf+9YlOOq61mq/YVhsHy9gifKR
9C4i/pJyeGekawKaVk+rWQ2jPPrM83UMRV4DtEhhWd6Ma4W6hmuXSDt7OSUIKFE/
YUiv/KzRYG6kJZDXOiYO8SFah2/HSj7b7mTKcAepIoVAcMfhGU3tToTbSh+sSseE
8C17q0BPra1w4o5PFpxZ3HDAPbYB7MlL3vMPQvkIL/TGY9eeA7jDpe8IN1BVMluR
6KVUpqGahiApkoUy8YtcjRn4IMh1T6kjfbeqXxELJLedfflUbOurYVW8Vpe0GCOu
NBEu/SBubxhnFO4NJrEQxZb5HBR8wLGMFFrPtijh0UhVMSnaDD0Yyl8sV/fwp2qW
uR1vTRlxdxm4SqPHQm61uOBJDTyAUEWrCadfMDaNfcFdl61cCVbh8PM9rL1AeGn2
jYFwwhpv0jEmRSlg3JIRKwBNCrdNx2KA1gN51JhXRaF9NH3TOOMqMXCpE/s9ZL8B
pCVPV9MVkpuHJ8+eq1jhh/D8GT1HK8h9PYTaM06cmkouUk4r45+Gjwc4YTOWtQLX
wxWCeMt/bwAyF7dPyOfkp3l3w+XWFQIdWiHCNsT6uVpDruVh3S8iHVtsa8hWAZZe
6T2fLj3aKpWfmQO8Tx5jF1EvBwtP8SVbdU9dgAM2NC8Pno1N6ar4IHDMDjy5AR6x
yGm7hO4ubUjo4hdJp+zMrfcMZEucLZB1wjYDTmL7QlnxRlfFgNd4UJt+4xOADxt1
pyyHeC1buCY8VkyKA5BulpzmUUWt6axSxsjjqI9arox6aRpTfC+k0AOr3O6xn8Om
2zi4bTa2VT3BtsCdrQizGmuzra7pMa/WKKgg0ng9f1PSceMHWqQm5XC7tV+ott8r
uhIp/xIJsRgBIJLtd3zsWrHsQ9rhyV4HSjj6n8Wzn+dIi+jps8z5oUPGzyrCfiDc
Tn3DH2oWETsHrh9ZNGpsBL547TddjDprcs96Nr/9rWtSe9jeswV86NP1+F+V0Rrg
uH1sTMbbh6wBva31n/2chXB1SxFX3j5egV1jitK6cHo2YPs8zsHaAUsLLcN++vtB
7X0YbaQuoCHVl8GZ34DFldo2sWptkL3IYAdeJkk4N8pn2gYTYrqH7o7fDClNJbu1
rFJd4Cn2b1lu2m8OmCHbvAJeuBC7DqJnwzg4caGR3JBKTJyx0mQBpAiH+0ZZJwAk
IwS9RkDagf7poVypOT4ylkvGVlalAVI7/Cg15Lb2ntYtNG0W448j4StdVQZn/qNd
Fa282vOZwMZQiGOAdMP2qHLXhAQZ4SImg3pt4lFS6DrfHNBqEuVyzKtjIXH2Z6t7
vTBV09i26pbE0OHqKgY+gFejvVrNaBTPs+AV3hf97HbEACD5R8BxMl/7x74dn2VP
i7/b5hfBTyl3fnV0/w76ocygXL+PkjXJwlzJnuGh0mXZPwVRspOLFINqy9c0g8P1
lRFBUFSJ+vlcMFtRvnzqx+46ZM+GdLkYsTPkORyhD5BkSG7OOlsS+Px9CcHsktEe
USR2QL8KE2PGSGBOHq/z37Pff59r7Yf7Naw2VCFnBlNBsJGSf4b9GkxhRPSV7VkY
Vcnj3uP6j/3nE557irmqHO2cddOIEmrTAEuLvWTw+qyQnpjiO2ZIHZnKEoJZAILD
BMN7O+HdyDqeZ8dsBDUa2j5xpcoQd1qodLiE0K6R+pAurVBAFzBMJxDQjn90kXqb
s7UdFWPFbh1RY1LfGavT70Vwc2JYLjXO7Pl+jdQwtpD7B20S5N8pkfp++6Ss+i3+
8GAerblPaq0Ex1nl9XwdvR+vA5yHmGrPIpPIfdhIfYlNo+tw4oRvL/GtecmMKXMK
Nu5/gbarA9fmUpahljzDFqXis0FARz+jO+wAhn3LK2A/v/wrYCp3Nsaph6SYjVUa
BDXodT6AwHJ+6hdMn412cVrijBROzV1VJq4v/Zqg9Q8ClHjeUsplQnBbdr1vjBxM
J3dDxqifZXII0a6afAxjKiOmLs58qpaIsAu5mHHC4xGmpSpBWTVJXzudY0NO3EzK
1Up46vZ5NQTmDeyqrBH/VOTB07dmcVKKUq9MgDg7duDytkkcs2TTZ1EE/dqMmjwM
j8cFWSEYqSjlHY++avNLA1L286062eD/A49PeMBJvvY0bXtxCMMhx/T0dGCugl1O
ensd/v9wCIFywAhz8xlmwo/ECOKWs8YMmON+fH9U47GzydeYt2/BkJkpDZfQ1miA
UUMKA4ZQfxDGRH/ik7YoPL6w/eoppVKEEgkd1q0TuIHWBfq2xiqmogJfLtcZ2HyL
`pragma protect end_protected
