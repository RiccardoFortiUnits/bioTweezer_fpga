`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Mbw1TnOrFb8y0FpqzmVW/THu21wN6ugLOtWVSLg+qQfSFlOTRMdf6f6ufKWyzgXr
jstPU4yPsWmsVWKCOPvdWOPaotyRhyZPmzvCERWXQzYmSQVMlgJzymT89hd4FWs7
E463jMFzee3tWZdn6ooX1cQJ+piDaa0vhRiBXeY2Gmo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
5yviqkDheaTiw2K8NKnMDLtj6j5yyqbTEOcUBWyHGmbaM48TltcCudAnyVE/k6jr
ZTjTwFMH0TimwqxvvUA6ACNxS+iciMGHLSUzi0LMtdDH5CYeiTzPFO0+/Om0Nqzx
WffZ4G9+KysZo3c/ZA3LWExWfLfvFxLZ5mmJ2ckJ8feQNtS4fA0MFr4mfMMFSHxq
uAjicd0ns+6afnU8nrAubcWF4qt+hu8Oe7hfzZEToEbjgMWTwdN3sK2p6lsVPNnT
9+QKW/+ts4BIFSunuHW7fbgEAe9te6tLgSlJo33EJLEnZhF91sqV5q3FLvR49Pgf
SGa0OQw49dn//nU45TMsjIk5Qmr8WHoKg/Qw9iM2ez9I3wXZu7UMI8Pbdee3VsDv
aW3E5tdR3EiZHg4vYNg5vQKaWW2E0U7s84NQvLk4Bh3/IhoOz1PGPNRjBwVShKw+
EU1KEuMr/YdBDGJ0IXyryX/V9b5HaYxxvz30x8rLeHURs9leIgDIb6zfgrEoqq8N
DsxoqnwbmRLd9P5VhxqbtHOC+vE+UYGGXCxfS+g2U+d6Xtt8hfuu6/BCbGFcRJR7
OWcH+Pb9x4yG8j/+IWGuqr2PkovUdfBqquEVRUq76optSK4iZgrxjc3TxpPn7nOw
gMwpiXeBUGH1FJb7qTeC928KA4fcneCsHO+XXUm9CQuPiEc2m7EepPlFWd2MDsuf
lzsAXO6DUQgj6RFwIEO3LTXVVWAGn1LEPt9kUEjIO5iud4rrgvTyE9NaDcCCZstd
Y1JR5VHPT9tB8HMvMZzWA8av1XdtZQYHJrNdqcobXLP+GCVKn9NB3YCO4por/5jy
fOsThglyTSaIlGHLgBmNzGJKgujmnivjeUyNty0DLYYuPgPyuRbbec7XmNq0KS4+
sfPXDrP8XJT5h+0wCmTvJnGa1MLXTfujvAyysM+u+JySXLVg+7kzpP4UWHrBTUqK
gT7LqxiWiOJEF0ywTKEul1qC+uytb3IbpbJLPmE76ZoWUVufM/rww71b1NBAauW0
Akn4F5NOo46f3k1eAJoQJRCn8SdJFuyW8QEZfl4aZPPW+nTYdjVUOfr1ySXZYdvb
QM+CuGYUgxRisE+0DvF5p2N3dD9X1Xr2TOz2HoI2XUPkpzkrh87ndX0yBUh00PRG
BajGmIC7H6b7egpTzJJW0U/bYmSYedv6mg9RBTmADMx81xGHdPQXTHv4yD2wubSa
G+lOSAsJxaL/4GFJqy+lepA9WnQM0DpUZ3LLpYAqSK/HJwS5PWJ4W7xWzrJg4CU1
/dDxp+WO5bPY7BMsDYreL7P/1LS9px7zYPtgHZGiPElPH3E9bKj818EWPTswNtmz
aZI/iSKJR5oudK4v4V+aTF2tTe9m04TAO1/o3pOKB0CNI8cu5Ua6iCXd/hkqhmo+
YBvT4uJXSHzV4P/DH15kcBj30Etp4MTHNvLDlIuLDhqeyUMvMTgoQ2Mq2Ba9scMj
Xav1VQpn4jPPzPdShnkDgcOpXyWx2VXmYbFiw0B8nczVolAQZvrLYyNFNQ7kjXFy
C8Pz0apUL1Vl7KMvfATt2uWgGM+fEKbjxWc2TyirxJwSStjd0GZh6yC8J7MZJMcI
yHB5tHMilk/QmLKObvpNW0zbxsZFuRHA5X+8hBkgBdcZkUUjQEC6jEfQWuQyDy8d
IWJvaD5DA0Z1kEGl1lVjQ8+VV1aJqLsQ3gMIc39+tbTVSpf0BOJ16oNiywdr9w4O
Q67QKt6SlI5YOv7fVnLAta8H/penTaZDGkuRv4BssX3En7CjysV/m4uzBLZG8GQw
I/kttYrQNalFDYs3RDdc/AQ40SjrYXzGZfYNfaOYBRHHrAkDFJmPRbSlu+uyOlIV
xOAp0l1vQFaueY5uzgSydBqkiayixZ+sLJnXPl2Vzu2RB+TXIFGX8J9trNcjM0YE
E2r10FL6+nTLDuvoWz3xy/mWl0gb5eC07GjNE2FAEpcumDN+sl6tU+qbgVP/E7wD
3UrhdewxkNv5bfbLjI+N4qFxR6/35PcUg5Ydm9wsrYV5A0eX4jO1eImzb9dozsj2
MuS5qdEHI4lc/NJN+w7IuEqgPZNZjOWGA7omUDTm7jFtz3tPUVJyVf+BtR3pQCOT
8roeI+FPDLMLyus77CZwjbnLhhHvHsVXnyDCg3+S7Tts4+XjuJF/GztqgG1HmflA
m559pJ7t8OcdW5r/XEyX25fObAP7akheMzcJutSXplHee/L3+BgIeJVFUXSS+XZT
L1mTEoy3jfApcBp6svjNcm1t49Xxxq4QuIatFXCOclpXtPJ3N1sRG8P2WF2+tDol
L8SKW9WgUzNmV+OiyBwsiP0AJcNUXdx9vnwP1HUDP2UhATSCX3Ka/Rz9Z/UIGD26
coUkgSwit3iivnvzR4yEabPOyLymEsSTwj7lEVvNqwOySbYZQPws0w+mu/rnvc+o
AI93ijIXzlWBgy6gTpQAvrTWn30TJ664Kh14hh9Key46GL1X0l4izcxgLAWZyNQL
MCTT13O+xgiR9vKYZ2cyJKMhQJtwkZaIO4PvDeP7UMaX/bcE0lyjzRtF2b43wtil
r6RMsVeU22+Jo3cw3v1Qtsma77yNuaBCudjityrvn/0N2K2COOXUtjQWNBfe5laq
pRf6YkePvjQN6OzFYEBdwHWBZNnwJ9hGLCFzsoC27smfiAqoz8tZ9doekNO7lzWk
9ZhsQ4LXkPnpZeT1HLQlBYjFm100A4PpVKPGa4jADgp5KRnh2wRr6/IjCCC7AMtk
v0csDNdgJYVAslt6oTdZl61fm9BdqTfFN6SPLx2iC/A5SKoXp4/Z4EIt0AFVAcQd
47rk4PfIPEsZTtx6g64tFrRJu1D+huZ8aK832VXFyajHDor3dKCmklA1LjZrYlSO
5VflX1e72NtciqlnNY4Vj3Y2gQk7+Kv7a7Dtxq9tl9mLw3cP1wc0nGAa0z0J37lE
HJsRBGKDYuEUpEUiu7SLl541L8OKYtCovWaltYqW0Uv9/y2G3qQ93ar5SjaZyRCz
985pZ38cWgOkwELwQsCS7VFMYB5JQseEb2nO8IlgUbewTjpPLX5+qktre/m4VsnF
kCTfFSt1dN+ROxSJ6CCHlBH4It8v5JIXQjshVPZ5WVC+6Wpuwi89FwU+MeO7TZaO
Qi9XWWwEAS32qYNeC+eYAj6q2uP+YpFa/x4ZERG/SI71hDNszUAalyNNLy23yz0e
o5H0LxNlCaxFkGbNBUu5bzbBOmYr1Bm32J955zP10nqDHwXtlSDfVtY03NwjYGuK
aFTdRiPCAmckxaMyDM5XPYh6e0hU3qOZdnZXcombyo34ywpWflI9Jf6Y1XVByQuk
7zK+1Sv5thsNJ0EdhciOOblX/+sQHVQGDtbonbnMMIfVCiTtKSia8EzkgpSa95Nv
EAJ00Q3bY+NVI4th4oaMQYO4KL6shVM/Dggyc/TADT599ebsBEyJIeb3vxjvec66
9FJutGVCyjRMRWrogS8/xhcp2QqO9uX/rOdGLRRed9pToeG+YzbBFDn8Qr8vt4Db
c0tuTbYRcTzR8Q+goDE69VfJiC/xVRsXeLMxbqMPicc8Uff1jtMBRJgLDbHlTlkN
+UNJmWC4nwLRJXrWkHiCfzvUrtplQ26DE6zOb4H/DDmotteea+4IdVTCxsxy8s0W
NzEEbvTuRRBW9Ekcp8pE+4u7lTBPtEkas3SGAeN74SifU1i3TnkLGSWE2qFkk60w
+cfpbiB/n3Qjl6JtY7guhHUHS7vLaLiGecLsy9/RjLwhL7O+B2UHFTS1fytlr8R2
FcG9SqiNbVLPxlrQZdTcfkg5gQxfQyslxbr7Wxei2C6Unn6Ihr8JmGqjnT9T4zDM
oTgIJlInL9Rp2hqsA7aYe+Ot9FsoBFfTrKzMcV6rbdotkW8n2ZjdmpTa+46KTKaV
u5iMuFRUGKrkIXn2Ygq/8V91HZoTCgwZEz325KeU9haYYDdEN6pn2SEot0+zZU7r
OkHdMQA8KPPUO9KYTAT0+4s6Mirky1JaS8SP4Pr1NVR6Rupt6sRZDowDTfsdUE3q
fpp4xa0HldHZhUPWII/Geg==
`pragma protect end_protected
