`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z6jKinzw7Rg7zbJ9IFN3fCP8MeYJzERaEAWe7Lg8OrH/mfguDJoghvFIg4RW+jOf
r3sK23PhZ5c58MKPqJpzoxwUNAQyy8vDPHhdVQWIeAtTHzz48GZ5b9/Y2spUlbT3
csmcGqDzTaH10K81SrqJTTg4dnsBCV8Av98fPuiuBPc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28208)
gX4yGdprKEIXeGLqrTAYk0LkKaBIBmgIwaoRET3PDfI050UDFZfecmEJozh+ppb5
ZXPa3O4seSmMipprfxMnijLaiReUWjH2k0FhRyoXy3k0TcJXdSRSe9rkJXws5bRV
RRfDF9raBHj7HO7WCsardbnVJFEMJpVcoMJ97sWX6YGSeEA+KmhDCO5r4yPFxo7w
adKNuuXML0XSjNuGTkg6bFIULZ7PGHhRjG4GtXHIw6J36hS+B5C12fvrxWIQEjbG
eZKQpvQIPEY21LhIpn+uH0kbahiPr22wYbquYtODoej3QgqupRiqT1Ync/7xLN77
O5Glub24bKblNbe1MhAN6juPmPN5hZQRIYjhU7Vs1PufpXZKKmuW1Jv9IRYFI2Dh
7M5+XpOtaKTghpZeeW6kswZ4Fz7iuidF6kmTei/ENdmHaZdiQkMP2/3Tgp6V4hft
UPaeRJntpVMDpVM0hN7D2d8XzuX/w17emNkLaTaG0JtHpZc0pk1Ez6D9+c9ueZxe
pdwLzYnicEhaz86ib/lwDQ+EFALK85F/meL5NJDYQHY7llrJPhk/fa50jxZQzs2w
Lf952aZuMl6zuqPXExVDDEmOxG3qA9OnlAr1kKAsV3xu4lnYvF+yCzUjlxz4LzwQ
Bqq/bhsUA2NBPHCGc/K2Btitey/yGHkBxSJbJ01GUinRP26nooXodSKYyvIw+QCe
xHVt/FH1T1O4jiZP848ds4k9TQ1JOm+0gsH82aH6ugsXs+wFr+T8VOOdtn/fm7K1
SdcE335MPu45laILGhvmKJzG6wcLLV/DvNtfPCQosGkH0ro2frGBaekSCH8Jltd0
QY5ogElQIdWd7qEvriayU5/Svvky6D4aT5p3BZzjzSVmRnaeLiW+CF3CTeoQ4sOS
aP31+auzDrsKv29vzieTG8MPyGCB37a5bIRUSM4AvLEngeG/Rr+qyZtlOpwoi99+
BhxL+35vdcXZVLPhIO6guGhUnM1XFkErXOHdV/UCNc2BIlkXUhQhPqUJsgb81uze
kNYhhFbNktqU18FQHg2SsxreFYH5c4CqgengnTeMBlB5VkKhDL5XGoS259v9bhqE
m19aCXJUPdQHjeT6uDKJBvMYR3wqWMRnqyl0RsE8RlsCzb6KNO2IQrzcDdwV/8YT
HVrcdJv6GbdPrp2p9rejvII/eOE/hsiBASIgYGR7LaoiDWOA3lsrn/yvmJHuH4xo
bDARp2sdwQGzXNQ5c/VCmSprtgcx+V7up4SJGqA6XFTf2rPbr4OHJ3mBzBjYJkwz
ZRGcGyaJdlBv2hijiigUmBrxJfaEeEi4aPoaIq/S7Ph04dvob9/4MdSPc1xYAFlD
VwZ3gFEzx2c6H/Xi/+unfAvvVKIpwg3M88wEAi2W4dgKXpZfg4E603Jffn10hAuH
JdWdsvS5hneB8dgALaW9dqLdBTxvfLuL98lRepvfVs2sviR0dOo7AOGsafDnezNP
IrlnU0gDbtY/Q9ZpTWlCELfmHXMCY6TAQLhM48vX5oP73YYnnhWIyf0+0q7UbL4h
YnMSbh8885BWuZXWBQrXDYyPLQFVwl2bYVkEiHMnOw8nLDLotWprkRSyl/56hkov
/5GgXeDYzzyGVaF6wWf4VcrDW8+LKbqJpAxKPOvC+D3rzY/rPuqpyp+Pq3rfRJf2
A0543Fadhz0LbPv04PfW8soErz5tdRpcyXK+tkAosq6fSKLtM3tVwQixMCItkTtv
E7nTDcm8WiDRA2ZGKh1kXv/ruMQnAxLHNtStLaCb75IHEnMRqu+FeobjYpkR18Or
K1kAdUgaSa+2W4lL/YiMa7WI6w0sM4CHmZYwxWuElZ7zW84glMZhXIhHVKs2ML8k
DWXQSf67iHfDfFAEZHUwNLDX6Pj5c+AviXhEOk0PLW+TCx5S4Nv4y9yOCKpPc4de
kL1qNrVhGbeGIHIKAsHwCouUji8mvRVmU5/qLSXQq09vdrA+zxCDFeez7GSS5Dld
r2iXssKduOvolTCThx8g5pHQ+EYFrWNQnK4WVyl37nnWEHtXOjShEIFXjB4NLQjD
63fvUTS17rdy8R8c7qfJg0gI7HL4VnzN5nkjgTIjMSNTb41SJ2BJ5w/gD8DM74Bs
JEJkEuY+M1c0G3moMszphm/nNFJGPFHF8KtZonl2wsL0Jv9UWlDEux9fSNN21uic
FzyHtEyaGbxuM1xXbxpQhaa/+kUggLEXioGjzYmOkue26jNOOlxe3MztjeXmiDL3
N+FfCWNzY1NtakhgoVg3iOPMDTbQQsfl8ubVDMlbSLA6aOFXCz6Au0/Zt+eYKD2P
gzLENxATzjYDF7tcej3dhhmPJ/hVLq2rea63D66vVgW6V3WCIZmSd9dXoWF//vfa
IH+6Lyo8O0uqkxHL7LKaMjfG2ylDE2r8Hvucm5DUO6VP/ZTGzNKuqG5NEfSB9mOF
IFxdnq8ylSG4KN0Nx7MGGFdmuEys/6fUsogCn91s0WcLyELvEi5X2hqjNzfXpZR9
JwBawTHv8oi7Ex/MIgqKmojduxhU3ulX09G6T/9J/xbVSTRnsQIKwi2AvHxipfB6
caUHsPryY7DMgvfTWM0b+J+9yBV0QaSSMXYML63o+E+ejDf8/GH+cTyJo0kMBY3I
9Q/HdRcSHa9pSP25Y2W3uzd4voX2lClFdstA9F7+1OAfNasyBfBGX7KFTBbhr8XW
X6oXY58Ah3Io2BLO0b1ia3M88iKS6/5w3pgQGM3ILV4q3Io5ocLwpeVhXNM1WLlf
pOz916SqO4L8SMDe2uVI6FfFH21Z4T1U8qi0sTFktMF/cL13om+gsQcs+djD/fxN
HR8hf+K50P1M6dOcdOQ6JcG7c5GIlXAWaVQTxXy1axeQsX8wqtk55JfCpff/iSl8
ycfiMOYmuMwoKgD1JCDZOeCW9dHz+IXjEfnA8ON5q4PLOGRMWthOhm5tO4GIH00R
IBwo1wHodHhht2N5rUSr+kItZMB+Z2OHJeG/hZ0wbk+FcCM/f+6x7UoC4XfdsDU7
EGPwyRka02olYTbAE6A2PDhNqs35QSezN7B5uPf/BxYG/AllRSZwTi+58FPjLN8n
Wsy2T4cQBxjjZ4ak+8Dh5zZ01tRvSjdFSqrLawFx7MFbX+i/Km3v4ANMfA/tEBX7
Kn9HkMDpLwEuyXfc/s832u+Ce3ZYyD3Q9Jifo/acDFMut8RkYwHnE3I0kewGrm43
/FUG1meS9FpehjgGk/Sn8X9Tu+N77DfiScbZDxZh5gP3MndGsDQQ/X6Wo51N1XiM
LaQC8i80MoGhcDVIwdTh+HkfK3y4a9Ujk+Y6LRcqTzmpnWIAyQDu7tOnD4O9LX7h
Se8dSVIVXt4JyjJoDK3D5tNGx2ootKlM/19An82DctxDsQ/3mfGHyDsliiuuBd3v
BkoOBGoFtOMWIf9X7ICJhf1WcE4XYrJByUdcJ5JCAjKjlM1YlnVBBkLuoLs4qDLo
NC0v7rzoFbpM6PzTtA9HDVL9juiZ7oq4vkBNgWITvoyUhoAqfQMaz3EPH6qI4Bnd
qXsUloRMM3M4OTRuGzC75YIf9DiH2exqTyCj3ZMp9JUtZ3URmA8CVB7cQPoel+tG
+hiWxN4/v3DNaQaERUY11Uw3KqYZxdr1n9jusTKBKKBb+Xz0KYmoYz5Uy4cDuAKn
2YpMCYuj9IFxdcyW2OFoo7iFBbTERPdP8leyV8+7/Wx9ZcjL510l7kutN2FVab0c
lEILDpzPN7Nw4Wh80obZa/NEKIZp1J+DbHZQWq96WfSI2KB/VL+cLroxsfV4dHRM
RlXa2L+xW62eiPXry2hQEMfk/vsTOAYy9XRCidL3Krt1x+7YTXKl7CiNddXyhWaG
znIKEmcavf/xavMMxkbLTYfQ7zx1GvALDozh5ghiqWm1IBSnP/IzkH/Gnk9STuSA
o7GZataXdYxZpKAG2uqI9zVf48U2dnIVW7KjAFQh2SW3qCEo1bI63ZHXzFxvnQ3s
JlmwqSN0uRG7E2l/iEJ/HkVcNdKRsT/pLMMn8KaqT63eiPKkBaVY3gHp8AOqk4aA
BQaLst3l6Ky9b8AgtKBwDCPNn87NMOntkvbhKbEpaWNAP4u6gh5ftwj1uVfcu6tS
O4OdIGxsAFEeA5GLluUsr/TdKIhrXDCyOKdFHeTZN2zDqibWqN74EXl+xwnxK9Sd
s0aBhEMwQw/bQ9QrA4LTxh1AJtNmcwhaLGCBoWFazouUNY0N7uErFUtKAPmVRrQN
Dvrk5/DWVexSfV2WDkNE4OBLKb+lPGhtdl4li9kiGdHLWDRNVm3D7mQm37zo6iIp
n6wEOQyq7kNnJ44JG3o1B/W+Ebb1A617kvsSJFL2KD27Wigb6rvONdeUflFtQmxd
80MM/MpZzq/bvFd6234z7V2GTRMLd6Tm5SpBL5gqc1bpc4kJPQTSngmPtflUd8oB
nX7HGn9nNdKG1AwmPaEwNiHwrWeUWHWSGcS0wywZ/8+5T0TUTUA77wq+EHy7qQi5
Yl4hg2wuP9DwTxGHYXRohVkAYlXaoZi0QKfezEtrHMeadfgpwCFa7IXrZsYruFd8
PFJ/nPLwjNFDQS6Sbo/qe+DglRk3hGGbb3Y8T9PKqZPzdi8gC5GDZYbYVKBl+BGk
O3EaRLR0R9JNki/ROeOK+ezxq9FUoACB5asuX+zWfsqZ+r+uQ2gs2eEHVMNhrg8I
1tdZX5HQNghis8+ZbrdIVTG2stjgnfRCFdVgDA/LCAeFRcw7XiTXZzb8POe5f2GT
uBBWB7XS32fmd4l/pi5CCJI7fz9KQDjliaGS+5T6CwHcdvM7/9xJex8OBKfpvIQP
T9dtFYFceqKLDcj/lxAdkTjUtNKKhiHXITdbfOWgmEAhKB7O2TaASi596/dIgqSc
nSiT02+hoPIzafWWCiSKdi1uDUDZAf5RgS0r9qSBWh9bXgUDCbBgdWsX0syBIJvD
LLmnZRnQG7f3XP6zfpboAfIoQxeAJdP4nyAI2Sk39Pue4xd6ceaBgB2tNuZj2rJQ
fiqDy/gokXJmI+KjcO7Ga3vX8udd7pwPF8JfEBhspDC9fokf24Z4xNzYbnIbgHwh
x39Domw7KIRWPb0Kn/WBTP66CW+yu7k3wjv1QA0ecYx2OfNvz6SxDb7Gpjj5i1cs
2tLh833P6euS/qMaWzddNT8GojH4FEPXxs/RLXE/ovB5Yft31exQnCRgBb1C1HiO
G1ELav1xpFklRHdu9I4vbcaolHtzsn+9kAGuuXJWjbHMPcuxgisIBYLDI8Zh5xgr
2NzmK9UwX6//chcLA92RiinFe3fl8IG7KXGkzH/qA3PSCMbTS5aBxK/bFNW7R0MU
R2QLeOwLRi+D8wY80FefEdi6K4ivsGsJuJsMlK0bAc6nbYDoljbPvIFY6mdJA5+j
fGL5HmlWJOCFN6FKDbQ0fFLKGFhnKAQfw/oAd7Xe0j+BTTXTGz8p2l3KRzczZLSu
58RQdhP+4PH8fGz1QUTB7rEKSwomPtuSidASqVBunnNn+cCOvoHewrl49IKOedzn
7YTwGMamVqJfjhNYLA1K8kuzqqk3rFbaF/HQ+ro8LrbPtjeSzWOlWk+w8WOcivfJ
1pIe0CPWe/gKizYy5rQdSvlNW6DMYtGdWWN/JvF7UQD6TPsX4y4bKUgMkcQi3xYn
lsywNVBe0+mTP8Zt+EYfDZmwj0oRQUlxa+5UUe57z5KDbi8U8nRttHLZz+cyAFcz
Iv77j7NavEEjF9vowrmWl4GTRKWp8FLSU0PUfDNz7UAWOCUzWaCsxhYZOc/SFdC8
l4jUyFAmpNvibHjOYo78BU9MR4GDeYYrex0mXGatgwaZY+Vckl+lhtpGjd8gdHxI
KBNoLAzM8P/o6LKMw7COdbHIijY1Vo7rJjPLkOqC135FkhmYpLOcXMn2JFdcWBu9
iXRaLyZyQrPpWtkh55aLkh1VAiZx6078ZBJYjbmBSl5IUOXYkUzaDGUeW3yMhN/k
daQOAAYu6P6ZO6fyu+x1Qxu7DNTKSvBBNvJTlDMnZ/qcjLLKfV6QQb7Zztr4GVdg
YVPQaIy3JAu1ZF07Wwz7mr3dQ2QgbkWpNB0ptIju1sUHSkSsSBbZ2r2YCVEbHoYL
qla5zXvWusHUsmR2BwwADBcXTxVjlAWAYdoaw9VevT1Xlex2fKeuCj5VXwnxamFr
uKYpKtGDQu/PJMjtFJtW+maj9yIP9tulQIn/UE4br3kFu7NcVfrf39bxloI0NOxb
mlMrxSf2a0xS8Ail3C+scfaCpLp8s13LNpjpicv16WODK8Y+egc7RFy1gl8yCviD
YmqoHn+7SRPJmgtvzcRQQBDtoiqnozBYj1NpYZXCwH33grMmA8IEH0CHWdzhw9MH
7yUTDxLpvoyzSoXY+97ZCjQMhvG7bum9f8nH7w+Jj4GwyryskbNm+RS+OZghnXuz
6LSsnbBupuquutFMh08tQZvKxq0Ks6nyu60crVw/d+FD88y90ZEwC+eo3bX1Lb6C
tns/XkwvBsmt7lCvM55H0IWymWqieAd4HHiR+fhuiZgTTfcjrduy5uLtUx/D/ARd
GRoefKfVs3YBif5wXgQn+2BOHzeOMiFKUbXj2oLjWn0rZsJr8BtPwWMfTpu+yrSS
6cjKoRTkVxig3P1Eg0cMHbd5QEzqDJpGVxvWVwNXg+/n3K/XgzUxDkYJxvPf8pkh
QzCwqpiwD5LF1QiKmwlcxEOalMie/np1hKmw99Xssf4TAkmwh6ByNbamGXKuU03V
NhT5Db1TZvLKCgJVfaCPMGjePJAPlWivjgUf4jsW97DdmD8WMJMHhF/x35PFM5Ft
fnwsSofSFnRLb9nzLqnFqSJeZBSTNvCfa4VIyaR2y+PRs9u8M5ux7sAt9WIB6olb
aZ/flds6ltE1nqPPbZ5oNiBsiiQxnsApQNgwjL3sY+PZ37Vd8OHYF9DrLFZc/o78
KaykHDkUmIgzWRMNcJ7eitH/taJubettk9a5YlItuSKqhQMSRyJ0D0aOK0NGnRDV
r4xnmeKcaf3A6uodq5vj1bnuFIcS1HygdzMS0lGtsroEWkwGZJUukUXXgPQo2CaQ
P60CUS4iqEeIVKNfrvK7lltW3xWqLaYT17DFktlw6KebWZKTcJVnIg9OVW9hAE3b
U8ph/3rH6QE8AqgobqQ0WMRNwF41WEsLt0p+5m2Mijn6jWeYsnk9yITbiK64QAIJ
LijnLqfGYeyGak5PkiFCZPbb4aDGBSDIFsWMAFwEADCrqW1edIG0n7rzAlE80MVX
I0JtipmoMzq0f+mWbzCvZdJDEAlrSPQLOMCqAuabBNRUxDFvdEi7HzYjDXiH4TBP
R2Q1c2aJgH+U/zXXjYxYIGVRgj+N4P2+1cA5blgtZh3BJ1SD5Drnf6i3DeRs9upW
1v8F6p1ZH+BJnyybSRKp1J7uTk7WQ6H+wgfA5BBH2t+SSXaZdtknrUyq2n9TtJYr
rC43Ea7gGxC0lNyuL+6UK+L9qKW1ToO2I/gua2F8otlTp7sMbyEFk2z4L2ehOqPE
fIjXpMXmQ0owmmkXs56rgYoJBtWChWrLVU7TmSciyiDRCcb+X4Ov0zmyu+H4wvXC
KTod2RO1fklEXRbI+aCj1B28wGsZh5Npejbkc0lYZ8Jiur6KJSlAAbB2907F8ATO
tNVf0wiPg9wNBmAE4f3H8TN51catRH5LWnCPq8BkKo8ovueAK29AN6K9ggqUOWa0
RZQf0keqlKG6nB0fDCeliE/SZMtj6F0H3NoIjsFhIkukVXPZgj/fEPHB7bxPHrZW
u9zKQLvKnkQP9W+/yNNO2r5Lz1j0Wpj9VLtjW8JH4rio6gM633GZ9f70A6/14KIc
BpsPHSmPf+/DWB2R6t5ldymDrEzW7P6rZmLWagnitqve1rTpH1Ek1z6AN/YgbdhB
0omhwJg7jF0tT0nuRsaWn65eLL8HCvZ5Xz21Yh5GGVMBByH1cLZg4Op8VNuVXnXM
0yy7esU6UO/EnwZXivLCSpspWA415bzkvMti8OVoGsQQ+tOdEmFSsg+2wZrdGihb
hQb3jpzuqiApekALcfUj1U/WT8H3bWi5NzgIOVPqT9J9traJDyImp+BWieBLV5+Q
PrOfTMzMYYnshPNGl3eQQGdfGC8TOyviqOZhbGmavo1RuPVJskU8UhCDw/BeOmvk
Nm6+Lcss8v/KKoXv8cSyWVCA0yhVE/c4wEsRsklEy8BwgNdcPkvS0lfXJ3rckKE/
LFyR5PMbUmqN/wP2jgCGr0d+NC5jFBGGja5cfWodvnd7RTguevQ5QT4mhncVixE0
V6XuSQY1X9+mi4FNEwe+rpFsu67aG66RP3IQeBebv7O9jDhYymDrzr7KcBAG8b5F
vmWEzGg8eFZFfYlgS3HsXzARU6WuEcejs53uK0Wg/0SZ7rD8My2e14hZYtY37fzm
70afymDTQbkuMkPK9nUYIz18UwWNgiCEpqaqWXfoKqHDbNCKpFicEH0bf6gVGzI8
BW+RL86DkUMkkRSgb7eMEjuenKFhWWJI16rEnzdnnZ0TBYSxvxbTwseKw334MrKs
QwCW7hf6ZzM+djNxAS2MlK6eu01A8JHwScF7f99hkpU996+GRi10cRTVBXvEJB0L
bMwQkc+MI7McqXa67cNYsM5opHxG+AcGg43F6oYA4V3/m8z7tSIgZCuBY0JTQGxy
wUbHEDCfDGFbtJ2zha2xI3LfMCLrUAP9p09Vs+J/QgsVAdTf53r1z4ZSGobaZAsJ
AFqothEggwVDQivyY3poys4+xBEHe26QpMf3sSmduAc4A1pI3Q04i9JDMDUqoEQY
JisqhbVMu+9Q3XJ80bObgnTK44qXioRhCrGd3y9QtYAy0yGFQvZjZMWOi2OllAlB
VYAf04NSoCFt50mP6dfl5Tl+/6x11Wwnz7eXBh5IGA79h4Co1eYbcg+JkcwAl6Lv
GDcawsAKlr7oGq5UkpFXBpEG6PN7h4M8uX1aB1nB0wwlIMcx1CSm7lX9Wf+tPICi
VbCKYDZOfzHCpoDC+hBtvvZuOoVYKO9vBpysJS7y4Y89rXF1G7qw524OKJ39WRIn
I4XpHvsNwdGhhtZIJOY0knBmv0c8fJEF7ro16HC1drst8tVDBH14uD0V02IPxZn/
CJbzs3Jf9KkX48NxOAUkoZui2plNw3thW4L9KGWbT+i20sEsA5oyQaYKARaLCH8M
UTvrYoYej3/7Y2TrARD/RkR1pz/35COhcR1goRwbj6PY0997Ykn4Xt/Z9+5GkIiq
igzfm7MgNMW1MUL7+Jb71RH5wByyzoJQMsi/bit+uRqwKlLBSTKWjk15FhrgiTCF
JZsfbS5pwGlyJNr7SheeetjS+pDTOWVy56gc7K8vYaCaZSgOJBr/4fvDe7nJbiO4
aaTCVh5jiwLnebNj2qgcVQn53wWpmuYWcCr0ntJ1jbtwu/LjN0SfyV2GQVwcOF5r
rCHooTyF9J7Ta40aMWe4hqWxJEJeuYs06l8kgbgSgNogdIRFmzMM7WWVBcWSidAb
zzl50KASjOnct8S7K6y+kK+CdIg17MsPBxfe8nf2aij3SVrp0LDxlakRXxdR9x3y
jVxX2xPHuXdeQLq6aGziEMPRP1v4FDZ6GIF4aj4VtflXz3+OjEm3PxrM1ORhEv08
gpfu4o0FAqaDtGfzpDZYTBrHJ4008g0XMsLl99LcLbpHyZWbyZzshXEPDHwRSYBs
0XcOHtyFBxQodFU3bymYULx7YSpT2BDufN9bF23TduD6VhXsSaYOk2y40sqpnY02
WeZxJymz4IkdJXmeAypoV9hXMnDWU0eugXimfF0Q+t4HXafvXlJmSmKrgxfI0/dh
+KVxF/Kf+1q2XVU+Clg+YPzfGdFihQ0agEI5d8x8ExvG3+Ifm1QwY6OruhkrZBrZ
4cSP1w31DNwKZuNjVsauYvMjISKX9yE49edr4aa5ATDZlzYLO8vFxrZO72Lz3mTy
c7huSC4mcDFUxZT9wf37EkF9TSRPCvy0CvgCt1sFKsBt4jCm0KLlzO8U/fo0E+15
UYsJKKbJQBTe2yCK176dgLS22BXOxhC4EdQSXK2rlW6euAQKc8GX/nRgxqgc2mhT
MwbBs/+8SbV7T0K95IB7TzWoMFIdPoCQz1OJRLDQZs7/qPeRFk9Ryr5/3sorjuWs
Xy5+6zyL36HVuQNz7npRrcMj5pLHzZCJ1JL8h9Hftlv4bTrO+maRjz4Me5WdtUG1
dRwiip3/94i/lWhW3d3GnNwsgMW8YxqfwrLYZNi8OpZuZp+HzwNmY9wlzcAM5iuQ
O3HhFiJdLgsIAC2M0SykhH+BaAmTL6XY3+IYN96hFm32nkpqHbJI2yB3IX8WXnEE
vpmBTieBfWYDKRqusdvDtOjKlot7bdSrb+gJGeX0zIF6Vv1mOnrQPo9P13IAOvz2
ebXIIsTjDyROq60fyYao2WzeYx902jNcSOOfD81rEn2rYyJ8Inc4xZzCNUlZ+btN
iGSjd0FavsBKt9vDdnbGd5gj+iRc/ywqU+G97kaLTf6nzj/WnnUUtPUReSJ7wG1g
VHKoieQn3ciC0cj5xeB/J4pB+7QqL8egSWLwgPoJs88C4yCc5hU10axJcm2obioG
1w5b8sC4iiJJozZ0mjEDF5nbH5r9g+oZLsBCOTBWfuMUOOwDF1qhC6CNR8AkW2Gv
8intzgR+aIr8HE8uT0g7LXcutFjUYoB3AA335D2Rf8PN91csm2laJ6yjmh16gqsU
9WRbVk2fN1UIzCYJG5Xh6p2+Pu2OANrGMj91zXY7l/Ro5v8NAqsRqea47XAPfWES
RuC2l6ko3GgD3KgBJYVpa1egyV+AUTzp/AFC21jXl3/JLW4sj3FkOCa/HvjsuX1n
d08HoCPcEtxOBZBjTaEr8XrP79UQLVKlCKSDuIlxNeJgvdjqYk5beuanPLWc8HVd
meLks6GAE9kVZ9m8kPI/Kyh2kYeIbVKzN32MeCwpopib7+ML43ZNi9lIIy7v2w0r
VyUNoohalSsgoY2rzUTp8oUuH3QdaXPyz9fpnKgI9q8gqv740kog5EC+qs17jhfI
ffNAl+S/4+Qun3D/7zCSoL1mOiBNdzTEwpJhryY357Llp6Cdfylk4yzen4PsjE4v
ikKYGUqmgOcqMucqN1KRQuF/eS1ev9FlwwZzqTebOYvR3bgvUUclYUDD/6lA3apV
cXidEMfrrrO66ZPnuYiEn1ko/pqQlP7eY+Hlq673l9aRyziDRn7RXE86fAhnCIkm
v29DI9jJ1MgjPUecuKFj/vcHef++WABjOq65mnTtkK4EdPnQAEwTmaR5CXlDAzJm
RgpU9Qp2nfcqNz/lo+xpfF0WgGxvNYxXhhlvNY1n5HZFu5QyOHwdUDCdPO2YG+u1
X7dOwpa6dFLXPT8KCYzFE+k8OF8YaUI77ISUn59nQAOy9qnJc1Y/K62WSII2zdNq
Zmq3Tpz6uUkQ6wDqBrVaKqHk8wwxRuIDDfPtu2LHXvSCsOpfwPYEN7w2aW3p2T63
51zMD0AJbS/b68cVp55uMwBTMx+KDIwE0VATb94oE8orUPTFy441t4ueR6zQFev2
lh3zO2m6tQJgahY0CdBqjslBRbMhZN2nOCjhcg8JgeCWfjRSHtv1a0/EnR45cdW+
z4A9hbfS3/kFxhGI63AULmN6o6SRD7wmuoJqWrZlBnW6tJ559Be9BdEsBoVuPzdI
HR4im0dhVkNKkrL5H0KqsXJcEX4j60I3GwqI1hu5m8VYHS7DH6Aov/FxiW6cRbDX
CgzPwmhdSXvE8Qji6nHmEBF9wn/FdOghJS2k8tpg9aovfsvX28Bp5GUMEEBf38dS
tY6YBa5TWK98nmevIvSjPTsPJIw0nXt/2+VPHNgVAVuN/Zc1mE2XAOEP5aSKvTRY
U6jCl7FbON5HSKwHQqnSNctfyNlrYjPpwrUeYEWGnMx1x3A2wSQDzg2+xAXe6CNC
KmHsXfuwJ7GB22JoMksADdQ3h4TXxE5MadgHOK6SaAzmAXcFdfBj1ebxmmvXHeAl
3V8wicrlFpACkNfgs8ttXKab/RAniW5P7h7FbRqtVKkW/tjl32tym9Ot1/oJ9n8H
QqoOsYY5KgaC04KpJhuwzELk+/aD7id7QZID/Wz0IPl5ECvmG5tXT38KBYSMvJLl
k0m1MPTzVyYpo0WNMcuD4vLcaaRw7WqaA7ggVezFcQNT/PRvW3Glsr2qtM4nM11C
lFv91TtjzB4MtlNbQja3D7RKDeaOHEjJJoyjggh0yfuJBGZhLj0mhdjUuiAqolTH
EaEq+lRakOG4KiTy8/MVpdlZPlSczkryetew5Y3RQrGKPwh7djLChnf6m1BAEKCX
p8c0hhyD7e+HabIMPMI2npVcVN6BGlY7Jmn7xoUi84TPoEEBcmCgit/x6J09riP9
u/6/7zhXqejlqvcO1cWySIfooFnZETiv1RtGBVZgOgX94rFKQZ4djO3B8sqqlkP4
NnC+p+Qbfq5HfdFbmXWSgTuU5pvJhY6rFCikZyaxaV71INoteQSk2iFRMDcJatDJ
MgIvUlhN5JegL6aKmBuNmS1R47mLQLnaXAT+DR8Y7RWbrUwksmll1o5Q6GiUozZL
4+Mkf2Q+zvrH6UV3A3UNAs8SWCM42/pMDQ3V5LXZWeGFxH2aB1Y+1FjSy28hoAbx
fOmjbHC7NJCMIIkQKiL/W1Jkg+h/PcNNfRWVaqFzTlK0AzmlAWxr8V4QsXbHwBhx
wsAXLekcbx2K1/97ihlZexIBn9vhy1eaJnWmRl5k7tiiX6KTOh3sDPEaeEe4DGTI
W2xDH8PCmpyr4sO8GdlJSdmBHx2B0q5T8aWY6Gmrd+5OLyFAHcP8GRtaVsmf+llf
pq8fENx6DfpBUEV0N8LplVfKNec6+4bTYUcqtz+QvwWO9EYxTYueh8nUAySkTTak
XMwPD6quW6OYCpFw8MSLWeqsWj81TBX5JhRtq+NV5JbT+02D9SpcWIj40gKbVJml
zGn8k8VVw3xiJ5HY7vVrvJWwn0vFna6/zw4qy2jRuwpCMYh1nG3JYhyAN4L8f8t7
cA8ixgkX8geFf7JF6s3TU6UNRTKTmDfRfkyfYXhZyBf+rHLfZokQ2V5m5vmrpMEN
6VWICEBEbpzyBTeMTbs2bTNOpNUSVhpmYqBmbtnWuy6H8dQYeemN6/fLxTIv9DvW
rpLe3BJFABGJhLKYLZxzSXZ3SUOUL/O87ypN/3UksNTW8B1K1td1WqZYad90V1Zp
W1W6WmibWo5BsI5G9K5FyFNrFzR7oP+zTztGMB8q9fCu7tST5LnAqkM7KtJmQJeK
WOBmCnH/5RHlZh7iydsPPLUqQ8jJlGoP6/p9klCLSEdBW3D6grr6EBiWbqRP5SJh
NR6TKihAIbSPUrQd5yWqBk8kpHqbWdPSy6Vp4DUX8Ou5zjzyrdT+tLuyZSf2JILo
PXiQLVzfsO5euSR3okmnAHnlZYlsNqfGSjQrDyv/lAnm+bYBOeLF8uENlmQg7usn
pl4TBYi/5UlOtK7cBLq34wgTs/M0XDCCZBwAD1SbmpEzxCE+nD964SOmSepxPV+b
R/2p/+1ybY/aJ8gOgSdjiFZDdexkht4wFmy/8690iXbI/+n2hxOFpjrY4GzLDVV0
sDnXpmDNWV52aom4lFkzDmFK6PqyXnl/qPBdCz6+BftrH9V673B51Tsd6CSQTru1
BtJ4wsxxuok8QuBAfZLfwE9+5w2XCjNZEF29UVrf+JJTvMMeRrgXY2XXMA4v53NV
qSSlykMp1U2u3pn3QoPLsZONtz3jJ9HkS1K+MbTFZkqwTKWKyq7HoclOlCCs8SkA
TOiUoxw10NpcqGcxGTasxpabEobujhItedKHNfsmq1SjAyN58Hm9TWx+HzTJPizm
hQh5aQSoU7PGyERAwEosuehMPe969W02wP8M18wBgjVA/aIsaxfPLzCqfPmt4pXU
GwXKD8woE1OQzjN5DGPvobcFuRBnkSxfV2itlOMrrLqzIFxquJgQkzRSyyGKs1uq
LyvvvT9nXO711wF6AXYJ7yzTjS/PdHZVWfoO6pCQ7+czVXdt/JDfqyAuX7gC0i+v
D0fHFvcwoWNfklrP4/n/voyl4gIXvhG8BVNrAR1b0hoXWpqvis6Wwch1udJLnTvk
ex3EH9elnu9PjZt3by7Q0ZwmmC+GWLWiSuzpeKDhMGqDeMnCQO9+T4DOsHZ0uy32
IgIk8yj1juAzpV9m3VyrzFEMtPhxyLDXDDJEh0mTGyd0naK2Aps4TDwGDjqtBLzv
e1W0DGPTw9M5ANA1QwhN1u3/U3R8R7ZjBKN6PRmmVsJgAsdvjwo8BbVBbDEEMFir
Dx6kTYkg4d0eDPTgdHI+fyDzTT37rZ6yT9fWQmNo2L7DWuutBSAA5GgefjIaj/xE
v8fm4F8x4pO89bPpEqY7HReBHKMOCbNZjlS6tnXFrE7cClrmQ0FofuBiEr2Rl7Vy
d98E7av35e4pG5pdtzqsLg/ESS24XtWt9Q69Oft1S9rcrmTaPyIE4cBXb/eloa1S
qAYrELBFppKfIZhD58TXM95p/BxItQo2YQI9LUU6ywxhwGxcfyEjr1ZzrMxTcTIV
YVT9amQAe6XJYKm/O/LRy1KrVhKPPovra7vo/Ou2cL25e6kgc4giXb6pJN02cRaN
OKhZxsSJsZub7hLvzklQvNIbPjs34mQBmktoRQBnfr+2b5kVOKjc2STcrffxsOsl
puNayJ6+xD6LJqKddfqLylGOZgHz53bDzxpYYYB9y4vh4aRKdDp0iiXnttuHLjVM
UxnNG1etcbpJ6nzvsu781tEDjOEmi+qvJPW3MKUKuKMUXs4Ho41PHNiBeeAjBkwM
xO4G0b715wiruVx08rI7yD6M90kaCCaCF8C7hTf5xirOjLAyiRYmirASYl4AYF4T
Uo57aRlH5FmyesVjUthK2s3MEIREr7mLy4/xrdulrxSstm2eyc2+nJXoTQpArsyV
hV8XO0fcCZiH1kDtqsbVlyf+d5Z7XvhkC7YivUZtaF5k3TZntegTO0Zu0xCNBOhV
HlYpr8ZK4dw6508R8ETiUvSt1f2hmVPZygjnfB8DuwZoD4Gxc2lJ/v/8JIs38gi5
HD6p7zw5ehtslrTb8qWY6la0ossZLGU3+rpUKurCpYvmNM2+riWbgcBptzqMeqVc
J95b6weYNijdAsi+4YYoeUQUAZTSktSrw8B6/Yhb3QIaQYjDWlOypaNnOgtYwIpb
PDOmSfMFznRATpGqi7Bwsy5oeF01/q/ZKCB8Y03qHqjemVl1n2lPPHHrWx/u1o9D
wKBXozdVyLQfdBd7f0KGvGG+gzvBCEDZxx2kta8NA0yZykAg41l7rL1CZkaWJAUY
3FTFffeXHc/0vmolo72C4QaiYu77wAwI0ebmfImlFbno/sZNBPUs8bITXg4zHfsz
zTfiaDC0xgDm6kuyQksXUhlMlz1kGuhISws795vZ9YfbqwP6Asa6/16H9OQzxxo4
eOFAY9JEvGcwMhlbIq2uezyPvmFfKJUJPDN+3ev6Ek9Xqsy7DJYz4RXIWCnP3ZjL
UNqxVRJfBiF/e4FIwBOTpZkYQEaSrOcGpQhwm9Gr5ll77dyRvTL4oKg4g40IW+O/
PF4+YXdhyxgUf8Tr+3M+DrcMV6CpTTyGx55s+U16v76vNuwZHGmtbPQNf8GT2xJP
qKOcZGUStQ27RFouyyFKANImi78f07NRs3fPb+L+AQZ+L5k4SEUi75Ua0i51eS8j
Z7GlTG+9wBxKgzSbp80Onk/ajiTxHIZEVcgKFIm83Vo5+eD8Xc8Fh4pgnOKozNgz
rVkC8Fmn5nc4OTmVF71h4zemygexpvsIxEYY0+nVcFABhLMV42IpGoiweJfFJmLI
5O6TpHtuqiq0C5O9DxVAC2g2WzQQRSBxyR5KiiEi5rAqWNHxFfeMvXlybJ+cAnT+
wbkVBUDS6mpWM/fIsHNxmaatBKzbP1l0lM15PT5NKMV2Xqa3bLS2O1GPrVn2pMpa
hgP9CaXWybywcmy1VrmXMhq6Z5o60w5Dxd9XxDUasUAKqa7mHuwrYVpyKUMzVU+W
m6WaXgTEaMpsAjje2MLQUcwrh3Ps4zsR8rbTvPvnMTnm7dyZFBsAv18VJDA8kgJB
zuig1jx37gd+9k/eTjJcFizkMR3ds45cvKXcawXNxdumYY/LjRuDxNrRTwKnmT3s
H3t1lHL8wUwN3wPAfb1P+x8R7UaVFP7kv3eGJzotMPcSpUAzEOOMtJfUYGw20dB4
jjWxMNJoVOaCZEur0kAoe+wqHUzXrv7PyN6CawyekgepdExWe8Ck+fYmvNeH2wfU
0DywuULS4DyFcWhC+/rDlfnv18pAuUTQhkVRsrMm0Sj9RSPg8x7URfeZXEkAwS88
bSS/LAg5prTe03Nh6YRqpO6Yuz1+CsMqjo3qZLXozWSAfRGkXrbxtRc10OIoolgv
G6NGKkVk+qynuVIjgyX5JyWIkyktIDQUWu5GOmU4lIwIDXJr87+bZQuEogC7QB28
aL1RYfdN7LVsavx52Nrfam9w96++ej/zxuPoUshn1LFp09mrtj6eZbE0eAXpQ70O
fDhKf2f3JsuyE5APnn4L9hjFbDUVfN9Y/fhxc0ka+u9G8sRCpjUMTX6aT/48o9k5
gXSgzYYL3Ao9sy01RIrTw1ZasR1kf0bZIdRqkiQW3HzN5UlsL5+suqsm1KS6I1Ul
h/n+fOKCgQ8e/OZEl7VCPEP+Ks60GBcQWYXXHpUWFI8+RNR9H9QIa+NMzQaTs44X
LaIAODx8wpzvj5khxLt1NTbrnbHaITmqS1GDJUjUCt0VhAzm4atIyASTfBwKxBtR
tzGtr23V4i9Bcmp5r2TMg1QD8U+7hm2Wq98BiV/TbOq0zEyNf9O/BgWC4CxYeSF5
npZa7awdiLFP7GjyLlZO7ctuPh3sr/WEwLloCW4lDeSi3Ohpf64QiN4Pt3TkfLXL
v4BDvc3gVoKK2KqZcFJStCkfBja0RXYEkT8KoMcbyG+Pgv1yG52XA1erQcLLtMDH
pSt/P7xXPI2Fi3J0a+8SB/dCEhc9xXevaBLygdV6LPFgULA+7tiHyQNYQFY+Y0gq
jDy1dQWsh25AGSMdETHU8h5icIXAxRbF7+BA8QA6MfTq+IbhbSi5BG82zCh9kk8J
mqPoB67XspjWNRKXF9D9zwEBDgL0zzZMNcI+gNqQCyPQ3X+Nr28EyfDO9JHk9m48
y4RV0USCQyXUOwyRIFrlZPnGYG6nC2mrdVyeSRtIIbCjdKDgANCpzzPofT3uBK90
2YvP5ZBrL/OtSbcEJmpBGheF8CVz8KHhFeOsCUPxEV81F60yjI5xkzliaOUgCf/M
E4/TlsCfmTipcmvrWO/O2vxFMunWvRukB2W8kskirHsdqIB7JXIFOdmRAQR/g/tV
IjJagBXI74uEmfIYdjdBIrxdw0rwp5Rk/EMRMtDp0jC2aXKeW9zgNBGu8toy7vkp
OmfPi7+2GOzKKndnRliL8LnQKRMZ3LYTNYA8lESLQei3I+FVvg8AJqRN0C9p7sa0
P04aIbcJU9VAwZSWLdMb48zwRIM7lx/+VZ/ii3SZ1nDyxAlvCDx4n6QhahYnSaBj
g7wyER1sFaM2gNzmZq+wfpe9+btvj8KfDNvjaSSuWRQty1PfHYQSD4jzhBOz8ywU
leO2anMhbo2ugdi68SQx37gNQXDwfiX5aU5np0kLYbTotbquYKoRC1IzYwSdIOjj
jN4vjrzh7I16NBwLsU8VCSKnR3A6E79z+s3sYzT14AFfdE5OG7PlEDn/HhFzWO5K
MYFDtXbQYT5+xxYScLTRxXZ4oAj09ZrVO4qWuFINXdLphdp98N1RqDQPviQlZQo6
KRlAyPJ5vYrn54f/heDedK0IXaX8MIaD96cJ5mar5OVPKCE+cv+YKXp0XAm/TDm3
lxDSqn9ryB4c1TOrQ+mSVE89KJxJHkSEEbcZC9qQVUzuFZaARK1dNibn2amCprdz
zV9rBge3zhW6HSNVfPcTfrTCgkKELUr+XCre422XSKvG/wuqxhskNDfvAQYaHmk9
uGcd91fFmx1pPnQY2lUIdEIqPCOEAnGxZP5u1RdkYCrNEOV+tcwcIKmv8mfj6Dsp
EUqak297RzmI9WubE1EFIPfx5r2sHKuz+nGxbruUHC5na1zjf73diVHeAtvnDSop
wZmEMStSZn0aalYkhSaRbI/5yLu/948Rj/4DbLk6SIii7d3YrRs91WVbIBE1MjvF
FKxe4wlX4BcwQ+p8HdzY+PcVcAgY7QckboNb9rUiRgrxqj7maAlc5hKdjc9pTTNm
khx/h7aBSYTLfPuVshz64VZKAUM+Aayja5H7Qb7AJxwNJCGt7ACnLhNONQXoY0m+
v6VmfzqygWf1+cETTJJwcFukv+GA2luZro+gQUpPefOW96Vg/7lks8KyrH3Yav5n
v0wMjlOmi9ARkQsky0l5SGcPpO7nDYxO94Kygj2lfmrUeK0cZDT0ZWF3vflzDlEK
m8vzMT+6fY7jK5WDQxoGVS6IUYi9KPGEE2B+8dywoY4MY+XzgIOJqIKsDamJagNP
kzi1XWWoSakQ5oWjYYwDnuV1/AnsJiwuQZK75r4oRaD7Q0QtJSe3dNfrN6amBJWB
9QkZV54lxtfj/kc/N55rLQ5MBCxyjtJ5I0BMScX75nbEcnud1GcpqEzUi/AQKHYx
LMW86mkuvguvfHpq50l0s/ZBJ2O177HkeJ6hgtqiQYOaeWRhtxdext3hokaLEw8P
jWWusUaP+AtSf5v2LoRMmd/Lhb972YkaeAWT0bYDvjaGTnn0xR/rLoeqELbmYL14
yZxcbNr09cJgNxRWhZ7sNlYjpyoRbZShr23mVpTJariOFv9jSNeuVyMHWk7gZMF/
k1gU0/SUH291iSNnCP5CZd8T8tVtdT2JB3cIoyuITa4DdRdSqlZFN9Aw4uED91DJ
EhZhKSeD40dUOXfykg3VzFfQkx1Auudp7W6qBUT4I+1mi+SWQVE7o3wY8hY4Fn+4
qcravnyJuARW+CWMBrFgxi7YEH5yoL8a8K3diH75ZhntzuTeS6SVvTUEIiioifq3
pS9KMpY5QLjOA2wkUaHQd61DhR8S7oewWOS8sSgPOYmMRYE4goZ0T8ozscb81Cw8
5Y/H09zL+aEk4dr6u4c6oXFLxFJs1LVQhZlMwmVDANNOT78udxHv+We31fqq1jJE
+AloRMgVVEgD8/wi/iqVSfW+rbQnnZB/eSBciNd6cSraHyIw3WVU3q5E1i+cqPbB
60NZzkZ+CAdiiVbgtvPi8B2uPboowFzRI6rdCLUA+NKk2iarku8OI7l0Wi4E7Ypj
Rb2ONhy6uS9B7MrJBN+T7idenOoeWPEk+wlfb4dz+HQ8LhRmJ5YHgsyZNtdMO/QX
PC8oHELn2hSlisiH/mhdinkA9zlSoeo9OMrM9Os/Fb5VOkWnGMuE9Z8bpxQy2K8Y
qws4NdG5kgSvtg9Oh3/O2C3+NTJGJRAuKhjGgE6RaOw4w8jAEXZajrt1wLnlvXMR
HmAb0L6mgOnJy6x7hLyKLdILxJ2cD399lFcEsEL/pGFnFltxaPZapQ6F2pMava/y
IRLgxnF3Pvtcbpi2CYU93JD66hcHlKcw+UbTvi+XtabH8kuTWiBs389feYfLDFg9
wGOrWiHClEsuHwumlfEDR15XfY+wEfj8k+aXEdkerX18pqvp1Juy6GiwHoQ5v2z0
sZzpKGD6X6a9RYwymOBZR8bQZWkXPPXYaNCgf7zN1hwAothUkF8KQh8ra73zbEBx
/WVjpoiNDlO75GCSgQkySUEvn85SaiEcPpNQz8ONN4SQrwHBVecZ5qSKVmlE3biN
+tjLpQ5F0E5VwnhnIFHYtP5EahGr/7DpkjgEkUP2Px2xkAw0EbSCFV0vkRHFKLXo
YA7eID7K7THkk9LjJOYJux96j+SYYAj68bjp8GPkv17TMPcX4irmUNL+wRyDqx/5
My81qPa0dw6IAfivAM5TvK4zvI5DM5oMWae/iKR3sZNl5aQ82aa0AyBe1Kontp9o
8uDyO3m7Hb0KKHPDBDWn+vC10mWNZ0yYgogGyPXJwGCPVnNs7IUbE9Try+Dm57U2
SuT4t876RFoh/Ah89IkkQrboGzdsOUa9dLyuJrSY6zyuaxuTK73r1o23rmErNDw3
xdDxgoAG2/z4GxVS2NyVKuNVMP/kK9CzprvJch7bdQ6Zx6LEwSpHxo/Tgt3c7j3d
YTWC0sPJZ/58EY2twlTBhxXFEE8u8sI130IEiDuhCkYOLBEZvxFPpC15gN2Q9G0Q
K8LdVx7qeJkj9qRiNW9BHs9AGWWhLVZutZDqnqlYxgSQ+U8oxu44vtMMIqd9oxJE
ErWSgbD1Ftxwpury0XIljKizKbHPIvwtkTVWxxvyK84xStroIslosJU9APE98cdi
qLgv13msqyO5+cL195AkhOiHXmvzu/++NT+shGAKEuUShoRxek7Ls8ugOI6iVRpB
SB9BzhxtIdwoa6At751c6iJoD6ZeE/z1rvcfT7TNuB2UmRhSFWnIrIl7GfZCYQYg
N0P4v2N/Sk8SAHt8/66aSATzbJRp1LoqOjqzZbqlYpABB8VkkRSD7aXzQ0ByDFz/
0s0XZMXQW2rQffW07+3lxbHESXYmjGgIYBnwhob+WURm073p9eectgj94/WgGZKk
w5xJlwevfMtYKG1CWPJhmd9KsO7jsxCCspm/qMKn937AM3hHNThTCE0cTD5bLULK
F7p467f6R/pFLoMTGCyF2blkFe+KhrbXQ0V6jCR6gWLwYsM7qZbwcgFOwGtIn0pY
wFCBBaO/PGfC09HI3oHqpQx+4zEPD5IrsG6Di6i5N+27bu/SbSsUqMqx/NCpw5+d
Eb7hxTGnAz5gf7QEU9AtvjHRM+Wsp8XxV/HAPSdgZwN6Ci12AFCvTi/PVtQFPjJ8
fTzAY0tqaYtM/Gcfas9cM6fkhJvty4sSAVAOjLsAp1EvZjclcHSN3YGKchGI7piQ
mCKQ/ABmEkJ/HiR+plwe8erNHihfEAX9tiny0cTIu6jwLVwxybT53vtIx15mHwgA
8LR2iyxxklyoX4SMH6qbPNCuEl/9zZsDr6I3vUuo8bjjzwalSvd4oAXIDOP0skbk
v1y/9Q2MdIUDRZrV4/PloQ9I/wiDbn0AjAF/aw22N/VsmU4tjqfk3lm1HaBl004i
CampsG896JlDJaBE672KWipB/tBcE7DJWAfWZO7jOigoIoOT0UcFt/AFq/KOnclv
rfFmRL+Zo5zHQXGC2qKaj4BRHqk2Pwg/CP3bQGrat/jAUbIXhMK23ph1XB/X6nU1
PUcWt++9RGyGpHyjVaOpbKOjNvSKu7mwC8J5soH4PQzs2ktecvBEVcJUa1H9jV2T
Jz9NbhSKMZoF2uBNC4o7UERmTZTm7JSVDeZDDNwllJhsXET9gGPkFpovGkcjI9Ic
3kbUCK7GgHfh3tssuAN6sS90BstNcvpOvq3dVEl6Lw8YusEcssPxlvk4fMi9D/s2
kJrs81HTukXfredl04mO0QX4JXZ2lC4MR/PjgrIq8R0FcNE8+L7jEnblHf9D5TlO
mPGPKIIwHBNjbz7E3ZEnUQFs3UORIm9KrD0rKOh+1GsHjJI5Qz72W1k5+J9x9I68
KrAGDrsFxLth+s+vcKBXW7v0XfyfTc+Psj0XKGoLXOWeuoibo2H2SJCLZOHHjM9n
DPtVyU7sVE69AXS5uLyLc1FvWWzz44aRpwFCJXb1I9Q/8uSdEL/N7JmWyglGrzNB
qJwWG87ncSrnpLL5CKpD5pOPBDvEzy1XhWAeB+mEWfArYDch2Ya1Pv9tW8p63vXC
U6xZe0R5vE/LHdhEqCmG03Fhq/SxzIaybdPYQfDW/ZBzsdfXyAcwfkbhHBLo4oSc
bwwAkbT5btGx/N2B7/8/JtmVRkDoM8ANapX3KXtBigYVv0HZfH15431lVm+IbKk+
TA3Y0KnIzno0PAQUaw84wn1CI/jlYD70QRG4R6ylVak3TLDwnvORfrYhcCo93GRt
/NZghkUxxu5SJl54p9QhCZXYonJfWiqjUcdZhLKXqhrdqRjxl3oE8DIHfIgvbIdK
PKw5E4nZnZB6bFqQ3Ydx61/YN3ASt82jXsF0rAqVo8/3mB4m77azDtPibSbZ18Zt
AAcxKqxItornyVO6GYLBRVFlPf6l4fUy5mQfaO9g78BX0VbI3N4a5aLBlSlXPQpr
s9FDMAzDqpQdajCwxWG6uRahCVk/jC3z6lVm0fhYN58N1XPhoLnFMqgmg4WvZIKV
0EvWGnQ+vlduYHuXdY6ri1tGnblXhgon4tY01JqH8/NUvtbLF5dy/niE2H5FWAzw
jtsFGm/g6y0aU9M2Il9Xj2kgRvnXxKR4UyTHvnHE9YgKoxQ5/RsjXZS0To9Usfrp
2t3jIylr4W/XrUhXDNWua9yRbBI+wZyIOfAMrptlg5q26ClQtsG5EOL5T0knzlb7
HgyxQS34Ec0yI+JnAuY3AV8naxb3GIewhkvr/9Xds+BqQzczSPaY9+qegxboQvaN
9JllWWjCK4AgA/WHyKv69xqSnWBJlBBptM7eenqW16avfPX7KMeipqtJxl1CJwgt
dXKG0BOS3o2HbJijMYKPdt+Pyck9vLZqHgDUva+7TO4Q4hjw4z5Hj48VppGWYA0C
TF6CuJNgZ1d+Ak65wlMaIC0IsWqZQP787+y8zyEx3peLjrE5UmS5sD+7FW7CM1v6
dYMZgthpWmtfSBanN2G0r8i+z2N10d0fZZXG7KKOP52GxULk9xC1GKMLr1DxwSSs
/6+QfIgxRBGkJyASm6E7uo04h6OwViofiJ2TjoSjNMtaX3cJ22agFo04VntYGB0L
/u3wLdddtQeCOURdYceHv+oTFOHryYLIeOJ9GGL7m0E3xyFLvi7QCLqnusGK3chc
uRhZu8lqmBBmoxOLJ7aIK3gPfFZqTr1iC+ikUiijf86w3984vUFs1Ort5XgqVith
i2xXGanriuRYeu4WhnfID+J9DGshFKZ09DIWgNLzedF1ubyqWDNgEV9GXfDkWhfw
HPFFGAcDF9Ag5/is9Qq6H3DUzWeLLPzx2uTOTepRSPzByhKD+NWg9qnsnDlzyKdV
5tKdHVfu6xNm390gOXRqCuu6MsMdZsswQSd5XzP+N48eBvmg5bwfLc4GPowYleCQ
7hyVDOtsTE3HTmS2grLjQ6PMKuwoAJmJKaKRQPOdCx3GkCONYJFLkzp6EOHu2m3Q
SXmFUU3ZS3fCX/os1Qs+/2jw+il8kPOywTjk5EPCrpLYQEhs1+IC1mlqv13DX3mh
eLJwGczVPYvly4akupiaqUFsP8X5/QkYvMvC4bRMbAlbMDvhYtMQA0W+foN0b+/d
mpGE/TuxSN16AENL6beo7lEoVLziWkKnQYf2T5VDQFcvaJHKTmvaGC9Xl9U+xW65
ENX1jjLYRohDQw5rLXqFNSwFaPxz5RvxMBpWI6ikwhseG8zEVoHJ9Mky1G7Z+H7u
nsSvnFDLwqmGHxBvEKxpAcX5JL/KMyBI5vKuMT9oMQA7gHZsg+nOZaZlmh5ZlTf0
PYZmRGvJLFgFOVlBxHNoGA9oLhthKOpF7Z1kS0Sqs266EqrpxXQIHDa+uCetY85A
dk8XRnYnGJr+nxycNLysSQSgpztX4ymC5t78/Qp0+Wws70etaKjiAo0LCC/XmUmQ
ZSRhjDMpduNAwLCVR+w0W4CzJWlW8lubIUcbVXxv8nQ8dzQcatdK/4tRsXjt4PI2
CsdAQsKj3Xa60dHcz1DZiyuLfoI7wO5FJWv9Zai1SP1WyGHIF7RUbRbo8O5QEDJl
phe4jx/RGTbT23ABb7gUcGw+nCt9ALyAAhyqeHHKe99rYBmhf7ljYfE8DRH1duXk
+Na2TqP/W23R6RXQRfSYPwpQf0g3aWFDIESKChbTzTP9fleNlnf9ac+8fW4hAIg5
iAF+Rm/Wa2/qPDPFWqwnm4F+ghudAlJgpe9on895qU+gpmx0Zl9EWd6hubE1BFTQ
sbMYsniewD/G6sSrUSPRGizOULujOrfGizqxT4N5agMLnjnyQJ3bxlLG5ZLKBki7
dHpHh3ojdECBcHGZtVE+So2wMso/ss8+z7D5UaAY70UTITj+jVumy+E/gcXYNj91
/KLeTOrD5S3Jppd9VFNatEjIMYaR9AoH6xFCPlrX5GjXpodjTRU5saZYj9vWkUNo
T4EJ3S1EjqGz7uYvY1W7RJoDOoISk3iceGHP1gkbp1bMgEMmjDb+iGNLIwOm9o6c
lzqrf1KbF8mHjy84ZWiIOCnFA6gIReCQFOBYEnVyPvPIO5NaTnJqqr6EICsyU1hM
Bcix8QSbGg80zE3LkyOAPoFh6EHv7VjOmUouVufkOeVbJU2QBymxFOQvd4WAvhm9
G+p5jaCYxk4ow2V4BDehB422lt9jAUxI/sE6Vu19kkjECMa5Y9URy/SG2y8Txj/L
1ogKtXH9kCNzWDZ9Wx2amCI+U8aLAjQFD9Fz5HANoUa538PvcIMdixNP8FfBrMzW
v3XgYrlnQ3GrodNJTi23Zff1iguCowWMnuaFeNwQzHVvbApS8YipPWg1eRRF8MMc
QTWC+fpZBzBC/QNjsL5TL2CjZaXzJwjQWrrds2VC+QUn8Y2AOced6ZgFLFYYaeRe
+zOGu869CHcOujPolfLGVkOUvvIPJTO+n1FamyIwoPolXLCuf4wkDlO8KQE56euA
cuBOn5ZfO/Y4PCzufcQKkaNp65hxYoiVn/pGrUlAAljcxebERyAv0YaJ+/H/O8iQ
orHgmun35sCwrQRaL7iPPKFYLXqoFhMwT1f0lWUy6TdLw4OIe0sKqmemTJAQRPOO
4fMFt1z05BTAZtaFvdyakei3PrsSDW6BDSje3NMzcVbZrbRUueaiiCcahrBYXKI2
/ROnqqImXG+yy5SgDy1jdWjlS1b8N57TKJTM4P62Qevx+eaqgzMjdevq90fmV9BK
oEQDyO9dosEVW6J1nqOtR3xBN2gOlXfrfvU3yU+NTqqTfv2oObW2uAhM9eZDVI8V
XvUZ5yKhHbtK4ohe9WS44TVHdLmFpH2I4IyaEbaiRQlJcw9yFPDaymmFAPnL5HpN
Q32uIXBjjnobHYozeomAarCIbXWY/3ZAZWT8E8F3auzkh7QqKBjvNF+3v3RBfp1f
sFSMYyAmTIOvLl87+mn+J2UWEmHjC5ugMWoEZw42gjX0H0yStMUXAwlum/GFW3xl
Q2HtoRzZUta/D3HNpPOIB41hHN16BA7wQVDaAxYFrc93Gihi1ozbktbc2uX7HVjG
SaQSwj3ukRvXtCQYT/kp6bF1768drZFvkFiNZ+ZvJi/AOgvNWkRSNGPy0ZICgu1b
faJWGwJdQ2HTuDG7ZirhifrbG19yAqvx37Nlqebn9pPL6d5BqJXyYDEiv90jyJOu
zkx/OCrzMokvDgKZAUmQAXxDHpb/o0bFJsKMf9nr5A0pVlkuAbTdHoffE7/2teIK
YSt3BJkorNEpPxjGEXNvZJmsd+fkBUnnYmX64Kz+oWsuKXNVCkLTbmteiaCZDNOe
LJgHpd9JEfrJ3aj7Irnya+SYKHrzixmWdxICb/yh7W0HlYvKFNXdULlqqbql+Wa0
njqEL6fCtGTefeN8FPW4AYNJoSemByoWUiqz01uOwkGlk5n1gKpU3AhcivZgpWNl
ApnTB3B3lfhHCeQcohGwmrrUeA2O+FAKL9IaNNTVIxrH0+9RnsPsb6AM19RSc6pf
UHVyN2ULWsHj7zmIc4RTaySH0gV1fKr5bsN/iHtTMFq0/0Nl5iqR6VuWTmW+yWHn
6dLQW6vp4PtT+KtPIsOwGBs9eBWU+QRaAVUzXxsCSw/U5iMXS83Nv0jvI+2vLo62
DnO8qxJVsEsO/1a7P9egeux8cqP0Kp+jPJIZ/8be2qV21R+z3djHv3GhyPp4/XzV
6ilSVnGmCE5ufEOkrnADmy24DfPCUDUU1H1EzhiFZiImHFmKCGjqsEGRHNWkPas+
Hpzno3p4oUXz6lq1fIPRaKdlqFrsv3z6xKh2gisIfsSRBrvsS9ZZkkS8Yly+Nori
0ZtnKBWzSjpuZ6RiS/k0TG6HMW3mxhtT0/uhLUTq2nXXmMgYoDa2Df0rFApmfTJ5
7MYAd2cFKHTW9oDonaUvrSjkzHr+AC02cjMONUhfFM2LmU9COtcYeBqkNGgCAzof
TarngDbzMf8b6xaIPQZk3ola7Gv6l7AE59k5kMPnTEgLjDjR2w4X8GfkNRkltui1
1Myines+iUG55YD9OpOzUT/6lBV9hMTamloq3A7RdDxII143VLUaNm/jUasdWoBU
q72n8s2NDOxbKmoDRT+DJA2nFGx0PmEsr3vIczxnm06UVIowaPsKSwFj7LQbHgib
H3Ah6p4/7lf2PdhVGxqR/eosKl+U0M2J9COz0VW8RVsotITsEaVLJM0qCQ0z2HUn
UFPlDNNf6Zr+g5rpREWEvKAEGl8LTycJ/z41QQLMXLejB5Kgf0A0NnvgTRGR4YJ1
uOIS9akypUKEKlyOQGAbSJiSVzhAJQTtHzBioitudcKY/Oqx8s6B1cbSjcVFy/kL
jTR1CbpuGabwodi4VbtK/ORuouBCv4kF4pQKPKkbq1rS+g9ZPJRshvULN+DvDb+I
IGFmBL1f2MyNsPrxGmgkQBcwRreussrmBASvmAt7xAIiHXbnZBonw3B9NIn5nI6h
RHcKLiE47RXzOoyLj0NWZHVY07jKgSBsNcgEn6bKNv10gZ19DCrJd9PnRbqw6Iw/
JgkADF6Zyl1/0t5A8DSswUzIGq41Ia4fwNMPNZfw7HwEOTAjHWpOh5Pk+kQxEV3M
L6BiTysAqWTg2m5sQezvM33zMiG9E/CBeWofCwHTluf+xW54hnPtvDZOzaO46OrN
00LqMGiB+AJEiuU0rutq79sa8c3t70ZsHNdWp89xCzq9Q1j4kDynIWQlxO9x2Sd6
lzMw8fgUfaIkzi/ibd+D2g4whNHSfzy8laKr9GLXFgrx0Jinyt2hIpRky9DGD/FD
kQHYZqXjq4sQzf3XAlvmf4Kz1M4cB2DYzNbkNK4U/+OgAxmYg/zeru4H90IFVw6W
kBIIAcVsnc7bu5/4fRWGH/5MRlbSq54qo3fZ0XhJsUq7daZkeLDBsLkqNNnvqr+3
fdC1sXu9ZqcDYltHZ8mvpZTLFi7Libee/uCv47I69o1hx/xxcAs3TySRdgpHmV8t
cwfYaSYzZxJFyNG2T8Dnlb0+plnLrcqrpAhJn3e5GHGWLx+KRg0iYmk5ZkWKSuzV
HvHjiDiWgTC8XDW29sMvY19XhzEn4UOs4cbxYHmtBUVB4oqX1wrW1+0ONktfJ9WN
trItx5NhGJABDnL3lyP1sP679TttGiogIrwGNvYbUrE0XNl7Ff3fSkZqI3YJi356
D4SXotZjMr6O0gZiqghPLQrFH5jX8rsjMIortxLwvuquFYvnMi6qKM/s6ysnVfJZ
F1qjX3UEc21gufaGT+N8Cgn0O2i0vALnsEKmFI0cQ5rLUHLS6YfNMf+Ho1qgoFRq
/aDyxJ6+0V4SevP57I66FfBYOWz4+wynxLqww/DX4sj3mpDTcIPd7oSud4MRW1hZ
VyLcledaLnshzxqg6z7aSTl5Amxq/FjYwOfrNflSWU5EoSjsIQQd76WAwgVJoapu
Ckvy34MHBdmNEzC/iKEtTOyzF4g5qeOv/PJWU2HZV4BKHOB3eidjcmHh49WlwDT9
xepnrOuV4PqSUZMPHPKNL9gD5BiE6dhL0e/7NrcvaAOaYTdNXFtBBW05ougYoham
uXtdAH1Q1p6blObEFZVBG8GoxuEWRQr+vj/IT9XAJ3G76XwAiP9xrd5Ci2nePQno
N872P2EpkJXoVkc9xjkCAUiylbWHXBU3cEQyiA8aRcCkc0ThMs0QY6h08JtBghsp
heir1TTjE4ruyLB6te04GaRXagySehvJDVAStNUrCPCqSU6nprVc8ioOEUNuamxX
yUy1yreSE+v/lKsdr3Ca+fb8uDDOnBxrIJeDtvWo83IqOTUE89kJz7kxHzwam0+m
deE1aalxOxBirhLukrz23gSGovCINU8KR8iAwg7D4kaBWfG7l27CuW+D0qaRJ5UE
eBoQdc3+FzsE+fSBZJ0HZu/ioMzGo1WT3ind604HjG848J1eGlirZcite1Dun+nL
6Z+6DEC0qHLtBdVU8PVjUsgGlbHlm3nf+7UWh6/1JmDfmQSfOahrWlzz5t+JzfPX
wnPr5ZFoHQp7KMdAAWmpeefUI/8qz7TTrkhqzuRCPqoResXGJ6vVAAjU+4VYmgfQ
DYk/Bq0UskScbnPwFOD/0QqV0I1rVYSmwzsjy/bRN98EkUtM6CeskHgbicEAgRKw
mhZ1lrhpaCfTlGzCdfnb+GgKDNt/SQ3RAJ7rGUcjbiUYfO1g0g+QleGIFWfwYeSM
VwLhtsDKQsU6F6XwyeVGm77C3AmltXlZdtlfvX/oWL/0nIDOAHgts0DMvm7I5RuH
tyhJShNOnWkFHpo5xB48tFT9+c8JyTqkTSN41DsncS4xnasdz0N/BsvgykPW9tJq
zsgU0ylPsSuHX/NdWNO7drcuBx9k3+dMzm3upOOZ4WBU871PpkGWlCbYYUut2XYs
9gB5743L7QyqN17XJOy5doJYAbAr91KQTtZ+kQDGCa/UmYyUl7nku2a4nb08EO8X
UyBCJUK0Vta8Ac5Izc2pQehiCxJC5cFPz41bL99ypnZX8SvUIqFhg/28MybG17/Y
VIYYlDTok4grgC4oWuv5Y7tmTyXhK8A7a+V/+iDVBZl5OtQWzWQpTcO8/AVPTSwo
E+/3Un8S6P5qgTSidrlNurGMgbbKI2R2w8/e4k5/syXfXP3plrJnF/p7CZ6T45uB
PV0qKfyeEETlHnBPODjEUNcWjkVBWV+tvMqQ1BRtIj4Mj48IXzoTloA/MO8lmTUE
sbjJac6Cn8aIia8bA9x/uMdAlgO47gtMcvj6U99BEepAVUgou5+sbTLaAgSNcKbm
nDSCHwKXfpnzh82vQaG1ayqzn9uCdVr/TXhZBcP587uqV0VxJcgwurOo35Xa8Ued
sYBm9xfDQpWky6tT5aMapVyDf/lE8pLVGH0H49gthK9BqStDD20/2Ad19dS34KBn
4in4qer72RqDkbu7jutq+Qyqd7LGxaxgS+kBnz3q8UGaoPfUtvKAGBdKA8L4yO5T
Olk3trw6IcIfYvxAd4mfAZNpayKyPtrA/4ct+2Bg+XKrtNR6IFUv7QG/8RPU3srp
nYgFxEWbopInFw5mvRRJjUVhpSG3swUMmI9hqqbTqzT5CQflH2iDAXviqW8rzjct
CjAPSNlmIquS+Q7axDgPa+Wn/fA3e/3LrRC2wXP4EbnLYHOt6OPMyOH5La6k2JmU
Z7DvJD9+nnRpYzETTENVINUOjoif8/resNKffpApW8L8l0w+/dQXGoChusxGTYXQ
m7MX9Pk7vZ/xlOCCowFq57TbbLfvzyZHHdSTy1vDqqRBhgf5au4/wMgFstOdRU/6
8k36P2PgS9mPtsxQc5RVwyzb42oD6Q45yNdntLLJ30QoxMbGYKZ3J7Zp7cIpps/u
GtcKjwarftmfdXF+8LbONPiX6Zj3zdyyE7ypoXqwbx4O47wsbXpJ2ZriToVZk7ma
2gDJdeLL9yr/2tCJoKB0HfTPtEJ/QWY4bNkegWXRFwp0GrDqqCmGhRHqf/seVvdi
ESQFYFbnIPzDsLxg9/3qG7+XFbz/FK3kB8VSGSxtxOpFu/iS48wbhc+12aG6pK+N
S8fNbpklvJdXnHIihQbBVoRa2PW0xQuUsqzG5DsMbY83vEIoVmhZW/ET6KvxsoHQ
KVkbo4CA5Pa3ByDuEpZWMQfCCq9qqUZ1EbXC/NDkOfEHpH8G9NwfUUbxg+3o3i21
v5WHYdmIeXih8gAU/aSpRibaEAmxTD1+DRz4wwXli27Ym1zs/TRsRMEgxVbWAc2i
oL9K+MhcvyuwIy9/lINJvHpj47+9oUBem5QBs9qgE9az+rVjDasAezBJF0lbD+Hm
ssP5q4uXwAq+uHk6P9kLnTs0p+mBV7pj0dhRflOKV3xnKtJRi/pc/GjUXhcq4mX2
FTlQjqmclmV1wIwpXTemrQs+mY/LcM2L+HxM2CgtD/NQVUuYADIsOPDATMpQ+A8x
UMG5UWHVl7NuCHO6fKP7XBd6yDPFl7WMeHMKtRRr/I9dWiXqVv6SImo6vlhbAtQJ
FIFLYMh9RCYS0qGRV2ATF0Kw1Nsc0yBSOiAT3jmoShVXpqE5+8PtBWMXF78xskCg
fXhkO2PZFHFgKGk9PpUTnrxc2JSoBSmciljngkEtAS7Hb2V5QHGqcGbm7K02VwDd
P+H+6PdgJaHr1D3cSGwz0qRJpGSD4zjxKeu/42gD3UDyxzu4R1KOC+rZWFkRJ+WT
Y6okc5i7nW55wVAFPzKwWPIJsnxv/C0bFtZ6678G22o3aDCGYXRutw5WyReYNGXM
TypEddblpfFZI6wErAyXuX7vRrO91q8WW/SVblqHcNDr/Q+KjDFuoL+oinDsyG4i
IOGd7sxCGZ/V3jBxnXpYaitnNhmHwczHWPYreYoRw//q21DTVlnJmiqq1ofBWdfD
CF4ftKAH34JkHbP2N3rcjgdWdM2ZvARYpk4T6ysJCJKVKUixovTHx4wdrX6Zk3ky
5wNG15Katv/8W67oFAsW/vB2rgKlpKQAmHnmzcNSe65F5GaSLuSv8A9YHV2y92dp
o5BQKzp0/0IEXGPlNPUJ+aWDOutH0qcjeYLo/8/qJmoBkCSLtSMTqI+kMqUfqHgP
z5PiYNnR4xLwu0hz7Ukt+QLAF17NgElNxcELeEQ6z2NQl64MuWnAEGRxauBoMRlx
Phr1vg0TpPXn7QNm/GybVUDSDCIEYgRpZAPxrmfbp1+wB7QC/KFWRBDhWyxwviqc
reoE05YHcDehw2+kEB4J53rJxjPLugj5JYj8dBKBbxGuw5Pli0amZeQtLlUuwa7F
kaQJqkYokUiVENru0UfRk7D30dZRzQJOCd8xWfjViEIJgWpdiHa/hq+Qp9NFoAzu
PTc6E0e9RpMY6MFm1DTznt239/0iVH3FBwXcWMRvmzEVA8VdXMRb/MGljIUfD/aT
5dJlAPiQ0MXTsSvi4ohZ/ISRp3l/MwjyAeH+UyOg9X5UI/mjpILX5VI1SqZMv4cN
xPiasPXpqi2fDMitsrFCCtp4BConcWs5mYWbQlJkt+FKA1NpuYEl106qiTt3PByl
OIjJ+/DVJ1sRfbAwt35fsfVNAR1OH5ThHUfhmN6Hh/pOFtcSDDGFtuznbF6Ct8rB
8odUj3yoQZely+DQIqGjkbDLAkyliVuog09b/FU+MNlIfH+oDgXVAbiQvPepg/rf
QTorOo9Qfxx30Ii0RXsM7w8iSjo3yGJmmTccLyFR9Sj7ef1OWLsyfNWOhRXGsKd6
vNwLgTgk9O5HZheRI5cE7R/yQ2oziYaok8I/cVuh9OZk/lRKG27DqMXtN7mFRK4X
ZzWT+pMzhfosKZfCHdd6iWaBYCmVgvTc+gupmWgs3ffoSS+FuuF5l2/3jNvfT8ii
2YdcI32Qxtj2CpmLR4Tqrs7R1rw57wmjJOC0j8BP4TPzE1D9cPskr2kcH0s5fYw3
NYpJLZ93SJjsxBrj6ohC5h0xgba4+oKWPD659oUZO6yjRVL949tv2QoWBgMWh8yB
HRXAN8pickCk9s+QzB9kC6Y40PZ5Wzs14CEiLd7NqYoICs8+80KdHwivHlK2Zzfj
eu9za6DYG3PhrC/YVC9Bh4R4gHcD9l4aShIs2ExxnsAhTXhf3S8TKdcVntfptDvc
L4NwdC+dNwNeqs9gGxqzU+KYBUI0G+8a6fjB3fYbcMeVe/7CrzCzie5JdqfJiMbs
2hJPXPrmGvxAajwbkF+Hg4hWOVpWTdZhQWOwCd8QCmxQ23fp5B3ID1pwiKPvfgLO
BLJlib1yZxkthXxaBwzRAc2TF8LX4zN0MykLdW3U4qnLuAt9mJTaxMi11Da4DyyW
OPpnX65q+jPi25Qh0QwLsX33h6T+NuJ2Ft4UDSUOkxy2Fz3ux7DG1PmovfZYWCcl
cUlsxduoAVbnZl26L75tTDZfw8+MkoHFPeT4S0YAZHC3iFzIslgqJHB5oFEXQWFd
bn3H/mtv8UT+Z2KFiRU9OXNe2nVRRSazMeC9J26zgfrqtQd9Gz+dLM9AvVDoVHX9
7dgwxB6gR5GFPA2pYRlkyQGe54+G1yRXEYKcLC6jIceEnEV2JYvfQQGivSBFq9Sb
Vo9tS2XGu5C0Emd8zwk4/sy7qJn/PIwrDUmPIe9xJXy5kU7DpzdkfKEjyaq+etNY
QKHCzAaEuUBKRNnZdVJpdOfHm0VAZK2vtOAfFzV6wOSQElr6oM4HuYWxjoyuI884
wr58aUPadGw0Pj2n7chAnMikFja2N79EqG+OrJfBP9OG3+h/2qUsJciTrXkDlrb6
0VyBStS6ymQ8kERbSYAJQSCAj0MYgtGCvmB7JCq/uD/MZgvnlBKskfJMZkfurZYt
6Hz2HNGzZTEIc3Z4ttMQilknz8R6u4w9Yo2A+D8hOZXfNGEMyXbjSgZ2TfxAYPTh
H966D6J+ZIOmLYOZgrWfq5OB1CfIZ9Ql0CcV+9MtU7SondkClefXdFeIn+nGvYis
8rSbZ85L0FvJEoSvErJOlJufQyZkF8cIQsixSdUdBORrd32MZ3MBHU00fKmnATgL
Vnp89niNzJ+RiZuZfhezeBshTBDModfOW8amqHN/LUxcwuhIhDj5t+Ilz8bcOUFf
pNrjlnmw+QAu9EQvjDTUtiiTvdLPwPaBx2hk+MTpdegnfoNXS4L7JPikCyzk7VDD
/MU2O/mswkizW11OJPhTe5c+tErdajk5wd5dzYpmLhmN99SNUr0o6OilN9UBRtHG
CXFWAA1UzujsopyP2aAX/jK8F3qAasesfbzJ/wmWI9C3/RpQ+2X8q/JfwmTv/1by
PJyzRcw3PlZhG+h2uYmgjQj/jvseUl54qCCtiwvY9+k/RqfMOcS9BhKarJBn3BSr
rIE3l7Go2i1K8R4F2KC1B13P0Sg0YyaOlcZS3x7jCxwLaIZBRO61M470sK7kOPKe
lT2nB5ej4BT8OmwXu2VfRWqqywn+x7+hW8TT0G+AuWebv7ez8aqNVJIuWLqkRaQy
Xan8KGv383C7D/XjECRxNwZPfzc0yP+Z2gGdOlh8RebyM53sdxomBNdMp/7dAd2q
o3OmSZ6q9Un757bjp1TAF/xnjHw7gWvKLVTbpiWAy94ytbcVj+Y9vjqQmlk4EgSp
L4NB1fFRIN5exMiKPEmrGnk3v8F0njCgpqSToe5XN3euLdNrbZD8p4FZONlHTkLM
zIjvAmkstjykDv/LogBNUhqx1hOaqSGbgBwtnqbzMgaiBLQMUc2/9dEGmYCxjaAp
zmif2nt4yxHsGaj0yxQkua7hQKKV5UNKdVAi8EY5BzG5SyfKA1tjdKEcgLINCIVT
76esUdsgZrOph5lwgcrgEtAizpSNxCzSohHmupg03hrfmyIqucZimGTCLAJWt5Ei
SZlmhkmavNeQ4WR0KZ0O0bcJIYnY+2u+UOhelrLvHU7sC/WYuMPJn3pW6Gmk1mYJ
e0m7ogwecaFV8LkA74KMATriQSzd6H1hZDI9gChN1R4kF9JYxx1jKin18DkAUN52
N8wr1EFdcT6fxdVKp8iSJd74XHMCdWiRI3sR3fy2yJRiHZAn1LVUEHa430wPL8am
jkICQWvhL49ahKyEa4icmFoHgeB30p9DX9saTwOqXJa5pUAWAsCdDwFmi1Thu44z
PPLTcepcqiK8+uMqrX+Ch/Cpbhc4KjXCm+BgzionaV2VBw4pHYbx231CJUe/OlWL
HWuTJxMuHXSTbNR4rwY1BgwaH21+6DLidj2LrT8kel9iczxFE2hs/hB7KAksJXAg
P5K+HrsaScjtTd78LbgIvL2cWP3WwVa7P8TxOfFEyIFrZyc42hbw0x5Zzgfx6xSz
p14NMPWU32AdRNVo9qHosEhcsPyX0dQ6wFsbgCMtZI0+RsFbcah7XUGGwyuz7i5H
IP8am3JJZHqOAttxKkJX+/C8U0kWlhnLeTni9P8B16z4Ew/ugj553O0AyoiRO+w9
82AvszncvlKuFd4dhDHobZmfzYOYk0QrzjYFiDKpLalD0yhah0wdEAEH/Yf5D6Ke
1nbYMRpptfmPd5GfTZ4jYjbgZhY2F6U5jrqQjyCaSIQZ6j6EaGTXDKmyXkDdssVV
NO0PZyWJAoDQo/vFRNcRkS8Q8fGSpNQOh5dT5/wxf/aRTR1PSAohFp6tB70qs8s3
TZpDa03rbg0myp+7xLOmqfmQLvr6S/EOyTQiKzx3wqapEzVBcUI7RqPqAWXpH7dR
rbnLPXMUjOz77oKGBXgAUIep4hsER9PdUUVGZZzGLO6KYxjVPswdwEu80uwikxyW
SjI+QqGMGl76PrsWnt9W++v0zESDj8G6/SgMrfpm7IQcHc01lzrIkJ4TI4OrfO0Y
rRjMVNduiidpdyNmulfgXFt5SEbUC/d3hBqanVdpcEluiauwDEirDikoaEnYYgw7
6/mqwlGaOT6iPhJY5QNZAmKyH5ccshZfStj3xoV3ABJTolwuMX3uX2tWjL452kcd
/Gj+wKcF7alBA42hFVzVcN/T7M0sEHPi6eTbeSQz2r5wRPrYaqBd9wfA/4iJdBMn
mo8HmTxEfgL6OeSuSe1Zz6wHqHyoAFn0eleaVnHTEliXtJU1e8IsyZN/daEG2ynj
abiJprUGATcy/FtfRsXoj4uW7X/O1Sdjr4dny6gZ2MhfqXV0klGSAtDFBh7lqJ7u
Vor2owDjTmdWawNv+fBTcuAE1tIo+eHRDQJND7tm24BAOfvaGZYTMP3sp1kGVcgk
Qut97TVoK27rcDLtd4Jp+lk0CDDXi1VXFVoyQjmaYQxWGYKFlWPbZeEYJHVr1D9K
hbTM5GyMM3e2dpD/WcaoLDcGOMXnIItOL/fL7e69ZaBoERZjol3lPavTb5b7slAQ
ZdXzdbAL21F6mB6GEZmXe+e4pXn4S6jFnjaHt5nvJkVHv8OGYlFikd2BLBFwwqBc
Hq8JdGxPXF7RTIr5HtpJaRVuapmntYEggpVj+SE0x4q4RCwSQ4l08zveGBvm2efz
5DF83qVQdKnjGyyOCSzk6NgHyZN9S3YBgAskU+taKL605Q1eKNyaSiFmtTJxe8AV
i8CIy+NemGoyeXMeN+oeDgULVBJwiBvjXhmyuEXC8ssXIrpjAWOasnUNA47NxfqI
Z4H9wsrXOBStUff2klwsXPe83E6j5pEnaYw+fljaVyn1fOd4k4jVJRS8zynbzhZ5
g4mLUwYe5+WXP/TDX4hFHTVmfGEXOCNUairaE7JNpP9ClW5qCp9SjpQsqnMZwCw0
bAib9F9sx9fnY3RT0JfWEuCceeV4/LaLueaik+GqxMrhnMomIRvb6PEkWZjPxAtG
+4+EZxrFLx0sBR+jnSiDD9Glckhux3d8t7+ZamDBANpSpoz9bgIwSZQfHEbE/7QN
OC0Ksc00kbBgF0pxWeshTQcnsMmKBhebrbmDKvbtVnZxhoTiHvNS98K5Jf0v0URc
JA4p9Dp6O4VbwVJ2zjdZPUBlvhMzV0FbF07zYJx5rR2SVGxFfOvab66g0dLyrqlh
FS/D/ku3AckukQkxpZHJuTS1CWd+wMTBYBf1fbmBnT47wZeTMNdVjhspSEH2SrQ1
Z+DGerAPikA4oBbNEEn/RgV8aDimKtT6MGYJDWdN+h/4FKrn3/jZJXKWTq+WCK3G
iqyLUBNVaxkKbX9pC52ZvCrts+WcyGR8NKaQOQDBRpi0SdaKPNM2kYycTKb+4CDC
asp+O5/y4rQJ3hYLc9qTqDiYYzm7HZO/phvAoRHQxROl2G5ZGQATfsD4jFgIqhOQ
iUcWc9XGRQaDQldI5lnRMPPlCa0pvlRbYm2r7NwLHVLj7H3qEHUeTizs8ZJ1Ao7e
5cy4wkv5V9dgnwpcKC86uBYS9Vx9homS0e+n0amnf3PdLFvSAsb/gPUF2j2IE5Sb
/YmjJavZKphoKyEPds6koeeXCVR4+IcGHHEfxqZag1l92SEcFe8kUTO8BX+CEdD0
w8qLLtiA63TI5pEKTrtw6iC7CsAoK+5qTHKxzpCZv4nWxco8blwihyT8JRgE1AVB
VdZ7V3AoU1eKLCmaHGCENET0gL58WWwuG/zQfoHKxBxg1xya3J/q3koSJb7FZSWZ
hp7WxOsEIXvL1xBYOqK60SmQBJkY1Iavu5edC7d2QKrymwHqyhW0DJr7SHF46V7D
JGlflK70Q1Rbf7WUq/CYsZyIg7MIMdEXcdOdisq0qYIwM7/YsWOqqgl24CuXUTxk
vEIeco5KknILnZ0FLO8YUoAdhV8VbvmLP2Wj13MwpxsSErcHoDiBZ5sRmZTtFVFk
CtfxLJo18QHCupY/+idIjEe0jK4EOFaGaDhjAvisTp+qqyh+PpT37e/AYu8XZjQw
XZ4xfBdKTQVjJrhfTyFb8Qu+XU6+7aXYJosCjsEygXoGCzlWSWEfmUAecx+2KOpR
g+lpSiz+bLvf55QHT1eAkZISgY3C25bKxiYk3A1IbdImmQ8Zs3hISWaadbhf3Ulh
wK6atKi8ZRqtJp0jxIyzXxWyC+jgo716IOM/8eW+tO2P9rNO9yYC6o+o8MCxCyUR
DT40igFh1iedVKTfxKY7aY6nBabmHvKsLhzarM8vbgdxuwJMkwP76Y5TvoJzCsOI
MuC7Yh5kBy6gMYQ7DHLlrqohYg0JYLVuNel6CMeNoNnb5RjPfrxL+1yp6he9jg30
PvuX9NjsJlv5UN6D0nzwFBG7EyrrDvdSkQuqRvPusaflWePPc914dpwaUY2qOmip
P5E20KqKgSvlRc7pHwvu5Uy0n56fRs7BsIWX2eF2GXyy3cYHF/CVOLBeLY82flC4
rGqN1uJDolGPtxQ2vD/SSfylnltTQ6rmd79RE4Kw4rFTkKzvUCx0anra/Cl98y2B
WbTle6HnXvDJru21Vtfqm9uuguhk7Yd7Pq/Hsitjtpy80r0PvlVNcEHJOSuU5+ph
oUkt/4I1tRGrGgTh9KEnAUqhGnZ3Sih6C8Mddiyp0gI/CeC6JJozTqwCl6ny2GLQ
eG7kHCePh36rXXOg/VVdC6cY3zgPnIK9xrhxeQPfNaue8a2TVIrfrrKDFCVZer7l
h46mOzH+9hi6AoJkURU4YeipaHwzHwqEE+yqA/4wXtqVjTGC5iORA8n0txGJ8ALg
eZkHhUEwDS0bQHkqyOyTuIXUx86iobdDQwIbJsmjsnUl9lqwgVZMede0mqhzGurj
Cgo2kn3M+e6Q3NelSLWz5OHifXGV4EbHMtahLi7FZOT52SbBYkKwsV4se2wLvmtt
ai+mNdb0zeiXIlqDNcfEvrKan0Q4+TCrZB+UN0M66BbAKg+uwRs0NwFC2up1szSD
tQKX0GmK7aFJY/4kiT3zeL0PpIMFBpdCLFWUx9ljODljmC+KjRdSfqgxs3ysDvfT
CEQpul3hTusZYH7M7c3E07HynV6VbnsmrWAUm9jrYas0TqV5F29AkFyr2cGH713v
DCQX6yHTEhR9vlO7JI48jU5jPV1dN/taCCOy3YHpK0O6e5rEJNlDgOeY9jAP+su9
JRAY5TGbvJAG2OmgaFXPd+Vm4kMq0N8CsBshgu7KkhE=
`pragma protect end_protected
