`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oV8DM1BKca60L/5epa2AdeloewIqUi0Q0miHgaCBjh0jSr4cHZtngaA795sg8rW2
ychS0rQMq6Y6xsUoeTu5wirn136D6I1mXMH3VUVA2A+Saz2r0jkIi4jEFzZXDvFm
NT/Z/EkUPmH2ChK26NUUemUjaLRof19v19OsCda1p5Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33696)
eTdO9pHNh7lbaY8bch1PkOpsHmKbQhI+27d0F3kwGkx7UhJy0VTdM3oTA/horSaZ
8AwBKkeKWgoGhnGGVWWaUT53kab84KmYI2BCuAO6x5qhUQ/VEsvPfhaq2BbBytK+
/KhngSztHh5kFJvr3HUlVE7HHPzbqiKSA0vABlN8PITH6DF6dBP8h2ciZiZBXh61
i4/CcCnbT8+7BQ5RDfBCqnlkQaXqUa0vLSWlADWE6Fh6dhKklBDW5DLrQOCSKkGw
JYY0rjZY3G3cAYYXshi6QhCUqKuWMcTRcEGgRp5prsRp5AQLU8Dtp6ysg9TscFlU
oRVqPVgTNs1d+5uSAw8rLa4NVvgYGY9dfJ5gks1Uap+yCN4qUTt6WkjpDx7J54gG
Xy2cf2cUFCI9Um6KOWHOZR3SpDEYF3pWZFXwVKs9cX/8fdHLn6TQUaqcBpQElZM/
PNbQn6Ya0w19Li8PGjpaQQvC+Fg/RvwGClhRZKkS92MYAt1U8HWhBaOAryxaTePE
ILx6JrH9b/VSTrjfDsrM3TWlM09eELr4BeavQ3gtV1eolKc9qqoHJcUg0zEHBsLY
RX/y2rkXFyWAgs89nOkmX8fYwCYCk4SRQkcX1yk0laGYJF16gzozFuwlWLFP4uNH
sr/dcugHJn6PQmGH190shRfSZ3u6Stda+3HYk3hHOLHk3zEWMakwJ9InFfWjqvDm
zR5usyocCsmDS94lwG14JWOvcbpFCdPQ9IWDVJwbxAFmhHMV9zjgPc0z3mHJjc6F
mjmwDxgkPsGHlC/vPHKFXrTpBsz9HajJbGWOJANt9eno3yoc/289IsvxyJlmxZyC
jfltqygzJm2ojEqO4ZE0MmAwn/34n6GxOfYbwF92l7w/u/35Gfa2pnSwpI+OTiOG
Dk4sCar9YSpVYFDx2VkRph666JFPx9POmruZZPzj+aVQA0N4Kxm3tE0zdjZGlDpw
ppJ9nf3PI21697JBMlzSBrIQ0vdmfpAznU/+5AaAGEp8ZC4LXVtpQMaMerEb9G2x
OIlWLV/dKw9G90KueSTeuVTGMgKCa3SHJ1GaB16v3jXlaX0S8jx6khgruiukChrY
DB5jQIZHJqgZlRjPexmY3aMnqpExauH/qEKpBkPjrMB3xrvf5cbP+QKjvy3eYX4D
OM8tYsz3WH/Bg+g4uojJVJinvEJLc2hQ+Cudo2JSDr0hGbUp2vt/rbXBqII9RHO+
9nSlB7/CDDCIhc3o+XAiaataB0Z3NIRQZ/eZisNE/3jSZTj9wVj8s1Q2Pj92xVBh
nDS10/GkSJ3Dxu100P17R8XOS6v0c3L02p31WJbrq1eYSDBHLhgLJwdpNR1sJGn5
dFs+fw+FM5Q19UHReu5RP+6rrd3ZDkZqGGXhTVx4gA2Wwpej4BdMmL3UydpRMd25
w6j203vyXCKJq8w9vw3IN782YO4/fsn6lZMBpIlRGTmp5dwhiU3uXRtV7LYvF75b
qyGV4FRU88ZVNI77KE40my1I553sRoX+wMRtnYTwHxF2JZTUMYfCTflcbIQV/5W/
QPlA2f+Mz2+UTXIf2/OM78SWDKv4Z2Ozdw4Iz11ZNRG1cu5+hDHgvVfajw1nvUP7
NrbKKQutjfyctq3pIil7T6JjTvqvlEroGXZZwhW6fb6CVbogQaD7RAM9pR7EK5IN
ZAEiETVLWwiQ8U/RQs7ZNQk5/nSA0BN9/IHz/ji7uYA+pf8taDzL0pFIxkXZyNQg
oCKlTO26gB6a6b+THLgnTC6Tn3xpJ2uOdndAAQY01PBqJEigL3IRPhcamxAl0MNk
VHCB08T0JBu4pMTcvo3B8xbYJc5flgNBYjhKalQCYuuVpz9ftdWfzU1TA1MR5b9R
9IeNS2dqNf5rdn3OOhd47U7Ds9srq8rah2eAtPJehXTv8KQ7gZ67ceh7wGF7Gb6O
zTvOiBL+DXdEcYt9/VRiuj5bTAf323apFias/crzUrBIrx4s3IaNEKdhJ6RLgpo0
6f/0+lpDhlnkp2WLehBl/TK3mkcYFYE62PeV7dVlD1QfD3NsiLJreJs3L7skWglH
h8bys/fVPxKJPviKrku9QW3hDw7GTJO7Htm4le1il526YENsB2JJ8akP0X0/Iar3
Mi2/6NnhLSaSOV8q5PuIDW0dd+UqKqEDvus/v3uOy2ECnqMXr1ean1Jes2yIPpRh
aVvRxgpchd55pqYJVeuG10rCn7VIOE1FbOvlmwH+LvrB6XgNVYZJNGGIpFfc1OR7
PFsSU5Lh0weyWK6qppaG0TR5r0twt9jck7yRQDN+8dzVNFVytKcLyL2NCKbqzhdm
GfioNjneKnKSHiV4SvTmKChtM6tfFxUkd98FHHEkZEKkP1JosLK8h1BfhazYUBj4
Lec8KHmQRb9zPyaW9Cg9TOdAqnPom6+UL0XMgxei6glBh+RHI0Mq/1NCvvEIHhqj
Wij1T8U8O1LiO7n6ct6kgQRMBFcoZTFIUfXhymg2wkreAPfkVatvqQzyBNFEFUQL
cPfarZJVX0N5yoPtaHZDFu+Mqa3H8zdTXX4AWOzmINcle/4czH1crGjotqLFYX86
tLMW74Zi1OFL31nwhuX4FEsccW20XSwC1v1N9yRaNHzS012FCrqFq6WZtqckhbmD
MO0+OOmhXqYVqKKKGIIIyHrZoHJmIeK/zSoqotzIGxUAvT0gUcYIOZ90jgRIzRpO
ItmIi86/cpQZK0/Rfv6wSgGlEffNPynMHv8UUwZdXEc+U3iTZPBTm7fOWZ78aN9H
TJYP8FIbMx94bkGbEN+tUdK8txS3daAJ1Vre+b3eG2Ea5a4V4YhFKePOQJZ59aHe
vIhgMYDsPIdM/dZm38SEkRi4Zl2LEddW7A7WdbXI/BnEbjLwtDcvX3skfL18E469
Z052MWuThuaiOZVl/Z4G6b8DTwJgPp8SjC0dxGBgHbQ4qYkbnpgHMboy5liF5V52
7bK5tQ/14FoUoFfCAyRqPP4lBDhkblyaAMf7EjVZhSn1rNUqGNzG66a9a8JvB0ty
la32/xTZhJZkhcqi1KvXPzrrpzHZIEyegj5sBwTsubzTvRGgEYgiUM5JLO8hKncr
+p9OE88T75PDisljIBo1jTupvGgqYHMUssQdaS85sfqEtJcnjac5y+v3YryQLUB9
A5e6AbAXQEgBjhmpq2uwpqGLfz4/vquJfL7JM21cYzrNBT+d0FQ/of5qoB/Nc+80
qgO16Gwrw46In4f2xTT9jziufSFT2b805WbsQ3pkVnuEcDL5yQunINimDQXjIaze
8M4LhG99yrx4O0KUedGB0MsLRc0ccI50N3F8RhdEw8VNOS8g2N+jhicT+HW2veXA
YEZ/QSh/8MIXP9pvVx/XCjC99kmUNuzU+7CvYQhudSL547qb3qlHKmBK6XyKblCg
pvXifUVLTnsx565hDDFw/z0KVEaXpAN52NtDP661D4UDNO8gie1bmxKy9Y9QIpKI
G+JcSZxLXkR4f2QVAX7mnxg3XnNsRhNB+yvQyi2i6NtV/CLi9koifIH49F3DD+XQ
UZoKZR1bgzm4+dKiujTl0Pt5qMCyIj01Kfo/JxpQ2jAyRnrPCx8MUpPwYmdPlEFL
qfR6qDXSzX6JoeOK2/I2NTGGBWGCPlSng2eot7C+xIwbb2OYR0qgpUpH7OMh3oBJ
DxqjqHtmh/APF8cj+ATz+STVvl0fO0TnQkWLZd+mBcTxRBGD8sgYP3j12oHpX+IE
VzLpj2CfdoANQGNfReYpb/FPNqQTHAFeeJYpk4VP76Lp6GsECTUYsWUzt9YbaefO
I/nnmGR2wfMRV5IBu+fDBFa0UW/P3rj28lfRJAr+kZ86tOGliz1+I++r4Wf43edf
1U90sML8ip9Tn2cNYIdGB/ouI7qQtDciLvWDo8HBEFLQtZob+CGHtvnZZdniagP2
ni9BG7l9cylebW+3W9z5q2VLllFb9B5VzXwwzhUEG35++YJmCDApLRMTocUdZcfi
f/jdPQOzhFfa1MQsQWBQ6unPIZJB7cdtTyEFP6kbVOITRuB+B12J/OVCHHVAZ+sL
eTq+f7hoDKqLDwQwITBA6kJ+02fWykoTlxeqJtVhbTSFFzlC/HVzhg6hC+Um51VD
HP0fkvMJ42YPy/2sKk8UyLSwV5SzWoFWzg33Fy3djLsxrbgFgahLmu2Vq6qR9eBB
AFED3qL0ZHHm89BeopBKsI+kWPV6OrswazTiijbrGQ+ec9Rxj5FiA+YZ3ktRkpom
OPMWR1wlsb4gwPvTbdHAtET5wlUwv+VfKasFj575hKaqIT+zKqG3eqgf6IK9cDts
koIJHLgncRxdUteei8lT3G33RFkEekyk4D5w9Z5ds47uaSRyC18D/NMaZYDntLW4
251NKuATOeqFCmK5JbAZ9C+kJBff6XVlpwnP8Bx3RDjDILZfBsYZ4Vr7AWILUN6U
eHKD5AJjbx1/rfcHnbbB944/TOhBqoANqfeuZH0IYLZ363KbCdgTRIz28HI3XzRY
hYQ1GsbXljA7Iz+H8jY3K+eExvhdzAFQA3g/22VIFXc2Q0EqRKWoYlqaedUrQPzS
6bgyijbPmfqJVHdDte26RqZApGNYnRTAUGuuHs0RLZiBpRpZYxnqiWPPXjOE/DTI
poe3uF4uur7kH/0mKDXyIUdbtXcctTKAHhuRZ+9QEFk5psPiqaUEf/kPOqNQgFsC
ETUfa5LBg4lgjbd3KaDg6gqNYAV2GadHv3oPNqtPe0LUwrTHq8TxyQwKmB/e2eq9
IKNuIxEHv6kQ5gh7CZBovc9wvR8sr6b+Ev+Xv/vr13mCqhbALAW154j3gx3mWTtl
f/08vo7mZ0wqkuDsRaG6+RRaFAjNecvw/6ahy/A67dY9n3dsdmpPG4RUPwaPU7SL
X2VXc08cBE83wm5hNaw+jFTzjvzonOMJjycUkUs6bYMyDs4EGJMBWb74959QulQw
Cyv6P+Zr7SHrhgnjT0j63/mAZkEcfMTBAjpdeIdp/TLER3I1SL1tORC8z+gnQVRc
WnSjOv4YQ5r7XPyF5zvWhvZdJG9Em1S78N1lVxw2tE4Cwb7EJNIeaa7YneaPrj5s
Or4Jo3LdlqXVvbtVck/TlF9nq9M/PquO3DGOLDvfXm/5RRWo0gEMg42V+u2f6t1l
NB2Ztnxf5LTlgwBnGpOiH5sl0mTaQukvj37+HEui8jMT8dc2awR8B/DEcdRMnIcb
t+v3KqK53C1J+Vi3C/kcaNZUB4Cft0uPJyBtElj4bp9uJhU9ppvyTp29RKCVZG1M
XrBsLPrr2iRcIFc+2NhyP6ZPBup1fhNzBajeaD//U23bt4Z32tGsi5Ctck9SX22Y
ZqVFqgjJyg7AlcWfIHC/Bbjf3V+Y+UP3taLIG7sMyDlNiGx0SclCvL20Uj71wC2t
Mjzd8jxT/ZBenDhPY/auMfalB+eQJHpGT68rGywOvBK95NasbbnuL8HsL/qjlwHK
8akvNLCFX0bGlYWevdKYeshDRgyC2MTGKR+09EMljKuFBFNlyNZqmOcipCOaxMbu
U05fTOEGElAz+WiPGADPQtYxN6SMy76J8kunNCqDAHkfobtNww+iPcxnUr4JHddJ
kKfvGBT0Eri1YzsvsEqRmTuy0kmW+ZrheQIGfxib6U6yHkgHesGyFsFqOvTduM9m
UjUrf/wunqEiK7xFJ2atlbA9PtEUN+ct+UHjZ4ap0+o8NKCEtVSiuGl7Qes6za0s
Ka5PcY6uFZw091ua1r9ususBk93cqgDM5IzI2+fygohMpB9c9nDa0U7kokJDUS1/
WvP/TAecLlZAbZ8pt4bzpAImJfsO6Y3zNDuLWwp0wvDHBavN4+WfnAZgPgEw3vA5
PW3cSx+3JwP2PH09mdCTQh0GtBvTqvYEf5ksZCZpsg94sfQQOmfFouNgHE+XwAKE
LkqcPH/9przX6Cvz9+/bE5QlTZOxT9fxrAY7eVBJUkvipjyM/fytMttDk90ep2o1
90WARix5m9p4fNKXh+v7BxG5uhj56D0zOwOs3KOCYGA056lgcroblM3elh0zFzfr
4xqpsX+k0rvQr3qqq4vn1zeF5XoaVIVV96b/rt985qRDM8medi0YMTxB4RlVvile
/ZpKxxqQ0cujl/1hJnmUT/eK8to8aTLAwmJi1XbgukoJ1e5Q6deWcM9p9MbEs96R
gSUz0JzC0MMmqj0aGAhUZKSHlpfzgggdg3cmvLilQZMrZ8WwkBDB3O8iRQmAYbP7
rYGm82LVutl4RykT0qrGehtGMaySaGKnL/f8bUbP4YVO8PndtDqs2HMGEfwdFli0
hfIg8hZAvoOjEUYtaXTkhiBP8k8dAoTmGDcb080mVMZQ9hbO+GkWNYVYX6eD618y
uau1+4K5gdlX8NEaGsnFjfQAkbS90md4x6T5JEgJkqL9s5qUZZuNUVyQ4/igbFVI
cFprxEC83AjjaUJVKqDT5CCkXLr3Whr8ymTDZS+auparDHgRvz2JEnHUdsnTgeNB
F3CXsKUZ1WywPzMjUx75h0ToMU+EihohN3ATmstlODhg7J0HJs1efTWa9P7suN+R
ltkxLelSytXpa+MmcmgWruCvs+dW5nLtgh/fOpHajQ5tC8uJ8QC29oLum6gEqvM9
np2byZOji02R9OZ/7c0xuItPT2v9vMopQ/LVKYRGfU3lRjaasDajH24IYCqQE9mB
WsSkZ8Yi2l1wgBH2WPeG94gx8vCyr5PEgj1XzGT+2fd5+/bYEYWRJH5Reu36lrU9
l4uQ+yx8bqFpwQUwmz5gsXYNFAkoFEs0ZFBVGYL4iBDDW3PzZcu0X4vyK9T2oXBB
K7880BbsZ+icYAkUuZRJipEOmboeOcm7WoOXjt9y6RX5moXB+DdY/aztVKJDwZ6F
vmyJYoZsIbOMm93VLqC/o+qTUwlr7sCovR3vv+6bksyJ6eGDpEOY1vJ05e5IqdiW
mS4lRsJ967J0C90UKhqnesphXTI30S5cWFjhzsqtWKGXBnVPHI5smJ3Q65IhLwz6
5rgZRAjq0dPCtGUnqk8fnjpRffXfd2/l8wB4GRFQJILaLYHjbUX6NrjJsOCs5KNu
W+HYQGjySogLIBYt5Jf0Znm00ZjcqH2If4uuBe+wGFYE4auG+9yT9+Gl6B/Q5/B6
P0D2OUaI4vB2Ch4k6H6G2IaUuQLSczn8aAGL6EDE0ShPz/Bw2d9pS2zFD8/u95D2
UQi8EtCHnzyni2BUGZ+AhN3wpgIBf2oTl08ZJ9CY0m4i/9EKtMwSENAawgK9ffVh
7N6WMIxy2NFpILYScHsLBUBqjOVpk1A+VqKebASW7F8SOPoXJY0rCCy8/mH6A1Q8
kKuLXNGAdFkYw52XqxK0H69+h8jSpYcObbjLgkRYRktbGd8gGJ8XZSHZiHqgexxy
Arh7NxTHaIFVnkQVwjroC/AE+Hkqv57zvxxiFa89Pz1E2+NqIpz6iYEk8HONo0xq
eyjwZUDMtxxnpJr3kkCa3jmigFgb+HaqBXsbH6yxkANSLM196ogMaEXtprKM4rUn
nsu9P8/pUlWqug7kBiNGCr16DDY5KkZnWZtQLUY/hG+x2LSypA2cO7pzl0FARGqZ
wSw6ly8fFhaVC3V8mmn1mGkUhu7W+Fu8ePdf7HENZBR+3Kdci7nrkLz5t/JNr20W
yLyl5Y8prix7tAUDXqCKrG/oP6UrQdW8oqFReyemsEZdTRVBDqhGAal7OT146IJC
LsR0dUWBRM1TI39rrWMqkKNVAwyvvwS4jwfccp4Kar1Ru68m0az6uMb7aUUWBWRG
zpx5aYfbq6+U+CD6M7jZlV6rpkYDyFa8vqlhZf7annYKXmceqvg4IG3wofFIrMUA
c/4f0hBf8hhZ6Jgx5/EHWx31FIRnYltvOOWy1XYHU1aTnrpJVl0jWpM/Uyezcare
rs8/N2HsPBWLdceFUu3128dSi59ePLEF6Zj4cMpSuUCT7GGKfeqcyiG/ytHHae6F
sZMtUDU9eCc/twqfNqMHrEnTM9mMciMU900er6KcGuELkukT6hKU4JlMl2XWbrKU
MKvCsIylSgOFSAQ5758ttRplYqm1RhDcV0VOovfg0sxD8zUl6JLcI24LAOHg634q
piur7+hYlyic1WgGt12rSo0n9zv9LXGkugJjm6qMsCrKaunEe7iHHc41IwxfgA+X
nvvh1YNvkjKMP040iuM534olVzl5mblf/MbOZeUfnxD9o0mbUSD6jYUCRS/qLvtr
kxhEWUK0VrcHFK0jqAvqKDwUPzQ7j3KjxXOkG+Dgd7iu9j2kcP4IN74q5143TZtk
1m5nnelsAzEww6YOEBGUVevkq6NmU/6qCv4308F3GsWXDDcBvHm5Xi3Khd9CjYYw
4d5ynHkMkFtuimwZPhvEIshmxHO4/ypTeex4UG/+3Z8ZKx9a95vCWECT2IOr6/Hc
EI9NcaF/wi3+L6IZ8EBG1I8fIsqsCiIAcD7SRZyBa9WhMSvX+jetI0zTbmQ/2cvA
MV22HScpfSnJm/plvdn9LsoAz/DTa2E0jtbPP9GEiESdKBNqZc/mwcakDwsBHwPa
ay1/nYvhfnUmC0Yc7dX9uWcL/ru/32OZeCwnt+IC0iH2Zs1XZYERjGBNeMmCLZ7X
TYNSUANUFUE/uCpqJ2B1Jja02uMaslRmxL4CcjAnMhQedBFLMFxEsF4OuAmYxgmz
tTOyVJI5fHUz/XamwGbLn4gmtZ9NEImj/TSAgRHcI7mVpxY50nJfESCqjVPkVwPG
WZpiV2aHR2Jl59cwYmlyzklcHJcpNZVqX9H9EpjzS5r6PyzBicidTqS3py4LOVzA
lCM0mVltB4C79FePnw46Q5epfuIJ8yf2YbZSvbxX9yxiLyKQwzLrNxIVs5MGJ8gr
KmCwYu3H3inYLLyz0xipr6GvAxfj6Bep3sL2bNTvuTMko9F3s+ekpsairP021811
fvx/ZGdFr/p13pcpasm51eq+aNGTsKMJPtZpzU0RmC+H2ESH/OeqMj7qxzWNq7/K
tZFMCTTAL3McR+nGSqodqJqj0Nrah2JpcCgP/S7qCOcPe8dX6LJN079wu+nLYvBH
gabyxzacFwvuSRxZ4E3VTtDJPVyIvuc/XhQHgiwXJYIfFMWsxfFmVJihWiuoLn3F
x+/Yb22NPWbaFhhmXTUp4Wnv0kS4IGF4lNqoHAiwsQMiMkmg0W5HONRlCS0esZ2O
7nk6ZCIaqiL/hfCUAcnYtULrlfCNa62VshfdlgYW+UtsUdZE6Ka+nU47FrVs2QQp
XV+cJzCBer3EIBw9bGhy+qRf+43BsPhI6uRwpbuntuRYsCjOT4xQzgeGH8R0v0fZ
2NvwpkvuSQDMCNY+AvNBFlG/gZaeCMyOcs6qZlAvzLDjOw+g1STaHlzTyaPIouuS
q/fhyoa88T3UlqtF1U+DnQAAWZoUKl73NIO/EN+RftFsVxt0lhGH6SNNqquggEKM
i+X7cM9L0uewhNMFW7+LBYuGmcYI9r/ORek7/Lhd+aXpNHk8z5rrk+RM1ZHGurbK
D0oMiQuz2Wgkc1VRIf3TRHVtkJ1KqkKrrMlimejt0QHOsqeHO75gkPom+YHueMf5
HJhZs29zczGcPOpN5yTiAz9DM4lu5c92tdYU8wAChmn3KdnVq08zoXBf83WZ4G3R
hWJhhJwhJ8Eq8wrqFiSRlkNzJv73tBwZxVA7FBqHjU0K+7molvJVKt4VQFmughKG
yLkUiTAjX2kC6vZHhbsnKM0j85bj63zVbubl606TO6OzQ3UZNBytEkTiiX7F3lSS
k/fzklU9k18Dj3FdGySm7/f3ARFLWOcn5ejXgheL3LNMM571zZTLApz/FExA30dt
jl2X++9Plc09dVZPhZ8RPRithdpuvT3BgvsWq2mF1gFF/7TSN2/fTe1PG5Z87pai
ok8BK25rgScf4CxNhMXlc1by85l6Cmu/RZYWvnT2Ip+6vKsCxefF2yHTacWcuSba
JDfXWqfunIgyOxBtpRrXs76z7IplyY7jEvMbVRUHta9lYqUZ/sFLFzFyBS/CPwsj
S1nQpjYlCqMIkW1YRj+9LYB8CDMvqXL5kKPRqPjsSrmY4IKu8HeHdHLdxrkK1pPH
+Lv1y/638IQttn9X5VhwtCduvDKuwn8qqhZtYKVYgNSyOb1UExDFr9ECT1G4POrC
LOAFUUdZMlXDor3KCo/UZXPwzCoJF7/E8geURvJA5530nJkOgfOTwt1RztJQHZz0
ThxlxowGGNu0+cOColjl28JYlbLs9AbThfC5tNfZ2bP617Gj/70KnLfTwOXOS/5k
7Eb4wFjAZ3U+I+Nh1JWwdN6l8eCFRLE94I+wSdLJlF3VGD2HARefHIy0RumExY/Q
nPbz3EJzNjy5KeIC5VsYc1tGwzK21XLOQmovvSD9arpvtOD+l4dnrDtT4b7bD6ic
DrOC4dQmesSH7vm+FuGUlLLATubjeW7beQVNRwZPEKbCYK8vVuSebqyFZJN41Qqu
Rr7a5Zzx8d1A03WWWpIKm7RCWY3CTCjCLFOLS/cQGJ7tYyHB80S78ElWoyifEDNw
nbvrXTyIxjm3cJBFyflPjtVro80nC/0cTphDhRU2GL1mt3g57tGR0AZdQvt6dkae
2BwRJbjDrmTPK9wjhrAmMC+J5OS/HcAXsX8cCfpk1MG8hFQnYEzHDckkJ36KM897
jWUNO1myMwvPkG5VflcoCqAoB3jq8d3yB4klzRSJY0ygJ7ltP8tRuuUAnXRaudH6
kSO/l3cHg8v7jXyMjS7XgeFj72iM6yrV5XH8CW/zZ0CVTZatBHJLj4Y83e4hoswo
pCuJUKmoufnbeDL1LPkXSRnFqsSmS264upWA6C9Kz0F/mCp6AGgzUwHzSie6jPHd
wPL1kItLzMlv4JGnRzx3sxV84d6f0H2T73MnmVFe4lkzwL/vxrvhaNDEyN8/q5Ig
BheHm8qfd01POeOf+bQsJGNSv2xBMqIiUIE11KqNh+OBak4N18Lxqy6hIqk7MM79
cCJdC3VIs3e1zJuOXLStF08IqsEgEnPl0jEKB1fE8Bew5wte51WpITuCWei7sdo4
bRKKEOIZVk/vdbM7cKujjFCz7DPF4+0pXWDRQZdmnTfKuOkasxHqs4kraipDhjFD
I3YML1jAIPNq/R3V3uZIkGHZCvQD2cuS4eerwl871ybS4FiyhBJeo8q6AwoTiNjw
sAkLpytLGiPGQ4YvuPkxb3xaLtVoH3B4R9ObxsXfSK8N8ip5NAdHPTZGCiwJhj4y
eeNSMh+lyVPeDnEoBfxtW8zmOe2PgMapcFXJNzS6r+6T4J167lGtXHBGSEM2n7vh
btmE8nmzGRf4HHKfdl5pCylYWG9r1cXOWcf0jitxy5ZYkDHr+k5rvmJwxOGTgH/4
9dXBh03FOmAZ9x+EKyQ/yxRroy1vBN6PNZDc9czbMUq8bo68qlYGiiHYBeQ0CThy
kBXqyaSJPuqIMzWHHvLuWvh0sIeW3ybX+eL9lFTlpBUs2JIXW4jETqx5grMGCveD
5KTuzM8DKNLYUQThDSOo9jr+D3znva8km4uSRJEKAXF+CXyk5jcCNbkmcMLDj0vA
8e1IleDTsxhVP/N7fcwqMXd3LL2nIOH5lmLnRuucmXHDlUdi7tGqJ/IrJ7XlBfch
eFJcTww/Yeqwz/Lr3Dx7bPxMii7xpJwRy5GbTkzxa9JSdf4M+qWxBx2SWmnwT8rm
zlF2kVVjhE/GAFcTZsRne3qL707xcUwo1Y8kKY6UnXjfR8LMcerNiU03vVlK+fER
V49NEikkrtj0sZmAjnqiqMMyE4HiXTQLAdvmkLkEWH6hKuddqort4h588Z2u2S9O
VBPF+Yh0NCczobupBwGegYkhypcmK+9vpRPyT6lB3JyIDvODOFA616Kp24l6YbN/
QsQc67A8HspEbTOXjTm5lL6viQFi6q2KIlxeT5I5kiW4DkSTV9vElV6px4of+gC7
moQN6weUiPovzJZRdGbDMLBEjHqEFe1VdnE6GQtcbAjtIgDna6BZ77V3W4NMxTvH
ou6AvQKu1vf9FZFow585DdCOIhvJFFtRUFId2M6OfFMQdmW54L9e+aPVTcMpCaqW
LW2dxZ0d1d+mp0V9FMP3NWQZ3yf85nuTNffuKMJ8ObHv2veUvkfb5pqgaboO7h4f
agdb9YsFCSgRyjQsjsk+5JUMhLRNY4Kg/4N52/6QZfFpWTFSKerda8vpRHjXLMXv
fmP2EOzvYL8GlOjX2JQ5Vvx9QRIWpwYMT/Leqw5yb7417pQYNgtj+78zMDdKubG+
yumou/DLeW6BIToR60vebRKNTUDWRHl13NOiwknKjSq4AKyMJJS4Zqfx3LbnM4nY
Azlclp+OHm1VxBl9+q0Ygwe6rd8K5VrH48CfUsH6qOv35AqsY+u//iyTTXy3Rz8L
2EGYaYBntksnFVNi8rYd9Xf4lH4zdWee70yG0kSJbREght8DBLtRKzeEPdudxitK
k86hhFCfQr2aTnEkxb4Pn+kbMkfMJrAm9WKF2ogqVEuJ4iHVwhmHg1DYOC8Ak1ZA
8+wPRbKX+m1DFC164WQ3/LpDL/QqIsITNYTGOHZZjS8q6ivWUIsa0Ku6lhDjj8wW
HjjKSbvcd3RxPHWiht2V7NCxvtgYVy3ZySdFRgMlpKXyz0qp8JcJx3Cktgy6PCpZ
KTnf5Hx+MlT0dXGfjcg6RQT7/KbiIwCEkFCer1PiFosDrI5h/sK9pHN9BnwlD/xs
CHjg1LTIQjavVJszq8P4LTlLCnAAtEGIT/3LlOCT6ln1ffQ/Qmh6FHN2XqWpGnlh
qtJD5mg6z6qpK8vF3wIls9pVjAb+ywnv5gm7gQiPZOkZ4zck2VBWNIICakszhuf6
nmnpd4FzkLEPHknX6RQPLeQ9aBmFO9vm4YGq2zIaIyUFyou6w86JMHdswxuV7PZ8
uybIVa70zilJpJou2o0PRykfQOkGdaNPf1E5XZcIV5CPn7hCG26qd4dLSUu8iBBs
alK3WsyGIJHt30qfcSwITMZk67s6ty6d517MmOLtNmYwv1JvZauGjm7tgRwNBSqW
QWaDyXniVWruUpyRPCOaeKqu2TXYlETGX5P5tx5Jc9EQjtt3IdpU7LS+E1IwUjWc
O7BICzBPVGCQL2agtlOeFLtXglCVBUOeEGkN1rtBA9M/nlHypUUfTF9v8ACcjMDn
DLy/A4wXzRNMisl11yAqABIAeUyneGz3kvYW0OMkrGRzrU8WzGfYngnCAUrGehyC
k+yqAk+g/D28D9KzLy+mTIF41j7vlJhSKOXAY6RhFDOueDQMgSRoCCh0Dmc+BgXY
ipA5rJEIW01SaFAf1Qx3zVnqiB/EYOG3ndJdYXugzlZT2yQ1B3byvhttc4Mnmcv5
aE/ZRkUIBn6W4a0TKCdUQIAeQu3+WySXzJHA/sw9Oz9eJmDhYcjdqpkJhNc3wvIY
zlxaYeCctMSWDFxt4zBxBuRbg/V4/CWWNFR/YfgmrX+Koik4tZ7M6uiwdpcWHFwp
T42+UTe4OsI5JZNmEStbpvAU2d7RZsBiwaITFuekvcS1oyTdDJInxrCG9SASPenV
EUv1jqcITWncCf74ksXbPXEymTCSyHp/ztFrSK3Y+etp0yMl+7BYWJxZytpgo8dv
myGEY4ZU98Wo8Yar/IrnmBIyNFhup4z0932B4/3BmQrH7MKGQYZB9pAV7rVgsDiw
SCrew+1UxRcb/rIcWAQ+LQYWm8l4SBX/7RwlFwvEXSl6nckg+t3O9GdxbRRPyPb3
sRIK2lnTfQ3uoWq7bx4nltBOIwCgS+QCII7mCM3Gr6vM1E4ZWI59fZS90vZE9D2u
5M6tatJHA9pc6yHy6F/a8ZTMiJIdBTCf+caZW1hb6nfCcX43XzGUaHvdWtSeTMVJ
u0kjyZ8OYsZregEqy/auu+PAUJq8mp9A1h0ohDUsppLpoWdHwCeVUr0RNSALBV8v
iXRcayAhYF1Uko1C+X3EoZ8nsxQPfK4+X71q0+exoR9EL6Zz3RKLppuEJJZzcLPW
isik+R5rDuIDnoCgdMoyBp/ju3vqlwIn2a//Zar7Lb3gnTIYKuEQN2DhD87uetdJ
5OQYnNJwC1YvdDRzar5yiFNUMuagtoec0gpFJUbTRU0jAFXKEGwJN8L1TogPNp70
MpAX29zlsDK7QZHotHBmgTPtNkM+vqd69WNH6O89TyCpD6fgmn4spG/sjpAW/Ugf
EETdIrLe4bKP9fTE9Q5Ll9SGMMI7TYb/4vY3LGxCL/Pqmr6l5TiWIUaKleQkK4fu
/yIfMO3ca2JBoxsyovch1QRbuFniSAwVQGpzljzACZq3gZKOsrjgsnxxipuTOiw4
gaoEWaz/izOGpj7MWIgsishzPDfscbmDK+8Z9zuL6bk2O6WqRhC1+Yp2L14b3oRw
HXUAf91cxE3FEvIhdCU0n61f+0o/ZZMggEN6two56x9Pl0cMyp4iR5SD+1As0Asd
i+t25+WyTJ7ZzuvW8SPHzyLUjsDnosorBwJTd9iKOpu1Ski5L4J9BuwHUHxMUiLq
XsLxv/StDpTCDubExtzvE5OWbX9wbidciE9aflY9TMw0F4QBhZabKaRRJ+hs+qpb
FDr9EZSUzU2cFhb8GA/pr3v/Xi6Kfjr6UgtP9oAYzl8fteUahCn1JZYNpJBxCWeH
kA+bNNWU2IlIjHryrcQsswmwzMiLUONxM2Grb7N6AQKrpIyvDfLH5qv6djMymF5M
CNJpfnwGSpj9OBzCweo7U9BAFOIrtyj+4ZhK+F2xzf88XnlRcspwV/D2qp4wjsMo
AtAOdgX5Nt8Dugn16mGoF4tS9XKIx2NZifN7IL3az14CwdgeE/3tiDtqoOZxTDgA
RNPMvwm0eY5cWLLM+Cx4vPTmOxb/x/ESB4UpnLh+2psLO6nQBr/ON3JKDqRzFVtH
bJ4Vy0Bknaz6rPf6X2XLPzUpis7mo9BwhQMJQOC/9S5myYEeV+loxz8tJf5oeeoK
IggVaCi1tOnORvrfgvB8WYzJ0dCQV6GznfG9OQwk9GOuhotE3IYkNwQ7zRoieQPc
EiT5cgS5OoitFTit2yBpPFpV1ZkM7RlWkvar6OBzroM4HO1cB2l/ub/1xYENv6at
AAomTdzunuIoCRsOZPV3gspkPvra47WvjH7nHbc3KeRuDQwnkVKbmNBn2cuKuKvd
zksE4cAQq2XXryPH3Ca8JGzTko3AH4iZ+0MhxS7lU01p16MqvkjbJj8n0HRw7Mp1
e9puZdUIOj/szIVo/zCyj2/SsCDCnKAxBAH0nYXVJymiV0HxlASmc9d2YVITQsJ0
dBWIat3n4KhzKsG+G9GdWgUz70+5wjFXYAx4bUJP+quk3Qa2EXYyYmOQJneLrgNv
uCgDYXgRuwErex8bD72kHrsfaUrQQ8bs0vKsldOX46i4jYUbR1063AzYbx6LMkDV
gQJIQrr4VLUqpwCjCVBbu+sp3fYDlfjNBujnhXOimUucCWtOYScZH/AL8QGE68xf
Z1MryA9JSLNdrOI01V3g4qFhlo4j6zBZGA2GH+Ng+AB0Vx/M9za3sDHKLTpeufnr
Mkrnix01Hqdz8dinqH2KxGk5CT9FYcFEyV7ZnaksSsfroGREbsMkIdMg0xn67mlV
1sn0AJIrc/L711JlT7yhpLim1YgmAbjJvklKNS4V274WEtgFIY5QFO5L4zzHs6jF
KcWp9w7nvrAK6y/kPmEZrX3uD+tHaF9MrCpjO/b7runjfCyo6BYY/hgDxzzzAG+9
ecEFGEakVDHhrEV+kpePA4CApSQ2IBkgJBAi4JT93ouqxMptuLLiXqk8equHxsjR
ozwIdxr0D8iQ4Cir/6I3SyF5Lni2dmdeTrK71ZVHmSiHozLUTL4BXjD5kQgk9uBp
TkujsH3sBNjaDG3CwMHBjqey4nKqo0JsCTqlqWrZuyf9sPK/Ou+lxjsFVdbwEJ/l
cN/77AwZK+LUziriRUPGNihQv+Adle5+Bx66bjbUorFFbWXeUz0z/S4pQPi1LMJu
BG9AlpLBVPMaZGzT8JzRPjS0llbl9ruxWskDkhbmc1s1fZrYbYiVr88RBmZxzTk5
Y3rlbD9jIgPt4Akf0DpUzLRRYvK4w2Uv6FUy2cE4pou0UO2cLkxRz18BZdWWII1B
uTTI4BdPSyhz+XxPedSyll3w9jl0AaW/DUWeePG51qkrM6X3zZ/ZqU/zLJTqqn0t
qH7eV3lmUIz02S7FB+OrEwoXuw5+hhiwlQRrN4k7JgvcpqqzX9hKlgpPIhmBzCP4
OifQO8j1xystJTbKDH9ASw77SMnGDQDwpsrAUFWpVdqKjuI33c46sLGBhLYoffqw
wYwHSlRCJq0jTx+KUQEErZPeY8YusxE+qBoWfFbXptlpwAPaVZN0ftul70K/ToBE
aQ8cckIZ0ybpPtQxrm70YUvK+QEKmIPVYQIMnmljjJqQh9DH8TSw8myhZPmPFAhf
K7i7TeyJWTni2D78NNhNkxAOvTkI1Wg9ryRIAwhsq2f++ZXC2YUv6gLJBFUqv7UX
tGD88L3ORO8uWSMaE2C4U7I40ITfQkCZJnSg6JJTla6gNkU81oVT4DoeTgsxHYiH
53tl4HVfYoQdWnD25odpKva8A8yr5uQ2QPiPIJTJc/kiSN6Kc0ZoLFCk0vqe1eIi
jQI2X59sOjguXYsSOftBt3z+XlS4B03HbqdWy+jpeuaAz7M/eDFzO5jq+BH7n/rf
cfYJqqoHd8yOgqI1Xo1kVCj9GDBFRNuMYVuR6c/040D1iiEki6riADxaqVkU+PAh
lhtxkr2sP45YivOUE/TR/rqcIqZmCtUCkoYjJ/WwkrTFIJUMay1jFsaPWcf8i68m
YvSgMcLwmBSOI9d69YE/ujH++9OPm+kXjmUmh287MlKbSgWAxk2JVGH1mrnfxHHL
yczPnda10VhpimVm1B2ZHjhM3kv18yTGfRGzWVwHKDXh9qOBZV0V5QAL609juMut
v0gBrSFFUbjeFqInGVeQoutAXKQSjJCNnt+pKGSl8M55mirqi/OhM09wsu9r22d7
VZa5/kMhxZjqu8wK8tH6KSUFB2b6ELeaJDQAhGWmAwm9Mpl1K0of9S8us0z3nqkp
Q0GA2yLKjjQc3DG2hV8SpRcPcfQQ1LmWimRKTJ3/8Z59EPOt61Gw5n29x2zPBPpk
WsbDKXEppU30hThBfBYWprQrQduzza1+FOh3FF38YtuxX9A++MsQEiaxz0lwLObb
VNNmMKaDOnctsQuUJgrgY/g01OzQR19ndKEoC3FZ329x8gF0rlzrZ2ufe+xNOOH4
NHlQHulFDqY7WzpU7sb8c3t6a5+VJhB6mdondWqpBEXFrRJxc9ehVMy4Y7LLu8tJ
a2kMi8VF7Dx7rJt/Fn+cHpcA3ffGnxydh74EquH3D+pagbAQbI/BARqgzVhriup9
YXWwE8LiM8nnuIrh9Ye9BlbhoDLIGNQEYa1FJQJ2VIyC04JV1d9ztrrHkSDt/RPs
AAqZ3Dz5LPdqcSBIjv7y2NNpjnPDshU6otY7JSLcU33v5UkSbDoHy83Zb0Ijw4dM
2Rhff3IwBza8C4Sc/VkqnnuwsiNcX7XUpQy5z2Tn1LxmYrb3oa6jDDMJdEyXFUKZ
NCwDonsgnuILE1GiO6o2mJvgCjRFKXZM35jN9TVq+5eUbv2AJK28TdVW8MAJYHIW
/Rrqa6A5uJMdRTok39+JRyaCPtwz7vpu0pEDBqBHfPiKzNCRsHdMosKTmy1uIT94
FLSI/chO9NPhiNvXCOQjRFt3HSB7mpyWr/Iv+vO9FLuDOuhxC9RZzx1sO7pW+Rv6
ghrIxGEH/sqHcWC1sUfWMZ+qZfL6L7xXWL1rUgGQrYHB0f/jL8MGKEroSajCJBul
Ye6YjpwFTFve5Hz2x4/Qn8DoHx7ignWbfrXf0zH4eoUAiqyyT6YYhkybQN+LhSlr
wtwYiHSMlozyZ2UIsTwaHz9QW+79BQmlt58TERK3VwpQIo64y9QwlwCWk1uKE2bN
Rit2E8UjSQhUqLn99BG5g+jptrW4EYwX+BAM48o8PgitWUkORKLSznSAwVPZ6jHN
GKzEXjV3giS7o85cuPOxDZ70A4OqqJbL93J2y4M2+7NMwoZ+U381dDO7x0RieltJ
xlr364kf9XamgAivX9dNyDzcR4WHM9US3eOr/kBK9oYZkTWixcl6xHJhX4qvBS0i
7gYHRtj3sgrKhc1ps9hcrOSW9jQEtpGrGHaBJDEDtD+NeP2RhZ5i5WP2PbSRNe59
5oqvyfSE510MMRJptoNkTGYKNSH9+2a1Dh5R5HSgNrOP8h/k3NnRfYBshvzoJQAE
gUMABbVmy9+nXGYvoQnENC0n/3tNvcGkvRghQOO+tFcDDuGSNCQnsZqTSwIkfTMV
Eqf6AVgih6Cu6gJBnWb3HH4EDOpBPUmTGUXY6jNx5cX+HeM5cM8TQIaFf87NiIyT
R4Akr+mcvD7n6BhgZFZ4ZZt3FIDpH/8H92fKo5wASgeQQ+EiAh7XBzEHVfR5q3Z4
41gd1eoJZH+B4sCOGBpXL4ZV51uzG1D/vnUZLYFhQee14EqyMBQKi6v/m2J2HhhW
S26V1XIY9DlHPDyMWPZ/F6VCgyCx0JyVO/E3Iqpg9E1QvLqzh2RcWRdWdMRz/xux
xOYcfa6t7XqbsWwPB/F+ynKNvglHc5kyufBW//sFqryL3AAfUxofIEUXcRA53Rw3
Z4bydrcSIa4Vv0NmjXDT2Y9PMBjwgquQ38DZqKKowcAbpsd/cjg+nibg4bv/3UQZ
6cGYLQaE1uQDlT5m/DMAcuLditbF55ZLnMdmcBrBen1X4L6nEhUXi7vydDnrldlw
OwB1YZ1xNBbYQ3KZZELtrOdgkY0yY9edKSLiXJfd1NodM+EPqS42orueU6rhn1PT
Z9ggQ846FAYVyEt2luxBYSFocxdMrvd6O/iMJZ/TyANjtgfpOU3tk24rbR52C9kD
08D9VevR9HkURdzkwPY30CjRawuK9Pif4/AljrOnlhoNzjxmvhxt3i/Zd0vtoVYt
+E+fSF5Q01cbRpVZnVWIvGXzwlq7VJjzMxOMxEOQ9R9PxM+6fmBxP+ESNQUnIUdr
xYoVYZDO91HGW+/9Iyjb6U63yw/OtRCHvkKRGvrB2zqr36IT5Jq2Zo3vr3JTE2KF
Ycm32f76RCAXY6iXeJTcQ4mmTzpy0hN5/A+dQ0Lq/N3yy9eIZk6wAGmg5rG4Pnd8
R4uAfs557HPqGkg8HR9c+d37vxNmyZUH3EDAywoOV6bZfQdlr1E4DXUFcPL1uNvD
BzYH05G41P+l1PsdBmhuW/hM2mtotLz5nOLhGW52ybt7M0f8w34g7kktT2Eyuya1
Vtd3aXpqbcSxkryZtvffk5UXqrCz0bjSGt48o9rLrJ7ExMFwROxSbE8l3fFCb+uh
UdX1duXJeS8i+tF7xnyy89f7zEe6pVR2xhjTBd++QfXZKIcu4/yuiQ31/u32FAg0
HdfjU+8XvM/FMavsYlea0LBTUl/Wt0UuQvzPBoyCJo5b/8ASnJONvxjN+eg2vgWL
Ooo9l/IGpYH30qOM0BSLNtrv/cgJLYDQ0Bsp/bw5E3ovzm8eNNu1I5PISHSu1YtP
eQ4cQCTAljK0qwjm+3gA0K436a5Ak4dG7wHMCR80Hauc9PDvTJxTDbZiEPIScOqT
uah2I5tuLXMVCTdttc+BHL0tbfgJjsKqiDuY7Y1kx24czt8TPlXHaX6oEjfgE84d
f0OxrqIfb9KsAYr9oS8/5nFu1v9gQhYwJOkwILujYdWagK0s4PL2SYtTJDDizmpe
Cvh48cLOCoYqhtN7pY2M7yUaoWBITzWHVYqmtqxK/wAHXPt/lvIISoEhQA6F632V
Wwc41GlkEZHMAQD09qyvyh/l1Fqp8W9kBryXn+tLpxAweOF5XbwIHgVSe8u8FF/u
IkPDc8C2nyjzjPu60IeuuH5wixriM/EYj2jAInNqqoRiPP7tNGfHFKtQ9RdmQn09
vB0IL4jkLnIjyRgXzJr8vQmqvFV+iNasxL3WTRygr2IS+0g6/Ndfff/RPFm+FnCv
5KbLFo51OWa8HjXn5WftqrQj0+RPdUJwI8M0yH+mKSvxbHYvXrrKqSGY/+Nr5e56
YOD4eL9/Yjehg+11Z0hqm9rD98N3OyD0vqL/dVEUPWgKSfcDfCHlaWecNG74YEFc
KFf7PpHja/IiFa0AptkAJrJbj39uakPbPDaiRxhbfS0So9ZyuPcLhhpCXSQTDk8R
LfxnY3EMgj8HB+jo9vkURtMAG7PlbRK2kBdrEp5VICpK4BomtoOSdtNe3xsq9+00
uIJS69p247NyqDN/ckeUcZQpCVHuNRP6H6CJ5FXlj/nXhAtoqtgVGDoLo70AN6DA
Siwe2Hag17tCYc0znwoeJWUC9GduYu+72gYZNrtDOqNdlvWgT2qaOYlJAHntlPaL
8wHbDOSG64Ocm9pPIe2TWw56LtsZBo+wZwFsGT+p8uXZoAc/pTdenujwXw38W04S
0VqRKGPZeBKo/B80epXjWBVSXlRmwwqUqQhBWOETebfza7HLTFurI5wo2U/8Gipe
/p8/AgWvGXJ3EI+wg7RCdf8lN6PxtA+/L1Tz2V3jQmWp+j9tTCMMqbTe1kbJYPxv
ujecsUoS8JYOt8UrLJoWblStDsB49Xn4GsM43qGNeVV0EVArX9OyArbYLscRKsUa
BLpKi1pJMZUVBPxCsdFrPgjvIfTVcygr13uNpJD4WL7jXuQNc6Y3l+qs1ucE+rs7
h3Wn7qOKTZ4ug35K1Zi9U41QM/xH/0TZUrHhTIIIrEvKp+BIupNKwrueHgTUF2C4
KL12LHbiSTFs6kUVs9DPOwpVoJiwF6183R4tr9KmeQ7PBtEqLVcRK9AviVG6tuOk
a1J+QGeCIHYASiSDKTbRaHWkBLCTG6wl2pzrMvB/HP03D0wX3bWBPaly0DI641QS
ElfTMly7m08vqdWmUycDyV8VLqrHUJlQTMWZDdU1vOZ3auT7FmW7jWljzscM8xNR
tZ2MW3ARJFOJlaCDvgza9W7oUlkrXR9SckmrxtWf0Yr+dNvx4Nc7WJHXDFf7NoOb
8aPNHEPls9bVaZcCzuvHmOznehyXzcxa0xgn/TvAOiO5++ZunQLR38vmigfY8j8E
oayh0lRpbf020I78VBEtEbDyK8ABmlnLZoVkiORBRB0osLJ0IJKHeGdWMierLhws
6KRfsfrfNRib8+r7im+b3cy+IL8hsrjtq47sJ0sr7AToAkIe6Mjci/IqZ3ylPp7a
77GejbylgR29763vxeUUGjpxy2Kh1nCO6xOaPSakLA4JIKQGj7dsawRqpUoL5HE9
WkHpz1xP7In+pDfjV43KLxWGOCZw2/6S6Kz0ZmP5SrvVl+kKbsors+ZZ8yWpT7RW
SnRIgRWz0460a52nMti8C81Ps06ThpK8xgWkDfTnh/UYnYLEczzqufItG+T1yUaG
m+9R79tmWX0kasSidu9HaCQe2dySXI1IkvQa6+WS1LE8voR746OWMPVAQ0Mci7Ag
CWNVFAXIhhsaTlla2MgCQeEM1jBO5wZ5en+cEqZSxZQWaTWe/SHNuvApz6cGw5Zj
BkKEAOzpXsbPQuiGqAN4gQLL0lpV/D3Ch5obwwPSEfEximjOXHXV9xMJMsT0q1Wf
SHqtFipwHqAIuCS8XuObANqoJIZ0oPqMYaWI/xnYEkEIePZOH5bWmyM6JNfLEBQ5
h3yBjnODt2uNGzIPfbsMQl/L2aMGJtCMm4akHyZksPvWVdMrv122SyrEYz4ep8Re
emFr6PYcxzkSpt+HlXk9Hwot/ysUkR7fT7GTzaU9/QilN9K5qX5EzxZpeLGTqbHZ
8OJS3jSKWaSfmh/Bp9/lsKdgCXSYXDTwmmOpDqMfs3yUD6BEuhIyezKBl9mSiQzv
8njSdRZuKsSgDLligCvuve3OprO3LvW4VaHpIEPQ5TkO7ilGC4TiZTVrA8F9z+Ba
4J4SJ52ofbo6cWhCmapgZVgOsmL0D4SQUg3RRpCD8Brne19swA5DN9+o8lWUe+pu
qaZULDjCKvS/XOB7b7Ysn3A4V7cF2H+WGSVWcBczGpTZcUG8d6CRNchHSTp7Wp7N
gW5jXiYyS0irJnVp6fF0/r8VdwmFDp/Gs+jgiKSQct6Bd4xJ2NVhmmO+M68heTxf
WcGlT0nPBk2h8rjkL7Ln6Y14imheuoYH/tdTt+tR2UJdtLFuu38KNyf4xJVh29HX
i2SGPaesQtSpe//39pNJXbAtwkK3tUFIkoT8f49PRhGZIAUWAd8d5wzipUIQHE1A
AN29yPFsuF+f/PDeW8CuF0ZE3boUHf+a6Qz3O5TZk3gyYsOSxDEQJAuwxKlySfNX
kw8pvtxcWBEjUe0FMSVVw4ScJvrNCcJpmoAPw2qbOQHpWAQkmeLUq/oDqAicMHMS
+gsWqul73wbALYWvnPGGcFa367qlFfqGTNZGPuwhx95ACMc+EzGw6NjTq17Az+TF
bLYfJiV6ATrbV0js/KQHN9eSb/hVbFgXIlILVUTbarEM3MSgtqp562p7nPaNVMzw
+ZeedaAr07NnjPuIUK6XYu4kYaWs97v90eWmdi5fQOvQc82llBM3um2o/CLT5Z7/
cOguak3t5W5RPNm7X/jJZ/xff+3GrpZJsS5DlRju2A3MIgBBQ8viV/J97k5Ag9W/
eORyDnhZRYSqyXstQ25BHqp2RXKLcB2WBLPRkig6R9DlbqetnOtjJnbU5hWvXqzd
JOI2XSRpxM7tDpvLH1s928nZ5KqTlNybCTLJv2uOnoff4Lg0+PKBYuJet4vKZMn7
Q4I/5CkPlgCQKSv6p35PXn3wbrLGYAheeVEQfxKF2Tqqy3PgccpXxfuja+9dO+xI
U/t4Rom+r/rpvqs8ViCfjiXMbP+6Kk/n0+OktSOoWzinsfUI28nfsS3fO27RNZ+6
M6svu08oQKymoGkaRczRyu0kxfAPR38s3irU9IrBRAz0bhfel4rjsfTIOio6IVK5
4KmGpQftzqIteFvgy1IjhTXPW0PLPcZQvf2G1fX84lHSqEB5bDL31rf2UyvUfUJs
AZMkdqzpZi8r1XdxwUfEcU54gP0F/l5ju8hTqvcouv/UZAbqVlCaHSBbD2kIchQr
Mrv0G/YH2+oMxsTCpW3kdZ4hrPOHWXt6cCJLJjV1Dqojx5LF02AesTmFsZrSPv4L
/g7ks9HF0Ocn6EW9tgbZw1FlSNODmpdeiB7Rr52CKjem3sO0cBFJ00p5MJahUInO
vE+oLkrI3w5UMJOjQS6J6tU1U9to27sEo5/OlH8063WUJXtUCNPDfJIlmESLm0KZ
GsmTIpnqC0y5SW2EWp6F2+EHXI9sUaApbaNY1xC68pNfBH5ktFDZBWcIUwjQDHJe
6pJrNcvn3dzzkGo3+szl0dEtMdFIfNtXcLGF0u1OAvOPL7dxfjkq47H6AMgiYEeR
cU966DXRsotzWB6ksLJgCZI2VL0SqfOt9dl6N8csDTG9woiGVOeHSe9gvGDgQrXD
/V/vRiavDSFVhdhX7zL7DFuhdNAuvQEq914FdPUjcca4ML41fYYZLOCMuwINnGi4
/C2MBKrJ4sc5sPrlaSFIySVAOSIAvyDKrPpPI2FRu5eAo1eytz/HrXtWgnVbr0ex
X9OpJBTAAcJvU+jNH8zq6G/hFmtd9ABSbceyM2JSRBXqOoBpkjcnKUWdUHyOl1fF
6729u9w6vbMKSI1YJURoYpMcvWDNGCR25o1lBEDjJApsVYHCMOhPXc9k0PuniAHx
zLdyvG1qNtCmnKyqkfbx9whglNFCXO0BeY0yweVaHHxnx5VSKR4qRpl5uAdmg0lW
t++9rnu6yMtwZ6wtu4H0qzVSS7WQsBMmDG+C2HbFliW3ApwgIMq2xEsGLeUmwfHu
yXb/JMg9dX4dX5iogK4cu+Iks76igppRyVzMQSaRrmRh4N24+VgsiCIux6TpKKGP
G5sxVZLwdIDwTn1fgG2AO5wL/1xwzxmt37c5CiVd0L4OHsZCTur8H0TJ19mKQm+G
d9udvZRl/e9HQya0ciTPHojG8fu/mJ2avArUvNzDc1edYj9Vv14hwo/Q2TPoo4/D
Hb6aHO+ULCFkA3HL6HhQb/tfmq0hN3dilU0UME+Sm/rDJZt+VYGTIbrSz/hjjR+V
P819gwsZqtzMGH3sKdlozJgd7lynU9XFoFegDnYFBfrQlkFz6EugWeUYFAUiLYCX
qaWgIuRykAe4pS9ERrMHo1nyD4HcR3HMb+JPjI94Y1TSOW+gwj1bmNqAm38SJ1sR
2SndX2ujTBvc18vkfvah4o/wqSTBt85tI42v0c5kIoBlgkNwv64iuhV8NjuYolMu
Da+ZvnF2czG5SMct0LfsuMyPcTKnB+ETtTZf1HtAVziMntuCCmw1fSijqNxqhQWP
TUGY2JXqaTzGZjaBt9W2wyhaJRMb/EcONFRD6qtGaaM8jmP3dCs1mpNLViRwYs+V
u5+dr13rq8xhtGlKQaedZNHESdCMv1A44npkluGzGi5Vn1TQfIna9rBRyOX0qSL7
gT3CaxucbCnDAW3nNR68VBRPQ731ZCV3aTtfbEpRF5oP7RlUcDF29NO2OaOI9P+K
s7ARxSLcdj0TxjtCqWrzzxjrKHSd9AhQ7yXOxMKNBWl4ybykCMtNjDkuRnzj4G5f
II0BEtkgKv0Lt5vfT0WPC1oyqyVBToOe8bD1ZWTeP4hJYMs8FAHdOw0ELgx1vOx7
Ojx09TidNl7ges3fIZPLYvUL3/DOYUWuDKXI09Ugc3zsL5/GvIb/iTsfTIaZbM+w
kRPTSxSqx+QsAo9qr1wySOgVtpwIjm3yB+khborQnuv2CDRm0JOywUYEi/Q5a7Yo
h3nSYtr4CaBL1D0rqZyvbm0NHe90GRr5L5BgRsisvmVfDugDDob9TX/dduihMcl9
A2QWsDjXuZgp3teTT4RnR+O0ze77YQ7fqV5LbtWviqMAMKHQmqxLDzlPzVdNGAu5
doGy8nFMfZvYJzm5gk+tIh+fmib9HQrHko3fo5w7OQIN+f4/VX6b+E2ojiQWHL2d
NYQXFOcmGhsjbRi6xwNiryjy936fhbXOnusbXUaxAKcPFAD7djw44TZtG/LmH223
KEU32FcbQiBYYErhSxW1ynyyPnuqGqRRQsW0nBL2P8k3cjKyVqi96zwHwqUip7c/
FBLB77lly60EmmoipoqDRTo4gPkRtxVXvKgpQDz3t1NeOK0s5oaz5/V3mKvRS+G6
XfrUdL+5/Xa7kQrwrFwYo0kex+eusS1az2CGWmD0096SQsd2j8pF6PbNdY6q2ezl
gq4cRYdrOVt49pR741QzUUGIgzmzL7LTNhg54S66edDM3/bAXafAsm9gf9EEKEjf
TjLeAp7znn6yR+ugi2djQ/Z1aICf/86n3Of9Mod4W97owyFsTF43s93eD8+2kqEe
11IGKVZU2NOypguL46kqIOlhR3SbKv4+OlapUvvK0CFnlDlyFeEO6Ia6N6zijyW/
6VzW5agOUdP7zly6ZyxoQ49CMXEWLKm/qkCeRhWwuztdG7SoNpOt0JTE1mgGF51T
LUPhf2HPCn4Wralhx/QKD0JbcD0gNKcTi4o1gnaeBXZYFQHI1RY7NqnbrslkaJVT
TkZW0EIbpWv7TUAdieEEIRn8nsjrkb3KrKtYVmh5H8oBjjelxRi7QB0rZar4gtnk
qvHnC85bEzCi4kmucKzXy403xMnGus2dEg8K/dwwgU3A4BFrO85c95BRhiUrILKG
Yhif+vnECSiiPjUGcYHYjE/IZDKnWGwaMMs7ah/sxJfxhYfb5+3Q0b33oSNGJd5k
i41Zl1/ZUZ0ZFj2DYioqbeNMXrSg/m8pJy/TYOzoIrapjJ5ZEplBsBnLfiS4zthh
vbGR8X8MMaefGXHJlra+3lLMOS4lOIHcB4HtomFNXJTt53j5LAUMvrYuhZjJ6seK
wXJMQuyuqT8WQ8Tg8aOwPfdDMVpuRzS//6t9J0QVIJxhLHYu8Fw1pWetUAO94hzw
J9SCCXTrv5b2wLYKI3p1TmKLyNfLIzNkoAhY4KjGLRzSzHW9t8bdWGW9GcxpJA2q
S5LkgBvcGNX4rmA4jW++TEGEzCSYShK5Bz3wjCiYrf2Gq0nYvubNJFJ0zRN392k+
Ht2B43c1tDkpoU6lZu3K4jrjpy5xgghjDVx9xwELXTeFl2wgAtY5NrxiOtCIo7WC
MjMet9x2Dwp5xJTbzsEFuRHccsBsRY+6qKX61r5uDZqUkgefCGE/BFyCMEl59h8D
6T3XsJkgHbcJ9Tgnc4YD9i1Xtf+Ld+F2uZ0IAHRVbBwG8M1LosDWGCg/phrhioTb
TWIr1j9yToX5zvoqCb6yPw6EuowVFkGLdrwoNiovtXfTlBYOpIfq+V9+uWzxRNLI
+MS9SdW8DEyo7zBmllz0P+popNfxoOnMPrJa6u080X7v/XX1luoDULAFdtEAAMA+
Lbh+bQXXhI/s9pT5lmz82w9m7i4btWLYp0rwO1FyHUypDZVz0IcDou50GJQVbEG4
DwePr+2YUg1nTqIxbK+zP3o8UyPB8+5/grH4pYXp6T9FMQaFUgFa7QS7B69srmBP
zZv6/K/By0JF0l59IoVSdkcN/FvAXoBKiqNsA/Brn8fCsH7bvVY0wLwiLWYwgeDm
A2nLGO1pxOYN2Fj6d6kuGjGQyK6zfI7QgmzOVOdltzfHjxVZB8ViT612yL13C1PM
p3OSgnePiTXDqdiy9DHE7C9sM+3ejXHTeyMRqoVuaSwnRroRKEduJxb6YSjRTeHV
Cr1raudzVnM2LuC5+j/JFxAoO3ciYpjkwwstVCpbEb9pIRqL1eqQVjam0IxiIi/h
mle7Zctz0Rb8IeeMpAYxbqpUaoTkttjCQEOnJQHCIbIOmuBzaO4bptz7vy3/PHlL
JwlBTCRSRebpB8HveO4Z6eUn8t2iyRVdmc2VmJpPy8E4MKUo4I4uFjMja+xfyEV5
8d+257qM7w0/5eKPYNqW3IO/LEqD2d56a7FOPWxr6uDszFX6qDaeLsCBC4hJVFF0
94Ngma0ywiNwGqeqWKVD49gL3x2BIJrZl5/EYQnfNQL3CwcP7bnZxYzDWR7gT49r
5S38YonA/2jEBr3Va4VosiIgfUlw/R/jNwctF81qMmOdj5bumd+6trQQV7D314KA
ELW8sQ9X670tdbW2Q6VpFEp2WE6PO0MnFZ6tGeUi8abvfboGTK+ZBs/oWhJh2P/S
CpK8N1OpYfa3/kvb652f6hknJUuji9FPiuZTfYrcgbeG6jx32ACV5jL2uIv3pr8o
0feaD6DcMoTm2wdUOJNk6nBBD/Dk970YTT4U0C/n0oAB0NjANznnaEIJ2eOEE/Pp
Ienu7bmF1oueewUt+pvcNL/0cSvJy5kOls+iQ/BjwZlbJonEFCQH6lFj8RAFu3vQ
b3lwXpQX+G55eMsf22DzNLIehixKHDdIv1wcYyCLzbL6Pfponfyyn7SWtbv0WuHT
SY5oaGTksu3tDy7gqMbkWAogVCB+1TJaSgQdt19lTI1d44cINAsIi/qP1WEdHqDv
kv6Ahs12BFOB965PkXL/2QjS/b7TWm361MJzu9cXqzOOKowBwi1gPJABhsonQUFn
wzeHjvLKnJd8Nutyfa6scTCF4qReJBTo46JQgvTqSlEk3mP6A8MGk6yC/cGOdOp2
TD1gZzx1tv0XmNgo6fg5Ma0XHOQtdre++u4e9pOldsOXFyuwjMWr4WEb7Pvqz/sF
voB4I0WbTP/BzoBnpE66wY51J2IIiptpuLV/GdgZF4JDxCG6yLakC51CcCURcB8Q
BNfXxfgDAbtpgKPMIUo1oAEqmdtkUAWsESCFW2HafCjxzVLZaHOGn8SmJhtiDE4j
HrkF38OkMLQNHSr5SRb0QS0GHmrgbKG3apZCVe3lypmJyoMSc2kEw4y2YGcpHaQK
/U2FzZl9W7JaX3Em9t52KASAkOxbRgD17fsKsBwnkdRc7hlEYFVs7S/QNh6Q00GH
wDRnBUhdhAVuZQ1ohCVGeWKKRYzZoLts/0UK9eGaJDzKxhiJYFQYVHI3VmkGhNKb
a0iqAIlUeWh5wEIi3qVkAMfAFSpm2Xag5nKNOnKSY30JeepvOOzWGyv4pe0e1Rul
xOjes2hOYJuB1z/u1ZGyBSJRNiaxAp/JElHen4F4KvMLVDKAJV66+yMZCCB07psM
0p5tIrmYct10+hFoqkh9YzidtJ+OsTAUx/X6Lq2APmVeL3jFC63fNZRcHbKUtvYM
A4HA0QV1MoAv3evmY1QBRmqbPMr+vyEgOD9MvICg7ri0lLsx+5PhAWQs7I9La2s5
yDlXoSM8rXIx3dsD4Equn3emhMgl/W0InYkew8V3xMc4+kMLpd7QKZ1jB69O/XZt
rcs6owy86yKZ+2SnHZcWKsaz/txmFFMUmAb/ArndBFc7Az3ShC0+ZrlNAMRHMba5
bNuOdzrbvScjRM1PoEd7kOMpXLXtXSQH4jqt5JjsqO3Z9OxPkv3Zw8bkTtbmXTAX
Q9Bp+4dBLLPletRsL6V+h5oxtXEkOJmRAsxd+ApJqgXzHYz0UkfABQOVsBQ1hpAb
KQYb7Ubi0lM1yMtvJFoTmI28prHAUnXehA/gMDJq8Kk3V+s4P8ocPuXR3gmq2ugB
Cv4CsDoYIT974pOBFirWyGqo29yw6wfrbKeZ6JUKhsabWkc77nHvf70nEnLK9hGw
O/pwE1CY1ZZLGAlGo72U7i2HbRXJDt5X96Qi7TD+x1heuud0tFj8niDphp7J8Bzn
Z5XiuDTDIteshjoXXtxtgi04jpJymcH2Z0SBJWDAjMpPNvmDDseMHQe6Wp9LoUev
iZCnrR6zOZaYWVI4BcCh88tYEPtkMaLxdimFl2gXu4YyDxaOTiHqseFBB+1quwyf
+SrrOL7Ehvt4C4WMGWz0bcI6nB8NdoegmCGjWRokKmArGxjfz5DvlXjcywckdc+K
omNpI2rx8fzB/g2zrPnkbqBcjxTDvHuiE7+GtDWBzNxPUqQT7hoPpgpqVhYGFZrj
GG1Mh9XqWuvzj6fMjvL//GWJNNaJejxdSOXcNpnaYPUeHjgS5lQYWAto6Le2KFSA
m3fToHcEuFw7/0ga7I2B+1ooICNq0CU828Qfp2OCc635aK41LKde+388dlEUmB9V
J/IQgqK9l2St7MLpYid/X3mNaQrRdWYGgBzgeTZoCSf2LQvysLSKWuBQG5kaGYx2
iM15DRDGp7cp4SqrEMutP1tWOTTFi6qOK+fpXBMeT9jI91HZKkRMD6IYATyNM7aS
FOzpwSD2ltQhlusrsmfkgQEy+zrlTWFPUB77Oqr5HAcZK/8TtACRdp+N9WdjR/fa
Tgi3iVwimsyyuxEDiTGl1vkKW/9JaTDE4Mj+jinYllC26XB1SBWPmkmRw4eUFlXF
MezPpADEgy8L18PLpBKjfSYs16aQiI5SEA0yBvrEn9qVfM1oFfF9Y2dIrs4NcElI
C7RMTb8Eyp9N9ZfU+BdHcipiPiezHDSbzGEIk4J+KBEdUw0Jafo+hvuXMpRIc1XG
yIDNOWEkS2NXF2qFQ2sLg70AKv21DP0U4X4Nc+eVDR4kB2WP4Px3zyGWHJbkgHBR
qptXt5GxbtbJ4rkWVaie+42FHDV//LRFS5ofW6Up3VHvLrJLMRFSenXiqyW962a6
0IA3RvToVIzqVXj12x4I8IOkGuCeME6rdrExgF9YvJQGg9OYwNC/1KybBiEePJTc
CmHDBCPi68bLCcsKUkchVjIKS2jRITC2xef1wL9LvHJmR5Of18UoGAuBAw2ZvMJG
x6N5kVeG4IR+eq8y7DYv0l3sFSybo4ktzzSQj+wYVmVS366Jkb0pjBlJP8hIMGPc
qZ2UDzVidLHP9Om0DzLHPYiXmC72dn0QaxzpNN+9xZrPcljMghmWWXJoXfuUo/ok
ui5rYGAE7kvxWm1W9qmPu7cBsVkcBZG5EgmfRKR/c7Jjx3owkGGlB7AeCvGmK5Zw
wZJ7P2Bd/dpI2ruGix5w/ej93IWqVhyxK5oMK33aoO4luKmOwGEhVGE2PsZsM0Xu
5TjTopkUXoSp8MKdgigaZAsMl3uwfgQBPX2T01ktq4dOCTaQwQWFT2Dj005e9ZAw
XNSxRfR1Ww53ECOyofRbXS35mfycVAM0GeiAvf7ttQsiOR4NIrcIi2ApBWCBUTLA
9gq6/4z/3yhJWo3HVu6UlmRujMslGVQOyC8MIoe1uWjXTDVXA19FcxTuYlr/e2ad
It235yAPdnX9TLpHD22+7mwbTVq7B/xVvo0FrrRloSBFukjaMjItOAW2SoYcZgIO
9v2aSmdEZm6bf2b58J3Ht0XrEmR1rYvfdMGq6/szm3noqF/oLkKYXCQfqDFujw1J
I3SSmX80Cc94sJHQz8eziCC0G8AenMClSLDRWWyFTeNGkqwybJYBXh461U8UWfSJ
eE0uI2xU5V4aPD81XfdMmyxd4OkVVRdN6aifreAWqRnwdaNR+ofcOomSBVC74NZe
Um7uMhN4Lf0lIccoCy8MFmrwgwHrcGeTGL9J7muM4P7OqCwV/tjMWaLYyTuZYchS
nfC3jHBJU3J+30q/rZQUfqVyYI9NrYHcMn0ucZRrP6eIhKQo1FmEvndtTGOyiqmL
Mxs3oVFyHHV2fxgUw2Bnt9R6esVyHf12i5dkLksYBB3ywyKO4WTwnKkrXgM6zTC3
jZaevAYmC/3BYRl1vvOn5mVUD3+Hph9vyUHKXh15RizYkiXH5PBOXNPXcu6xH+fD
CPBW3dch5XC0MuCxOid6fXFTCFNVTtE0V79g2X3fK0N0LNI6xpuvJu2DapB/f8G5
0fyj32kmJUmmH/bZu7L1gwtJW/ydbnESReQRFNeImydYVhZqQ50kiqRnbAQT+gK4
fefwWSQJuBu5ZrUl9rrvrUJjJJvr/uCkJFRYnHehkD0DdqKGSMtjGylW/fZvtV0y
1ZGbAKAHGaS391LtBIgIn1E5vmJsuAwUuyiLRRvkpOHRTNHXUyGfp1nue8NWe/W+
rBX3mUye76TC2z4m68ZW8IpVMnG1HqI9lpPS2X11ekXa0xqG+AX+by+XZA4NU4DJ
sMz6/G8qI+EtFQb8Bz3U4tmPDvFBdzqVP8K9BSHRkhIIXhfzFESWz0NWjWKVjiyF
NaPeSMq9RWXMQv2y974CgauZK8yh5mPpc79s52aN6teZ1ls0BtV353X/YHEtD1vY
5feekWkuq9AYzqmZHGW+ZXRo4wuEqlGYJpfMevXah0X0u0CJIQcYfoVMpkibndko
iGcqLpl4/M5JdtL76x4r0JN2clgfIPzJi+arJWnpHS34SHqzWZJPsDB0hLS4jE/L
w9KpdnLSbG9QCFcabOCIg1OXwVpFMIymo6K96pj5dMLZ8z8e+Q4/YndixabvSiur
8Kqnu9/2/9GpnG24tna5Bt8TF4e8ypON4uBIrnPBBT4e8YqlVDjx6CLRBbUBkZtz
t588VJmUlO7IJl7YiP5LkLJkrctrm2UyJxgkvxxNNQDNNhHY6XmIKjpOHuXXhT/v
MQD/kXv3if4HwD3SDJ+pTAL08n2rikTUMuFS4/yExLEzizT+rgIhP4xV91Zj+VLZ
v4EjfnV4nOX2qEwaA3aRCzrRbGeht2Uyeoy/02NfIpyiAi309okfjwxgVGFUwMO6
srMR1qYvpeqfyKSluW0LVu0FFZvybLxfc1pWQpj6ese1gb2qPnC6JKvjg6fW2Lp6
TXUsRqW6uwWk3R/IVypKobwYiJ8x0Fe+4E7r/hxPUm2kZUkYtj4tbEZy5giieO1R
F4mTewuAix1m4A85us8WFibnwSYjCE0xbxD+DsuIVACKVPxyBqYUFhu+KFx1TVhN
yBAy7rbUnzyJnnouWVLnQaQfM7pJEd15ZJClPl9GbVlyuomfGKTusQtwoYYaOoIb
qC+s6OTu7Iv9BIafECeOFuPQEiCNw+YhR/q3yARDTGaUvfUqrsI9cvXQXrxbGhnm
tpK6OLFYveykm+cOqKp15PuzhxLccePPv3yr+nlNa+teif8ZMtqCqy5GQL2DUrvZ
UCWHM90wX1l71d4fSFPMRY6hh6nJfAt2gbpM8ci+bgbQBzjZkAQMIVzqpvXdKWcf
6PMZ6mkTUoh0CrBjLu2ST71d9wYpOrr/O9UzDRERUxGvEIMfmfigk+IYs6+k31Xy
PV4fYginI9oK26/bxSHF+pWKXGzqLLbCiOEQ1biXcOWUuKJn9N8lpAu+Kdl3mS0u
hRJ/Yic8G0bbPHntZb3iOPdnxETVNYWzkTSXfy7IUr6rvRaFvdsELWkdEzap6189
ui9rg7j8BxbuVJsn5jyVrclVq5x/+nyhGlZvOSlEDeLyyLLt4PjE0NEhoz/9Mzit
kugogz5aI2xEmSekJn7dMjPA8b9dXb9q5d/TPsoodyCZgmG0uNyCC35HzKJeqQ2y
jahNThNa1wy7QGAOMfYKH1N6eE3JIYztQZdhKDuQKBZVtQd1QvWQBMFaSwqhIoAv
OmuTAB/zzAFATEU31TjQLOdEotWMU6mGhCbHIjFkXiJ/Bs79Rzo9OD3F8pqFtZiC
DYqNrzbswKV9ufhBKihUQgYApw8IUWRr94zD6p7iH2jhTAtEOYteRZOKVOhpKko4
/EO+IZr0VJpeMlm7ZpeDJrysTTRkw41670xfcTl3OUUuP7hpeuHMu3Vy5C4BnFD8
i9Y2WxhU8BAt8MJAm9t1u7b4YzE2EDaYB7mNlUXw3OIX/UKE86YDOFqO9GuHVj2/
giBqruFwPc1K7ZzBImZP7zBtRSHSIEz5erdR+tKJPC5BjM6GAZBsksBhuC5Z+bma
fUEwJmiaz0mgHSHo3xWOxFRcEdJRvLQ0+XoKxqdXBa+yr0ov2QkdVk3TklmAQM8Y
RXSqSQUWj+zCzCE8CUcz6L015v4QFboC+DQLxE+SZFzTNSwfM0+Yz+KkU1Xi3S6J
JtXMpUFvAQ3Q/N7QeIfOtzR4wL2OEww3lAzNuXh0Igsegq3D44DZDW46DBURWA/M
gWQgjye3/RwEGuDsSEPBrWF29c7tTFZ4xfnTReA6tofKf4ToM4aWa7UsKHAhm8pE
YE7r0BVLe3YBXvYpq59CN+RKezFc1/pQ0euAHB6xyatcc7ukrBdSmld43pMUHAN8
kHKx6+hwsWr3Z74rJmPcuKfUaTVQsoUIDp5f0/xG7yVFyi2n1II/0MSu3pMmLE+k
R9Pz6ckHSSdlPOKr9s1Y7lisn7ZYuRJLJ1cDIyYOst5d22nAwYI0egmqNUTMwAgB
kmeruCYdueu466gbn1DdLuKoiEPsji8yLBGT8LAtFMUSyZKG82hhjz+bbMZWC7xg
IrgNSDH2ibPhxqhDHn3g7+NqeMklVYseioxrxhXpOcBEJxyHsiVO4b8mWmzNaX0q
Gl/FYazChBdL42G9E9c9+R3WjWPKomfSFJxz3xNG8ed3jc9l04fJhMfqkfuI2ase
OgJ3C4vUhHCA5zo5aUO8yvyXbaaWAkGObvL3DHxt6+hpNDFP9wSNPv3IlKmIV8p7
kQUYaCMwudKFW44gzA1Z6fYHWeguRlpxCr3DY1Kq6JwXwWSGCxxC7p6ZeAv1m9QA
gZh74A8UTjtHZjIfFoxXuAOsjO/o2YM5CxNnn0OcaTBCMZcx7jG6WAZGu750ks5M
Gan8uSwiUPsh8gMJ6MbiaXfiRX1G2HDoTKs65BvkfpvjndAYFskdL66D1ExEPCbJ
aLy9T2CdGbVeM5iUEhZvd1sXfy/+AlVg5zMJrvd5ktiXPwi4lb+arGag9xnNMyH4
zSjYeeokw4Lxu+GMReD386gpE3mL7lVD5oiH5f6WzdWMH4NtOvUOqV9tn8ivuIKr
qY/unYN+fGbJ7SrOUruGUzOMHb4BHdsH69Awe8QACMCfiImrtsUywRk7IWhwAUQT
ZFmRnC9+168+vsQYzazPZ/Ef/2O0K6k8rYtuT+Q4QvaTHS8s6nnjvQX6Pw6stWLw
OZwwPipxCSeFIk4Y8EvTCghC+z7GycxSXVboHdLmu/PYOcmYxJaZA2YDgJcTGHic
RuyBWp5Fgk5xziHZw6B4/TwjfMoPebB8eVn7oDoOH1iahWiM//pMmBlJFzUnjjSA
At5iykD5cMo3x4jjZWPOXqeMs27onUBK5WCH7tg0d0vJodDoFRXqDv1bxgpJjhi5
Ac/CTRnGxS9nQlj8kM31cVr4fI1WbVuXstciWU8/ETWfY6nazEdWjeXEuPGHsitl
diwhokIOfI0HsT0fRVt61TV6Yr96DdW6wJKQs3Sia15SepNDV26kma5WRpmczOca
yKoy7+G348RfU8/UHj34TPtlP2Dqpr9bOEXjBGhyAHzB6ze8yzhec5Y3HA2BPF5V
YD1tz0DKRNWc1i/hsIzmzOUbXfxBAB62aeUNMyc1nlaQ/ea8hOvCcmcyjNkvpn7n
icEtwh0i8Y70NUqkBRrHt1I5HsMgatCL9xe81tSsb5HMJ+kXZ2TRDrrzeVBBLGZI
cCSdwpuNZZ1Y8Am7OWoV84ynKpJNbu0JJGtJDP8CYaZFDEu/IiouGCdoj932EpB7
G8Dba4HxgPURe40+9S05R8IvJIqsHTuRNHjIKyYwzgaUJNM8Gd4DOxljnrNONcZD
rhBMQbXOM6sYzk5QconjtlYB5ZWEOTKUG+Q8iM7v6kjMlo9r3KEX59dJuX1P3DCA
KhmrRpVmxkFejbgCqz1LGaeKYBRX0AdHhp1j7qjVTUE6eatSbYzlOqY7aF9/VoT9
dKw+6slOr0HocztRtPZSBKnAldpWPudTNCEH1kN/I+g6CPtkLMt5czGThCTfSuUK
rg0CaWrHdjkGKK/OJXaucKkUHScmjJD9qf33Bf4wJdQNjW85Lo5dtvkDN0CI8NrT
Adp0UECIk2EVcQUfa40FL0IizV8r3DEzhOJDtHjRCA1pNk2hiYVZkL5aoebHxVse
CJoQnSbScrF38/qbfjJ8j6aG/KCK5WQP24evjU50wrewVFh5i2gBQIMMns9vlO9q
3lRenXF9ESVbYUbQkD+ib2XN+GYXf0s4nb3w9/GhSm4UvXKZK5/8fqPzCa+MCEK0
PtiaST5Agm+sZVyentj0LY9D9qkQ9fSPMAAS+zbrhEffp6l2zVNMqq9+D2OEEh/v
d1vJu2l+ZAg7Bt7b9XKm/vHddw6x//cnGYZInSS7g0/PbH6+BHzpxvoahqZftnZi
RtWtYmrYaCI8kx/RIfp/aoSyqkVSJVhXm+r7gi4VjkrAoj66jHXZ4Yue4Zy/DFjo
0lVPOJwRaLSlXHgaJyd/ljge+CgjTgTSTVKk8kmgMP5S4dYG9RculMmekac2HT/a
5zxEN2OsUs3/UZ9H5KSw/gLx8XQWc7pNSxvCu8tMEL7E9/u1CDGw67ANZY5qsOid
YJA24YKyyJayPz99hbybzGJt3vUjrJGwczCJW/i0dlVeNCp8aXJWGsoWLQ61WvAp
rbs/EqXElKg4j0AL3ZQIsapeQWhaDYqCmKD/ouvopuricFnn7mAyarGZSOdix1zm
fHI4Yzbk+/LKTZWKW2j4zN2bhGixZngAtQCEgsD0bVmnlDEwQMleSrM45fzVe6Mi
MUNh8CCN3ys+X4ac+9SDQrNFHKc/7r9Eo8oAnBd+acv8EEJFBFqHF/xK2hbhoD6W
jxGHKQYFfpin+tS5W9o54mmXtgOvExfSHwE42YAk6kVmPQosuaMK5X+js1jACUlG
b8A2GoyAMPC5xEXYIOdJqZ3nZ30lyyU66HRbqgS57SO86ScFnDHg2XYu58H1vf+m
/k0b4RZo7wSGH/raX9UeG0k7ScF1s5kX/dD/IWWc1X8g5HOP8xVb/XWtzudjLQE3
YP26KoEpLwDRlHSAJCpnBQvTfcoEka09OrPM7cqvjjHKSHoA6s7e7gLiqXx+6nwn
ZegIr49BRgY4CcQFR9Ytu+HsddmUrPSuZJ9n/e0d8iVFrplOh/5THwqicXll4lhm
c2XE/svGT5+cRCwSg452DqrrtzZfdxkp7nJS0XyemKHPldOcaRkPwwSxwUEWj8gF
/k8oAz+l00OT+F/CR+SFe+8baxibumb0QBcI8U+T0SsyU0tiXLlB/SjhbYcQyPZF
XZn+p3qzhmyz9qEKU/ePAEg7ppLT6WE4snMge2gvOI5jLLOwr/rojUzrw1276KXh
kc6IyCczFathL85RkckTEtpxhOFt/78yogINH/22D1oUxlSb/kSqqIlpEpe1FZl7
uyk9IytLIfU/aT0LoDNztl9fh0hiT1Qu1YF5bFx6tXnO8iSCbISKaX8XK2jSI/w7
ffRwkmXmRZiloQ3zco4ktkaPBlzG3GtWqMYGGMQ+bbfa2TH62fOivNN/XibOt/yY
JgA2aGjaicZLWK5NaDKdhOWNkb2qyvBAa6SrBHuQvdgXLgr4UiL2lLr7VjkBhYZM
WGLAeSOCnD8QOLBCbEbkJKqXjDciUFuxoXCGwJ2uJtyR6eVDS3LvGjMb8ca3Jiex
3jrCFTnBI+fJHrNFeW43sa0cLXCJ11uA1RreCu5dOOfs0uM8lGC+1BM1aO7uGUWc
UpdbpsAlJj3rn+ukDrf+Q09/iYp8gNW/uFnu+xuvn4OA1TPbyRUTLBvi0uFi0YBK
xJOty5QfxEAYVBQwxZEs/thlFMcHuTIMmLJCkaFLrkMyv/oTO2Gu9eSAgP1m9GOV
Kj1r8zcl6/w1oOJbDAkErpVZ4sYfUngHg5TokNyR2MeAtjp2THtJm1kfrtDc2J9d
Ci/8nsmT1l9FOzZT5XN0qEzqhzHQQLfNr1rCnb5a45wMUJAyzC0KKc4ca60M5MTR
Qb4fXBuX7A4zvzUQ0MBu50dc/kaqCXj9k6QA66iVdlWs65JYUyxDm7K2O6i4Rvo+
Aq8o6AMS70YYdeSYhyqPSK0lfvnu6LpseEl2aNFh+kIIQhE0t1nh0Dd7LG0cDZ9j
zjUppJwRWtnMnJYWuPX5zYEAAUQObHgNe/whUDy19RNwRsHok7yZjUTPOFwVZPof
wl8vBPGWycLxIVoe8tyoXVdHcIqsN97h6fesz1xY0S5H/SDW3C6bxa5tba0KbCfO
l+zhSURmkPlMsPoTCQzIi0eKRcD0fQtGqpV69iFIqkjaM8GtoKok43UreoCJLpjK
/syq3PxxB2yC2JTZeKEFcbEDiLCAEw++TzFkIGvBbfPqNF6GFtSmffzbYPkrusjA
dtOPv/Vc87EuTN7ADGD0u5DFjzXFPHBd7M4NZIGECVM0K/uWTnUs4V0Rc1Uzk+5z
VFxg1djzyi9sDJoU4Qr/WBuwsDIrC93OIo5GzNJuqM2NVaOhjLyInGBiKmQGmcSD
Zjw5dt/XA8U3pfEMrPkYUPOoLwbe0nv0uWhmL1m9GpuNN4p43NQFvx92vp18MyUt
QWpUfIGLhJcwSfNMLCAiKiXifKfFN5BRbAIQ9RCsLkE/T682gnFx+wfe7uakaQsN
JaM1Y+DaIgZjn7U1srkxTjrY+eDDypF6MA142BWu3iHYTUfmkw712rhRZybUSxUU
3UfiUSwzQ4iByI1UOxX2Ts9WNhVo0iWaW/2t9gL23T8OLk+WPLdWb3rtZYZ98mFd
1b6C69hyPWKTZ/dlrZ1FW5Zir/QuNHNwfZCU80QxeF3rAUT8HlJOTzmMsUZ645Pk
i8m0Ivh0wSIERyyuW2em3v757TWxzVNNtpOwSTua2JjxwpGzh5hySKjNyUh/mbTy
WV4ME0UVLrgMcCjJvd7KRa/L69GDzPnNeSqXSPnkJJ6QVJgEaiB9XRtjcgxoZdwp
iDQNhbfUI3LZAVl2JiyLIFnluG7jxCyWlrjJMKW89YG3hi1BgNuKzBjGwGaYM1Qe
tNffNTwV/9mOiD0l/CruvaSUigdeRzvD4En16dz+okizt4oW704h8Dt552EGxR5/
CYHXOPfJGrJ3ehisWwaT/4rit72NcO7tHZG6/armz41+5p2zfZUT3GpoSPZxCP0H
GIdIB75cJJ8Ejo319nv/VAi9fdrAnQgsHFOTEuJWv1IYNb0UIH9AhxKrNt4rf7u9
8EMi87c1Nd216n8kOmiiZqJy1iDeiWir3tYJtXB9cmRSXl0pN4aUvc9DUrrAYiFl
XuhRF7tAqzzE/dRGeb12FQHbL4XWOhpmEA1QdkWBUm48bKlQ+gih4fbKAtW33Jcn
ua9SnmjVgls0JccnVAtJcrGAoWIbQ05+eRimOBSynw0sqMz9VXKlehuCac2NYk1z
tgjRrx3PmQObxjsXsuL5mh4hdaKs//oeBg5/AMt9vnyPfS0+uABW7eMc4BZ7r7X6
weL/7L6vTAa0XZ66Lkh+YALsoj3I/KNPdZ4TffKF8J8LsIpO6jQHZOQWKzeWJzNt
s+oulssciTYhSIXJxcAKFgwX8UQX9AjT8BQ3dSuEFLhrWhmAL6UDpPc6mg10n2QF
qu/LWMyZRCG+3mKNXUORUtfmU2N5WiDAWNzEfX2KkxNVEomx0Qy13FlN7+UhMRBr
NJ7Q6kvnADShE7v7GgmQ9R65EPDgzbAA4gXSGdK2J9tbYlF9sLw2TBV9SYUaFtK6
OPs9G1PEjyz3299WSasOFh+fZH/GatL2qgtWNuHgbQZgnpzvNy3aIiazpAShfPn4
XG/5/YaCF/iDdHNclNpfwDx5hi5c5bwm7fFYECLIq4l0ChCA3e0G0nOFotWZpKgz
lHyKglsBGWPi4xxHRXJydhhqFDuEHQfdQjLifcX++t/gFQyOdutNFzAruKI3CcRh
6h6NZ7jICGaM1X7/7ih4DUQLFlawq/fZ+6RQxSfmUN8pTnJ4+8pOxhIYrMiW7/lg
SLLlYUOhJ5LytPNO/Q9TXxlS/2mkYmR2bsn6mkz86s3AftIGVmHE7kJex7dwnTFH
+xiWJaUI8511e3jlKigpP29b8FRwEMQZWSOeh75Y3gXf+GAUTTA3cg4wGx4C1OKf
dlMz3OeSKelFTg2OXTWqDR6ua4hhM8e8aKBOwnO2N5S/HWcF0PcZiSvcJL2SclPe
UrrLSvzDx+yGg3V3iXEbbcbT1FcvnIgGRvPmKXgIutkCEspW7/6+dmAEq0fVt1su
IE06ZhpYNrQNCdFKTBAzyayyCguvE07+mL1+EGoGnCTasj0XxQfvDLEU2dlbscxW
0szXygxWn+78o/33Xi6oaJ9ReHkGYVnldTfdmz+Dcu2hyFgcMH+F/eAYFs+apOsc
8OKgKoxg/hYoq3PBYrOPynHN9WAPFopqvHdCrwz5kea2xLOM9iZSCfPI30w90leo
9A3lwzDq/JrZndSwuT1G1ELtTCixC+1T6G2l0awQebhYb3AXgTo3MtYNRx+EljOf
dqfQbuY5lmch0Y2cbBuW7v0ZexwGMISYhi1yXiitO6w3bziRNRC+LTtvubv//Vhe
ObTCTIjkM/I8k6+ckII05nnR4lQClZegbqH/os/ss05a7i2tp5POta1leiRKvFT0
3Fjan9OijnNy4PKGo3BsnZ3v0Co6COqJ0t0mja2T42rDJw9v3mogjCRcKUvFwar8
Fpso9eXWsa9Mxmo9DkmCxonjrPxsAH9Ifs39k1kr8281xGyIdoJzbwvURZUq3/jf
rAoXdbiB3NCbT8NLGbFMEN00k8ZC+w+p5ag9+s/P+sbbch+0kkOdl1VG9s4PSg5u
RqhixmA9BZeU6dJgOrrzFrOYso2fKfcPLah83f/qao+5QEQ8KAPSL2g9zIU55H29
4Som5jlF9J1h8NXkyMStrSLCMZDONGqXRFNEdDK8dkNuXro2UBjnX3x52qGQNe79
2ucMnqUnknUZSxvGDnFZvxUkqJp/o52eFHwkK3OS594KtYWOb/syDAyj2LXIHiTS
ScKl6tPNCQIR0xA5p+8YR6vS/QdP2IB39hQrHgjNnL1ntaazqVFv4Pb/CtfZ9gmD
gTbw51RrcZTRRvtZDasmLCP+1OlPCl3ftntmfPp/k53nmIplWlcOlG7JkGXQ+ZPC
x0h3tFm9GKMA16VmNuBeWWq+CKNP4lBH524HlnC1AMsk2HiaXPHTqa+h7XRBfFqe
KpFsQltMXEAovT/sKPxTh+VaR2skPfwzB3PbJIrwRbtf/m/7sBEeE7WcXcNbjU2Q
bpRQ6itKbiz6efXLkakzW2GpCMRNTXemrAHmVd4P/hUjmaUDd5syaDPnKH2etL8t
fN9U8i1x/SkfLGmqUi0NCjIa2q4RCB/+ZHwseeMrRGEjnIgH4Xt8yM2cXy1cQ1Nn
IYuR4PWTSXbzqeWNo9aMa16n9AMwKLgNDne6VZMXO4VhmeT922OwHJR+Jh/FRL3m
/CGeHpR0A27Rhu0CRh9cZnN9R3kqrBm/TSbhqbnQBk7vLV9T+fD/TLBe5OvQwXDf
rTWv1QUHjx1MRTjrSsLZKSLKovnuwFK2hnqvHNmX+jR10Uo6gR3A8CrrEaIzYwoV
c+I/gR1PvQlP9hKDhBFS4PcDHndZjn03sTLC+HB4cCMMB4WdGe5icqo8h53rOqA/
O/ifz3PVvpyQrKy+QBvxE0YfT6PP85yTybBGq2fZgykmuTEiUggMCfaiakCZFKpl
YRUwZO+bYU8467d0O7NJVMdnYlNsaLF81nq1V3drntOG0QlcvgOmp/pYw9HhfXo1
/1LRjvdQFaaGTZxXHADnN4xCBHTa5FApzu04JJVCJDaaPN+kuiKi4cxkbqzsRVr8
43KZgDdSugSWroOuPYOm+9ggwB6xz3BrzMnxvw8RxkrjIRKAXL/s2mD9/QKw3Aqg
twKKExGRzqfHUIxzJCXXBSlhrIUVmWKIWdabsw5ogquHz+uTOiUU9wV3ziS11ECQ
7LUgKe+yXjQNkLwy6Y/F4FsmI6aSxhI9sLHy4HdFcJuamI/MB6iqaf+Gh/jJuOmF
UmM6ZwNIqGHpoGcyBzOCgBkdwZVs11olDviuPkbtVdPIFxD258FGWEhyA+TlcmG5
B6iw2VkepE+iARPItaGu2hwATKA2uyeJO6YXiTfa/GhlUd3X1OtfeTcfRI9gCuP/
W04brAK9M0ofoOkn4YNK1ZUQzM6mCA2cov0ltcsI6+PV77U0ankADma/cYyH22u9
hEDPezMSx5OgON+qHZW7foU92NXmAtdofwvhn6UtEvFYzdZEHtPwqEVyB8vImjYq
P7A3E+GyIP7r4CcUogRqwxKY2WlOoOgzPWJtbAckY7bygYJUQVvGPHj1/bhBhuYU
RsQro/2mjLWM7fFsEBcQjPRPEnBsi1QH0qg0sOPoVcKMaUJJCV1QY6R3Gr+5LvNd
8eBOmNmzO3PbRuc15OEeB59krB10EkKRxAxgHH3C61pDa4suC2yKyUeAhfneaefP
eXRf6w5EpeKE+XiDrnS4dwbnaM3cfRaw/WD8Q67gfndN1cgL7fBYo6Dalx425jpE
5w4YPBxdC9ByC/OLk9XgW+x2fN3pvMljed7lqNhvfTxCT+n5sn0eeDvLebLLBmO+
OABjncM4uG4bXNGH7GkPuQ2hJPF2gO6aSIaDu6gBhDugA3+1hjhHlxzhOxISz+f8
s1btMn0P4ABIeOTtL38kl73isRI68pDmfNjZJbXv8iwg4uLMqXG5S9OGU37zm0gu
j8pRZGSsxmoE43DSK9uQ3lmpoB/lpyDxIISMllTIdkx8mzdXc1C9GmqENGLXQCZY
7p+rE5m31emuAFNut41mi1+pH3Ke4I8/k8rJShu6gUMMm1J1ZPUwxxwt2u2c3aI7
gFI/tpWitmgZtehuhnILU4umUWJATEXJI9ZB/MXwZGea5Tto4TgvD40MYx5tNLuV
gojnnovBqFkjsuBzdvsoT7HPjYxu+driYserhLvgEPll5v6ZJpR+slpOET5bfBY/
c7gposGc/TKGJydvN1kFrKJnQdPfLYmSqcGfabp8OPPrBafjVEmCXwuvI+pst9dp
WVMx0SOXLUvxNM5OLJMwSI3MpZDS6HrpWkZ4QZp1pe2mKoWbPT8acz+80jD3YV38
0+2XZ7cPmEdIiWtazs30eliwD/TYHRnpKUAeCgL1gZIshZt9/8sInkPJzhSflpB9
KZa+jxD2VTIIKCp6A77ob2+ARO4etojO19/BeoYd1qsJ+XnjXWyvv26nC6bsC9uZ
hi0OnK3rM5wWkFX/VVj+CGSHY9pRew/RTSod2lSwY+sbU79OIps0OdTjmbLUO2U5
NWLfVZBydlCwOfuHQPlpbkKN9tzu/Gf35MbEoZwlJkY3LjP81ok2Zzf8qrExC81o
iDndxK8N7mPw7bE6Bs38CjbZMRU4mRu5MzoCpdgkpgzim+54u1ORk6VQj7rM2Lx1
rz1NKKGk8EhKNogwmnPWD5FMpSE2LXQZPjAJTVjd3AcU5EXmXdh1+yiw3y+pGq7j
cpe3+YYqF3aK+SjYogtl9VQFvc6NGAhJV+5UaG7dj1LBpaarsxdAqvt4VD9qazJF
gZ1c6C7gL90xEvwN7leWUzAIuv3uxooDwSEkBY44P9oRFgmQjL0vtv51SMHMTL4k
pDu8K4MHjfWh1ja+1xZFO10JdDyyew2GDuyL7Q07Yg6zh/tU4TCZDDjHikxepex2
X1m6fhUhRt6o6uE/7yBxMDYudiS9P+FVyGcSkpTss709U01GCszzzRAWXnps4rhr
yJsLGLEV/qzbxczuHz7y2UVEw3VtkqGFozrk0CsOQ4TXKwyzhvZEksOVwMRmqlNa
Ve0jaPc7PBgy3Sgpf81NcURRVPdKHihFLj02QD/OArhkooXaMnof7eoW6I6Stly/
BnBHoOMJAvxPuTaoZc/jJMLLiVocOxnFqhbom7NWGFsUI/6Whv4OIHDxmiXWW8Sm
2K+pUvw/XaVJYYpsm45lKwMdw6ej/u16XUBLZl6RByiYdgofycd9ijbDdtRfBcbv
dcKMcIoPeq89leSWLQoL5+AYfrI51N4M26TFM/fU+fmSV5WU8ag/qy7ZMqQO8bIh
oeOVg/vyf9+lENeHeMwGYWQ9d1Sklkr/YSUdh6cLUmIyVBDablygklS4HzM9vyCu
krvzG15Ky2R1Fkx/aBgFo7F9+FtyzcY3NnuotfAnqIlhvT3bbrZVW6CqNOZ+0Ef5
koND5M26jFaMtYzPZiNpvV86q2synEThsEZfFOEVfyByGDUrmv2L/fZpTNjfjM/+
WgQC16HDT4iK+HMjLjP6BDWRi9CvN4159d52m/lv4nH9re8HT+X4Jx4+ILWyOgir
QcPDBrSgl3ewHe2dPKIEPYF6G7eqiUZbqh4GqTyBqnPM6CcQKBrwaQh1JkGCfXn2
DGWfLcTNZdYCknGAEYROG4gwLVnKpeJVZVNuJLhLRZ6JN46o+Xu1iueBrTgEzsRp
XbwJbXA9SEmA+pSVkPVoZUoiRQ8oNVxCXGEscUwrhACaYWH/w7tETQLDUzGQKrUq
UwIztScB41BeNKQZPo7Y1JaCGuThbmyVkbktWdmWTK+So2pnChb2AwmKDgB3etpz
8bu3vMXl11YG0zDqDQKPoNRL8KYc59//c2ycIJNgz74i0NCV6o/VWct9BUoUE9Ws
9AFuG/mOduXV2oJEaJf9bmiKdUz/B7TxGZTgM6r0ZzwJQ20cTVdj6jRNVCsjW8hQ
LAZft5oXyRt5aLq0o/3S2cz/rU5scyMSicr7yvsdGmZIaQvGLd7u34ZFLFqIj4Mp
QVecpfDhYFy2/RUV6UVj4+K4lOsGrC/e0NUWrL1PcGV4tfJFdh7VGyjJzKfQST3u
7i3d2rvH2Rk5I+PC6FfKDeESG6Ygf1kZ2R3pqyxsCu+ocdPiOG5chDnYcdcbob5V
dJ5J63CccWJLzy/EuxCA0hotYNNaEHlHeuU9kRGkD4VC0igwwshQEpc3Spg00JFd
HWyZf3sEYt2zUSXxaGkJWiFVc+G+uhlBbTZp7lDW2fI2XazEqXYfB7+o+UoJsfRh
5RmAvqiT5hJAlrS68sKvy3ySGRuNj/wHOX0Tbm5/8KCJDetgb8jbCQMShiF6fCtI
O9QSvvK1iNZQNduyOUEdXPnu7ZH8JQXsF/sbNwA2+H646ogtEwn/PMFC9i9XZMgN
54oOB5wgsstMzREgLfSrHbohyGk442eyFL0NzR9rd8gS89g7I7s0LM6VBB6ZIEs1
7R8DR6HJP14xlfVMXqf2wIOychDrZgCEw0uFAjHWuMfCeVR0SKx5WYTKTsFi6OOK
sc0rS+e/7bJVXbYAgFsXXRxHCM0j6sVt5XSR/wg/aJlQ5/pSxBUF9i6fqUp0hyGn
PCHDZoIRcKhn0yVtNgTz2rHWx7G4bUPJ52khDxn567ubai5PC3fDizSmzKbpxq9x
vTldiBwt7M1h8pmsZCNNBSOzaWxlmWC6Q3XVtQH/EdVRQ6ZFPj/UAgDpE6CxZJbv
U2bQcqBsjqbWO4lFyKgz50JRPr3zcSFbX78XUsjscEEfFEqmJfpg8Yl/6fA4VXqQ
mqN7IK18wi4DUyVEFBmrhOG/cpUTJ2l0bBr4+8AsBW4nw35jHxk2yDYkeIzSLQuC
8bF/0j9DUKMUodtWyKs4zSfGS2TUCDI5Hb5P/Z40cOVWLzuuQrg+enVa6GWVnHfg
XaV25SQx5YBIrqjwJtSzEFvSg/F1u4oJ0zCqGmm5mEu3nhzSzv2JcvYCdpXmXmht
9QqQqpW7U2YlfpTxeSLaKNzSOM0GO+OGG2myQS8Hu7gQ8nmS8Ir5ESAHgyqNElt5
hC+FGUeArE1Om72An1F3ssU5LeDCmli4bu1yttoKIR4WuAg/qqRWCkcaF13r1hYH
6whYlb8tjgPKwEPRvGbLOH02qhbGtp5+XbASz1HvEZXaYTDb61t5bKY1Yvqo+Ovo
uzCMl4ura+2nedLnAyoPNCDjOqrfXMmRdONPhFU1Cro5ZwbTyaUDDwoaS07fV+g8
U3Vw1lMHXw6GN0SSEvvs+xdOjLhhdrtlUNRH0o9ykts4ZZWWZf9CtBIctItRCTNJ
einiHaHPoqNzEM+UUJbtvRrnM7ZUyNjlbRuCuNo/Y0a+nU3Fw5h6f/Y6n1Bf9Qjt
9ExM1S90rCtWdugBXMwUoBI9HsJob1ar3Yo6kPzk9SisUxVRjbOZdBjO27eGPgk0
vt08vMM3HCSQxItOALDmfRXzUeVoLd1aDfF4Ednu9l76tbnw47utoPhlCrxHqUWj
`pragma protect end_protected
