`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PSlov+SqS/TF5amcdSkf2aPwA/m+FjRHfu8IrdwQXY6eQhRdeGuUH8rX1aXKsoFU
agtb8mS1sflo8F+Azv8jMpo1HphA1B0TP/qaefD/PJjChnMlH4r7gINeEqQnJc6G
7+pt36JTs99X8/FLLMoL4K2RrwjDSBH7jTm9IU8jaig=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
w3FPQPmKzrZ5j2lDz4FvPZmFXnrclKIbWFlocVPn4bBA2DtLQkUts73Fke61sZ7z
UlY82qpNXVPZk5I2o/UTW+1g2NF7+LP8mZT2kCnTCtrZ3e7ALGUhxPxMP6NKa3M9
kvmjCTPIUpJtA7WdWbG7e/q2UwI/f8VVxLYjWKzZWz8VG/NDGf/iR5AJ7iNLA7H9
eCFAjT87flhqX/Wtab20HblTim8Jv3zoMEbkdTNo/yxkxQyxgkRHwVtyxlJugdeC
P6MEv7ygkkb+05evlWWefG63/FP0Dh0LPgzc8YKEBCdNzVsKKMKhnx41aeZmJ4AA
TS7tnxmbnLBZOVcWM50DL+7QNx5JhppDanweKbRFUYGRsp/2ZC986lOsmjO3SRQC
CtGSZqMmuJI/n7uxuDR/eMcpPmpJrJkexbhxtczPIMoVgJTsYv/w4/WYweOkSm2Z
PDb1W4QS2TNgLt1jvb4/yzacGhhLxEbbbB+L4js+bh4lnOfeUnM49+6pRS/ZRNWj
MiQ1ux8Ogo61hxSuKf0nGAmgrutY7g1Vf9cneRqREbBHuZwq4M0WEdh7IwCfhAao
BRNa1EqjlR6oIxM88GYUx2QUEDXzx2RzMcgMR3CI884NursoTemFNmyBsHGTSbmA
Bv5i23RDBqWqCS1hI2n/rUob6OqTV8sNaE1pmj8o8Zcdq7VduJQlQD1yD/+J42VP
HG3WsUbqrqoQ+9bfHzXbMcuNLKGlwuxh12+E4sP/6hdpI7xArwIl1JZD2IIEbYxP
eVXtC6av6/xqyUnt9drLvs7vwS3kzP9c5NiYo5nCkD46VBQVkccLfov0wAyInK0u
IXfzS1fSY2pw8V2a/Tmp+IHI1FrwhCXPvrbxE/uM/WnpzdMUCHpLylo0ThB90jG2
FOfACQ3OAIuKlqpIn9YpnU67R+RsnizVbSTvqjtjgZlgHiYTXeBDcIM2X071DMfZ
aChqstkfItp4eMU107Emd9zq+WEV71wY5A/bjY21P0fChLkfu4VbPYhGVNbkF5Q1
a/KGHgrq4Q6exMPyOKyy0vFYDO9+gijICC9eqGTejLeaHcwwHZ6wcfUM3gcbsAvX
YRNGSMc0u75tBjMaPBXcm4kzqu8HvPPSGbCtGMB7cPuVoAMXTm+oc5VSFyQHKT7y
jn7QuPFSzGPCTaAxU1T7kTXPorpX9gkiYQFv79s4YahA4PxYApVPCQAbH90eGk26
KzI+GealDn8I3YbDOvpMLBrmZ41SDwMvKe+3HDT2s23oRlrvGFxmoVuyBcnSocZU
D7Www1km6WNi95GvtJD6gy85/VL8PInA03yIsNj+C8cS1wK0cpl2OQsADW4QI4JR
MIm5NEuPovgHPQRmuUWXkLjZ1gwcwQfBQewew/nC4FnQiGagYDarZAGDB4YXqY8i
LdEs2/BxHvD7F9/ynvr7Mr0rnwA4G795rL+BoPbvAFciTX1C8ohB78Lr2oG8rvLu
Xv+0n4cLzGkcOxDp2QNUu57zb7XoicaP4Anj+HQjnx39rOhmnz1Jqxy+F7LnDgtd
57RuK3ZGAHHbNdgKjfqfJK0NrFeBDjZY5PrDgsqhtqvARKpL0JSUF377UzKr5HK9
eyFAOSAe1ua2XjepTuda93YiIjFBsP2ESDToTBfFQcKYXbWLkn534cVYpcgbBPAt
Ljm9x1b93cB9fY+ax/KK9OaMkDxUCD0da3wWkRS1lM4ZL72Pw08NllBdxN80RlRx
ATYxHE/mzwQoOcGUYi3RyN1GAOUHTJP4/vjZ1IjiB6I8mcopxZwa+o87R/b5mk3b
cY4HqXTGvLdc1fmwRk+CxVEgOts3ECYNOMjDrKDEFvZenRaC90CE3HmLofNCW5zA
qrVUI6I6MxRMvWS3cG+cvB3NryE/CpVxaJe2HGhiWc+7yRbuCI/MMTVFkobt9/61
HQN4Vsbhk2Xq7+fZb3dYiCa4eOLx3o0jffkXOvAc4Gf36vscEKez6UXA4xOWrskN
z6ylIm/R9gux/ED6pIHwucPhUDnzILP3fY2Obmrbdhw54/MsWCvaKmfzUv6w7uWE
oLPzAJ35xThy9QH1pFii7/dkdKCQ+jTZpylyc+IROPHGfUkjbzBNqGyKcTkJr6zB
zirKc1G1ifUXvsHDMdT/C9+j7fFHeJ7U2uMUvYoVode8KuNlGXX+g8COMLU1uv69
BmB4xH4sKB9Os/XaZvbh7lwTXDw5Uy+m2eA2jua8BRK9YPulJUExLJooa3O01Qfc
ncbXzH65E4pmyWrkNRQXpCjaRll3TYP8C8r4bAQTz3yZAwnqefsaoMDV9sqIHg1h
H9uMB3DNdkpZCFhNY0y6xtbk6SwCtoDiVp5kWSf738vWcFoiFIerYCLSCA8MUHw0
dMO86IfO1PQZP8nXPr9RSKqCqwFH4o9Q2RwGcjkWALIPzyZVFKHscvIgjT0KXEoY
Ld+Se4o7eMolUTVLJ4cR1ehdtuJLQWmJzKNNQCK1Suah/fWuIKUTTbOrUE8rCfwq
EfqN7Glx4nVzOEmZtg2xZGsyUI4G01om7SfqXcGB1PUdGdlFDQFzS8kj6H4FYc6Q
rJ1OgjEmI6D/MJ/Z9dGvVOwbpI6mSglcwmRdzGfSIqpr/6bcqbcI1h7tFpoluIFH
9l+atJfCB6JLvQJe6UgCoLk8A10gjhe6ggsFyl1bMg1jNA4Wjvaz3VpbclLGkvfi
BOz/TxnnWck/fnRoMCG5CoELSBkK/v4G/CiXxwNBg2fm5MAEeQRSorciiwCU0FVi
HCiWqo7jD6KnKoX30iiYo5a1CSCnewqVgsbCrZIot2/ljdKi8qAYZRequYu7U9fb
Da3H+2nzt6tVzTkfGvQVyy+hSbGXE8BmZOLNQtLT8/y6b+FAPtovWT+MKzx3UoGl
V3LD9Ay+A2iyx6wyh5CyuW/uCuNl7PphOonZB+L8EuGOfPjjiSCuvqvJDzb8AUJl
n1dpN3aBiOcunnD50/2M+ZZvnHbtZwlukqVzA5UEUL1t9gBp01iDPj9KOp2d4mgn
YAyaRZThlPMKDuXoRKg4eCCCAbnwR4pxBIiqrS+720SvGgRsFg1dmKdyGe1scGDB
QDmPhbmTqJbIqPAtROp7gwA2AdGt9bXTEOV3HORcmYzmlpSi7O6SPDvgXpNH8LU1
LjwtE8q80Z7AiJ/KXXKO5ZZ0aevSk85+rWa9RoZYCvGvEszpY1l+Wvr/lnALfqC5
x6tp0Tae6DfaX6K8NfkGPrfeA9nmNC5AyRyntFi8Y8iYmmoe6JP8SeLrMnHA7ZUC
x+Yo5z6BPadTblbFthRE5MFJzKxONT2qacRYq0XYJ325ryGJ1SWbOD6AM0eLvTL/
wlu7IVztVjlof+gjBydgmmRIXQo6xE5LasZ0iiDGfGIlsDLNns1xcfLwAueTs8Sp
Y+DRyhD84XBIG1tFVobL4zTac4l9nGbwFn+j9uk6oth82o20NV/lTRKwrN0JDLHj
ZXNJhrIASOJP6Wj3SqOLtya/m7FpyzMFZiB0eLg4ZVJViLbmCihCzyjhKPkN0OSw
LxJqI9KdTgwxIImYkzoWTBVXvT4Gq9kiSQysHj07PsMrmIVZRpxzsoNlFl4ohSkO
dH/zZBcYULL7N2ShTVhbVxzEFPOHJNx6zqKGaKHE4PKbFJwCozMB/Zb+F6uU/oXy
HbFdKXKyZhFrbysCjd7Ztnzyi0lr38swB9BflJwo6vd1LloAJLfzH+L4Hcw9a2A+
CFV/xEFuFMUi/B5i4TAkJKLXSeaoOIgPooEDCEX8r4QS+Zb8k68ctKQ6iast3uTk
XuhOQKqbhGvJG6ONsmni5NLPEytwWPter8aPpHoTlixDQjZcmdLaNKcTMWGF9MkQ
JlDl3p6HT8+aIsOMf3RdXsrgcyuTxJZh9GasezaVchnomdUOcDBh++v/ZVV42Tvi
rNINOQOoXDyKDl8eUyCmOHjcjkA+cvj+w5SEWJ0QNBwMW8LFvW8DJDDt9EU0CNU7
0RdbEse2seK+P4lhqXzfD64b21Wpn3hlFYgXHxVpovjRBbIWX5KaZPH04VhQvVKA
47TlCj9IV7Ovj2pMY+o5MoLMROER0bqlMBEDX/Y1s55jo+UJU/0Z0MpbsJoIr9Ch
LVBh8CNy4Kgy8TV0H/E1bWBsmWbtUzOTlbioMyKIR6a2hHRPOu/PgjSYcq5PUBTk
korWxaM1DFYR4MWyU9IiiW+If/6VufqNmJA9uvhiXmcOpr8DbR6B3jRDdYeIvxKv
DI8oJRYih6XKYCSXonwb/9GTa/0JgS47Aok2oEFsJCX6NV+VeDSaaFyflX4Pi0lv
cAXAeUWg724Os05ZsI1ShEmfhMJ75PYY8SGeSPOcburvLn+lPY8uHS1waPwwX5DK
kXnO1qR36OQBR83vRwq4YXqH0r+9SBgq+UN1ix363x5K4DR8S+OL534Qwrc1POim
j9/sjh0xO2aS2+0JXdCIA4cnh5BJcjDd3ATCjdS8D5H/spclYJnlB26oZVaQAK1+
0x6TkJytbtLfBHOa5auA8dXXVY9xdFpr4FwJcdmIWheTqtm1RsczTOKmoHNMQXq7
Wb47C6oVUR2TqeskbjPstaFhqHkZIkXXTXGEmbH0/mUNmNZU68tghsfjVevJStz9
8g67i2NTXkogxXp3K+2ffh8YawyVtNriq8xOnab/lpKVge15lld2HnN9BdH0PBLB
2pZOC12EvXUR5FYYRHQYugsk0i/R+Tqp4xklMpQR7l9O+m38A9/7GXonoxSey8YQ
pRteYap08oOXQSzbFaJKJEutnCDwliHxissxRhEfnyr7OYNMKWx29iE7310PWYEX
ElTMvysQZ/OuPS4URy51hymOWjaT4FNCFfkoXj4SsfR83JOKewFXMloRy2xF7z53
apsKVadDetis0HqlWpSD/urey0hIjS8lP98gsOA/HXkYuS2MJzZ+GMeNM9KxTiHH
U/Tfz0AnxLmN7V/K0ULO+869qCJBP1ezSeDp77RTg6rcVUcaZJjNBoeX6YzBh1Yt
P3yck44hGSh41e7peqQZCKDO0eqxGop31O/EjRhBewWFGc9MXuhMXsCvCEK76y20
y38M3gLw3Rcz8qAwFN7FE4sc49kvOhrUGz+gPTqEpwb2pe1JovAnzfo8S9DS13Xm
kY4I6NOISBQROIArdwcV/dizF/0yiy310tOwLLY3c2MKkEakPld1DBgcLk12S/rO
JEn5OKu4CThqSzjojXVZ9cGGfSmY3RL7k3oXbgxa4B4S6KNaZb4T159p27RR1rcJ
HlE8x9dCiHqRGMquV+bKh6rEbp9u4+WvZirMzwQdfigBl4exrgnp0W745oAmIijX
F2559DBfqoGpiKeRtrFLB+W7UwiN1JL+reveI8yx/HNx0CC1ri50d8PEVm20Ystq
vav5KCGhwKRvAptNf+fcOa5WCPpFUWZMQGqsylTXY6WkfauWUVU8awayp9xTgBtP
QAy49eiicEP9rbIW0gLZVBZIRbr3vSsFKtxGBIKrzCI3IVvvCIHZfBWxVgwzyYpl
7LCr94MhmyouCL4EYDdAKYHMtXzE0Ay8fIKar1fOI0czb5xN6Y8J1OJYIgZdLPtL
x8b7ki1x+phXAHwhsiDE2v98iUoNsMU87MZIQtuI5FjnP7tsFB9CJkIj7Jo/4nOF
7TCqCTr+wk91nLnjX+i8HNDNATcKc/6RH7JpZMYKq7lKPcvwjyS8o6awH+jLVLJZ
aRUmOUxfEsJhpYHYCgajCmiAL7SSqrEe6eWPpoKlKlFLJD+e723uPZbdIV5ZvKfb
UlI8huO/BEtmCZGnVSL6ow6CjsJWHqAui+HpeUdg/OSlrtMS2/5KgPlU+iF9Uvce
axPYxrQiWv1sp1uX1wtSsis8y3A4ISyNMxruSQKpt3A03I6c7DfW/eBvJStbtjub
T3l+kpdG3jfce6gmUPsy8jRN79D67JRi9csHG6aw1SeCFME/K2UMKq8DzbgFO4a8
TtqTnO8KbHpkpmsYmsqZLGGF/jx7AYp0ZndBvJOWjCK1tRzMPtLvNlMF3pK5cY7l
axV/fiCE7YBXMq85P4kpGoiISbm0U/SfUJfVs1IDk8tNTKPCb2NI2xoQ8+RlWhko
pmRx074FVWdD1XM6zx6r2X4XGQ4bNmBXWnaukZdYxbFEj6Rc2W17ED1j1Z40pXSg
ZR5gdnbNZUz09n+knTTkOu4BvNa2ffyI82UIZnVzytoorcT6T7HhKjDWL2L/CaGU
07TFpgSyugY4oD5plxAY8KDj3M1hx3d2ZuwFCJA2R27xQ8h0DJOuxkxNSuVXjR1T
l9HA1s1XZAWddPLbdLe7EGw28bqwPKwrgIupESkEmcGRx+0IAtGCmjNJmqjYlUjm
ZXbaW1MZaZABjFIJjorIIFZeDdzcKObbhuvRBHcVKIvB6IEs32fO5DRdQAYs8v8N
rz9YExuat5NV78iAItCiDxbHk+1WOno6xb+OwpwGyKaK5/sgFr27KDq1rnOj0Plr
4A8UE30UhfvcAuT3o/5GgsYuQwJNQYZXHVx9yNVJwTc1IBTbijj3shgfV6LF9ztm
c7i5MR7A5DyBzfzbdcPXRr142+nqtoT0FaBatHFoNTMTBntoxcX5B77e3I8uRefD
eR4k+CErrV4tqmDOqR8vx33M+k08ttDS401lLkxJPx1bP9k0yD2+iaAi00VkG6Qa
ff++RB524Dha4oezRPxdaJzchnlhOGVPIEFKKVh7zAp++TQOHc6h/P4q2FrE5LR2
JDcAyESYo55ZZJIUU5S/YOV0u4WM6c7ejdCS2fcRH+q2rdZ7Se0T/yI1/1Hf031n
/en3FXKiWyuWaQqbWIrsDLz2jMvOIwxFXZ8mdRPYdVRjx7e5MccDOcwWGf0c7ZZG
eZ68TIgP4+QLx3I4psM4Ip9shCGyrgZg6k4FQt/IgAo7gfBK57iAhVpBOGEfgMRw
`pragma protect end_protected
