`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bDNCKbTclf6lzyJ64Jy6ydzbFEFYljHU4x97+nEd1mgj3kXTCyyBRrQKYs0v7ZO/
MFjOaqzhUEn3VL4QDiUQktzlnRmrnWtoak8233jDN1XjhJo0Qi2treSUjCc0tUV9
oWBhWQ+cgeutWE9oUAedplBrXeCu0WoZeyQrX+Osg5Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
dmiUsWFmiXOl1DPaQtOsgLmB5wDqOhAm6fvvR4JEY7ySApw6NmrMrHZtT2odbAdG
iQfCrejFbpr0BiKvtJWPTLGNnxUmknPsMtVY0sG6LgJjBVKOch1Wv5+Cyk3AcwkT
9bubPcQFAanH4rUhLmT1a9sQu6tlKNj10nbUOn08XigRrqyJfjz2iT9LhZ9jQC5A
fUc8wxfKNQyPaQHGphhZZnmeBJdrHta4Qg2VE9pCGCEvpE6Mwm1F0lIYnCE+crKb
DNAtUi/yo9DI2wwAcyNjwbL2BPMat0zDCrJXcSpTS7Xrgme18Fn9jaIDf0RoXof3
YlN5J+e4moSquhxHcu2puQDJvuARhvc/vpJmCUKry+nV3leIM/pwceCAOxAUbdw3
jmdoO/zfsNFoxyDRqawQa6rTpb0fP5nLZiwL8PGdNxVTA2xjyGWkj8Rwh1YJjBUd
o61UgNFTlN3WRu/9z6MUG95hzplSvY51b7QT9eNtHiTbCAxmwsMvc3NDhZy1HTKG
2L9xfIS71p/xk4Y65u9wQWNbLy7AtMdXxnJh5cBR+q5qJTksnyMkVhzt0PK0OZ6L
NLz5o1JQG6BmVuA2fQyu6MJiwEyNI3ivNiaAFUd50XomT5WF/0fD8BdG7qPZbbp0
pbax81K5Gzf3Rar8YRJa8NVvS4Wx5VP3N+6dYZT2GJ6LM2aVefc0L/aREWmRfii3
8yEWLE14k58WTb6DI7R8qYB/iuUDICv/2OPVlOBPhQHSGaPk7G5t+bB+0XBxEnaJ
7DCBew2J4EZtVR3V6GSB56CkiI9IezxIyKb98yB9lg7uA3G0l/O32HKV+mTsfrVg
a0RxzsvBbZas5Ze6wEGaFIaJ4S2Ekwnfd+2VQvRfA1WrEMM4xqKuh6BRbXuwmF0X
rCzTcLIJN7A4hclN0bWMtgiha949O9VHdGtLHBIp/NtIIGlGpobB2WFwfKIPyjUY
5CT1jOditCSJ1UC9eQWUV6WcDycHBMd4vUhAQmEcD0iCdXcEBLX8iVceyOMe5oT/
DXcdrL0bR5vrDPJzJfxyROHcElgi2WNCgINZMfDNlqvfBN0AtlTXSgqbBXMh99Aw
15YfsE8vDpyi6niVcOOWbLQvdISxSOsXUC69F4MTATl9EZzypjnwLS4DsCmFwm6n
fUPT6+o1/7GvEUFmlG5cCLMHiZM7Xw84rASaLL3n1V8LHeNg0cqeZeftzti4HntA
u2f6BkcaqUvxob9EaitcDup7CTuDypAAQOBzkAv5KxfRAD1Pn0zpJlGYrkZnz/1q
dh5F+OGYvGd3u3x1o3W98KpLbeEFeA5FlBqAOxKi83pMspUxOrNv2qzupey8o09G
NydGtZ99bRjA4TptmcO9mxEz8E8jj+mgw/F/6yPCcn7IzydwNz5yPeRNAHuLOrz0
MGYyXxFVUnhC7zLzzy7hGSrXCSR9wPk2db28vk+mr9g5hWto6PJ+jKKFdRMAWgLV
ATa37Y2FrixYsWVr+TanHmzHDxZzbFaSIgYx4zY+e+wdhtRySIBjCzDHWPkJpgF6
LfoxkQz5qDqWgK2dZ1ssYCnCBudoK2CMkbN+VsWHKmXUTpAX38U1KGwz7LWnrUfE
wkihi5xQ28uQObgMjp3McYhE+eqxqec5ALN0pghDfUQQmeYoc7UzCfomCTVNCk6e
YB9NVqKIwI8+Ikrcpmo4jazsbdUl0KFgABuYZq+b6CJm5VONnSNYi8aRVFQvISO+
lv2eQ6sRpTtjF/evRK2qkH3FifHd7qRdqVG+1Ri2eDx6uffgePEckonXjcuyOo3B
C7i/mazDhobbzNxwzZgDfMvz92OOQwT59Qonk9oCp2kpVyNEtf8x4SYsl69svVzf
Vg9ir4aKPgtWMvJyFkIIvpag7EIhXJOKndjv660aa+2i+MULHzZ0tX0/8C7mx/zO
2MNpl+TOU9usEsUwQtoWWojzslJzQCfZ73tHAR4C3jU1za0jBFDGsXpF4KamW+vX
0c05fYV7JmcVaAXTkJrBpWwgqeLH0vA9LBRdMtc0rQwb7NzGk6qAMem19VvSGEBN
zRerI/9i3IuNEqODOsnnAqcOKcuoi4N7H2acQht+u3zR+DT3af36t5psllbuCmuB
Ym1LjSxkamQLXaM/heQs0uoVbW+9LDVxTtbMgOwQYBbpX7wAetRhr1YXWYU7ElSV
9tOZJWd0FLr5OmmN2rbFxzKj31446JgdR/+SxVNV+jZi//k3KLnMsMGhL7Mwla6Q
qB2WxsnGf8sW9j4veXdkbraCwRFoak/KSs9TORxm5FVAHo/cSU/x/ruJuXKS9T0p
sx1nf8hI3oMBNusXWsnqyCzo4uNXzkRxF1snw6NQEZMAImP2kJK6y6/ZC74GpZk2
c2b6/Eg0s2bWkXKplOXlukw//7FB4DPhBxltmtsiVVWh8L2dBOi9kC5uUvxa9+lB
QCqCv6PETryyAILM4lKktboUjx84vBa0snyQSjD21ssOzSvw1soJUBdqi/JUkD/P
Xec1yASMgMY5dJqxl8ujgqY+1Chggzm6GHL4p+E9PtEWVN11Xd5//YT5qo5ltdSl
V2sw2HJkwxVff59XrtvvVTvhN1GCn7byLlCLKl8MwnuKK1psG9+VW91BQS4zMWmk
ZakqAieJxNVfbBDhMek4mxHMwSeBwXLQW0iTXrAbhgiaYi8a4eIFTXFJdQF+J90H
yVJSsxg1x9pl/FqfXQyKHIMBUnatzwQpuR+p7XyQnG8xD8b7MbV1vXwzPLjaD5H5
2uevB1ET6LAaAWICBA8gPEoBAXJ5UVzi6yN3t0GZk4Pnf2Y2RleD5JC13pdf2ckC
lo/eHPFjrhI3FuxWVGJvhbTXfhubXi5xOyC76SnXGeJf7vJ6InVecsC0L31QjCVG
yTsGWQ4ySJQl/QhUnIohpW0DtPQqaGTAQUwQ/QLJ3n2IcgTO8r+f7yBm5uz26gFI
n4uUfS0wx47G/e6HPbBAglM1pwQVt/oFEVRK4vc8CnSqoRyTwzy5AzIJFYjHh3iW
c93RLqFhyIqszHJcCBc49IuurPbYHVRT6Xu6KQjCY5ehO29TfnZlR4wREI/sdonA
eNFWbo+NCf7O0P+Yfa/5L0D2JAlknKN1hDtI2nNKcO3lpef5zgd8wthO+f5/6prX
NZkBQNBsrJUgjjjfUVFMdvD7D8tFlqSV6fTyh4AZUPoORkG/Wtj21PTzpI2Y7Oyf
LUgzhfdHFaZhLfPvzDjrao8Tc3bcZNR3nHrQPipEQNpnToRiFeojoNVppJXTYE5P
dMy/Zuu8Qav7BtLwVPQQpVwrUgYedggX4Hw5vycm6ICYonPTiiJoG0KZeyVtRgE7
Kb5LbkL95PRFvyD0LvuVhVL0JKxghBIT991lsaqMrFCL0295xKa66yfxiY1R80O4
4paQqebxNqMeOrdGh17WReMyyTVK05sU2rXjv+A+w40Ii1S7RPdpPAXDLdTdUJhk
dU6xiTlCPIpeopXzYJaXVSDI71wJyzCgyRw19zYWLzRWD+fdKBoululrQVm3Zgr6
saJ3fSSkeXsltHU64Mrn5EOXXCIuwojy0WyoDhBrb9fXIKA8pFNIs+lqIhtwaqcq
kSTz7XGIxVtxFkANEnSYZaixd+U+hoRvRVu+vF2am+lXzt6GSfZMkey8mq+oHFlb
MiUcoeVHiMF4rH8q6WQyN1tjijjA3VRn8C3VrMT2ovtdLprVj8/xu+bNK7A6Snfw
5wS9bCBpG6ZEjdZNZ4tgurRa8BlTaxCM32zPTpbLg97ILP1VvQXN1ee6AbkHwLlR
NSlURZ6POpcyp117Uk7+K8SWniXOgUOnrjVph6MEjO397kfUEacovyrcVMwBjZm6
PN+4kp1XkNsgW+aMvMDVdy2u2B2uApr8QYPm7WbCZizsPLw2bM9UBlvD/ikh2v8F
B2OKbWgqN0bIA/oUrFZ/hQh3LWS47XAjIffsDBDqi+GLgMGFtfMC0x5mSjiLqVf1
rUCuTbagxvYZ6BQiUYXNKSLutm7+1bkHCsVT9Q+Wavpstnd2rYo9mXVkzGa68UD9
93cIZYnWIaD5k0Y1qM0bOnPrnWoswC5+vVM+L8iI5Di8Q9HmAV/T6R1hoLipISSV
L4GlZyFMhivbhlgF0J62wTM9R5kIPWrDe4Y8w0dIFKs=
`pragma protect end_protected
