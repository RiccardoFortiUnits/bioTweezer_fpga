`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
S7Y8XL345pPJA2teiquDXtY0jAWM8Qh7I6IXYi8jvUtv+MlgPjKLeU9V90v9d6xY
8A2RT/CC9Qd+MeBqzLMNPcuOEvAz073jbR8DPI84yxxWiq3RI+M0rVN65UTL+dMS
UmLboJ7hTIh6YnCztrcbJVPBz1OIbbyKgWxthdatmlU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8400)
P5/qrnxFk7AIgm0sC/jUVWwr6VriV9aT3WEGN1feBiQjFMFZWBRvn9jJJM3DCOQb
el/Ksd1vSYAVA+QfIASmiVckQKzryg9DDon5vB0uhR6Sv2ercSb3fw9w2kw/1vEb
FgYQVIEZMMeFo5IKO6Iv0Hmv+zgo1WFtJFuaV06JO9w+nqrsOeOknV7olvninlBC
9fpkb/66wqRga3dhSz/d6OxB2KBo3UDesGauUFKSLZZf6yWepDTSEVmZZrbHFZ1k
hy8SELdzjCesFwmz/gB0XRdNejhMUS6EFkij/tmhGRWoaUBlzx/OWsj15gKO7sNJ
UkcHW2oMreCBQEL7ALrJMpqM25BWYzDXPnAFcEAueTgVHQTa/mHG9R/onAVGRW6M
yG2Rpc3jcwiYfBRf7AJQY0KJqdRjaadtPbAdtB0JZtaMMCcscDoogpZZSdJ38kPI
F1B8g6hMVWarETp0crd2coLr2ypFUWUoBzN6WVtIbR6ef8+2KlA7Kmv4Z4VJi58z
vGPTrKAmllGDIy/3B6R/UWVNAJZ5tQr0u9uJxF2ZnKgr0sGBCzm3nEYwND+6ciYw
4wPqXEOc/fImXzFhdF5sfEwKARgOB85ejfs2qLGlf6JQnUkxhfzOmvRb6w/aVzxH
6fLEUT0stw1vVea4n1Uk+Iiw7S1gLY5EhNa1HP7MjfSCiaHkvvnaHfNq28BIW1g4
/urmGXB5JxjHIAIU6iJOyODttNLCPAhLcL3cpNm2/iI8gi9YK5musLlGsVa8oGuI
mGYLx2q0udjcGR1hu59INDiEYMokKBvNDPFsI8xGVmFJCe9Hp8ZapMhZcID86uII
JYXetENqaKwzypLA2VPJggaQT8K6fR0AxrzVGn285RYkZiMRsnaJLgpY5KnGGfdY
DoSOtycWTBmaOFngElaMRcrOwJFHHKZopEUCaXFxGBE7vH7VeADp3BW0TW+WAUlJ
fqcfdR0i31zCVeRkZILKNZ/QfEi9NlUaQwEQWRLmwDEcAYveHez7bTFir5Cy01ew
zwjT1PXQQxTk2/kl1Fjbk8TUp0PFCuaN8c0N6HJQyTAQ/QI6Z44isGy0ZCc/LB92
J3DfYmiV7XYNVQUZeptDSl1F6PlSpQCvjBzm7UFZ59Luz0bYdG/gouuhzjVSqonM
YZDrQPAWEF1pFLfCDa6MbN92qRJMPsPmOj74Q4zaXoKDg8enm29fRRJO4Gc2zSaU
Wxf0BcHhZMY0ZsL9QAI8FN/wHuvqjwiKngO+e/CKKf5ltiMIcJdsid3pWDDXJANu
l6qTnvXkOg4kQZnek/GSaXoiBTIjyimo8kXDzNKGPXOTXVN2ESgDz7hp355gfbc4
T0YWYcnMSP4XCxq/t/DAHcgIbGWI+vij+hlDPfD/a2e9AxoFPGCr48ytpXZW3y6a
U0x1MsCZeTKjghSDCbo+CxpcmYKHxX2g3u2R1h0WQ82koT3BFSmn5LC5pb+yrQDb
avQAeuku+VoD7WNvdm7RJoqa2XKhAS0sv69eCVgEKTyYQtpnuEh7WTFxMdmvRS75
IAa7Nr5UXXPkKUx5PykSZbtl/vOlDO8InxTbIGISSnPzWuCbFpf1HMPEDuK7VZKA
OoeZgpdNQjQBJzln0muLnp+vtGP4zZBXS2G9BmxPxuLroQfI3TAdhumczSUU2aiq
VQ00OxAV2z3cjeGxjQ/u4eYhvVJLAB7qQoX5Dogeuuj+j1qqcOf+6DXZg+OSG4H6
bvLaZDUtOnw4tiTEHzd2MOFSufhuXnrVhkOTXqmUzHv+cT2uYb4Sb7Wp3KsWZpgT
18bONvbYNYal6QzJ2OG83sEDeaq0qXubY+BsqT/juQSKuu+sIgv2ZfItN0q+mDna
g3tJUBQs2z2I6aYug+E7Z9uxTfjMuWyiJCtq6UpEB6sw+X0B/G+d9PnQz+2Sk78u
wR83o0uS/l3S90GVnbMCR/yUSsA+NZuA8FD7VVihzhgjRCe8j28T7aOeHh0kWjay
xQF9eeOHTa1oAA3/foussc50Ha0Rzz6OXBmwmD3+oxPH93nIL+HS/teak3r8UVV5
pU7JImVckTojv0biY0o0nk5RmxSr3gWCGfgmgtFmLjyygMly/kPv4PvAGHd4Werr
TKvgegUQzYLPDuFFFuJDvyLII97PNxvwwrWhOPeWXqqmjCm0inMtjqXbkLq5zmrQ
MKp+Y6O2omJYh6P9vFKOwjvQIIhXd3aAkuvQL54yEUgTfp7FGciyO5gDrBe2TFal
F7Z6wiiKkRoWdLV/PHIUkuwqw5b+KvK+aZND3ITV8EL12OT/8VJ4KqU+sARQbZg1
Ft/xKBrFYyWYy+bYrxNzWp6w5ibNWvLirwhPfmyr9c4TbtiC5sPYEi98pXhCUzaX
hji5/S3s2kLInG+YzQ9QCdjbn+K148YNp0JiiH6Az+K9eyGUvLLZR3cgVVtPL4zN
68DhsqBQsbscERaWIsB0l5D0jtyqCW3bVxy2E51ewfxACY61z8vAqVgbdDnyPdn+
DL8djQOYZA0o/b+xhWNw2Bz33LR8KNjDwtDFG/0CxT9lbjqQpElw4Qf1/QMtVnLf
QWiYk8oG//ibhy8BEAw3hO0XfjCJeEwqx74Jl2lWmARVewc8JxS0X9PSgAwBmwmt
8xR2oVoZZWQfP8Cndo+YFBpZoGTv8wCZBVFPec8Pb/8W4ETQ+OiHsFX5/POKwz2O
Pc5Wxa42f5XjwZASRJ3BDR0YRgxXlZLl8EMIJX1pwZ7st0JF942M8TqHyRKiug9I
sq0ff9fV/rIEyTqBpOypEEg4gYCWskmW12zuPECxZN5g+IJYWQ4MjUmhnACBhZKi
uzWUhN1ZPmpHtIttLL7WciO2k2bcTwK0SQ7WUVSDzzT6Z42AqyhRLjICwo/D/s9k
qjTxXXONdDkMTA+MOMV8s4M3v1vBqOCtsksSHUHLV+lvi0wqMoOdg0FAWnfZ1RUv
eHcXmQYOHdX5GNOJkO1pnlcrX48VyqGrCI6oiZMqaH4NB0vOgXqs/3muvcjDP6s/
/WIkVO4BCC4NMxKbHgemqAmH2s1V9c2CdR5hswik4mR7+n15oZnBODiYHiavIfnM
HAYdSsoiHXGhrUd+FsQjJnIiwIo0Qux+5XDI17K44l4L1PRjT3DFughWIFe/k+Yq
F4lTmQ3n5tvUALhtUUusE+vlMMAWi+oUZZdle59c8BtdEODnN1mV1Fcg/vvzGBVV
2+h6mTTMjA8E3/7aKRLwZhnAItxcBikmvdn2XGWqe2wWEt9n127W6wSS2QjdQcSv
CvSzDnH281qNuYRg4q0CEa6c4Qbaa5aAPFMe4yeGMzfG2zOUALPkk/P+8ABH8JcV
C+qSbx8bsSTad7iWLfodt0+6bLyhf6a3Ga5+kQ8YsX0pQp8QR4g/e90diGgGocI5
iJq9yOtE+ZxVKBEuqBvvTr1PhaoJBzXOxG7nV7gnMEsLvCLlnGQ4xFFqxt7cb3ej
p4NtH56gfy/SvbodbGoHrHKCRb+38TyBwPfQiqKXEw9T5Q1GJBvNt6FpF5Io7d41
A188a9GQdIry8Vdd0FH4CQxsYqrkK0I7dblsdae3mglegXljTXtgq7smndDV/MQq
mW/XizxQVUXXxzikHhhH/cm1IniyxRAJt9dyZnMRIM798gm8+yTHvOa/dNdg+nDL
zq4emNjXbJi3Gs3eo0UeBsq8RCRHfc794+921eNF0NAFaTZ7mRHZBLtlMu4ct9wu
zf+GIfmg4y+SBUh5FhL5F1Aoypo1AnXxhQ4g/zt5rpMzEV1jkslpMAGY2/xXydKK
cjsvNcSBjStabyrCN+dLwEsE8Z1l3GVTMrt3CxwdlEWDQJByR0r7P3pkt7PfG9fz
zdXx5/l7w84JLvNhWosq8tn2Jfz1CDWZ0lZImOFONCpa9NxJCY+4vL+LlefXs+rl
g1oxetxVedBaqP4oKwA6UwsIHSJfadVegWLCW6KGODuR0XEsuFpVtxSWMN0xIeSW
UBgxBJdTRo6y2u6BTlhH7T08SbBnbSb87WKYNGvmqtrs0XBK8KeBBQu0TAZiTPtd
TVS8tMVsS0PIcCKO4UDSxh5x+CT77jFOKARUpJsdypyGles6w6jTgEUV9dUBk059
0gBSkpolyKGlHa8m7BVzDq3+239KJAIB+2XtW8GPVQUEk5ZS8EK4C3yffHp60r9F
YhA5GWccXnLaMkts2DY5JEw08KGKhpgNcXkyhiTAd7z+//5xVnvluhd8DiJItlPE
tvV0lk6Vu5JAD9kd3fBCsmFDIg6DM9M4/jYRztVWwPcLy2ZExU53k5GrS9tOZtai
+FgNr8q0dSwcYE7qmvIg4L6PdOxoCiry9ocngUM41JVS/s/Q96Iyq7YmzmWolTIO
dwYGAItgxcPHPGz7SqQsPS59ruA4YH0LmnCt++TEN5rMpeUQxIWxQGTr+c+voPvq
X7Z8U48atVIG3xGw78JISLBG9ivRMv6zTCbtBVYXLXxX770SkTlx2aTbTs6TsFQz
h64xie+OIWzpyell3nZqd/XYqXYJbbV7uXCB1gGZwfcxSnrDN1l0zMU+eQo0LDcj
lCi5/U6n8xDJajd3mABffHkwI2DCzQTTOlsSdb7eTQBh4LiPZ95pwqCetknGymkE
aIoknkEOuMcemgMuYBMIhHcYOO7s8xllbijkYHY9KQrkY8rn35tbq5sR9LEKmIbq
n9cf2bdnmKfeB2L3J7+aaVEj+zLPSAicgBZ3bFt8eNMIfTKualteMo8AmvnKexTQ
RxoOPQf6C+UeOmARSlHxo9OaFYMOkECatr/kVnViL6guY+VJZZnz3gH3ii5DvFqE
xjJ+7VBCvYjCayA1RTWP7HL1NLZ5lqaUkScyOI1EZlI4QtFX9PIOO0a+K8SyydGF
0Av7pAVKMsYWPqz4M5D6PCFej4/GzjhJMsFkgF9zS+0jND3H3d32DgKZyy9xUMCY
/ZW2gcfu+qKQ5L7cK4zPBPX/lVD2r7fv7S0pW/bJi5fdWpCEgRsmukbhThY67Dqe
r1pyK6nTfRgGwz//u1Mfb2w+Xqum6nhJRnLLZFPawzGvm7IYbM4+1RDkFbkkn3g4
8U+zojDy9zQN8nPI9ZzhCJ9xbCKfWco4sGQ7nA/29mM6MsSPa7FFEni+ww/DiTbb
ovaOFV+F7FhayWXD5yyA5J9LeKKc6j2JImm7UOFKXTEIeazyBB3NssVfXPB8zY5U
5RE6ND4FRGhmlpz1njFijlRjTHBUB6cDAeBAA22gtu7NYAY904lq07fkA4xXpslZ
klSnc5WOz1Z3liZ7Igj9bjWVTgAI9AZAImdZoDyKlR9VYD81Fx+JatHPiVU72obL
qqwp6PnPf0OAQf0M7QGGhd0rYxzpZMQzFt6PMEISm2qfdJth52GljN8hRuX10Hgz
HYM3FkJjPOX42lAm6oSOCTW86gHf7SoP7KgDfX1qokyqLQGF+XyrlX2JXN/9CV5X
qooFb5W7Dcq32m+cV/gapzCw8QVefZlv6dKhiE7fMgl55b8QcWyfrmLs5CArMh0g
9XG9lNj3WtGZwktjQaOZHSI1+d6zsHaaL733N9BtKmcaNtrEARW4m+macDrBUrdH
TTDTTXe85gaW7QddyWQIDG0duTui/EnEvEm3T9KPpDLUaJ3nz6HHd9HPYhnmUNN1
SGS2YXvJM27k8F4khfrpkPzc3VOkGDVB6jzT0t+5qQnVbE3IrLllwUtHYxw0cJKl
6WEU80XBzYp4Y/XoF1BhcGVnIqmQ6pCuaxSc/qPjUCsZc3ZS7J+LtKVm4eoDYxl2
C1sLyoY2Zp1f5LsTrGigEdZe7GL8CDHWtI2j0MJHqlE9FTP2U6yTVfI4pcZtEHn4
Ha4NUovIGc9+kTmqbyVTXIt0mXJBAdLbTk9igyJ2dGE49Yd5NhmQgIUqdjscH3h2
mbGQovC//rL35ftIy5jIAdabK0ZDK+vqmlbNfQ2jD+h7ORgNEcJN6e+hWiJKkNeo
uVWMiSNFnzNWl9qtYtzdNJ6kusl5YXnwpQgTv5QayjKMe8b64Fj5vsY351VFy3Xc
YwluyZdqlgLjrFV6/BS1aeyqRXcWew/nGIBu6bFrpU79sTVtae4WzswsYLpxOYVP
ngsbcn+4+GHUyPrXPSUfLQgW8gFywNofQPtRGWv0EA7XnHpywJ69Pn9TwYL+VAAJ
5nOUD80ccS5W+eT8XFayYNKbhN8w0WGiargIIXwbYEel6eO0hlHX1IZ5NVlvDfnE
9nqPUAbPTwJGcKw7XOGEM6OdOCUVKD31ioKm885ObQHf0FwkE/QIRymQLS97HgK+
ejQrU32gLMl+EyrYbS6CMn3EbV/m/ope3YFgf74blapMfPpbfSEyk0tZ+PCKSqlr
NS4+0CtXd+TDg5Y2jLaGER1QH5BnQBPhKtHpDHS2VBi9WH8qaEh0KrqGZFrGbseZ
EJx4ajMDkwhjnx+4NvV0pkgI00g4wbDmvdIFW8FBlUlsrgoKDvJuanF5g8g0/JiV
gXc1n8eo7Ua1f3gn/FR/LqRwUTfGWqpTWhuJTu+AnOwqkcN22mfdH0QnjvKDJZET
1XlaXomnkem45OlYU+Q0+bHgVAJrmWIX2Vv514z471MIL5mKSGjT3wPEJg2K8/V2
voezCjJ0aL0mBxGnhkVpFqeXjrOemTFUaCRH8VNxH9e4BAZkF5au8pIjLKGZJ2Tf
MQqlDyXZYhAS/AcR8cT9G7ru43jWxfXYihk1ldKNuFexMVGxrhgiHB8PGV12aFAS
0iaCItqrG6xZt9/aYtbrVqtIpdkDArLOaGkAFZfcPT0ZFcNRQNa9A83tWKjzLkSz
kTQbOfnB5LK1O/47EXCofGUSeFaM9BXJMt8e/RPjBsBgZr7YKmDb3EB4HpAiBlXf
YcaF2z4WY43+uI+RmcsW16Gx4LQglJFl37NoAcg2eUQPJxVo+PZgUtWiUsTxH0vQ
iJOoKw0mGnFZ+SnTx+Qi0B1F2KJ0hV4c4h+aUir9/EMHkXPokg+ZtRrQX3UPznYe
ccKjQH4ySZKhvX2sFzSPf3RFVZAIE61oPY65i59HBe+VPvg5ymyLsPldChIZCX/K
hg1QIeul6sRI28Zc5MJnhF5ThBsGWh7wkb/pIpykvCPDOwNmyWKxl1tKUY24dNk8
ZU/EIenduJY8iHAAZjZTe6fTEJOWK4HdfOOIbyf44hW2nyqqUf0aoevkatE8QZ1o
qLnUGDLzIiPaRpDmgiNbJx+4RoCQmrE9sTpjXqP41HE5PIudNTUVzgZls3ilof7e
RBX3tJ6ODFRGvQIxl3T3dU4FHoGA5iIaodAH4FC/0DOUXQEUoQmafVEXIxUfb240
w4XZbIX/aGUMWblYKzIY2sHIUpItx4Srd4vs8lT7fJufQ0XWD20gl6TfhAJOrzTo
MaqL8vO84M4cZq1mlYAyL9abjEooOxrxY8UvGLJCNJjnMduwIFg0ObSug46uP2sG
ppuXDvpFbEKlRBMeoqL/Vmvz3mpkjx2nGm/7/cRGpLGBVZO5k7Cnl50pvm2hmQCT
Cdbe/dZ8+MDQPgBbvb8YHkJR+zdL5ClY7vNkWYXxNPvz3k+NtBYuQI6FLpC2jidR
K7ylqqnyRE6qdDrPorYX21RrUnKt7PYp77QlkmFesIgEu3Vgyw8Qr4A3N+qzbqYQ
BLV2sMoihnICdvJsqMBM/4WdiGfd1DBIyUpCpcxYn1NwKqNAkOUdv5V1vPKL2VDe
a/S2SWa5e2ZQtuEwLX6cCJSKRoBoOg3HYSg9z3h++WS4mb4BQ+nGgESXj8TZhKSC
zCKJmEaFx7PwWAHZZBIgnUR+te+FlMwGHJMf5jnrbyDkrSD9pthTX3srFNClWCvw
cMwT0eftRnn4RXEp/EvJEwHg4lfHzzbSbbvmsSiT5qkAiAtP2fpi5QJZkpNEEbFS
2guDFRoxtxwzR+BlfWQZSLwxZbme86SvIWm0R5jfn54lG/Xarc1bL8MELl9jJD4A
QQmiweo2ZswSQab+A0RqrfeAOVi3lCCMQBY5zBSGGyV6jwmJo6H5CAW9Zr/z0jIa
Bt9rzl/0n1xCZ0uWlWl/pEA/xc7yS0HB9/VxRqYEs+hSVM9TK/nL1PDcS5oiYoet
P6oDxksk/qJtaHhVkG4jrTrqI+ELi1o0Vimou7hr9vDtdL0Ei2EeZZxQqi/nzTZ4
yco8hSswdF52KX5Hjp7XNhUeNAb5xzTFz7tpyYRKtoxaowan/qhqrKIcCzkngI4h
a7un8gNPTzVkKymj4dgOdMKsS8RCkqmHYyRwhZ5c3m0B7mtTDE94QUmqEIRx6P46
poCk/UqYgzxxHJd1iNI/O8Y/REScIHV/lAd+upNOCUj4Mi/tzvefK0RDz3bWV8kv
Li1ex5VuqvQ1q/2lfmes65SlLVeHgBV+r2CEBTtKG861dwL34/i43YzzKz0DG774
Ib+f9TSN+5ZP4ueOnCSy9o6zVMWOPllnSahsJBid5BuG+m04Rdnrj3udYGIDgbS0
+hzysAQlf+XPbvqBJHhW9xTZNWLYBXynmB0hTXOCdqRMBV/Olgxh8mzz6VdgPAs1
upvS8piIEK/aJgx9/UW5pg+3VzJ0ZTs+NqYdmrwLfxM0VtfmZuMwdXyUcvqqiKU2
grMDTA16T3eVnvS9ldA+5EcHEEDXVfKZW+mc3AYUzcVlECPVbfQoaLoJWR7WI+1T
ohJvXw9a78kw9Hf6E/cfPSj1kucenav+kbpSoZQFCAQs+47KA8s64LryUs2hG6K9
Yn6EneuOkr6GRP9WIx4gICpiCtd6eTJmoHpU0zEY78znlve8FkWMfoO+753KsLf0
nIGV55rjmpmLNww1zhBBBszZ4MgMa6hLHtGFpDKrkGsiCLSbaaLgTyzLpJHJH6we
y3+47puxN7UFf356ZQ10ux5IKPDLOg1sRf1bOi1jOKY2JwUkwTISPeVGIYIuIEsd
fM/DV6hxD0XG47WAhzVY+TvoBKtFbUUggxW7+eMvugPc0zoekaHq7aJOsSs+B2Ui
TPlMQlF8e/IXMkjgGJF0j7EpxyPy2v11swK9USMTQbP+NpXn64X5okzCw8j9lYuV
VJSkVbK3gQ9R3sxTBtIKG1lRtNCGaJX5gPfXn1s64J/43zf9OqsxisA6yrqCiaOt
WScjYoa4/hEbNgPYMFMMHepbV91T4vKaSXDzLs1SN5q5dn4rP7RWATP+CmIzuJkf
jQvhHCTTctkd70uNc/Yu6S6dEDkWF/1zqsO8x9VGEeCYDlbKSC/LK0XdEs/N1irK
hCyh8YYe/hQQm9BCO5P/tbBXhvF8FFNrLNBH3SjLUy8CXiKjW3tyTAS068X2Hfjt
CjUsFUr9CBVm+lD+PFPRFw4J6NarE1jDwfJcFxhJlmUompcEepG/IvlCeo12Pqql
jL+4UQHCLTo4uPteKS0XCccn/AxNe+ZyaV8S+ueX0SBGHh6Rfu+ot/riIq0QOgdO
OLUVBTZ0b4wfwNRXB16khrFgycuwK/1ozIns6g+5rUrdNNlsdTCB984apPBDu/ZN
sm+drroM2UvrOAtx2PMeoso4055KlD863/gNJD5a9Z3DGAgmEXPfSSQD6pTSO+k7
Gk8h4lppwWilwyjZrOJdMxg0kFEJ+goQy7cOEj2GfGyftZwym9cpgopgosHrwaWd
YpeHVFUsQk1dAxNqOV5mYCAM7WBKYigRjqw+83if9jmzPRdAXaZX4s+G4lg3xnDe
oUePWgyO3eQ7a7Yrk4PATrxaPkEj+ZQJ/z5gCgT/7kU/I7C8JF9WkD+GQ+NTZMrx
kZzbRI9wCt+3rMyFlPo3svgVAAQYOFhxRF6GXJDbntF1iUWXeVnMqwrZCrXchsUN
h2hvHLWvnwTA6LSO/W8hZjxScKLm1E6nXBlEo1S9ESGpmOcQcNSYtniqfFFVjis1
XSda+3aFyHz/LCqF+TzMXLLE+L/3fV/mANyuRZzS7cgcyig8jSQHU7u4HWxrB9a+
z8neUKTcWnTQONpjaqXB1/YjmKqJkYJP+fzCSklVLNOSrDiBBCyYga3HXqxtuKvI
j49ClOCQKCkQPl+4uoGd5Oo0peCuEOrm0yJRBNx/accA+RPIvY6k7oUMyR+QhbFq
fduOfuCYyOYOOPAzp3bCuGqVo7Elr/KtzIhFGDjsd5XUaNvBDsYjD41oHp2LcKaR
1ld4wSOvd5jVzAclEX4Vi5WFfADCUS5D4VbAwohKSnGwOLwXm2PcQ/Hv3O5TcwOD
GPTVoD7H710zJ0MzVYFRe1MeZ0qznIFg4ioFScCQAv7kNVG6JsvXh9b1q1rxYpXm
YdQTs/nI2nYcCpoNyDcepnHzmlt+1icOdw4zSMShJ0zauiqDNlVlWS0lgszGqksq
doKoS2pVIdVvlBkY/y2CPCerbt4+Dc3S5dtRPbDQXOPuSomBiwFxRNtcsynWD37A
biZmMigpCg/se/IddQ2fvvqKgKehSgFuV9yNVPIFRrQngPlalCHd8FkSwMNC4gb2
66A9/4Na3pNaVN11FYZl+QCf1r8XYiGJfBBrMUPUZcSjR4e3eWbnVIVUtX2CjhUz
fXbnQWbsNH9O4jTYkqIANI8Q47gfhCHaEVJTYonNeacw6yXjJ0FngBLIkaV7Q4IS
XMxmclh0ZU2Qj46Dno8vhFdeml7mjGV758vJsI63T0Tpah0x91wqJ88ubW9JaPx7
D+xDwAOgmPzL4IKbd+M9HJnDN3Ghtpa995We4bYjfwZ8jBHCZCa0zOmL8Q+ERqAl
A6l/QH2bs4oZ9FVs1b7u6ucyhoE0FKkAawsBCPKeeSCWjQIfVqYbTBwAhORmyOP4
RWxhcoXrCp/z57z4lz0qj5ssc1fQKKQdGN+br9LdGXw5LdmLmqs6O3qRYAodXjlN
wAZfROQSPq4V9c4TxVImCnHeJa3AEwZLqj6hsb3cIAf/qa3luUMrkgfwc8nbqjbY
4zhpWpAtCvwGJtQK7cZ68Gns1jePDCTfpJLbsoXBltColGApr2sZsoVkw9j5unXp
NKIJygRqsz2HHcQouwXC0uwx1s076PlfZIaahxSyIXlB/dqQ81/LkpdipcT5+xTe
SpnexQdlmuNEApRt57ujT2CZSHUvaFW+UuN4CrB7TYMIYMGI70ovIopsCguaSt0y
pNqaWdEBk3wV/MDdLhf9oi/KN88dScWtCzOYEnNGTiRtRSTu02PuYQ0JN5vtf6KZ
p9+2vB4pN5WMCGl6IWfWsv7fl0kqr0tFdsZdHTqaDtSwby5VmS7189sfjA/IovNG
`pragma protect end_protected
