-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xY0TMEE7keu7C3QN5f+d89TO/7PG4Bfek3V1gE/x8wrmSisY/kZ5at7if1NAbQ/EXx2pj1BuGcZ2
Bl2YseTt857ycX3qzaZChS8Z6AX0j5AQsYiFV+hECsawCIumOyX4nV9VSyl3bcoAOwxSfU0U1S6m
PjnFoRqVduJFKyLeBoTwzMykQd9RfSv/jBktWBTJLsNdNSaonvw335CYpCe/UsZgDYttGJEXMNr3
Pg6jkxMgkSM0dyU4EXJX30CER4uaeWt+Ugjx9HgkAQPSZilHxZJZQJVC/AxbbJ1QuUW9aTv7SwzL
/trDxm3WV0LtMSDQbllVIQACC7FixGINkUy+iQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3616)
`protect data_block
eXPSsgqL3mPWAg5YatMolfPzh0/knTkUPVwwHl1bMsqA50DZp8bG8J1jk/YsLbFXUra6BxIJFJjd
agWlh/Cdw26LyWVymH1vgoaeLQjOsaHCrIH4O6l74s2R51+HDmx43YF3ENcviaIojGzzPg9xptSq
47JtmJ3ADmbD2DKFiYhV7R0U08fvR2Ce1/vYcb417ySHnWDv75TybGq/m2+OFagvEI1Em7OAouqL
8+3rw3iXaliU15SNJ8A0TKtNs2Qka+cD3Tb1zrJ/OHunibUNIRPOrx2KhIUOL6Yc9Dat++rTSch7
q0xDva4yVHa9TIg1lujhkCutDebpxBHnVlRgbmD80FamDG7ZYVVQOF5XU57L+jnmaXeRT9JG97uS
FmUQV/bnIzvcvJ5InQt33SrS65OVx5XOOeNdVAVBnESEHpDwaiVHMsf2iU8uDJ4y5e4hJjawEj32
2jF4w9zH6+QKI97zIhYZYsJ9hsJ1CyboMtRA3hcJuV3bMa1heldqN/Xf4B7ROGGbtO89oxfq/19P
XtByE4Ixq3/1GVG6qLF4of/3y3Xby9e4QK3xuIvk6P5AmpHm0llpwVB/kfvO9HaAeVFfHS5E3mZ9
QVM5qKXX5heOGbYKyc20uKyPpGyeYpti5xvf5MqZcP9z5I2/qBqIvNy4B9NUaKtnjyDvkKsM7ix4
NRRJd22YXTyKqAye7RpRNklSrUn1tDp0is7RSYbZtplGJEYSl0jGaQjj1p0NBdsrf0LKaFDmYGlL
UnTjVThDt3dM2W1sGym+MmeYOn9wWgOMm9F8AniDFV7VOtwWqG0y4p8Fo5oIQICVxGdQVixy/Qnd
E/CESQFeQz4pFHBp4jEdhhTeiHaaUHWBfIYPgNMqQp+FHAfg9HFk9JveQAH0J0rMQ3NM2+N/oH6b
0EsWrGPcwKzvbFGMNxv7CeFEs4DQzf6ZI4U/5axram9G+5EywrqJ5PVZrVAfG77aHHGMP6Ishsit
kWJYiK/OWGN9kNd+Bkyt21MnG+Z/oluuB4DAjyE91Rs9oE8kmRPMJgCJenc+6J5FIRWy3ogkomTN
Ft6d31Ck8JKoDcvWXXClYPmQw6bZkfbm/m921mDYNl44PRs8R+W9+xr01XKfygkZ7CY8j4RQvej1
Sfep5hs+kKaBvCkbU4EdIdn1GqiyBi/VTeK3GNpa5x5HzUeaMXc9z57aA/1hST+LFBnWvFH34XBz
xW3ob5oQymIF7USjSjGW3KBhdT2sHMbRKGGtO3slslb0yI4IN+HQ94m2NoN5ChlmiLhA1ghiAjJK
x4tujwTx39sAcLyugytgyTTas+xkawi3vdQEhM/uu3Ls+TTOAVzHf8OhfibshFRaobxEAM03LonV
B7leLf1zAX3RNNGd0mWViAfmbLLpR3RGz2yjN+1Ph4wbZITSvBHTLK01gjz5cJUka57uccG3hF+L
GFXBZwqK/Tav3psCSpkfW7VrOTuDYAGkDLfqOwZ/EXzvML6mSV/s0vHVGPp8ZevREUZIwT/cRvn9
lEEjGFaaPQJLge0lRQEkUM/mb6ZO0+RwzttExDJn/sO7yq0jU52jnS53Tn56AZd2OEcM87NINfum
Wr7XWcjbRDiYpkRJu3QMmBrUqOcNVoA323knVosQn5Pv6C8TsRf0+O6UHdtVk45nXMSNs0juSMic
la9ubBpgI+psO1QJCPDeXQa8iFwYRq1+imeIjve9XF0cHfb00oK4uGzif9jH1pmnny5C9V0a6e2f
pCFXtYqz9TiaMtT10F3GgNATTH3U8nET3SYO2yH4N3jluThW6MkfXnii2H30veyoufyX7i6ugR0Y
5tekAZ6K0augAAKo6yDakBrNU3ghDRm3zoJUinzn2Go3YStTyCLfsPzoBThkuSMrhEo6cTSJj7HQ
DiqsPazFhzPGNSoX+MqL5GT3L5HK66Qw/JfPhNfx45dCF/fEBfLbTnV8l+RdMJt4akw6QlINahkU
umNek3N8zybCbCDmBoCo1rN2WWzeu7Y1Fn/8p5ZvkMOUHg3R838+WJBr/N10FL/Oxfzq6bfPQEk6
Z1rFQ1kzB0cAWtIRThG6Tl7QNlsCKEaPNwCjjOPe1SudIrwV78PLnUP6iBwW7aaaBFHTtV48geva
5v2NxYhvc34X5TkhtTdRSUvlinsX0C+cQ6VnkuJdHTlSiGG3u88hgLLbhsh86yB8CojySR0W5mIO
TECUjli1UM9Q+FPc15YZafu4okCk9xZGbv2gW2hqnz+Fo8u24t8S5sRclY4ANFQdnlK/Vs9Crg4G
nmq/N5DnE+5sDsziIr/+P/jFTXgrsAk1Tni1H04oexQkXcXAnTvUyzydmxGZ8S+7keKQ5E25JAxT
01sJgo2RDYRJZYBJsgzbhOEsUwqkh9YYF8lyxfAgim6mWiqIWrdN0nMn0TL9ZPlqqBrekacj9vnL
s9zZZNgcxN5neNQneB5KUxF1PBDJzrM2AP5RcoMNIlfB5t+9DwaxNfCEp/arJekM4ySyibE6oSUr
FAyfbXdVfiKZOo92EQ37GFG2e1T2IstxZxcXQrZiBCaTJZtqplbimMy+Q10eMzlQa/JJKcrhYmr4
+WKn+vZnGRX/ez20eWvHN04JEIkrnPiHaWhelNAyiHzYYEvZnZHKfr5LCCF6H0Xe4oyEN1EzVLjC
fc9ON9Yeil9FxdlxaSKkASLuFFzGa48kBHdbTcnXI5xX2yswZjn7JOotm1oxge28xdExavqimr2K
3vl0PeihTvSePsRRB8hcX0fDLj23XgnZVciZX1Msvq5KKW+y1l3xe2+wqVWLLvvYyTtDa1HIDcht
gRKk/k/Oha5/6luj6OTJ8xIOSVxw0+IkzPP8T6xKZcXC2rPW3tKDmJyD+nG+T0BnHhI+8WS74Bdt
/ggfDleaX30e+t6VuGL5Pv2yOch66MLPbN4BxEn4ZBMmoCO1uXMoU04drA/yB8ejTVVgfK9MMBQ+
5YpCgiJeSebQPGYjp6OoFgLSy1ika/zbW3MWJo9J8S3nhVZ1i8IahYbln7+QCXmlejKQIy3TZ57x
UOgU2rVFsVcPtjJewvI+xhC+0Ge+v+ntEJ0ZO2ujlGDcxCOS7thfv69rgwGjmSh56KBSlmHxfSvZ
v4/4doYXGnFYSuCcrBLNJIIEjvsG3mhmVAVEMSBTdBBl99W9Ut+Q0+VrqGiO11/8D+ygy98Bbjk4
6r747sTOpBawKmP9YF2ledY4N3t2MBk2cyMLSbVxoZyx8ekrWR8x/nbpLgnrd56od4BHTPUSu0mF
p/SgcF1D7PJdEIETn9EqzpXGgIcAwRuSjI/Jcgj8B/vQrvhP5uluhlAtb5Jutu+zGuzl6GMuSyPT
/bXSa0OO2g+FVmTThZ9R0D8iMh/qAP9UlXsAYR7uGEz/zoZ9WIQH8IlfAOvQRIkSC5+eEJlIKMRC
uK8aVHCp0EZs+30IIzJbioQci3zm9Dk57CcVfyi6sAAHe+Tw56ARrVbXVO62qfsWjeudt4fsWeJX
VDS4Plp2SZ7s9YisD0tcRfvV9yDNuv+RkyBYOW/K3Vhi3kNinnuF9e9jgcHrJFa774Uulb9o1vzv
OlXBOGvLX8A0F354HtHwhAfgCxZBoPXLT6d3G75v6aQqJIow1AaXTx5LXT2TTF0bjiEX2GVKpEeI
TKYCldR3FLVekXNoK0Rpy21NunG7SzDyrO4a4bgZcdQtdhxG75+MBBEHQGALh0bSVyaAYni8tIqf
gi9+Mn0KqIKncVNU3AnLLlDsJZ25MSMKKhdjX71jwNIBgoETu74dNEsE23jyuwVVEBhfZxEwYZln
ns46Nm1qCPHenbb6jzmwMRTT7hzGR24bZQ+9JfFKG5CReLkW6pYkOH1D4oO8kQqAo8uhn0jDwe8o
e+UK6/bcSdN1HtUag/deE3HhYMlWr8pccwo7F0j3P0ZEKJIBfuwLopoKHUwVU8y6HYUH3iFO0LNA
f9p/z4cLpNNqG7yxr+yV2Je4XMyxrQKJd2VuKdxY8L/HAt2FpeEC55dI02DfWIZ5ao/SESSlxy4U
nyLYRpZL43vRp78VfIGKOId+qCZYhyhsdhw5gYFcuafJSTJ5mGj3tvp4QorVzdLy2KAvOJ4OZz6M
q2H0qurNUPAvrpiCjmbRRIfm8Ibs0DU1hGZjvL5XSkuiP/l8huAG5O/E1exKURTfXtf0zTwmq3OI
drgZWNbu40+fgylyB2TrQAE7Y/FB03aOey07vdhqnPyfbK3RlL7sZBA/vdHPo8rsNEduiiid3BQb
KczcDp61JAFkMDECuil1xuK5ltYGaQ/TU1pQm3VaCxzAJnQDeCtCepWAqUe/i4wjISgB2uvkO+sm
lihkTQ/USCI5z+xikbxhcbLljXZFbwF4OuicYeB1qCuxFLrIYsyRWAAvPKdetZBVoBtNJ81YKt6M
R+/zmr1xISdlcsDWNcfsk/TdNed/MGiE0K/m8+XuvtgqleNR0N9dlhvBHYoySZSdE1v0SUD/URGy
2xYXuIUih6AHgfIovUQN0t/9vL66yooEydRLTptvBUk/y13uW3APpUGhEeJjCB47GsFKNqLevRyP
q8hyMR8q5hQU4BwJ0CbJW4lUlT6/0ev1/gkNA4IXdFPgLwGWlwZRqtmZV/nWtw9dJ7WB/uSc+zaR
OMU9l2BM872+FuA5xuWXSVn2dg3NMLNxFMfWo9aOQVkdqGnu3M2Ls2X29fbdlbUB22tcuVWkBrgm
qabWSUC2DC0GdHlOKYtr6JPEa+cQudo+1314Vf3Ut+L0/xt+mUgvbUbgU6Hhh4WeB0Ra/CAsh/bF
7CkP7E98cv4GjpGJ8iRP4Pe7UFY8Va0YRA==
`protect end_protected
