// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
k4/wg6rATQXg738jTzwdb/qhBTat++oIe103SlMgXkxCC0L6P0n7EeUChl2Wc4SUAiN29WaMkwd9
fbfNJzEZIj6M/Wr0Su0lF92NdWso0T3HzwM0e2S4RF1sTHsmwXtYbg50+/q6H9kQDJ6FFvoXcR7q
Zxz7mNfw/DkGXQKPmcFlrfZhnAgXGJkoRJ4LSa0UbanQOaugIAtuYdWFezWi9SETv0GrdjEKt99p
7pR86W+UQYBUW9FsskMklMq2JRPFbSsv+1r2WVjIHnwpo8y2nJXVgUq/wItves5fh1xyXb9pYiPF
XUTc+vDYsoiELy/OIRAw2AbQJ9FcsUK3kauPsg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9440)
JUdi5qHYtOj+2CyyeB4ntO5wtmYwAFraX946sidYjIwmCa8kebVUs/kXdo2ed7sFJAgM+TlSQFg0
0cF4TkS/tHtUoGIiQxkhCeA4gJ0R1B8P1AD+OXjd2x49gbnpISsaMvY5smrG1lY/nxqPlfJOT22N
kjXWIdMp8JkRM91G2riVIeurzbJSQS0iVQFCC0n0MRmZvdamcnKE3BqWzdL4YcXLz9EB0LGcdtfa
oKn/NjVnJORfWotjUJlHNYRlVluoMwHsz9Ws+EFGIwvzNe2MPZm0h1rR+rpYbwnnmKluOLQF3doq
rTrLsaiY3sbClpBE4WWSWx5ifcpkhIZHc6n3stko9MqWOyEFDITTWDX/wSJ/QXuyQdNMdshUTsam
xIy4uT8K5wPwPf0trKOi2S6DoqVti2JW/6/se8i7H3BCXufFBslDfdbyVyniA1oinCIRmrDT+fmD
2R6OZMBvtv15wc0i1tQLLP4DwFsu6+VWDXdVIZHkfSO1ewpVo4beG9FZMg++eDv4yBZVeICIvfiL
u4chxpuvtr7UAqiHk/xaO8QVWBg/wX+usIXDeswyP+ho6pAIBjWbS5gMH+rRiTdmN+ud9xFFCva1
6tpi84yhtakB6WWdg99/08tq8ENEfknNH5DmEhl6VqYJ5WzA59SBrB5IFblO1bReBpIJKtul6Z/8
pbfKVDqmw1/OkbovO0SbURisajCfRP697Ch2ryJNjHjDveh0Fwistg0geebUQRb04YmOsj7hzj1u
HKyo4pnDgUAexHcpscSZnb5JOTtBHF0+Wngr/WTVI8w1WupTQSe8oiLL6QLUdicP8Tp+ushWY/Zt
njCkunxJxYaKkHtxeb7Ms1yAkijWIBjxyb9RReq5kGUZCijEkyK7LgVgbRr/iXBJRky2pVeLC6ym
QYR5yWI+GT3SlPiAokpPDJAe7Rrjzhpz+uMz8cIAiI91cEQmyDZ/UVEIz80DYXp5Qw0RRi48fsoJ
YNOEyhrurBGiKD11NfyHuHJdyV4OHCfIXViqiBJyygmW+w7w12m8x4p0SHVVpi3jqNUY9U5b0rDY
LSW/yHw72418M1JTAWbQNr3gQ/V/JnkDRZqCdSmTxHnKr9ktWqDT9XKxhEfH5H6TrSMnolmsMZVC
hhmgIHewbLnHRxMscE0UzKeJl/8qaiLubF+p7vad5W0uA3uib+HWVXeTUr6J3PnbQYpxH4XVsBLu
txNmFg1wBBZqQ94QvDwHPUYZ+LziIGNtcH/lWcdAy0tDkp+6ah2QzfSmh6jP8O3x1JkLbs01pxer
/DxqANyYzBF+oG8bl5zGQ/PPqG+cOgvhmMsysp3KZTFgX1zCRFem/zddkfCmJFgHjSvG3rDlRZqx
eKibGVY6Lt/8xkhy6i9pGFPoIc4qtDE3oTYOQVv/IkW+jxu1YDHwZqIeU9uiKOTxACrAxPlKZoZ8
7Q5NiT0k+Qz4irLvkQwYjeU6scpM03MGoyJF8Lefi8Byru6fs4qahOHcztAL2IMEHodW5MYHl0F+
mUiQR01UVSi5MBm8GNkwSkb0e4KnO2S+Kf8P4Or/bljhqiwjLR8kry58umph0JpsmISW++VoWYwH
JBCfX4NRJaIzkND7Rr2deMaGBqma88F8O/RDpbGOzB+L6HePUckRtbkIxt7vCoBGROZE0v2EtNKu
rbpcOgMuvYct4TNWt0dIw89DVbxoGCuuh9aUnC4irnowZ0dN8v+gc38DEsQGABOQ1ONL6XqrrhU1
6ucV3k54JqGjjn2K8WWPzDvw9b0/rBkqBwaUkvybN+o7GUsaDIpaICE7Bl/ODlBKqOL/ExjNq1oy
vHEF1tMD9wU++fFz6XiWT5BXNkWGCd9Rk5UG5Q+yzblmacLsjctJPJfHJxbvm3fALNnL3ctZyaY2
cWdlnFCZl17MKhnHodzgyGjXn9KiLbiHdSkbSBg0jWJ0SltqHnjOBwtPN9fbsbHGhZ0ODrMvco7b
AqOkAF8mUyLYKp55WsjFdnWoJ5TrkO8bymz686TT5cEDFWD25ETuz+MZUmum3xfZ9CNZxlg7DWOM
u2kR8F8a+cuAtj5jHzMMA/OfpMx6bSCatPeK2QBMtz6/miRjyktcTqaN0rLdZvbloTY5FD9fjQ8u
PfWkpRQ5huvpkzVlAALnJlRhqAZYNV6OPbYEeOVojHOScDAYhW7Ny1AuIvh7xEeT92n+ZXejdlGi
Rfssc57dVirxuWSevPonihTIb04+hjU+OsvkVARfAYLmoX7c/eztDqXK1UWk5uYiZm7VaYvUjTMh
kUa8dVjdBWhXXUiRfWYENmO27LZ3STUJ51A++A3F0A13AQrR0kJArCCztl/ixqfs0LhlW6/iuQ9K
Eg6j9xQOuNctNBvSmgQNMUByO5KTC76ZYpVq8XqEoUzgoxGNquT7O057EVk5asA9oiSd8Yxz1tHc
tHLhb5Ax5LY4Jg9qFSjYhWTt7sg/hT72Qx2cWGTHukbkxdkwhMo0XPzl/AcjmzjOzXwbAhNJaRo3
nXueahwg3AOJ15smoD5DVnQbHIo990ZnHOFMadvYqzUBcIVDH/tkpq+gToLOcj0++HAuB1YVxrhg
lS/mlD+hNHkMNH5L2tKPJekAi2rMLNirpEFeB8rKSomNI8EnSPXbRIzb38EHDWVOEqHl/GSBFfgr
sIBl2eiV/Gn3Qg3xrfAmAKPB7elCi7rTqWZPCB/LdTIifQeJV13rVg5EaY+jr7wfxwty1nKm33mi
dAVR5hV6qa/yrumSp8NEeW3KOPEZgsAhQnrsAhmQd6HUOEpW1ogW2i9hLk8DF3uTWQzuchnS1fS+
IT1PNSVaQRZhnMHLfYnlSXzbAvrCyMCRqW49IMj7xMtQZVrMuNCINGcF0rRa1cNODH9ayPuBNI4m
YP7s+gyUNKcSHIMRVVpEowToiZjtt6q9xxiKbm67Gz5NMdxI55yJe+XW5fmsy94/A+O2uk1hrDoC
5OAUHK11T0ioE2E3fKEx6qhLSaY3xMXQrf/mvjCXGp26YPIwoA9uUGd0bmuOTmRDXFLgxVowDS08
xDIbBoNbthpxxZrigTcfyDWlwTRvchYntIliQrZlCy37gypiRDnX2LSkH4YKpkHOy0kilurkpzZg
4JvTSCIuNeooPGGZeQoI03QOcp7c2g1zV3iI6orUdth1pVjzfUSox6dOkuPBvdGSJnJcfxrXPmA4
W2nWhYtjeEf+n3N+UMRaQUYIMzsxX5AMc68FcC//51rRLPL7RXofVKbnAaVhaBFPMXC3eJK4khuy
NFo+rG+TXDQNs2Z5V30n2Pqhft+L4IBQZIGmo69hvMVkuUyRvuxoYO8lJRnwhS1evNRwOzQfDR9e
NxHfAI/a8PXhzHaU7uSyG0MccT0WE78mLNznGC+yowAq18XAV4hdpibLIURGzmoQ7igc0de3UmB5
jyEi0ZhdkZBbkI04WqsjjC4rc0WWXgYtka2Od7kVUUp1Cwj1Y31kKZlS83A6eLrnMKnIZCXaj2FM
s5tf0jV/uikZ/X+ozkcx4lFtwD8Vl/9AP7Io36E2iUfm9e0MefT+bk+vMicciimURj7U5mRNuptG
XEvkaJX1JKJkWeIryuiZG40dWotbBUpaNQhzTiI+g0qgXEfVfXpjThn7Oi9abf/KzrTPjghg+WW6
6D+EgKwy30cPxO8FDQiVV3KlDVkb+XMakUB6poDtKt1Q+B2iuEKyxxHGh7WQmLHDC1bRICVWXbsG
RM7lgpc2Qx1EX7kUpPGP6UL+g+UAyXjOhojySn+prM+1ALpUQOtMRqWOiGldfHVnPTlCgqr+/06P
TrVj5goUZDIR6VAnfkuCMPJmZdy3yApPYdkB26waTxB/hOSQXqCJwNzpQtsjFOuAhqe5zD2WVbHx
o196s80/TuTrcf6Ti97EBTvRHGQ5nLTtMviG9BsKmZF56fk/Av/hmqxYnQ8CP2uSBYKQTMbMuXXV
KQhLHPErPFKGFqKOOt7gdxiKbSWbaPvx9ZrJD2jfp4pXrbHzCnxsrSnzCDhaq6+pusTi7LLHestA
vGqsMAw+WxcY1yuT/EoClfGtMZx/KZhANB5QfR28nK5OzsYYv1tDpHY8sUJCmqfk/Nl2BjKPuKJt
Q6rqOYsMR5unzzp/7bxlBTdrXtyMU1Fj5FQGKJQgmi1DHnLuc8qlEcuNnamLT3FtEESKQ8mrSycN
3mDJ9Z/o/EWz224ovPVLRsdvgL3A8aAPsLEEOTlJqhi82Vc307Qlq2/WS8tQruXU87wBQpK1DXF2
k+/WbxLYNHNwPwwTYrPZxCLZ42o/uwjBFhwK6OV437TI9C2f7maPj0/tkRKeLpqWb8NPjAGGeIF+
tlXdsYKot15uAbMLepXwEaqcaeAIXLXcmcD4GVH0TkA23hFgsllFPpW1/ZuUk9TXxynDMQawknmU
dEmcdAYLictqdT/qpgAT0VuZNaUhzxNMbimQsv/ArMS8KxvnB32ZLCjC8nWu6ZpVnJ2xTdm53o7J
nXCdJrRjCEBslSR8LVXe7AgpJrFZJ3xwasixhs9sGDUv83dY97FO5/zi83Aaqn2PKovBUhFbpcn4
dJCEN+1kwfyYbPWCICFdBHloxKIMG5TKE1E/VauAdtKWB4BGxUo33ndX3OwbhCcwaEIHIDE/+irR
0lHeDARy3jLXbVacYW2IZognWOs2Y7kcpsvbpAAZhckaSCmJU9vZx6T+G/YUj7XttBmsn6LyoOvr
6lJXscO4m+9xL8qJ2IO1DMFgukNvJ0TBse2HWap/vAu6je6jryiYh8HNTtknQlwdfGXp8xeHvA4j
p64ksekVRcBjDlCFmSznYR9dchSWKjunHdcp2ey17Ui+Y2kHtOmhfwoTjh+evNoRKw0AOjVw8Ca9
gOc6Vag3hAdm12U4PzvREWxw/7Tja8kfSmi4AD1a1SK9N2Gu568YWbcfdme/DMosd3cMgQr2bpgL
UfB0oPFE23TF0HgX2kX9B9oo06QcErsIMYdxKv67DFnyBKlLyLli5Oo1YJC+OKbV/9qw4Ec23SIp
ctVNoLqAn9Ko6Ck+/eSSdlRcpHskiBErRIGsN8iDS4e1UF4KV42c8+Dn8A4xGsVuCjEKa5v6YwPy
LzS/Uv6VoaEIWFMW3H4JWLHwoLXlCqzQ/DIh0oEHpYuFL2Q4AI6iez+WmEF7CcFcmQ//inSqQV87
kxsrZI1imtel55EeAJozMSZJbI/CJ8caZS58oLuJIvjRmAhpxFnuEBmmODCMwGxoxvhVpkL6ls2y
skXtayTtzK0dqJ6L/BOQMfcNUt1//Al4iPzfMlpDyXG2vGRd6BwfiNbqSQihKIJtBssJPYHx0Y2W
qMvKsyECOtYNHjoEnHGpQiNeaWIRgRODcPkDYt1g/asDaDDZA8UrsVI4mi0V6LZtKOb3gnfVnPL1
2d4EQ10vwndodUnV+yEVfHAaRZ/QYsGS3DLhnsd2G2ZnWvcf2PcLKCdoWn5x/F8mPpBQUOqZ6ZHR
jcb+fH3gRsHaQa10w1lMo7yUcRF+tnvc0kAcq130SzMXUl+nXymqh5lWyrW9LYdl+8x2UJ868Tud
h3mFpJRNZZPEkY7gtFBzw4Av+srdEH9rVE2qz4Nm6R0h3jZSiKDK+ukcRAf/QxX9W7Epbx080c3s
S/QXgBoQwSdn2h0401VFraeNR6ry1PpyOkLp0zB4pgirco/FmSyX8p4Vwy59dwIVc1JySJKbgZSW
y8XszAZiKuF0NK42QukP/PTYQf0PyIdxUYfoxY9K0husjeAKUpKW7RjjQgDEYzDi2Ft5ugH69+cl
kQZsF4tZQZXZ6bIqia4/d987k03RHxfBCoTOd4O62yVtJt1z1jIKd0XEm0LLugqxsQ894cWY8zlS
QjZ56dQV0ZCAYNidyDP5NYPCtOZwxydwZ7980I+LVax42w51DKK9t81hBcAPWwNzLRbchja0VcvC
BF2p2AucC6M8ou2Y27MYRYxdJ1w/ri8wtZ6im0ZV7zirEif2v1IMS6HGdz+8LlwM92yHwrPqrxDp
52a1/6SjE+JskgywUbFB8bPW5FqXACXDWYWOmajRe9xRuRL4O1wXk/DuWWHAcZIzziWO397vVXR+
GkgxHzmpBlBWzoI9AglbUIfhf2yg5bPRFiIildXY7YZuZK4dHvrJCH8imFHOnJWfnUy6vEmAE8mM
3pV0R/bs7gZ4MA0EZYRVoixfWo0CvTWrPjkfzHw1uIAFWPpMVZcr2cwW14dEsb1qBz0oay4YnQyz
ZbfHX5yL7UGE9kvBM5L4rRSXqSC1phwcvHxtQYK5zbKIrdZUjW5huqiLdh6X021yEcerfK/a0tKv
IIinZ/veFmrgfBzhPJJ8WoCrNitrcx3a46eHx7R6yGGnUECdABtd2H1Pge8oOCqct3xvGmwoEhzY
X6Po/QvH45J6K+rJ0Tdn4Q3+fL2j/Bz0oHX1yzPhiZ1tShA5edpc20hkAargK7o8Q5W/+OAPD099
xYHtnSEev4dXG11MWERqrd5dVEoYD92WhdVms44YTIixsX03Uuu+Wm/uvD1PiJxjncO+IuW8vy2m
ShX/j/3XMMtDRjfra3u2E+rlBY1YqMn7krZEIynl3WVwU9DyND1FrcnnWCmmfo+uEBnR0KVs9m4F
75pNbItOBsrTIXJd6+j9kqiHwAnsmT9gfsmMHJ1iJFtSp+aqxArBGWAnrotqTuFDCbfD2+cKjMLu
0oIjTs2EljuGEkTZEcHRYuzfWoJFPgq3xVq5n1p5271tXgivpcyFJ2LbHUxjZwNCL2HxGGJoUHin
lfDDJZyJQDhJRtyR5yLm59U2r3OWtdKCIk67L0JqWEuP8bocmjkmx/yDyq41uksjuCL/HogvMCVv
ihr5UGreqlzS4HVEWijYjur6ayxQK3EyKDY9H6G5uOJLUVdppH+i6UhqZ5fy8EbP1MtC6kumV1QL
cMG8w9fnBCyh8BHpuFmi4bIAYCI4PkPA6DO1pxfkcdR08lHHCjosNNvH4H/P/xrxU28ebMZsF6TG
94lNfwJm6hRh3GDmJyQUu0Kh7VC3RH8Noc4GTCUevsOvgiGk+x8NevOgAuDmfw+rN15Pn0HYZP5Y
k7pAMBlZRZkOGDNB60M2mHSY5dUfWJ8Dz5LfBw0wzUv4Y0bTBlntw/PfIY751QsKGQ09HZABfr6V
cw31Cpu8UwekbSuPpXXQ3y+KBea2aGnwfb6PAzQ3w1H/rxSOvfaxMxASshcvVuG3ThLZzLsuTEiT
EStAqlQbtiJ2enMze6gYU1wbfn3nS1ZwfNiM6wVQB3McIXEPEnN4xO2qBsmWqRi/x6EraJMZNUd6
RG+JHpDLM/5AlkVej/4xDRCmghPUSaARFO7j4xoCA7WjlAaT0RT/sGgE7ha3Y4a/7/wPFXuAdVEV
jRhckAoxEBTaI6nlQGpFta5iiVT1n7FzasDeQI8c+J2v/EWg/VMICdHgLQa57QHBjNgggoJ/JgiA
z3lx5TX5NJfTYVLt8cSZPnf0NWzYNco6fMyq0K+cFlqgEVWfSg6ir6wuGPKkUERXIWwqvynRKxzn
D29WOhkBjOTrROGT3pI9eJGNDqYOJ/vgGSTiKawQw/QZ4caPTxtUkMwlPbK/dNylra+daT3NbyeV
euob9LN89LBbAOhxrgzc/CBGLpEL+lpQiK10kPpsyEsPk28a4jwGlCe5iVABSC9ajnJMuC9Z1mC7
+Ke9dSxv7Prm6A59ScXytoHLKbuSRskVayxe+fTLsaCsYSlDasnwGPLAjD4731FzwugKufkILRfg
+ltSaJJNZ9E1bf4MI0Yr8a59IkjucREJdC2je0a1KF/m7+iTu9FD7hMe6XZLPZD6qcISQHQrcFI/
mTDC2ss0USkgM4l0L0pIPhPCgCRKxLU4V4cvwlxrWHoRxizHF8DwoDpruRJyBYBL1/Rf60puJCiC
yCob7EY3kQudWVu9tfq2qcbSGMowkUl+g92z1AATN+xfNLyPRalBwTaBfaCLfftFVn5VhF0PLIpI
e2oDpvkgbS7FZBDW5GJsU/KrrU6y7VQEj1hj0H6xl7o2q345ch0F0ChLTZWjPrbP1K0TEY4arFr6
HVKWn2t6eZnqph+vt9CEkCq2c2ofdRC4hLc2DZkXWFWNHUxZQmrpshxipalfqILwNq/zMBt1o1as
nHHiwpnsDw40Fmqa8JrzoteYJ88x970tnxCpuPluMRdjIaKP0jHYTtewhmr4fMLE4DpsQxknc+CU
sQrazfLnXSsFaQ/sjl/Gh2PgzqjBRXbQftGDEOs/peK1Z5ZHMtDtEcV0s3rGf0N2kJ1+V4eu3evL
XnKY4THxqLTHyCjbKP4PleIHaQo9w7O0UhkoSlqNXGTodiAfaWRDnTW1aj/IQXUMdKeN/8eliwNx
Ee111I3EJLSL9kredHYSt347tp66N3Z5rI0ABnRvoSPVSk18lnpsUvKuo3/gEM/x6aQ0GfLFcYCj
6wO8wkXI42Wm3IMMX0a/ixCvWo+At1OFIDNN/1BQxiwlvgq1/FFk4dpLzSq4tFoM/E7it0ycFka7
z1uZDjEr8SSe4P50/JdqHaM52+0u1ighLF+MsU8bzXnT0z1vWB0lkTzKGLtQIpivqdCHnz/LRM5W
gwokRkMNF3To7K9fwsVPM1dNsgSStPfwTZLOV+nZs8ER8aAoUHomcbeUl1NUqd1DWtfGhNbOEWgm
9MqGB1NDCpSLyApVYl74VjnDIVIvvAOmVijghUAkipJbI96m9kVwy0iFYCKpg73Jaf2TdSyZUT+w
bc1foesF6iIyCMcoJkUSvGfNjb5PzH7GzX9khdlrMe5jFE0jU7gbgJnrMZQqNK20rnJbEyHsioUv
VCNAGGMG6Hbk6LSzsAJ4uT0H8lKHm+VZh5sCibfb43jgyM7FN88b8Pi+gtpU4X6fhidxLqzr5jrq
ywPcOH0WfGE+f/pojyfR2vWkV/cipt/Iax9D4xspAItxkuqxhl/w5R/K4MkyDAAu/3ok/afqc5nC
NVNsShuK4QmaDbkkE3lNAvAugaRzZ1KJtotRI2CNvF7mnkJExhqXumuTC+YtZPU6yl+lk/9U8Map
T320MxY8imm3A7LZ8cxLZOQCf3nFZnFq6InMfVC35o8PXW3FyDkRi09LIy4dhCkNLnYZBS+s/UpU
t1djAgxTYJyOdMAo8G6zfm8X03ssh9QV1Ti0WwrFfAwt3VgioWGyKJHNI91m+BE7rT9U8mqvuzP7
Nc0joJpWCY49DLf66WbpMDF5mzpnkdCbNyPCze1VpHzMEaU472EW2vc0xwAxaZSaVc1Ys/fY6tZp
3yLBDDNvBj6L5xW7VKcOwVFSAZTQRNOHAPEEU2a9LfU2zXRquxrJISJo/UQJ/l9eIYQV2vncZao1
kD3Dja2yEpaQJRUJhoQmMwartC79YVTtnrCXVdKLnbIuPzIvu5Tr5msxgv+2Yp8kP5p6LMWN24zO
ai0txmzndMKB9HvwAczsMjFO0o6KNmChzLRhuM2kgCg0PXsw1gFVsDNcB8DIWWCBmedvHPZUc2Rx
jHBQ2rNy3+Q1X/yCgEtSacglTQtidkqacbQ6Lt9/vlOQL3hI0P/NK6SdINMC2IBN5EXGA/dQnRO9
8LcHhnOpmdwS2/cQTXU1ZxI/OTP0ujSX2MG56fV98dl1Dmr7p23uRksjQzXtqUvcox0aAsNR3HX0
ku4H9WTgz5ljsYPO0YGw49bGmltXCguzL5ekD23EKN+jzuQm4P8xYZfS9t9jt5/ZNOGRCOe7xQBE
o2vWBTVL3+dY87+3BzDypjyUpE/hIR8J2Cj2p85dX4JoGdv6Sl3zRFoBwj0x3QRJUz8HoRH5GXYM
YY4ps2kcViJjmCCsVCB0jvcndJWLZwJ65QqaHXNFe3dQ8igP0e95xVMPMjkGIexGUJmTRdbwilYL
VUo6o2Tsz5YYtVM4GRV4Bwiy4uJBTgFhseYzVDleLr3aByMYTRe7XhRtR+8nJvebRdNzJ1pn/yBW
liBe3rREW8lBlyZ4UseYJ60s6jms+u8rsKAwTcXtUlYaRWOmCiAe6uoj/oY2y7h/u60/87GkRIGs
4tPxygW0xFO9k0qhCsCaQnq20GZ7X2/1DUrrMMqWJYNvZs+dg+T+LgCceBkMUOoxEcnbUS2D8mhR
gvx4mGMvCrLSfPTL0Jz48pIxUwEM1l9bBbfe+vJD8WVVR9aX9hjkcNk3B7f1wxGFphgOMFbBb5C4
VqraVT/f2lHbaGU+gU6YbLYzmifkO+FOzEfAO+bhItos6c2OutxPwdPg1wlP/i8gJzwM19qN3boq
MjSF8esVdPyVH0Hoq3b90NMee4JmJ/LY8QIyl+pVpLqUWrAHVe8y01DN+Xd+xK4BwMDajp8ZvS08
iazyFAiumGkR9W5Iqko+u5TrGCplP0Brw3kNUQ19mDdaj/VjHbR3QIGxrhD2jgwSORHsdCSKidF8
aqLXZXqXNfx8leXsqXBZENBJHwElCH6QJNNjRzpwQQTlVPFsN4s+5gDEjd2N6n+cvhC+rSntgG4Z
pcaVIhvkMCfAAcaEKeRVSNX8QQ/Js2sSuFQDaPfTKBcdVXeWEM8nYCxF3iyUCIFVch8ciWQV5aVh
qSwjF3TTpH4BMLpccBgxRYKPm3ndMmBGF1hI93HRxdP2uLfIFmUph8vXT76Z/1NplbD4W0Sk4Z+F
oxOi/UR4RTE5QM+8TlPUYjIWK7wsoirciBxsKT/y0jiR6soZiBrCWrM6IHt1zXsAa6MzXLs92ppA
NIbjlEv2qsyX9if5xUSH7fp8N0+qW5BOStleXvYvoImRCcZnPXtCm86b1T2mXE4NldcEyCWGlWze
oDCGWeKnsZcuwwEh9w6Q+m6O9OLuNDDYb2iTuKknXnOVnckF7QzCww+M3z1yEuqSfrXwWsHqfNM/
/PIaMrMbcu+536PCFBa0qWG0RhKfBn6wZgQ0Ns+SdBwJqKVYJS67ZIGLSrtN7arumV4NWvIGqFZM
0A5NGRd9rBEKHgoUdAMLNpiPVs3bn4xOcYnyaVrFZOvwekwwgnkWcWwJtNxFcHNwauYNh5vCsl+x
cqBkzH1KRFAePXBz6Ie/qGOEsXxWsyA4r/9ABICNzyx7qsT6KlPvb6hvGsSKyxYPvmQe1sjk2vHP
2SvIkUuig1//kumFn/WLP/rZnD2/7E3l/PNDHMg2MlzebD3twwMeshVryM/IRUTownLI43xOLnYZ
MuyK5vlqfCoWshJN+WskRThgS5qwdF0XaBH9n0MRb9+2qPjVUmZjHAOebINLvkB9cFuQOkit3dIq
n6MSOtLUywPnn79gDGAVLfiSpO01Zir1WprhA30vi1Q06M0Yd1cW1G/kMaAbQdrkqxNSKe4ERxkd
lBcop6gHNGu0gZXZNbTFWRDC5YUch+5lDPgSUOKKr3ficRz5owIo4bpmiVL/yZt1Lq94ILt1bBOD
L4szIkX+yveRdPZet2lIRUXJ0lZltK5O6U2bs0eDuN1yvM1YUO66e8XyG7EJrKK5vHYDgsUC3i9W
b9p6TiWkgo0RyA5g6amVlDQoh9kmJHpM8hsFnyywhDZKPZlxBpK15t+rJw+2t7ABWLA1bYArtmtS
EDCOUrNj2GKKeeAOOWMVdDXz69ufSBi2pM/qcvSjlAsv5KnC7qEAaD2HfMFtz/3ZRV4S+J8dKqjL
rZN6pXkZWuYSuI7sE/pOOEJKMi08HMZrB0c84kEP/IHxtnFxh5voSaao/3FDH0Uz3n8ZJra6e3XS
KdS1BjqhrLCwdAnTK7n4o63EQ7FNeZQDeVOFxKGv0WKy0SXbXEflVsGDFx8zGI/l5CoDKiEp+8oW
Wb/FoUExk3jwk7NE3PUtD+I564tLjfT/p1bfyfl1GtKR4obGAH8ugM1Zn0+Apj8PF8WI4ntYZ3md
dlCdXy3CcA4MZw4JelUHjNYY8T8g5QWGwqqPojRmf+mSqVPX9vKTIJ4bPqS67tnaCyrY2K6NZ9sk
QrB3NL086odAWMx+o2p7VSS6tzF+lfM9o0pcHKgU0C9P2SC1O+y6HTCzB/a4Yqo7qo28fp/lB5sF
I36Rw8N5A7BYSmKA4cjTfb4dxSLSvHNkHpPJ7bBDtRDI+MCjFhXSm++4t0IzHtVoH1VfukQFzRID
BZnuwCc3/H0DS6b5lFmuW5o/kbgPuME2xpDAZTuZgHIJrAEy76621cQnzkEregr/oltKYm/0FX9d
SQny7oDP3SuYMQsJ2mu+iXHZj7r+ii0X7uOYX1Hw/VPxe09y1a40cowb1JQ7SUs8CB351XBd25gd
rcGk9hDUF2wRPmyK9w6c+bxihEko1lRnaVqmPILcOultkpuv/xEzytfqOXxDr9M2koA15N0HW8Xk
YhgAqn3gszBcLEWz+7zRhjKyjiQYGYGJDWksH0dcsHfKVnRpiaVady1CGaVen2/90se7hNepf6dp
j9onC/Ae3plNwQ7Inn7T9XWbRJljTtfNJwKg6dQZDeTIoj7DsmAuAmSXO/3kOts2Yjazd1/fu92m
atFAmmEvnS6ivsUYKxDvQHIxBzbJkA+fVm8kcx+px9j91ZXyJNeDac06f9K/3Ov+fdHyJtFEVbOp
UvnYSTOEK0ADwg8r59LxD68R7KK/BeKTlFn5Nx54r+ksMj0=
`pragma protect end_protected
