`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MT2R6c20OvmsgB/H/cSiEA9rb8Gvab7dHgfWM6wkZnDgrySOlTeeE38TggXDG5xW
K5KXZDk0kVWQ+J1Jkx8GhUvOJVrp/DDN1APWCnC1s6rx2OFfOgHkfX3jYd+30zhW
ve7J8nIiE7oiBZ7S09mflcHNcovXkUW/1T7JpKdbhAE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5776)
gwV4psyx9/8jzscO4WD/d3+ww2k8o2Pe2qXQiZvCCLtAcOqetM0sVjjCrAI828gm
nrjmUwqjFlVXIr+sk+4W2rWfd3r8w/C6iKvecpJCuA9xTHHsfzhN2433JIB4ufj1
juzKt4uxP5C1tmXqGTA1zpzxUEYHI2NJcfPZqiK4r5AMbSDq8wp1rMGB8HdEXeqa
LUV0VLGm0aJP1j7/8j1pHqT8eCFB/Y2VQeFigq1UtwYXKHzki1TMsPbE9+GOOrCN
lQa7JTqjxRgEAlSlYvPA3SelMI3bcSUYdnlk++A65VAHmdvlSRH0Sr8aOE7OhPxs
5JYAQJhXKDFODcuGFX5OP7DrMjpE923FCBf+G9LeGStE6t3rODaTjYu427i9ay1w
Fen5eOM+ljRHjWC+A0eV6x9xYOmqfq1nIuo+JGo10hoopUpaQEdx3R4KGlMhtduZ
+OG+qZzsX0TxEO+Wg1Wpc+GVT/HV7Ovjb8XHR1prUC8L/qmuw5ia6+bJHQiLk41t
71bcemElri0MGdLueyw/nmFEyRmjITlcc/YP5Kgb3BxVQ46U9evIhl+J57PgXSSq
hAYAcgbCxx+53G0aCgdg+rOYjbsHizUU9WA1innlR5uE0NMrklilHFTf10v4qhxH
hXc3u5H2g9NVH4abwXaxGTZL7HlgAZGosjSJM6csMxJaXUGnkbYkfXn/ZYjKuZli
Y54NoeloTrH6Aoj2CRDtPAa1TJiyRm1AWMSjeTkua3NFcRAdds/afIc7n3zigUas
1MmN7hbUYIUsXFviThqNRsu3TkAqqRpOKGGgKwzHK4Wh+M0lUiOT3buwyeo33gR8
0byN2tbQIf1trlhsvcAzWhvXTXsfx9hSyXGKTOeHNIp8mXMoThZMYAaEBZw0n+L3
9rYP4J6iNoWxGAb1dakepJ5pQ8xryiw8F32ir2iv1yN6sAPAkHUyNSGF1z3o3Xnk
ej36yaZBK+dmJPQvqG6dhU6ApNACw/PbbSvqfSdWHTGCkhfdte1bU9JjBvxRaCZb
bW76w35kNUHwujBhzCAeXRpOuMvCLcoN5xsee7TwwL8j/E/ZmB6xiu7UZClybdz1
wqrP4fr3qO6Nzeo6OsXGuehGTG5oIsJHEyw8TSMOAolPHHxWf1wnqnTGV2XFnoJj
bw56KXKla656JSrmoTRS5A7EFC7QzXSo/IQHgm7vQJ74RnV0xbgxGzjmI0i0xP2u
vUq4cgn0OH2vhGa3OZ31b4tK9/wjzsW6ba6I1fp3duqF5xS8rC8sy7YGGFl0NFbz
t+0/ficGQlzkZzPsc1Y62CrPs5I9Tl8Jq4Uohul7xTA3NDvhKYquU8pmlhLSjqfi
579oRCImE34y/qvjYVnZMmK8J/lQ42EwfzaRuDrRcMiVzp+bCFOeJfBc5VjTOrWx
sQzMwN/7tADvz5MrKVqIAYSoQ80dKTn3ImXU9FVYnayiTEJAR70uun1mFmCRdtYK
PFLzbKaYg1+B92gZCzljtlaOB6gZ/geRfREPohlPZCjV2jIGx0R3+jvQzgj0MoDt
kttouKq3wB38Q1mZ8uZBFIr6pFFqSwIN/6mMhJR9TjXNHMfrbDu9PIWv/aG8EpHc
UEz4ikQ9sOCswupgXL4bB1Dmc+I+VaiqoklMkXSqTY5c0P5Z+DdW4JICWyOza4if
pC8rSFwZoAzh1I9ErX1VTyUg6B0V9L8Px0pEXop0zT8cw/IqxrbcquUvYwPekB+z
TtGnbv9NSwwIFiyL33R8X0nyzhpstG59BWdUpTW95cNn2uKZQfOAWA+pFX5umqhL
DfQmUr4oupRRBf0sSZNroSdS4u9iOLK6/cgfglFUS5vfz3wBmw5xdzU+cOL3wU0Z
IPHqlNlg2HYM1fyjvdJvZeFQW07BOmTbVd64OscJaNB3Mr5D6bhb+4rtHih1YThb
FTu5ICwFNdSFWLaPlTjB80dUE5af5ns1er3/h5uqg5P5ce8LDkV02Va/4FJ9Xqvl
tgctxQ4PQrnjXAoLkCAZCDPI4LRzUUXzBS3cNZmluMDFd71Cyp6Hu0hxoAhDso5w
Ivj7wVN9Z3Al4muAIi+FDATgcOiZZxWRDuTc0OaC/WC/cON+gcnMc6sE/l4k5e2j
GXd07V7A32pl1/pyejXkfdwyM5ZfjyQ6q0AlFgohn7+CbNHuoZDcEmJ1b8Llt8jZ
rEuTjdANxishn8F0kq5d3k7jVt5n9+6NzlExIJcG2O5pvV5EacLt64CdgurhAaIy
VxC4Y6xcLtDLCUo/wM2E/oirQbxCbR4acD8pAzk9bfNGhMtm99oqX18zm2cEchrd
XRcdU/Uq2rvNi/rB9z2gtdEzGQkvM4LY5w68HSU6C//6kdbjT+gM6xXPc4/g4hUL
7u5kw1WDx9GrqZ2qZEPZqjrPDVf/wXMlu8b38zbltbIwEMwo0YH71twFgU2/6jhi
/fhOVCFlj35JREmEbrcZua3YrMsZZ2GaIwoaBpOd26/yb6gjuiPedMxP2vvXnfqA
a9HTj2ms5tbKTFn5eewv/Iukp+440hOt7RokuButP0bi3bxj7LWzweH80UqgGBqd
h+FSyhsvx4IDheLR9mZrv2QBLOwwZuqdiAVcoEZ9wVDPc2VuNJbUYmO70gLU3aYH
TZRgNv/3p4Va5u6Co+WbE6EElkSM9EVKzmrM9vcyaM5TkP+O9Xmo9W8Se1zjvPP5
PpBKf/xCr05pLct7irs78HLsE7BmmvQUcqqIYSPKG9hoK3l+LEKlRj7VkO7tyfQm
RqNUNekRGxUzzIjHAX5coX8DP5HwDTIBAcdtUV0e4X+Lh9nGQ9PtAJpsBuR4MJw/
b43nc4E8h1dxi7GkmEpsyuG4LGQnDoe/h0x13vCLiG0QIYBO2AfkePsWmmDPBc8C
IIP0AWU4bzqoYJ0jKGR+L6VSG9A81eJ8p01o8m5umrNoYcosRx+rkTuAuQcwPC2f
81jAF8INfHyaiOyYU90CqFk3cS3Ci9NV+0tkNjpJex7QK13bt3wcFsSrH1ZJXveJ
p+0lhr1o6YZyHqQQnuREN11nnkZhsiCwv5xSC56p+bputC4MWE/tQhCYNqpYRMx9
3wqGoPVhVUl9+YDdg/CjYWFFdl9hUKvACV4G/BuVi3DLAPoWXCx3TdjfVRc8eytR
pzs1oyYl9g17ln3fq3OzYhykWCWrSSUTCSxvUQa++wd98vJfLc/ZefRGn7Kmo6zS
h0ZEiX1zH0dGlrtiHOLedsi96ZKjRPoHhhTU92jPPtf1WidmqNOQ+Sw+arDeOtaF
ZTSfTF0RtoUrN+Nmj6ShRfAHpNsl4NsKbWKm2obVskz64GmAK8nUJXSaJV7s5CsI
aRVKLaiafvFbQNWJLmvU/z6sa8Y8QMuewxuaOBPOzgf299UlgKLeWDE7szfMSgqq
JPVF55+QPit8OUFM5Ros5vAThCRFxCd3ExgN8FN5FWO4bcVZnbR91Dtr9n4PVjXX
OP7XZRaOABSf954JFuudD631zIVLBIGD2/bsPeClmPOh0yQK60uOJyszEUN8j7lF
Zz++O3Z7TIWLlrFnNP0+skiQYy8J9MY4O5yynaE59OAYS3pO6Wc23sSccHzIHEUE
Uz7lY6N+Ll4MCv6PWbA7BWFWSw3iz0L7ndN/cHUlE8uvra/WlekP/sLELIw4IbmV
57a9oC00ulf4jcZAM6Gkig5CSIKV/JIyKep96bj6QNDguzyxSbvYhLjOpyQWHCDD
K/1Q7AIikh6EzGGJy3i4uJ1eet33/R0AWe2iQCaq7Yye7fy4CyA0dfj/sJSrsJV6
j/9flBDLnt2ooKc0N77g+WCU8ZT89v2g8WvC7jcBiYX7IPoFD4mLU6L8ns4ksHs+
5CANAHwduatK0DkKVqq/zNbnTBNFdu+OsF/G4fWrgF+D1c4sNaU5jpzN8EmttMNM
KJx1qEdOOz5KbiE1oIQOUTdFxUMT92b4rz7rpnTagpukMo/n60moj5+xrDj5tVXz
E+sZNzTXo9LrCEg1TImeTcUtJYHj7t3Fyv95zZxnwoYsVbv7gsHHrOsvA0GP6xCL
/lKxCUx+Bdy2HxBq1Yf4Ip+Xv2b1GOIz63igmxJx/rT2rUxekd8DvDTqTlDh2soy
31ExFD10XLsOwyA8zPNnSYdZ0gJRS4m1210PvwKJm/nojXW7QSBDzRz/UOu8nhAl
Mc2KopV+HzpAeL+u8ONjpHbmBPs0M6tnr4abqnJHBmIgG92jUpb0gDGBeK1/jjYw
5Ye4D8FB6BFUb0J0W+RI2TOu4mtgxErTeNCmcnXaVhB8yTG7fmw0z7J3/HtgUPRT
ZbOKsqhcjLcKfP9/N3pRtv4OjqcMtLENQn0lnPOM4CTQV0Motsqk+TW1FAluBoI5
zCXYbFzAJePif6M+D27PgcW/+S5fE3b8Cld2Y23EMN4V/NGVoxDJnRbQotKilhE4
4PDH3ayQVWIdWTPcTxBfuCTdsLlXu0erg0qEkK0DR9HEWKWTa92xP5qwMaXyVGSj
dL5/8uox9pGX7pQFF4c/oE9lIeEr3VcIty7RQK3XnJBE0CPZqtKFnxriAkUw+1YT
9idZbnJlyAnu1HaVHJ6qlx1jWlFf1JRUccf7uQBTX89cubSCEujrBLrnl8x1LnmD
I9t11eHJHQhgngaenXfISsaKMaOPgJkh2u0RBwR5gMELhDMNiulG1X1O37pLDdON
iw7pRF/aTnjfYLLgqZF1ftFWYFeEVPU7mTIRWtraBAcl/ZjClb20UJiyUBlrMe+S
79vUsZL4WbHQgugImn/WGrB4/ANM2dpDdkaRhv2p91z4QF1tx9WWLJQAz12YAiK6
Z4yr5LoR5rQKqqWyKPCfJoq0YdO1hcI7EMBimG/8db57W9ezYToAutCqkUCzDrkX
nAZRPWRdNMflfU+2aEvpnqBAhBBC3/lJ5/kSBiK85EkTzBMfj/sIVQQuc/A5VSdQ
l4iiLr0l3n2Wh9oj0+zrZmIGGeQ/K5+4wReK6nUcFZ8C0hSXVEQ2+X0yO36xrHrW
Hb10WNxfb97vzddINMfi3ddIVC55tcJxuiBSJWXEo0E4Il5bXsW4S20Vs/pzVjfn
L40atC4NixWSHA29ATQ2xqJE0I/OXWtHLrOJGQPm1iMFPXkMB+/QQewCsZ7EhLJa
olDlfLegkm8VxJdkOObO4Oiv5RntsP9oW6Z1UN8YLTmmNHqW0D/keVcZZirn7FDW
Z7mlR4rNbUl0EeuzYp+nBdDlPFBG+L06vfRyaE5YO9QsaHes0wNs56Fz0ZC93Cyh
JLNoqI3s0Tq22CNC4J5CLEgtx4ETwXKWHD8HEeaaZ/sbZ7RA52aNxzKpgbCOtDtx
ht3rJQg+XqGQnymAd/p3mUvE56Lu6dJI1jCEY528AzT1/cZlFTnPxsVnemTQOyP4
O0ugEIJFQ3kgfgmbA7z4U3bHA9YNV+DEFmikyMM5m5QJStz5W30ypnvXdqK6Z9um
W8FfTvzf6eMhL6OHYB/oiBfa3e2HgCMnWezFyelYBDLsF7jGpu6SV1hdmHhuWTHc
xp4v1AsYOTde8R6w1KjALgORhnCtz9iuNpstjwmRB9c6SnbIjNbYW4f9kMUfzRkZ
rU33c/zcsOrlGp7y4bO73hmFM6r4Tvu2Ggaicf2vs2gwKpOkL1txnjVv5uKEGW9s
qvGB1Y7rp/R13+4RgmpOY6M30E/6NiM9THYqtiC17tbC5681Bi6xJSwtPE66abJn
41QxQPNUybIHfuP0hSi4N/7Tv/R3+nlUc/jGD1Jambt4OCUlNOiAlCvJrXB8wOVB
9NJQssrM/5nXZb4gVS8YlTCwMJAonQ2P4dPnCE4RDMZVos2ph3Ju89jJ6uKIBOla
x5Mi8JEIWpgnUNBH9hcYye8QgHeM7lBIcvefJCiuMAp2Vx/yLoVjQh94EDPBYeDJ
33P7T1RLabpAf18+sfraVkPLKsQmdU/aQEEOf+y05MEt3vHNdtEDfmdZIyZ1Hec9
N4PE0BUTWsNZH0w/K3ZuVyog9Nd8gW94ORHS7+bR+AHRuWZXpDYqkxFFldYfhfwW
bGvvCkcWsUnEjA5inbs6mRzWgx83D4gEbdcaCWxKKhAvvf/d8u2Yuky4oZpG8Y1F
HMGkAfkxnsNqHXQRIWALWtqIdtRyEy7V61nxZb17oSsij8vZX1HdzRU2kys7usXM
jabQrHwEDT7YNzqoC1InVLZimdyKnJXENYEs99sdHpj9yADYE47j30lKfsJnw97X
fLsU/eiJNOlCgYaSKCQpzZaAymQ4soWCWuqhP7XUfc96M67dtHQXhpB+M/ew0JJX
ukbfijJEkWacgT6qaFGBQ4Kp6yUfKNvhZv7EVVPlnJ70AOaj4meC067/pz4Hj3Sx
2TpPVmVxnicCERWL4XK08dLCWePVPssjVx1yGVXl4AvQxf1U1UGbh/UnPwhk+4AL
CQOlQriuM+jH+JFG6kcHuG6Hg4oTUR3uxikCpLaudkwNI+uw+7WGuFPCLmsqGbbr
0/MsAQ38dlZtHz7e4PGjfEDh/OldA1yAC+R6RU/yWFEG45w5lagKds6Q8k+K3Ozf
9jjjIUTWdrcO8dOSfRART9Q5cZbtQKizpqTYp2M+PUsc0G/s9HNcm0RvsiUSR+of
twf6ULInXcJzSMlLiWUfnOczHp79Y+mVp2UWwrRmH07NkFuvNDWPwDq3JE1RkuzV
7Fe25WqdAYmRYkEeifRtIS+umz7h+IRnPtAHJqkGFRPFCB6PrmHlfWibH0xPV7gV
Va7qesJ0ErOnmaIa7B/WlelTxi308cSsargooZGH8VTMURETXuppPcMUSCd7+1F3
ZR8bSPO9Qd5IZLfd1Kx2kSJQAfIb7GjEwDeUzGagfVIlwEHzk2NnJKNLE5RQWeQW
BFXMwk8oIAi8xE+z5WPrfmvtT8t0fR5uaEI0xvcAhFPPGEc+MQ44YfqEjZMlR5MO
Gnjxna8dmg78vc2V5eQ1IEpxVIvFuhLNVwx5ifVJApvKuGBkKjWVV+JRZhOdBZhC
aDsh1XOBzUTDZgIfspfYqZgYiSqlRYlCfTOMYH0uFj9iSWCRaltAIMR2tE5dA+tQ
zNDY3QEFd008aeNCAAvYsSj5cseAz6k0vDEkoNaYUugWlZk/IuW0BE1sWFvzhtcN
Xz5jzajls6D8SKic742DQhy104Ldx8dNJFEOx2N+HC0rpAghNjfasQ5xYbTjRpHG
aZbR9U+PPXt2IyceJuO6YBZOvDgT14gfa8HU5Ac2hKJdWxphcHI/z8pI+Z++Ff+r
nfvPvERAntI5X7c6TKfNpjWFu7CR4b1AYaVLi+EZlk2NbSxvH9znHZ7XRJBoNAEK
m3/gWD+oTlQk2TLF4slFrfnj40KGMKYw19itG4oKSI+kQk+70Qb1U7iH2tIII/wZ
aA2Q0XOpmCiCdtohzTnuesce/LvpLciKoebRJmOz16L8s5NglMoBVxuRu9WwU9S9
e2oBFI3DmBAx49hpyRkLZgXES/IlkjEr070N7zyLyTlFlRHEYDXMokgFXRqeN9Wl
Hpm8JFIilr8YBNuUJH+PeXxhBqtdPDNwokeVt8kvGx3FXqfp69Wf/qSbnRXlL1+n
bI5Ocw2BM3mm7STZ/8c6Coz30bKVn/FgTB2+e01ry8qmDJ9ZHPSvYWtXevQjmjKU
fSXYb5as/WH8yZAoT1udgaybaR3sVLaGLgxIVGg6envC9dMAyeKgEK4O50uRXfAG
Q/v+Ak1cy4S1N9YErMwHmg==
`pragma protect end_protected
