`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tBLn4zZ0Whzoel/cIrjumTltkSwfhNw0I/cSNkT16+Ne8LF3++hCga/1neaO3NGE
aRpHX/mqhnkERYvRsOCmG1xArWFb0t95T1b8s4pSw0v58EtCUQ9XudAXfoHwoTlg
jBsrSqp9u3VvtnD9XaqRNVU0c3r/o1wjArQON7EQEGE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8400)
awJNFnJ9NuQW4jjPiTg97xu5XdbGpzBb1MaX46pXNC2WsYUnPxSd9prnrQZQVxX4
BwJShnx5w0xrRrtPCe974JKpvr4WuvL/TPYWNAIOl0ipoagNAjD24D5HO+eXael5
CYRFFPwQzl1pICkV+GZpXtXEOA1uJyQIyi3WCXjKP7nRLm4vv24uaGTnbXycbynr
gIv4t6jTV5/Oa8LbhIsBlAXSCvJTKweMQwy158qBzKO540RFPn3MugEj2dIQ4qbx
o3fIHdTB8KmUhclb3ol4LXDOsMOh/0NrUWsAhRhIWumZC6FgHHHZ4Wvr95JwWbtZ
vQ8Bk9xE5lDl23uf5vhDqz3tbrz7L4adjNnXFFmbfKkEApebRyxQ9DEPNPoVsEHx
Ruz8KC7qgbUpAcu5YCoFb6Z86VG0Y/lHtnKOR1+XwCTUiidLuhAIhfEFOoDeREPg
aiUnwwgNjCGyCjIzjwx3XkZfOFWjVd4ygTv1DlXC4KRizYCt9iscu3OwBOJSOMD1
CZPP9crdl0ZJtRRVGLbU7nIPpoYDYBTJIYCvVDkEvH3zoAQy6IJFA67b6UfWZad6
WUiR7ctiKQj/Z54kUBTn2OTzJvNmOTrCutfuMqit86rAuzIMgAG3N7bLM2GtT64o
Ydkkt1MwDrPw9eOJpuRoJru0Tgt2zOfjmYUMe4UY8UVvlQZxXY5ekI6WwslpmU/V
xL09Um2VeK6Sxy1QkZOF+U3/Y9rQWQUnv5bn/XsyuX/tlzi9EtM0YGrH3qP46Ttq
mCGP3cwuLZKILXxN+uxM0zOEEMCuA1a5tqZ6+bdLp5YDYksw+6GY9/PPgCBlDkbP
pHL9rF3ER66gCqE6GPBz4GlsMcou6n58BxkB2xeiIvfRwdOuK9Ae98HuQd8iV2HI
4mYICLJr4Z1Yq6oW1TLhauiAM1zm1yBRu1ohulq0+vb90M5aGadyg5e3XOv+6mKD
7QiAwTLNDE05lJbVE39Z7j2bdhVlXKohTleXfLVG+/gfUtE44srjqJ5m+tH0Bi9E
MBsEUp0lulB1ZsIxNuDlCBLPgj3X5ZtyQbciwhc5Cl2BgDEB3yM/osuclYHRZQkm
9wrjHGrMf+KSh9MNcnkPQOv0U94Bvl7S50bP3M62Wl/gyGaFqToO62q1NI3HbI+N
KEcAn5cC9TqWJrbByVguWBBoIMAxS4pQr9PjbpgO8i3S+3tVkNIsbaOazjARFqTW
TX/ExCBbM7O09jYkApjbd3kamQwiVo4W0lCHyXqDPg+M5m5kn+Wp1Oo37UL+uO2h
pCfXZYEryBrqc6EVGo/CWTwjcSu6p+NP7J1voR9HjsEFJCtqbiwIkU3V5sxZSZ8I
Mhb1W2xwXrbdA2zOrzyfMBQLj3GwK3yKbkHCKVwuERWWddaktUJvrV0wH99h9R3k
4L+9j3pIe63L03MSdjjVS9/rB5Ie76zm9N730m3jNO5WHw3WjHzEiqV2wO1LR/nq
sof8Er9nDZm+l3dvvib1TbIsuMlKJXgLq/QCd/gZlwV8ip/LLZ+TUONKFnghqh9a
bgLWK1Y9NgzHBxbwifASRg817McMizw93s5EoDb6Yi8wiiHwCVK5/qrkCe9hNeCu
MeQSmj745edZdMvAJdhM7Bujdxmlw+GpC9Q/IJsqXBMpxmZumUXMmyVUdv8npeIH
T7i25ypkoRtdUpe4761ZQnxiAYgXNKPrhjFLFVXtPdDuxmyNVeA2m5oNqU2rjKvl
4Kozs/7wiED2VeKpKE/c6VBY0bxTVe3WKA+yV2xCcSkgKCm68TCIAIGbOC2kxHtA
VpHEGeTnI+alohoseJwJ0/pzHBcj1mkVxQh/cZN/a/+9SbBaNZrj1/NGpb3Qta+6
fH/M2LtAaHzRQTWwbU7K0zM2DC4Yt+BzMqBxc5f+n0K/Qg9cSMtKsQj0ziOnQdee
AG1ZZ7MAUd9BVQDIpXtWt7b3EKnMYewcB/9r3ImhLahATPjReArj4AoMzj0YPqES
q4CJJSRQRQaqO4MgAGURcKUVPH8YGRjN5uhsDyNbATlj75IMRVBd7eDROujjkhkl
1dRRR3/3PkB9k+D3LtLjxfvBZ2uP8YsULFpq02ANGV2kEk6aCs3a60BwsApZ3d/g
1+vuBFguBdf7tyF4Yu2X2PXyqNolZh4tNQyLy9VcDDVUm74jUoEK6TI71QRpHhpk
4ZKCSxbYRFfpEJBwh6GZyq9TZHlx88ry3NsnMUC/wA1V13q5H2AWEvsRdqTd86Cf
ItXnEI2xMnGObQcsWlTKN6wJWCFvN7iTl6vt03tT06gGWLdxlR2ciL7Ogsu2W1Ad
U48F6LgQO6M0gOVrEmUPnfvw/Qi/Xek342XDZbDpYqYdNiJTGHgPvdnMQkXFtrW3
sfmw/aLK+LmVFMKmzKV8GDJVmaTFnB1ZpHa/Sttfopl4Ifhyuah/5Z5xvmy7auud
zXMHf6/Uwj1oREwAE0rlQEW7NVyaQynN5huS/9J4S7NKpnKFFPCYk9NhATWTihEW
MkiYyeXg/WH0TUoAE/6m+oiOrqP7hgfFcH383aLZU4uRymp5uNBVklCtBH49bKzI
8Q7nRsr2o/XaBwxsi1cMRpD/4JzHjgb+yz+E/Rrnd1d0mQsXr/n1ijWPrzJI0056
lFfTQOttAlcQqp5NjmS5rxbLqxmS+ujnaiZxgQg/qncIpzljcZJGrX2z643rnOTS
IQ74TVHme13voK2iVrbXSOaRU8AEin4qmXXjwTCIAn92BMdjqO6zX4bhEKg4TChO
bwYWq3Kbywn3Sk+nl5wNun4kMy8p2w9CGWxRi/HLYn1xl8bHRsM8y5MGs9PvFUDP
uSgIBNSbkEhOWjMmQTeobBWFi4WK8Ailc8G7zNPTMaRKrgWVzZ1UAVY01jzOkcRh
5oh+Ngt5YGv8dLOeAadhvpCJ3u1bKpiMBOZsK+Ga2Invf/FMTeeb79s4HOKtpgfH
hTO107rIPs+lcKCGhSWzOUr4Vn8WQ0ZqbuWVQoMXPctPHjjxCoUAlEwuchJ32ICY
RRCN1pvizwE0GsScqPTtZqoAbriPujlHa6KTVHha+wbxuy3rA8g6mRKU0o/sP0Be
7+bc0ahZF5pMjOPS/QrXYvCpOSWsiBtu6287NDMu+aUyxB/09JGQE3aYTfgvXgja
I+CVCNFEHqp7PaA3u4Rby8VEo0L7h44FawsgW1MRLhl/PK4fcHBPnr9T9e4eaofY
etiu/g3zKRPkKjpUnmZiYG71OVWTwULDzmrU8mKt2Fw4cPvBA9xyRgCPGhP2U4VA
ODpBe1ecUDzYsFEv4o4ShF3XdKHtx55Yk3SwvvJOgUY6WWadaZWxp9bEWYkJkVCz
Z6G2wYNHVYAdJxe3qYJTWOjf6+/qxATfNrDCKLGFhIYMfovKHOpNVe6HzzJiXzT5
YQR/KuMaREi649bw2IG+GbgJQLtHPy3DEBfwq5lWGhVHEPwH/8qWIIqIfqXwtP2G
nrUY5adQAume3VNl0TWUmv8fjrDxXhGsJooMUfMMBcE+TQUJ2nLNUNGr9IindtxL
/8Xp1dafyyi8uHUCqIQXzXG6d4QA4Zbhfioi1nwYtbrJdIBStd854gao3m3iJ5Na
bbjNeJHL9cVl/+GoPqoDYnFswSAMFNyd3LJg+4E3aMelcvapzkk4CV27f+8HbJQw
Nq7ywyjUY394YLZjgq+bDe4Oh/4QxPzVTgFP/GB4Tk3O6I3MOXSPre9gEOh8y/eB
Ow5/BbO7f4EextiUkQpGgIz7HvmM1okp79kUjBQw7TH9sESUk/B0iKdHGsndCMAH
zjwRkFvFHLLc+VX/cj3ki5aYSAi/rc+jYx68wzDY5x1rfIE0QuK2qg2JDoHspkaX
mAI5GDCKxKm2nIZV2ExNExRYjMwsuEapaDJTv6cfpjv7a/1SOFxkgrfMbxaR/gBh
y0GLm2l4skD2q8LJEwqBxlNGap7j45ZzPWn7cuUFTLSdeIuj0IbLojbt5i8Tfw1b
NL4Ih3WsXR1VeTH2374QZCeabnmTHg9Va5EMTPp53U8zyJtv66P2kkv81qenNRut
jmYUXKlcr+pyrmWU7+P23muMYcReqIzbE2jltLS2l+Juh/LdbxkzY9yF2FKYBhnF
DaxZJLZ5/K8Jm6C1wzcJiBZsMcXLz8iSu1qilppV1w2V48+JkUhwiUCSTXlRud7J
3CnxFVnRIsN0+jqPZEFs5FkuqJs+1xwICEu6etPVF4bsIxbQESjeMbss0oxZTen9
2KLRTiLtetc3IuOKoKaaYAZ5qW/ht7zzuxQOETBIF+Ah72du0yMrJbrH4xf2yhhk
2lLexVILNuWKQHrA2UdITCqv2QknyNBBaQSF/ohiA40nyor+pp7AJ36s8XQ/CZrA
4DP/psdn3vVo2XiK11Of9xrWgAIlltEPfxT5tdghM/691BcBVcs3fnyJ/PTX4A52
ukOfmo7/vigs48DEw83n3Uj/VuBzhMJmiGXWBtbZ9fnEgZPC59N3o6SktcQGrP6Z
CZ3Qqpmarxf445jZ5xK029Gfg95jCABkKzhVRvvueeEVQ5g+JoPWf/gfGV54esY0
JNfYIW5ufGRCdnYGGR54/zF+YWSGUhAzO/zICxbO9h5XnoeiVaDjKrhoqQY+qDZF
w8l+GOOXyxfo8qeP0cVuecnzjkCeHZueBj84jn9RSVmOL6Jr+K/1LGUDbMMFgYUA
PVjcmYzqY/ZAvUeqZyuNx4z8FeCUTRqwJTN4DFRtUgzP091iaNE9GYVfTGUC733u
sAmqP670m6ugrTcgtSyA75JCgUUtwSXohsZXDsgHc5xenHSWzol7r6KtVa/hN9F8
ZGfmOg4eHipDzWYYBWrwXfKSlNHO3d36SUrIOd4z3c/MLNcHBkJn/lnqRXBFW8DX
Tmkr4X99D08Us4g9rPR1UdTeNvg/0qC3q6rTksgw2pFD+4M7gscRjqUtyCkQx1F3
SBcJkdJKyCCmjw5oUjMAYq8+RgHiefak0llYeX20Jok0ce378ANcwKI5jzjnXzR9
unDL1YVvoylnspLx/dt2/EQdko8XS7dxo55u4MHfAILz5E/rD9requiD5pZTebIx
/3lAatmlzU6B4o7RTQ85viq9s42Dd/dXu6rzSXoOJjkDw3d9i9PTWXYub/3pkcXY
UeQClbAR2YPUv/AEkS+tEhTIF0SQY1E7y/K0An+lLL1R/n6dTxUOwZG7lJ7pTgdQ
NPjCrwm9TnI8n0gse12X8WlbslukHfJJGLW7Bkm4Uu3EGikScp5Fh/tHKCrklPWO
s+3oaZtARYRsThCpk/CLBqUpGMIOMhykmcOFmCVWk7ZjxA8+rlvxygQL8x7hsJO2
s3G9jiCQKmEbaxWecq35wB0PSez81jDx63QbjXsN1AjV8l/qmdxXseuz8e9V3Wuj
QjjugflINB8fsnWin3TvlBYBzXxTyn1vsmwauCUNfj16o+zmidmFQJWvrGll9bSd
67CRzTz9XKK1C5/Z6CftetYaNuKf05my2DxFWz8HS86Ti/8igKr9h8OX44kYcVGS
WuH1zAsj26l0l+f3ANg07RHDXbhzu2oLbmWByawg1OFudkIc63ngT/I1WdkQOjeP
U/7JcQl0P4lI3CVMf1RxAv0v+suKo8i8dGdvq2BKeg4i0yCNg6SAPQnADvazoHas
jlTK3Y5tB0LeO++8Vi9DLLTNn2GB3v0ZfpXZyXRbWQFg4nr4RJOdkC+AjKXlBDu7
PFNzot75fd/L01D3eoYB7HFX84gbzInkHME+nG0Bci5w2FA41vXp4h/naudbm2rH
vJUHOwkJEtt32upI2d8omfAvOlu6YOhjBw6dtegsEdD/5X51FfcZl4nU2raDtzrp
A8nQZ8IcKUFqCdG56uVbceKjSPdDTKWPkAeA/HAoiXk7w4DS3r8Yxj8RDyJOaOmd
izAfJOAwykoRyFwcIzYFQl1lXnRwJwCtn60C0NluuJOY3K2IPgs6P0OI7wpWS4hF
S4pg45HfSqABmfYshmatVZ4ShIeYsElPhI6bznPbpNdYTcpY0CWLxxJnWsPOTSxG
gsTShsfUbp/rxEh6fWuunqu1G36KHrbKE6IFwWI2EfO4LY2HO+bCHoQRvSzdyEI5
8DLeegNoV4V23kdnqhAsW7q5hPlxlU9b04QlU1BGj44nhwjkxld2vXwRCTPGC93R
SAWd50XAQqtFc5zT3BGCYuN2fou4LJQ86oaZM+BJlxeKcFRCW3/96XJCiHWxqvX0
xJ8QNfyy2+9frVWJKzv73n1XS3zmQV9aaYHzQ1jp7+c72Dw/0MFhPJMJJQjN0L2F
USiCCmOxrwpRWOlYWYq0fk5ADu6bbeEk7Wd1vlDSuy2Ns5HMOW02kgiGZ41ApEwy
2gDX7TGIarzSWWCAsxN+/d7fPSFg9Qk+uypDiCQsDRLN8fED0lkHvKRYcZbmd2hY
7voWR30J34pwF1Ok6AbSzTFxNgNrlSErW8Xwi6m3HeuKt7eGu5uGqGUJBSJI5A1b
AcBiRqO5XwTXO1KlVPSOuoyb6kdwox5oFYrX1qzOpF/zmQknqIDVgTDy4tUdscDT
nHdqY0kVxHtXONGzMAcqJUsYbPzYn2+Vjo4U68KvuHkw4IOnpHDDA8f8iNX+LClo
n+4Q9AYLkbiliFi1MvyczK/B6X41gso1TyoDOB1AUzFSWTOq1OuPvhD2R7/1+vV8
Rc0C5EPhUOg1CtKNSSuWppbsdv5HZxSBpqiDX/EtMk8s4SPEmlhAAyD5lR9KQTBA
FmXs7oSVlbIhXdqt7iAyr0GYleJuMfNl0xBg9cCMToXdxVKyUxz3Dlg8mVxYyaxI
l6iNpamsjzY5XUwNeaci9K1V+K1GtlfQ5kZqb6ZBwvEv8E0ANvSEEwYaezmHF79f
Sa1ejFDnLvzgH1YW2Ju+JFUMM69fER/7blqbGOFCRVvdAGsVJpfhxb64tE7J2pQG
Bjx1kPWo6l4nObBN27NQDyBzdA+RjOxosZrW5coJv+Gax1lu0Z1a5npJ/aGWuybQ
eQc1Qqbd9Q8NxtNqObJx6I6BnvtJ5E/ZVc9oOAE8xy5Grb3v5fKjBGV95/vXyh2l
syMYiW2t2NYfbgaU6Tokvq5UE0xwqIILj69TF6FdLgApHjqhKrxNLVEdEkzZnS09
k4izcyWdVCe9ifE2pCTgQNN3uRHcKCrvbITe8BqwRtFASJeeJLMULZCmr2YmKF/7
NwSTQj8hRRpPIGlh3ivuaEEbT/CMadC8a+LoSpytMVrFPwOsCKb0+P4LLvUeCUVP
4GMGavhusGrwkssWElFOgquUwOXnH0Lsag0mfMqo7/gMgzjP3Jmo2+00lW9ZNt7j
L/jF70mHCPssI1ZkwGReCN2k4NYfvLeA5XWRpa3CuCoKQ/T4DH7uZbyxRnp47tho
zzb/wfLKKZ9mtTjkUCNbtxaHmp+VZ4v/woNo9nIPq0p78jx42lf3LD7xGsfVJEJw
Y53omwMpCAE9JN8+QkY0zyg5jP0ZN99kN0/0Kar+3EldZorqAKgcIcjj/IKnkJdZ
Ydm2gozGFlOBUoOu0wx/AhG2fh5+hQBEiNjS2Dtn/+U3FlazlbtZeDqld0jXGzFf
AeQvX2OK/H0h1MCdG5GM/ocRqMHskcgTCgmYyeUq1VSu5mLcdwM2Sc/sgyVzUDAy
0O23v/bAJxWi9TmOop/Q2Cr//u1uscHzA0tOz8M+P6G7oyOgwxZLRtQEAuvBsy86
RuCNfGFTyUarIScIvhRDai8rS8G6b6y5VZHqMPD5oDvuw3kPPDD4MFn/kmOpfld3
rAhPErEewKRiq5PtXx64KbIHRjBrGnGTf1dbbt7lJVkg8dXgCFJHuQr+JkG+7ut0
9T4fqaC7DH8V87SvVNSNuP4hhVKAmFwzWldQPaPqxipPTsS5T6itXaMERYI8QJo3
zuhyobluZaOebeJqm+qwheCFM0xOBKwpI969r8cG0q0SvYEc5bZ9AqmVDpw1YspU
LZ4BX4lXyR/5w3txAcVh6oIoAdnq0QAI1xziVJcA3vVU7A4UbxTi7ItYJBJ3roSA
jY9L7r6BjpiUOFz2Vlf23/E/mpV6fUdlB7sVThtv2+5Oo49XaR35VgcbwzBLot/D
ji+vCNZbyKyWrhIrQT17s/BESKVwqOEhm/WV8NHeo6UVcDlCx9kGyAGQiWogsI2+
TtE0M0rBEFNqG/Jih63knuX5OpxL2qF/mdzHAfN9G2H2yb4wQ2OQA8/xNvt98yp4
MbD5GdIM4jW6HbW92CN/OeIm9p+zKRN3x43PnLRvjgGe+vjdKyn2WNtdCczMe6yh
fdGX5k6NIu/u118l4WZ507UA1JjRxNWGu+/zZ77z75OsgHLvdoi4oC20TkGcwheI
sADR+7zeGqupBXfs4aLB2VfsVL48npASV2UATGJaHDynK0f560mOCsVIt4C7/I94
1C/EIC32CiRrnlyQCYIg3XWzn0L9rNLHO7fCi8bo82RUOAHW/qJAvEybJvIsjEDa
4xm6thCeAjd02G02T7cU7bQ6XNyXenod099u/4nzj3c81cknQygVOfBpXN+qlxya
MTEkLoHEJF12L0+jm2LD4MvybQ6lsO2aV8wU7bkrycxNYW9PFe6hkwuO9kqJgl+f
cDzgmPSq6DyKMrwHVGENHkvQ71ad56N3Fe0h5G13eMjQxlWApLUNqn6hdB6sJxQQ
KJ7/pQJwy2dmtzIRdi0K60gScQp8PphfTkCNyfshro+Ja7wVcwWmyk8BO7sqj2NA
+/Av2ikCvXp5AQ3xoRdrJcFnkXJu02cIGCTwhKlRdl+8/n4KzWi/0XxvxJ0ottmr
fCJkPDiKS4+DOqjvNeZtmUUXVpnUNCrfigFvZ8OJxKJw0mjMQ8y6ecGR6FqF9lZf
QbM6BijvWbGf9CAufB/5J3TwBElhbKD0ap/SdJSU+4McfwWqsKo7tUEowMFRGid+
ObeYk8tgkfoOh6cAuL67Zzjwo9E1WR4NO3UHWpAKRwj77KgrqJdc/T+0UpHchC3g
h+gSIyN0kQBXoT1jFeckhvCZ1H1JLEUoCMlXHWu102qgrbMZ6lH971N20egibSLI
JLXSq7c5KCNm2YtyVu5bouawte/IMM1aILqRXS8sjy8NvneHrSANysEMB2+pa333
lBQmQ9DIv1Zc7s7JeucgMpfv9djf50n7JY8nffV+6oOL0g7jMVDSxzb+Pt6ZgNyh
+Ub9CJ8bcnwgDiqaHEN3QcgjuCtwpNGICbDRpD/6yoCYIOTGdOSuzadjF9ntlTRl
U9go9QcO3Nm4blnSmDm5YsPGH/Z9Re2J6AR0mElca5+Y+xFHjmgtTpg6KII7M1Vr
uZqFJUwPkUctFKPshA6KXid6+JZrIGDCUrXLjxWmcCjPogxkU6LqhKS89K8GR05B
QMjoBlAEi36RpTvqwzom8J+qvkls4b3krdhUDM64we49tmXKTv1tal0ilQ2WaNmU
CXD9+KHDZ8mnLpHpgAXYiLgLeS9obxl+67FYuX5bg6W71WLym9P/laySMDXCuwXA
4QCUFt+IJmU8KJT3EaCvmoW8M2TPgw0LN6JnFAH+89juGpp391qsLVgAnH4xg2NB
d1g+4ZgZbjqrvIvyuUD21bFFMfes4u0kQzH0Gcb1PEdzvItOMjmbPdxtbIWxr+mx
4bc1y4Th6jOrvR+Lic6UUR0DXbPzOrND/SO2ynqxe1D6//oYG92O/fDaYdgqq3Nu
m2ErptMCn++EZ+FnwEIvqGJhQSLDissdxMhdTPMuQOXH1BBR7vAcDgRpmt/LMgGl
7oyQzD35RZM+IHft7QAdoaiVL9dAXwVt5MJckVnyv15jmbxe4QcSvvX0fHg2iHO8
gPDv5PNzIu584DmybmQC//gloqEPNT4avcMzXCEb34dfZqLAzeZ/U1Qh3u4uGc9Q
/pBCdAIVnS3RgkrvulJBs4vPaKC4s0fyx2pVPEMTvK0hbKA7E63CTK9VkzIxlTAT
vVApNUyfuWla9Ro8WgPxvgXUXfzQRNQREHWDlWbtNHeC6x+BbV4AujSatYy3ngcV
UBPmPVamKYjHSr4IywcBAuWpk2+BVf+x0AapZifrjEu2X4lA+/qvLwFgYuRMeEfG
3Gp0Kpq+f8IBKA4+DqObhi8lJIJbSooZNexWG8DBiGVSTlJinOIkzfYo8rK5RCHN
16+g5pl+eMK5sVEhU23xVoQ5rJjOOeQdIP0FfLkKt+loRKjgm7MrFrMA9MSkhViH
JA7QkXEL+moqCVLyYU1TbImK/X79lajinTsRWnBIo/VSIrM+TQ1E54OyO3Ihtr0r
aZwMOKBJI20e+/Ktxc3cHCHNYsmPRjsdhxoJmeqHUmz6287AwjNV/ud5eSHS+77d
Di6gZYKuMScb3S/t1+tBepc2p5ysqXdgAf/uKvKMxTkrix0Aqv+1QaEj8kGYCFVW
DbrXKY2k0bMpllsLbUF3s4fQNFYDmZgM6o6JsZEKP35RYhNcPctB+bZA79m4VAlF
XEgOlZc8BEdpMwFa+4zQ9A5c9cGDA7bOdKVWSlTjBgMjw4tZQigvJuCEL5FA9NY6
mltpxIQzfXExDNSysa6ybCNgfIkPWAq0ovC96aNEcfzbm2zxXbCfwF54E4aEl8oO
krglx9mL4XKtqWN+v8y6lFUCNIbhBcRvI5i2y92esbv8MgZgj413qi8wVHCBFEqn
aQvRlXHgWLQEaZ7piXwNEh9rIyN5KHHG3xa+K/osJNn1UTWmzwfiQ5BAMjNo7dV5
b9CrPnY/Wydp5AS0OG2TnV1M5S14ouPsBSrBpEZCwJTPEaKP7F49zFSY/CgbNswp
DFooez9e0RtnZgCchhydYRZBKv1YhPXZs7PDV+P4cS8z6GjzCpyqpT+1+RAvOPfS
BTNb2/WfForzURhngjhryO2EN8ugxrv+ysTdzqb1eq0cdWKTXrtiwCmcOhpUmtaB
wq45d66UyCbapDcFlhN2rjPcIp8KCz/syU2+NFr0ofdkVsaaW+9SszTgOYvHAN0U
EhS52F1a0KyVs+4pIUvOW2GBmQZ/VflFVj9tunwCtoaAZX66O33NbKqgYfbtRDcv
zOq60H/vsHLc1Fx6b6HP4PT3Yvy5bx8WvLfIsrznILzhcRsPZJF1Taj8bpmyJAyd
XVne5BhQmO/Pn4aVUom0qxMf/pYo0SaXgP9VJoWS1u0OrpupExYKGSrH0iV5mzGl
91ueEkVdcywuklFVnGCWKGg1gkcCifHT42m12ZnhbaMdlBepoK8PLO8EDw/YS4Is
`pragma protect end_protected
