-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JzndBq57IKWKdcFYhuee17yst+fbWu755fYd+dZoSpn07097dvvLgdIJIjEXiRAegmCtbxDQamw1
dDzZKhOPQ2VnRVT98I+1BslgPZJq8pegRHVMg9Ff0GM3+p53fXTsOLyZ+gnzcTtdcmVy6ur01aJ9
0VednLBzkV9p8xWi4/HxpknFNmwptQ23PN2ChX0qrgk3A6+nvrg1TLXK6bWNSGyGdG6N+jTpgdUP
ccvLxZccUHMpxNZce3DjDCicqkM8kPkkJyISpZnvR62061fyS9rmGa081ehTkUUvPxSX9HXDkWn/
oT0EjgkerJlGU4k+zm4CtNk5uB0+ZW8hHKEyng==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28736)
`protect data_block
kFQi7Uq/OPHfOT5QPvVNDPgp50qzwokFMvyAwCWF2IEqru5h/v8nS0+PCL6sI3kaeB/yf4IVNkma
e6NOfckMIX3YfqSBsi4nmuNE1wFPuaDClDZ2v50cwGFdJZ94uz+PispELErntVdw5zQuof7F2e9d
n7Frx0H+KW6Vi1rsAcJ3nLc4ET4PeKBbJjW/mXlZHRnY3q/xg9+q8tSYgzAl9hlnKriZJyC9MO79
si3HzH348R/4QRMvL9Hdzyj/hLwYBAmLjwJ42BPxSEhl0cUDdUsxfkk2rqI9i81xhsohi2QyCzpt
OyI9iLhBETfKASxVEi7D7ngCiemBfH3iH0cSZOnmK0rIvuhO4CK5/CNHyGQdLXEyf+N4YPQT0YIV
j42fGZrIcKa2JoOKwFwb1WpCTXg7rfC86mJJ28MwXp5c1R2CwioZ0za7RtlVhvRRe9dQYcYvE/m+
2p8+AYEmP9CkHKG9KErKi1YdS7eFYXJcHpOqgVX4MziDLoG9ZNaLXTOonEOKnK9zTnA37ZWdlvts
t+vnZSPqrLe7D+YfmhixaDk9Typ4UL4Q38LUcs68OLqrYy9bjSV3Nx9hhAteSohr/jJa8WAg3sN5
bc+EHg+iOxm8k6S1xdMPok+S7XtNHplA4HB4QApz2AmzxfuhINS6YcJwiUrH468H3ZKMOpKTMrMw
2i2xlFKW9jW+ytWz82LAyeO9bYP373G7Df8/YTSDiyGNVDkbu6vJC4XQZp0x5ypztJtEmni8Bwjd
wGH7Kd7aNmlMyOJUcW5BkSot77H+Ex509pmjDaA8IiNmSMHszLMnU6UHiTHkV6MP2w6Ogu/b6wGI
CL1DTJA8sSL88RqDeTJ13v22z0IlvckN3nUHLmb+VpgswPOC8h6W7LAe5ycSa0wOp7FL8cX66J48
tUis9y1B+hQ2vNN44bwvvB9tpj6WN/aZYQrf9Onwrh6QDC4MT1onZvvV5kJjYbFzlUAcQytk2xCx
J7yqPkynMVjZ7JK+QBNdiVFgqtjBX7E0xp42qMulw50pi3tt3pi78KJcJd3Ce+EaXZX0ux0k1Jh5
HzJyFaqNG5gAnOA15HTNTaPzX4LOw9v9J6w42j7C+RaIHVQtgkb5uAGE98OSz317ZOGg0svhKaGF
Hl9wmZCLxpQWkKLEue3j+utTTXKRy6p922tL76Tdb7A+GOqGWcEBYlbFzUQWUI3M1OeHPw+7RnSo
9DoCC24vhzO1vS+ZOW8ssrTYaRyjY3d6EeSLBEtnoDJc1YmTQT8x90yhnYyuBk5SpCHqmoJSucOI
Mzp8E1RfcK539riPyz1B2adGzMvPtf/O26TNp5bRBRimquU4zrT+NtFJnVwvhg0twD93LNDV9zkb
i6XLtaYbRsF3Qha3YTMNunOx0FFA6EPc2S4DJ8t8zC8Csx7drZiE01CStE+NWzCYY0/+74RiGQrm
aO7CZRUFMBrCqqT4puKaGWQjp0KdQ6UJGLc+IajhDNomN5zKxGiAhoJnI9ZevV6xUEciMVgzmOud
SF3DdGfmSL7baODXlaOzZSq74w/LXjpJHhujw7ys7vUBYlSE1tPkvR+kRWpTJGBFs3eRR1eWPK0C
TCgk2VB5lb55jPGUlYUhZ1+5SzeotHC8VKn3fx4lP415K4fjPeHXNTwyGPGli4s6P3qQrgH2j1us
vLi+3izdgf+I05QS4qVNtuAICuEaTRlGlakG2JLeC1a9FVFW9lCpgzFxl0NUkQ6YZTNqGdLoFksj
t6Mzj063h8+R8+QaQf3EWmrv97ynaiIF666hvyiZZ1iUtQHgX2cE1RvcVZbOUJfrBV1rpXfDwPam
a1qq5u5PdrHRcqyAFr2Pd55xQI6Heg/OpGJfAuYhEdsr65bSRhcIbDQy/O6boXpcJKsDNxEL4U3x
kHLTsu99/sgaQVMBu9W6g1/MNI1AARKv0kwdQQgFuLWhhs6OjwmtsW3vdlHCBBgS6y/ZPPsbn61+
hAJuLzjeh4wUuh6034q7kqU2ulYDXs5XYj0lMHVCqrmVNIhaTmhp6GfGfaC5jxx5isu394LJmwoE
sOVY+0WfC6AIWtZY7+uDki8xoQLMfH15iMUu8ZctFEZglpMHUjpfWtuYQyRUcmFVg+yerlXEMHOE
f+3aHhIaFk6Wq+G0SmGcmKHll++QUTqg015sh3a9xIlz40GMnjURluqQO+Ls3Ni3d11wL+nAfFCD
KNi6UIY6d6GKMnDe5iEDT71POF7feSV39PXBK7rIUymrgYznQ4HZGWZXDu6QYS3XXAmGwhZ92LtJ
z5Yk1YJL+qpFPfWS93JixRFdlfw3APdaBqu9LACI1KiPx4tlK2FYggwFXX0ckpcZRbCsnKO/qZ8F
ShvYcW79MBoUiIPJhJfI9h79QHCtyeaGSqGX6pQ1s2Fr+k/eUqa9jEejlP+RmnttYmfE4wqwzLdo
5qCn4aVBmPLPwIQmeAoKyrK57EtOAwCSmxLTgg8/qxQCo0pPVlvfsTsEPNY6TYOyCfL1us1+tHGI
I9SZutXVY5UKUMFlg1w/f4xIAyKzEclSS5OaW+bgvbhgngWEQk3yp6gcl8fKiRfx0nlNW5xv/go/
w+FLJpno9uCeCvb2d6CY43u1zTNslMl/I2qovbnbOIEFh6ys9Cr2863vqj/CFMM43EFhNLBJgcTC
9mid/PHs9rFsLvZpwxsrTheW6tnFwkIFpGoRsnv3pNvBMZfl8fHsxYOhJc1JfwBv1maEAJZ0Rmx2
f6vEqqb7V9/iv6b7iIrFklhBqeJxEYprG6jMDhUamtw4gSOxAa/5MLcl59uGRvncoAU2Z9UgzHfZ
njtGjcEjGu3X1ONBwYFuYFcZJVU6NjjyP99HmioNwCx02vEYJ8kSHctANOatwGPDugFuKuZMz4LG
b/CxUxzsrUOOWM1pMnzM//SmTzs4hpcUNoA9YEyY4Yg298aqKc1vj1cvCnomdMaY2DnFvFDLFHzc
V9xJs4/SpaZaEYg6sW3mcGxGaG1ktckSHc+m7cc9k1lhV2PdcI8N8Q+WCei41Ds9RmhRwNRwHQij
FylJMuyxkjA+3wyzt+EbbMW5QUL0cUN1akJV0M7BEyOJYRkUr/fuUzwH4VrFNB45Kq6DzmOqExV7
H2Eb1otqQ3J2VEvfHG8vc38R5cNbK9j9ujT+I0vdSRWmm1l6ttSWb8uutDm3gyx9Iw7wPvcUqPRa
ywsti2MP006D4bZDpQIExB3pG/iYjCyIJ4iFs1fO53xhidVlcs/A+NyqeCkvm7jc7DLgBE2/bOyG
Ohg09iMlr1DHWGCKWw/n7cn5IhufQiGj6XYSLbyVs1vXFyNtOXGPmQC9EMKm6mR8PZidOa5s3A1Q
KhTHQ8xO99nimQhtEQgyi9mR/j+rAz6QqUhWj4DWUDX5E8HjwsLr8gJmO5c99nVNExISv0rP6KjU
XBXumoDI5wXhaN9p8088uo5KXIvE2O0cghdXBu00abGODEGeMLH8CGKnurbqkKFlFtg76oyYEuTj
YbyaS+2TIvgd5hFuvB5qZvvi/MG8jOrp7kyq5eFYcJMH0dtsKXMvAEpFGGW3jrTt/TmeVKL9IOPW
1r0O2qBXu8QAAEmazEwPeiDk0dGp9EvjdNdqd6HY6SfRDPZRkM7b77U4udWjK1rooY0swXQ4CUwC
UL2cm7U3cmgK3V+7/ujPP8kMQZ/6k3zfOf6kgDQnk35AMBy6b3tSpX552q46nUql9/oPRXGHamMq
raVs/i+yh8vwPWljyWJhBNAsoFBObCo9eu19T/H7iouowtsHAmZqDcK726kAnF1FOQeIwXZ9CPnc
P0Pw1OhQAGrfJ4HiJh+i2k1CCTxEDxrely/xkI0+in4hEnt9IsRvS5RYH1K7yrFQRbs6YL8aQ9tg
++Z40leKR1ZteEOVO8dWzVle2werG7eA4hdqOs7XH9jnSUApkSBqkEaYKKITX1OIqVTByzKcA3HC
8RflmovnW0TtLutjiOayJuhDVhc5cjCNgi2Wb8NVRKpFGwkwWQtRvF089FRBbQ3/JX/mIvEmeJYF
MeeClb++legd8HsepFnyNOfSLaNvH9tndPRbuKaxnyvGVfGSOrpa3qTpxTNDudB8zaKjQneWFHfs
dzjUZvjH4yQBPk2+BHm3pX52q8uWiSbGJo2D3+Yj662dGQDjPx+A8knBcYsUREGJb/piff9PRN3P
lPr1TkLo1Z/daBj8FgHwFkJQxgT2OmzV9z3ylm8s+k1bigNZdsm4bjnBf4tqm/6Fz/zbgdbU0Iwe
kzR+ohFE7AKBBdDjfQWsfXUfCfUNRPvpGQct/rM+NPQU8NS+JagbRUARwlHZs3/WYs3cqK9lyPDl
NZyLXc4Sx1sdcQwLjUdPSBxIxhrEIHkceMtcfP2xMZZrFpdlNuU+eNVhDDIjnQEJRRZSdWuA6Gkl
TLX6veiDMz1yfZJURUKzUgk0Pu4RQ2leriatlQtgvCZg8RLMRpOFBSRK0eLHAW2qGLeq70GFDoGf
DQRQxHGXbVTH4LUgwFq8WuDJivs2cbcXYJQpzZ2SPnNZvmJ+sG6PZg4fCv44fhoyMPWJcB/qIjcQ
5wocnSUfw7PMzg05C6TqsyPqzbWqqBHCodf7IxdPrqzkTXZbAQ++4rsIvItjtE9NCmTOgGomJG7H
Ljn2rhYCx4yNPkZxjH/lz6gxKtE0txqhncMobGgNHy4H6Tr8h9QBZBbY9voRGZ28V9vAAIWKopE+
nbt2KMdAcplN9f7bDDRRTYBbsHrnmdePB8AF/vkkpTBuiN7sdUWkWPwBMvo5v2v/peOWpWamME6e
tQ9eqQTb8PXqIpEt0iaMOvxptKkJHx6kuqu24VjmC8gS/BpZMd8DVyO3GmvXOOu1M60oZdsCe0Iy
t+XVW6qQHbaVhZLBO3+IJ0GvBZx7qWXgdUIZV8p3W+xggjK1akBWh/+es6KNSpriacobxylw50jK
hF5IgGgqC8erWWFMIb35C90WtBScB3nMPbrzBOGVExyzVoHajv4cDXr4hDPH+31wvwMqtvi3ag+E
vXwDQxugFezn6NnMTYBeGmkRuKurobffr24i6JqPYsbGDOsZqHN3LxQCf87kW0JyNLuSBcDycX2Y
44Y9R6DsRLa4MnZvi7pNlJijjJptu3ggJEMqLIApyU6o9nzho2ByHd9zLryizsdZLRjh53z4d7XF
bKktQ5PP3/S/91Yf0fPwY2axPkaAtGe0GRTpozhnRFSfbl4gwjVuXNew4EpJlyhsoppIituVZAVZ
PfbDloiUzM9QXeU/t5x/nHj7AGyw/nPChmNZdb0sTAwhrh4POAjBrJBB1OmVyOF9+jTGe6k60/O6
81H6G2X318+UIDAE83zu5N05HZyBhFAgAMZOga0k+PpNuSGWFv2n6Uh7eF+Y/ocahb0/yiSbG1Dw
vP3eDZspVxRENAJjcqr60td671LvaE5L01/wMAIM1dFlUeaHg7j6jgrFZIhbX6JuDA9cCVz8cQAu
fy+gGmX2kUWPs3Mk1+Kmwvv/wwzVumclCUiRLlNxoW8kSWt9Fhswb21rj7XDkeOv7ZHJ50OSX0uY
O7gxSqJwIoqpFSB3s/sR64U5uG+dFlJo4PsSIGXv50y3rnK6qJSldm4HwBwXK5lRTPN+QVyzR/wF
Bb7p/zhqSHHJABbhcW5Wpq4LERD0j7XziA6lyYefMsVtjOZ/Bjj2SDQVgdVvwqwKu0BBMmX8SqZe
0QX8/aJNfpXXXgOf7LPpSbAMcgD2ZfdO4XvqZH/6B3Jbi8OUD2sxVNG/8o5BCnrMvTZbOHsZ2cv8
omQ3LXnK8qjfT9ggUKG+/366uI03FlyNF8/9n8FnU3yAoEfEEYIeeKBS8RhIEpvTU0V0Lt701rp3
avEfGDMKIZwhYf+l81RsdKVFCYmLzloyvprUjY3fPfHlNFknBW00sNNgjzI0HhKOvibZGjOqpfKz
qe6saTDcusZ68QUh3aAl1tQMMKvcarXRjqP7soTfQdhuvQWQ53Q/VorDD4ML0/Gob3zpmO+Ab1NE
DouuuysmJxp7C/ZHUqHYEphjNfVxvRqfao0RsLsmC51RmIqzBxUwcYWD0VZC3rDSrvrmsGCwt+Ex
5vKwK26lSljPLhfIkABuJkNIKWPQDe1LhZVfbZ+lyPasXP+vnKxeZLd7jkrzDEt+aNcctz4R6K7I
BVvT4EYMwRaAWz/XoN0qhpQCGihsx5MViWMauyDZo6lq0dljpBW0Y06U8O1tOqlVHDoH7Lja8OQQ
mEI6HmRXfaMbgbgsBTHWeYT+i9iuIvhoFEGTyL8GD7t0yMS50A/5f3NU7RjAnpcsiwKEn/DvSGgc
bImgzVAI6kc7uBDLnUQqmbZc9c6B9u1uciFMk8Fz5Pg94aU1f9zHSV1CpAlr7dedzu+6dLc7U3tR
qkBhgAH6PTirR2k7y65UgpE6r6nmqNm/iO8undbl7qS85kA8yzSCRKg2HAunMzzTp2EoV/ozITBp
4h1gBFKStfAO1MQc6H45e1ijdkwJc7Vc0rM79o37glF3k6TkxzlUSsYgstAvclVzoTb1vJeuaSL1
ZeqhTPnjNPvtLuSmYXwD3Hr2To/xiNMjGpsRxHzWJ/cPSw7OgPektAQvrk8dQAE3XOLlUszlhEXz
dP0GxFON6GymAleGgZ9fy+kxoKlPjtWHVBEjqHfRMeHa5M1KmSmMaUeKy/LJubkoXpnGWoX6WCtn
8ZT3pIlkVHr5j0W3uLXhMKuto3ybicA0TCHbV0RXtWmIXvn5voV1hN5T4DcgJvTYXoghV/dwdMKV
OAHYQK8HyNInX89mfZ17qkqhSv6rW8sYLz9l3nOknpO2CtxoXOvJd0NKzRQgz/tIJZ1gW3lxzWqg
uNR7Ge0/gWnvgSqky2AwCjB530+6junCBLtoX7WFQl2e1J3pgI3M68Cb7eSxLtw9+Y8lGKBNVR81
m4Prd/VzNYkBjv8q8VdVEqzs0ZwlOVmQ2KU43tnVRBWU39X06oCda3N2cxJ24ukz46aAcFN5mhii
A1/wk3Z2ApTYwa+5jKOOK43BwB1NqpJf0c2IbHNRI9U0Gt8KBpLOxth28Hb4c8dKRIe5m5hf8HKo
Ox6QYAOI48KOjmaL1NugHiZSJgU0LSw4VsW1D80fg9bAPpM8WkLd6rbNiP0mteMwLGbaX3BiiQj0
aJJ7Lv7+LTpSDFz8GlG1VpWW1qCuBYOJBOZTHD9CxwLZVatGy25LmDZmMlaQGiVOS5P8KQWhwe0V
L+YmkE/R3cZ7FyAm04nKT+jJIcZHrCZC1SSfcvxHyQpLxeene3S3mAOpkSfcCYLncbpGmYX2RTHj
q09618xraRDLAyhMfQvYkejPjp/nZ0hmgqCSsJWbH9VGZ2lIBYoeDqCGRJkrAbzb0uZDXMydjs8J
P1jaJ9Hr4wO30DMiJXlFPTL+U7iihwDcffUO0PvirQ8XWNUjuQdUwSy8gEkjTOFSDaYzb6dChYFA
EXAuu2skhOcxmS21Dqy9L47R/1hR++vkKJX8Fx5OlInvOINh2v2IUFURV5CzEeeYoBDS3HKkI32F
cABQIjwlK2DdnlyKPqAouI2lchv/o22lr8W4sWyeZvymBINLZXuSpZz7P3ar0zzgnctWqJEIJKcZ
jx7zxwIYQBe+pqRaDtr5Q0BPWqLO1pqty/v5lfKYZM3q8wXoNeVf7foDNvJ7uyu8Low7NCFY+EKL
7nYWOejRnsPdh5SQm9YqPwQX0sUfVYE2fyzTYq8l6xGuo9f9KPulUQN1cjy6TeduAV9TceU++rsP
7mqgCyMPcSv/p/X0NStjBeMml3wyBNZyCCqLsYoM/rbc2CqhLIQ6V1YSBu8+oAHcsaeRdiAWnv25
3MCP09Lr4CthrZ8THbv+Ey+MliqBAr70uihPFzgBFjx2RkHfKW+FPkSjrYIsqnrblktLFVVfJQRF
tcQh2vzv9skqcFsWCzGxXUyGYlA/Cdh6BGSB3MyvUvHANVffxVrUgjEdwHULL7vqz2Es1I/3I92F
MDZvRIXMa2pTrajPAeGFdUFviov66g8fpM2Gcz18SCPkhzdUICBCJ9G0eK+VOyjJ8TaLK481dA14
bYIHX3y6mwCg/lxLv9XebvEwRTWs9o+2DPEpZOdC7LCoVMqhlNBt37M1ccbsIWa83iBDXC1coNOB
JP0y5Jg5sPfFTC5/Sb+fFgQndoJXR3ncl87uVmmDTttDK4CSXQixpI4Ktf8DPA6TjzJrzm0eN3vD
NMMQeB9xgSCBSqkUzzjAZ/1kL2B9L+3lmdxi6NlT80Ohqodar9GzZ73OIS//+MhOHlRogjfPcuex
0BiMJa1PFnwljtLNtIW3MJRpZpWlIP3BZoEEIlX523m5j2cmQF/vZLxkCC7ApURmuOjaHWFRAfzj
iLj9J0jkMjWLMf+8qnWWdhAYaAZ3GMclUwPFeoozDl+FcmpfJQxpRcEH3I20po9WUBVse95IAk+4
eMSbskZu2tTe6EIr8m/5E7Fka5e5gxvrVPIpfp4fpbBaXUmgZcnqSZmWAkfOfOFJl8VecNN2/2Ja
qP+GrnR6w8e5853xvVSG2mV81vRanetyuccCiQUSVyA76Z59mCV/NrK97MH18/WtVbj2B1sW5BmH
SahHtxjrcmwf8X75QZGcc9YxC0CIPqEaWYk8zhtnst8wdfzXpdkHsQM38TjENZ2TZ4fAh/ZS1C3e
WQgagdC7cjUun8jG1mg1ho3bQ12XuH3NFguaBmplOjAWU4DvacIq+I5S1sSWZSeQzSnOKn8oxbn3
mQAJq+q+FZGSpIONV/yOys45Q9F6IP8h7RxUqUMiVEOfKP05dZ0yOzMJFi90Gr9xyxWm5z8bOCNS
bjX/3D46cnvRzCzZoNbyIYg7slm+awvzZXSxxI1+EAGd2HPjUEP0vDXbOUABFtBE42ikrvk+1Phb
kW+lt5VIFh9WHK1ebSDrAbWg1P8SxMAYtJaCZUlQB8HwbXtDKwOoiY6flDv3L29ZjZ3K2y2N4tcc
kslnmGvfNAF/xoMAIV+fywiCmxlrGdk84ToZoct04CiOjVdsLBJOrK8CqPAiqLF4YUlN2XPP7kaj
BCNZA3BGIKjg85Hm/eFiuGunrlrPQdqrnvEMejgP5OAoEx9dxPPIwasfrBSXAQ4+hACg4QY7yp1g
JmQgXwlhdRqGPAYw0aX5I+6fDrhaMGtzM0wz4j31U+tYXUbDkV5keioOJWbJdQyboFvnj9ncektQ
94aP/lVcbnyomG22u1gTlPQWYeW+hOsrnkA2Ghe9ABJK6fbUoe/NYh6MP3Z38Qa9olZE5z4utv5P
x8pdgqrmzA30K3pGveA43+39nNW3yHxhdcZOXaUtNw0vxXfOr5+7XJPg4/fFxUcVT92PNybTt2f7
z3TirrnAD+7ju/D9Ut/vSF/JsBVOS+iZoBW49v2NoPegs5T5AqF3HO1cjXokO64loCRGtlCh4C+a
KEUg1YBeuTnFuO0AVh1wAWsBZ/kazh0iH9uJY2stxDIcIBMimVIzac+ZKunABK6PDSEp0ashLWHD
AOl7UrKXpuwNMrE6lrt3hXNIqvq/2AgqwoaT/zZwu42H77X0Yyk6wqWxzKyhHVjuyqbGBp9/HTIz
o2T/Shb42LZUi0NfdZMsK0SzfwTF47HOG/uJYM3JggSeT3JRvO3pGs2eCMmPKOuWNo8LycIov+Cx
Z1gCmWOS+drT/ecr37CtzwZYSGT6BNu8VxsxYpIhysq24ai9M2mEeHz08WmxjLMAMfnRJhoVAL6q
BGPcBw15xMIQELVVXuV6E8PQl6sVKi/UlbPIpvuGKrcjsivt2JPn1JCMu1CvrE1Y0EWHt+uRvU6a
zy27gQEVAC4A7p0pfVah3CUPMdBu0h77wdoY27T8YsGHI+ONjRnB7dL0zEPDXDSCq+FmgIg7Vuvm
qXp1pjaNG5IXQcWfNfMyDG10+0ul87MGCw8GxmT26PACl4kGx33vZunKjio0sODby58VytvL4pGQ
sgwP6MpTgXI9Jjj47gj84yBLa+cOjijfpVd0/SFmIGePQzDeuU3IsAaHNaLgucRWxf8I+y1/Ge5S
/dM8c0VetlVWLT3eFs7DhQva22+DirPOmq1Lf8FZ1J3xoRRErABGRIpGuAhDlSAzN9BZTyZ4VC2W
7joCpcBFgY0J8/FtevZFLjj3DZXpq9EpF5yinpg8PfNxqEtBZlKYCexojYHuBJxnmNuoAiOJeSqD
36Bx5vZWTfT2uaNc068TeiTZu52hP8GHQtWchIlcD5y3toQmHSq+c+trXBmUTC/cl+HEorfBVcq0
YZV0ZHzHRKXLxpvXHwqk5wZd0j67V+6ZkqDwgM3cb+dTxL8H+Twm4mlVvlxx4KtgjE1OX8k3n096
Fph9ZHsyJ2X1HG/mTjgmDAU3XGVf/DS+kFrbmINLZhJXdpzJouPirOdNzpepDTukLWE2vtutFXA4
XDDD3SxfCEqXgCQHJZWTw7XlpFqnBjag5TISdwoScvgHo/BmCHWAPOZe7JlfIRaTJha765IeqHWQ
Lyz9+K7tzjFFB/qhgu4CO7HkYHKgwddipncb5HjAb0nDV3CmayesO1kWrwi64zhzLBDmoBUuGcHa
nc2234lcjoBHEaBGNSc4yON0cuGsugm4F77cHoKxI/3H+UbCm9O+ER97F8BJBFGnJSaT1TGMOmjh
VoirYCz8wsQ0b/5rU/eedk06qyZLFZYloVl1jKvkkyGXBW7U/qsbnfiH11h5lTXgKlDwQDgsPYbl
N3vDi64zpMFt9chartjlIiXEiIB6yCygjp0HqGqlJt7ZZu8mY+yHJ6DOwURcTCG1PJ0BFImz56w7
g3Ik3yNiCaPBHudUpGA4Svols9BrO1sTp542cl9ibCblFWYKPmpZrCrW0CvYrdNmLH896clZtJ6I
uQNVMqy9qG13lHj06AjEvDr1vYmedq/0oR/p5wlkguRRI/1jEuI2RL6p+XD8yi8gH1IwYJOo0rX+
LlCfrwe/T6WV5LK/tomp7fouhEEHZQaiKXc2UqYXAHGbCBnowFq1JvBhDkpxsGnmTN35pX1WHpRc
UjiYWdZzyilqUOYWN61Db1sln5xE/JKRFGO9Y7rdGDkSV+6/dZfX9paxZLOCSU5kHV9TZy0ew5RQ
VHDhss6X8Ojglx8QurnJgd9CwaxN+DokVcYOgWdpzgpWqhAkfHhmWofLfkGdA1nGpgzivkd7X8Q+
5pmYGVSwVpymwe6vPHDM37l+jqcUMPCSoqi6dwu89AapNS/cD928n+DO3PWsItWX1naCgTc2X2ah
t1FrCM/zzxMw4Z0WmXLrCMhw9OkBmbKxSizjYVJY2O+NUUAhr1pN6MvBlldq1YX036/Mfy6QdPHy
I5y1BpRSl6Ebkise/WMuWmTA4zX/XUESPaVyRVm3EnxBu4i5DyfgsiNSC2NFk3TMmn7lIlBRUDMJ
XtXRZ4Ub6bVRvdR4yfjcSFTRLy2KlEIPNgsJ3pYld2FWM2/hhOYRB9BNI9Pt6YA2z4WBHHOCafAZ
rPSA9qDxph+rY/pmKSlVBlnEXyU/Nzj642WYiaNPGsvhSQ0gFrlKp24WNqKV2YRYJeQ7mGCu9mFB
0aYbmMGJOSzy+ZuPDrgWbKJd3I7DaUeym3fFPXk0ypX9xpoQe5kiaLol+OmL5Am2yS8USCsorYwZ
rhPXHNWFG8nWMDUkO/73+vJqfv8k16huroSlxcFEC/48K0gPlhbvEzf7sxUFyfEtt2j4En815h1X
PlalP2Q/PbHtq58bWYLTfZkdz/sM5Y6ofA/z6fM3aVNyWVD+gVIEkYiq5kAfgwF2tFXbN5nWqs33
RNUM23qPOoVsRjffXNFUqMH6X8lrFdkiEuGgXRvAuz0k0Ne+sUu3Tx1yQ3uXdSD1Us4khD50KOxj
twQk9lUfp3Cx5ybhl/u0V6DBt+6HncwmmHJurhEhkWegk69u6MU30S/jrtVibv+cmQaUmcI0p6kc
CQE/63ekSipR6ElYmuWSJ1W1h2XqrCinWOP6qevJjSZNuO40yMRn7wZJZ5XxrauWdApIXeNCP8zL
rshM2SI6iF8TapqQplMyz5Ytwgo3BaMIbX5NyDoGRNtafSsxEZXE4PZpq/WBl894C3VnSEj9P+kZ
Wo+mzHW49O+sbk0A++CkWhvBVTxNKTCvYAK53IWhAHc9krtqINMwRlsiSFU694Z6A+TpqOu9i206
Sa7fP6e/UTb0WAOMcV/u9Cv2HuQS60Bilr79OO95Ucs+mmoTAz1B/cSY9Av+xbG9bYpggywJlXLd
vM9IOvS+exXElMzGRuEolVe4AAgxoqIjaEAUskNZv5M5zQMzyQOHyiPJVb0BtvbeK1oWeXTonjgq
liG/k2BMlFtHD5G/+GEc4ImyNRR4yRyEtqcF1V0PZFjIIf3Y3R3wnrzXA8+5a8Ruzm4JuQiEYEZW
woF6cLtIr95qg8e6SPZL+yhb30FYWS3ybbgHFx9QgPZn6MeS2fySP00hkyRKb5jV+mvnoVluAZ1K
aThwEiU91IMBRM4pNlyAIaqm0XFgqWtwEnRYxHo1qIpvPsmnuaCekB+1uX/wC17DJbyAnp29ffyA
aROEOGcq03oO2VFGkqeguigxeluPTx1UvOgkDS26peZqIuyQDkEgCf+Yhf67dNIx9BwSHgdUXuPC
qO6MUHiL6XqppR8jphAkqGinlRMdojtQwSYSVoiqXFsnDJcNrxKvvSIBJOI2Tqmf/cAeEHW/JDtD
3OwPeshpxMypZ1PnTLPSU35FduAVDa8/ViqVDdWzV4RI0FSmfWjgM60dNLVjlPHEtKOG2RQFnLTY
GM/UY2e+mwiTPG8buKJKV6OcaMdHoze/I0kZ0NnvhXEYuwoe3ger+fVYtYI8wzqk8kbJHoYCCuVB
jl7oGXQ8o+iAEr2HB+lr5l4pNn3zEhA90W85bIruZPcE28wqvBsDXP9r76wBMJsobkHW0nzsN5NH
emYPjA2S+z0iOAyA7YeKFxuRHI3vMr6QGWrCFOEs9OF3O9rqlCoZfUAgCQAKTkiu5+05Ec0/riwX
rz4TnFznTKqCNbHLhuWBCOlPzc0nqHr90H+0sZAemFsEPicgjfvMuQ3r5NAFoCjr+Y+6RjQ/sXsy
KeJ6B9upfc3bU0PIeyzCHOYjA6ZB2n8eesh7tjECXQmrnYl89IeQPu5FkvCfKDo4Ngsow1sfZfBw
cTkIm4IOIX1YMagBKPtw8n0KW5p7h0f7WVy2oo/PEAVIo2Cp7BU0OSLapB1+lYPdM4Jo/hlEwyI7
Y+hh9KhOY0M1oe37a2iMCScyXa7RC21ZiwDVBP4mxbrZQy2eFfKZdJlxgaZbKgyr4R2/7i+rJfMf
e2apL9MA+PTPJPhYRz1k5UGsAdffhPu89xUEhxf9tS5vM6geItdJz2+HpRd5K3+B4LVF9T2JKDfI
+6hFoREKi7e2soZPI0WEKQLlGSAJCkx42/h0JTfP53+kAWSgXYUr2c1ks+9x7pflhptmqy0pFOBI
YyYn29rigUfBlcUx5FoG7GJaWlGOOhg5qBhD1ToUgjAGjJ/1SuMXtFnol66qde2J89f3/dvLFfVH
njDOWxLIWhJ7LfvYDwpguEOQCEjrWWyMFagqVl1uhi8fHUDcApO7VLTB5g3wcMpJ0dZFt/6HboZW
BALdYFEBovYFoWcP2nN+uIAgHrOD1nfYxPCeYUpMpml5auix6uS4tsDSzg4RzNBBRA654smJwVAm
0Pqa125H7vUXtJa8rlISQXtvK0lHed2QGjlO4ZEwYwslRT2pz1mekPijhYGn4zFhzqqbZ7T9d+Ws
D4E/tD2FtomExGEiO3VYOvreIG+Ab6xjhVn3ZIAPhkpHCytoVEDbp4N6oUJoDO86hJ7oW489H5Xo
h2FFzzj8hERYgiyOBIHOcjNSjqLbazFHR67YKGYSwDdYOKQt5mjZzRO0WiKvJAYExIXu5dr4HN+F
5KPiZMT/xHS+Z3k85P8JPVDQ4/297q8sa+LCZ3jaGKFrP88nGxQ+Ju+NUXyaaBwyG52xVZ+CcroP
94UeAvGEWxxpM6xqIhRLUART/b94KNJ4Pa/wKg04GNA/F0rGmcC7rxdGdnQx22E6xq58nTnppMZ6
6A7vRZuWfIEnSwagZXPOWiD6xaPpo4FKv6ZCdP5j/HswZE4PchZeDjIOlmGpkfk2WhChsCEHobLv
dlV2jRQHXMsmf6bcczPviqPwjNUePWbXQV/0v/UPW7Fb86akau96saRZemxtPO4EDDcNmrRjdAlL
eV41vqhxJrnWI2JMdZJln6tMdkt2RQglyjTKxcK9CHX+/K7fUFQ8e3eTm6NnMA6Hl8KP8eZWv4ue
MG3y6aMEQkLEkUijCPNybgSF8GAxDh3iXOx4gwR4RWr6bqyRZa2XnFZeI5FVNEawYmBVkNmg+O4+
VkSHtb5KJcYaudQdBFZ8G2d4SCv2tZ/1nAz1xq4TrEVMeD0uxNvuY+ORA8gpGKeUTgiD8wV6qYPy
iHDExkElJ2NZYY5/Wq0FBCber/OEzPSvR0d/VB8oMXZ1qV0u3vwGyU8GHBIaXG5KRSbpk4aSHt2l
13+osGVRxUwl4NTJGbCfYZiUdn4XGhH8aFABmMZdcdoddbqf8yZgn0Z38eDMl8JKcI/yMewJHG6g
v0vCj5hWNaZKfZdoYr5LxU3M6LsS7wWEBj8CARENWHHQkWipmlvNWX2w7tu4/XEmFM4XR2/r9ZC7
wJ7UChvm/hvSZzi+IHl+sduEdXas3+oVqYpepVD/m7Gzdiv2Rh+mkpSCSEBPgxPvESVnQ3xWGo4R
raB2TieKFxo/6HeAFhx/QmiNnL0LtePvhrlsNlSLUh6sCZfBaj3W6aij4Mbj3veC+4lnhS21zJck
SQEcVOTzPOr/xdt+8dtTelHnpLjiYCrNzoRtFxPhUSQ/BKpu6MJgN11PqDZIfO3qFE0RlyemWXEz
r2TA/L0TbRZH+yaQSyiZ8UdrFgpcs40fVKfLGWn7lcf8ToTyl4h+brgjppmh+VR2bnyxdylbkwZk
CsnoGH+99ttJnljkcaibiWgvzT09qzO2qb57EasB4qCnDXJ9KqDBC4aoqtr32Sj4VASWR+5PV7oQ
+G1lg8bedukgpo4WmrUKBl5oDHKyN0BlnSQuj6+C6x7FG/064Z+siDtyniNNi1EIjrbs/AD5LVip
U5BUpaP/dcXkR5E4Dc/hTGMmH95FxJvsM4Vi7youMFGbhMAbFjluh754H5OKezFgxPOink3f5xr4
rbpiIMdVsTKvjJPGDgG/KLL45WBzqSfPfOg47YdgDwYBWHPhroTEQdNAP1jRNqyf9ZVbhRiIvDTN
g8rI7BjqVAev/Liprvk7sMDSc97WH5bwAmDAHVAl+WfvshZ3QJBh5EOibekHBIdqaNkUmeo2/ALF
cmTehMOp1kMjaARAE3TQkuA+j0MrSJpqh7E41Pnkio/HGSHR33y4paE7TgoxNWhHYW+m3uy0m/fP
fT/MqJEcu1QlmcrncNFuv7cxnrnnGwL1BbReCylDkyAJ4a64VBzXrV5d7sJuTmc9lVLbGYD9mzKF
ybVUFcYcmj0HEH+rK2XiuANRdPvReUU3XXd+QHvptf4NLtj9fCoQR1lyTnKiHiQlERbuO/1izWlj
hKtjX2qQ4ciHF5iKk2HkpJJakmAM1S0Oq/X8TV0oFVGE5mtI3G7c0Xsqs0JDKfQj9O/bYe5JwFJ2
go00eYymgcjPg6E/F5m9hU+pgEv6Uutlk/j5tqoP9cZNDeyeuTggkRUn0Gb+L1JJGFYn6Etchxnp
Mj2ryRX583dRyJBDJuv2mrYhUlNKBeJxoHVsiKBCufAjAOLk4FGMhyNOy7tYs00Ung+IOiB+T4ps
R9ViN1yogkOVKYvX1CKzV9HwJewH0bcW1lhp5C0uhTz6d7doQobOCzyCis8E63kQuhxEdAWEhwFH
SBMPU/dJXjvomnSYepd4fP5lWvcIm/I+NbWzamAs+aZ7MWsEpEydfJ+xbI+sF8Yee1KeoKBuRjKb
YPZD+JHXVhBXniR0ups/LQBBGU1SYGjpkKIjV3mA8q79fojXrS+0hqnm7BmlDDGD1rT9j8HuVVZl
yS30J5yG2Dgf9rpwNppvEw4ibJALcVV69uiVfpqGEQGDjWRtP8yauu5LLqLsv7eGEJRw0LCQ02Bw
ZlyQ/j4aRYt0B9XJvj1V0dqT1+L4B4EuzAw4kJF+MSRTkp5xOn4KIR0QdoC1AzUEZrKMqB5XmrVr
f8mG83uIcMxHQHaACpwdhGtEOrgxrHNZS4lE+c6EU9l0K23tJlxilvexETCgOQGdsbv6UP1cJ6T/
iFf/ENJzvs/XIbLy7mUzyLW2xu7pO44H7r2yvwDegQGCdS1ISoNdsFUryjrTxMfPVZf9qdEOi/qy
YLz3SPjmTygYu2a1cKhNW58zlP8J279zzXM3X4EXp+bR0w0tvN8zc66pgVF8kzGCeB6G5OKTe0uC
lym+Q2LlCopSpK5a/xdoOHZOVDVc2C2FZhSUroG0jpoSdDZO+CtnBc+UjgmkmNEhplvKD5Q3C38M
8VGPnazhBhNwsbcaKYrQF/s/yAyt5zK+PPJAKrnxDLoMt1fwGYqz/5HRgBbQhW4Yi0wZp/r6Lt1A
nJQny2xzXBdHi2gYVmsGIjmCdoEJUwfuvQs4aQOtXqOA5227WKC7S8lf6n2iUetW4DMNg/S/4kby
aR6XeQAmn1m8kO8dRSxgwkWQE1gKhb3hFnXnA/rlJdIMNvJbiC7a+UqesNRc0jyFPRiFRilFxCT0
9jUN1Ij3Uh/HoKrgd3q+B+qF71TrJQNHOT6UqIJuGSbnMPkwQ2khi7Wcx3th8l+nG5xtv7Jtkz4a
3Dr8uqtTGAiZOn5GyAcA3uWxuCip2UBPPQptXORMUM748uo1qMGE83Vkn5rT5+YqT1RxX0h/Ei+N
ergA61xZgLSU648lJYp4Gk/Sa7XT8YXB5z/iOJiDmbAgP+kDlTJqfLZL/nwpeneEieyuZWZoPdii
DKeE3+CWVKuHKtYZH5DDU+Eaa+WwY0hEjD+HkgQOpcJcL7ZSS2aR1j+3f2Iv3b1mBs7E+PBWH5XA
6RGioaFjWA+uLeXI/mUqmaWFJhUGLf+bV25qTcX9uBw2l7cBFcLfLkZWWot1DBtrnRKPSw/Y8aNL
eVRQLAeEBO3bA4fV4j7YJE8vxLu1p+xDrBFHnvgthNrS/4lWyn+1GcQGN/Uv5x4ORheJxBQt009b
Zf+mbQ5p/YxwPZyi+Yq7kNw0xmbhQZRqt32r32axTJ8eYtU2iQHhsI+GTvZNGc/mRpLqqbo6TRji
G9DogtAffPymrO+9LRv7NnJircKHgv2dn7QXKPtvxNhzayfhCwuAZG4ebBNxr30eXPzHlXudfYFE
anvhzlL/3MEuR2SLtbK8wP0XGuYsKRUpHEgEuzmVUjtLDKzjBxeDeBhur5gf7NebuzyJwf1+FYCA
+1FPFzj8SeROdQriArQVTuaAZqUtooqdI/4yF7dpgotQDBLvjeEPjmsaWXPZT1sFPlYua2qYDaR/
K8Jy2ihvo5utKfv2Uc8oI+aXfSq1qwIFK1bhW6BS9ys7OhFubqdIxgqjpAvS/pNmIQUbhCCHHVPs
/v7K8cE97jrtqnF2brtPWQf5lG9LlSWWdaUzHIPOunWdNu5Ozx7rfXz9gEVXBuP9pjby4kISgW4s
eng4RyQe6nm8xTQiXyH4bGC2K523CoH8jnl6n45B4JV1fi20VjPkc8XKCBIkIIZmkWuidJa/lO4D
bcbYG+pYDDNYDBToFt6OBXLJ26Kq7LDob2wMDQVQ4Y6/oprEbnXYBYOsPc1+lrG6iM28JHj/Qmec
dMorfwaK5wF3i5laGiIFbGfzC3wDMfRin1rfKLraCVK5lCJPBjh1W+NW3Bw2bgX0sS4GEeJKUO6A
ZtD7pQLo3ima0hxJRibKCtW/mB8Zs/9aiaxuKi/Q4VxBM4TBH16IojHFZelNxcbkXrK/Fi1rCcoa
uYB1V4YkWVhZucJy6bChctGbGfBC05o2sR4ep3bJFNX5d0eb/rpvLpiMyjRgD8xEHwDhTSbdo1n0
ivlHx8xv53c5y/WXPTFbEHoSoZIER4YUfN1Ea2OaqJs3s0VEs5VngFRDXteRUNcnOJ7+VT/s9Qux
0B2RYx5Mz77IS9ZyYHyYLAxdxbsREhATrnQvx5jJ7O7dkytFH+eyhy0iVQ8d9G1u/pfW6GguRHY+
m1buaZ9eOqt0JJQ8S5nArffFN/lYhIixikIpQGh4p0vSbNB2HLzpRGycvZBBDM49aIm0UoZIkyur
LndJs/jmGLO4jeRGL0CPwBAQPB/2sZXgxfarzMRSndxK6uistnEF9nw8FH4e32bvXvX4lJGrLnzS
W72hqREkF1HxADb6QIo2JMtoki5GyOa77NlLzpuqlPbIsFR2XrmQmSpJD24J7CVdLWNQjTTBqOpq
vCmmgSOOnjGKgDqvRDfYakza8DZn8Hq/u2c+mYxTyjX1bfkX9QsX0esRijzfI3/eP3ru1VainRBN
fL2r+vOC50pHdYW2+W4qO91oa0aMhgRfN+KzgjVt+xqSNHxYVUI0+mzE4oQXJf7Tvxvy/W9KW00v
EeqT5DDn9m7YlzDbyw8tvjE6MLymkpNXv0T49rNZ53uvPGHSxG6lcSeIsoXlVOq5weYk8cC8TCDr
KrjiwSIVs/86QafE6MWhA//tNO0HuQnaV7ESgdCT2zfbWRj1+YhtxduiUJ+3OBUf7PLuDauwVfBW
6F2C+JsnownqllGxNouLzPlpFDc8raVVbU/quFjVIY/w8h/hQRsrBT6+XlNegoNJOqygi2U9gzVQ
DLEG8YiEw98yP3++nkEIwQJZ9TnG1O1igoNHNSwuwmeyiQ4mGJkkOhtWSSM4gTQoZY1WAhZNzJ9e
lIl2xxJtzrE0ziwUFCwQ91ujpm7tWJRxQU0QbybQdMAINBl6wq3iBckDumudZ/6t5DCK2jso1vAj
/Rr1MpgKAnUB80XOg0+rux/y6VC75IaoYjI571HUpT3LP5nTIsj+Z0TYcl/5TvkXr3tgV/TrOLg/
2FoppMv23FVh7s5mYkoCMKS7G3g55uE4LqIW/bWP14hnZmb047exaIlzegWSBqnadOsUWqjndEkY
bn5lO295L2hM6T7vLueOISijLrTyPOvGg2tofPztj1mLNzTKJaqOM5hL+o1AKlyUcxg9VKfW7E+a
VUmbkouJEK8lXawsIKZaHrxuvNlEgNz4rtghHUSJlIxjS99qgjYc8JYMXBgS3mBvOazX0XCMEGHY
UVluH8t2XSPRLC9TDzJ2ZsKoysfyOEwyQonlp9BiEI6Sj6KLJICMWaGFZJt9TP1o459zu9lNBbwV
zl3lw/fY1wAM0StGPkJDbbyqE+J040haebJtyauTYaHa5lNyYiWogqvaAGjIKocqgsOhQEZyOiEr
ZczWLCmb/5HHWrfy8K1Kg+CzcsPeCfuPL6BMfTWQCfaAI0IzFPxd8YvRhjei3kUQXx8i8FywiyOR
ASMOEuCfgBHojCyDAJK83+EHHT58lRykg4bi3ZsYhNc/mmzfNhV2dnNITz4bvvnpPSdgujyevFgV
TXXCH6DYmdoObFv9Xx7rU99t/QBDul3UmvrWwpRLyopoIYuhBs/KZfX74MBdCP7X0SYpkF4VF3vw
LA1bFvAtUt31k20QPW617ni2LQde47i6CkyMVSR7ulCmKe8H2ZIZKJJRyKV2g8xOv+LDLTVYsiwu
sncDe5Z4r4DlxFI1vILva5rvfkd35YVt9LMP7y8CCoTiHufnuGyKSVy+YTTfTSnrBqkHLRm24Ocs
FqTSFW3n+br9wJS1eH9OEAnRrl7PHPlqZocAntmof4YgYT1gzUvhN/Jtbra7PKVewjTjo1riIYjY
qbP1zqQRUOqPtv2kOrX5I/1T3CBCK4YhLkMCFpVbfQ8bCDPTA19j1BDxuFoW3ULx355uyyemRtGq
LLtu2+zU9UwXne67tYsvN7jALOPOfblvW55JQfHXU8xAkU4LaIUw56M8NnN6QU+LQD6LxCF3I1Gb
jszukkA376+1lbBkt0+TJB5cvkPWEzqnIpqd/KUVRsesP0DpYzmqAPQQwT71uMHkP4yk8oAjnf0G
UPy3Snnda5TWZmPlrJvXqg6e5GLHAtEdTAJYwqs6MDnxNsBr4ATMHTyGMODUy0n6JFN301GdCjI5
77gmWkEr85/nxo2/IYR7iULcuSOmdaV8cMu8wGGE8NKIdEAZA0dk2jXIgTXzAGuSo3WKABvhhubV
hbTuJpEFn8Ev3tEp4FxHXFfQBr256s1KjU+VTwri1bS6cTRc5IuIZ3S+8MCJYLa7ThnEyYN7hpc5
QWtDg3ZCPAJay6h/3FQ4MwHuZw4G5LP9ayMiMsmmIVDTuxqaBRffMr6e6gN4biHVD6qSW0w91zXH
bdenq98Aipdmd0vYuo6PMWUQa8fOAoiF/+3VLg9Bva9X6wOG6QnFRFLxODFRhZ/gUtVT+AT+DNyo
6zCr3OM2hXtAUml9DGeg8N5qb/dsdqsOFPgOGT8PXiQIL7Cdjb4qREfgvNMKnfThTD48+LfjNpVU
W7Sk8FQnWI/7mqwAUQMrZbxnF87euZ2iZsX+1Uz5iXtAac5xNqhpjl6/Rr3E92c0NpMjcf8G4ZjD
CNHUozJWP5/P7TsS9J5oWO2a7rubiIO9rKF2YaF0bcT1b4RHJjXmER707xoqG4LAud3nkEBKAEhL
7kMMSEB/wsYI4sVZ0KceCGeGmNRLpmcUEoE6ii0caIGKiVZFcvVoSI6aTifR/SmFyk2ZbTbkpXdT
zXDo6pDY2Vqc/qr8lRz0hlU/yTm2gyEuPGPi3LJIyyO3lCDthYYt8QvezgNpaGfuclPh/8s0WWDH
eHjKy8TdAbfPJwwfsvLcjDWjHDAM/DHZn1NHkD5LoOrvZel6rsJc/jSabcJgwmHSEXGZxyiMQAuZ
8W5Z7NhgwFDg5W/G2f9jnSCtkkNFWAcXMvJ2XctPdGxD92CZM/pCH5Y5HRGp5agTVMoq3jav7gyU
sN3SFOlPlcngWehohFZJ3rgtC+mOWMjyFbhYlsFcD43u/R0o7g2AuG7lUKIoHCLNO2v0kBeod4Cx
5QIpZy+L6+sbh+Z66VxJHdsrDj4dIeAkH2j8vsag3C3VMn3IWryaIhO62HBYR2HsaTYylSQmhjD0
C9j3YMwcbGzI+1NOvMqXQZCJ4meU2inMeP7KqgvIiPRK6ga2ba1Hle4ZfdezkkQD48QjMSVCfuxE
WA+8U9QxBxbokQL7RYgUB4pXm8KA75jt29tPz9plw29fRiBZ6ZVRct/4i8YSnEZ4xgOzUswMPy7p
aJLmJstceWSB8WZdEI4KKKs9pmmcMt22q6pYh+Mp+j6eunQfSQxy8ujQVHO8hWgEQxCx8ae1zFWg
cbsGbPGCaf2fh5/9tMdMQM/sJXAzLPE9NVNd2GH6tMO4iTa2bgXCanvgxb3IW7Z9xOJcO1PD9HUF
hnS3PqywMOC9OFoogaZ4JOMznKvT11l4pMQ3OvEFow4tGZm++jlnLzsNhf8nk2k+ehv9z3BQbMAX
gbJyT8iniLCoOy7WQF88mtYjjDS0MP9rfX5B9BCfKT3U+BsisFkBVYz/qpsAg9UDfZxKzTyJzApu
DVA/dD1KidmRmuN0qOt/hPsEQ9ZrR56j9KnqL/XeJRJuyeFtnBBSmSTFi/GWb+eVghg3bYCXG4jh
gQB2d9M4e6Yu7FJU1NEG2XEdS0rktG4jmY+xs4jDhpQ6wGXHWLGUGDASNooHPqIal7pAxrOVIaPL
IoZgpnziBzd7lJ3CGSOovCIPmTNBjrSCwuzx3eUAzscoIXsPNoeWZ4PEZH1e8ZLwUXEo2O10deAh
L9utj5hbbeIpNOHSrDITtLcY+SOuajzOFbY7KXxJA8IG4L+olauVPNm/WWYS+Nncz/aw0XxDskLp
Q+VTZ6wg3DiOM1T/kzjNRKRztHJMoTnk8ceGZRwX6FZtDyA54c/22egwINz1tOZQTDm7YZWV6hLJ
oEo4lpzUuZ4ZnrFEyoiY4G3edGaC99PhPxRScb3xCurrrEKTNazmnecJB/y+Pzgzc55ox7/3Avfj
UmIVW506vWUEoS15wqWp+gw7Hi0Fz2s4IKgNkv206E/ULpHnBesrbiuQLVxfuc6z7gHetz2kbRYe
BiySWlLOcD+mgXjNbvte68f7X3m7qHGBBol/sBCFqBEG7L9+b4Q4tEQRvZXvzWXTJfuVq5+nWaBC
V9+I7zR+KhQC2/OPdTXRu8XrDkC+tsa8Ty1penREp1OAlY4JvWYx2t8oc2T+JLiGdf0iayCyJAxi
JhJNmk/iCbQXaB51ZjurlCzKGj+UDq0KB97jcRgwupIUos8H0/elNS0QEeUyv8iZQdPxRN9K3yE4
9tiBQoFitZJDx39P59TeJuntC/jvddM4r5xwmSf99SVPC/M2AIPuWXzEd+XeACZP1D1WwNG2cN4W
hFGUuURkLz25/l+otQMPGKlHF7lwUbG0hnjPtvOHVo9Z/Ibc1dmmbVyFxtJdUzKd78U1yFmGLnIR
V6N5FR97MvKH3kSJN/SvuLjQy8sJ86LZNaPSxx/MJbAKgzpGau0wL9aiZLt+YP1XKvuVr6YjUvwM
eIHdMbUdo9TNs6q8bitPu7ASLdiNAr9um0/uOPb5wTyvYfU7Cr4dL690Ex6yKd2LIEerwMrAzL78
NEgT81SAELfbIOW5CYl68wyj45CDzrBeEONbaOuE+JeYfP6JG6+oI2sSSvwpmluHUAebEjc6L4CD
fFVHc619DPykFtZOs8+4SfEKFSrbSJLxuitJc7KNPD6J4p7Vu2UtfI5NVbyYZd5Z/h7IolGgWkyT
63tjCIuU3BIOQzjaV/q+JeHpDdCReAm8JTUlQuMc97Ms8mZa8pjaJbrAB6PYxqAq2WaQ8OJdoway
ULmJDvm0mqa8gQv30IQslW00fa7VAFEAGkwDlI2m4Ju10TA5JiQqAfEdG+NQ8HTjJblp1r4hoqOO
0I79yxOt8Z6QEge585+46mayUQC0LXk0txOUf7AkRi5t3WAWJF4YOSa4DkgO6h7iqfB5ov5eXxrf
3rvUWoU3l3CXwdEyVyHP9VUoHkGuXCabehFBxLAi6zjdvl7jMYs0Vm7FLiS3LOuCqUoe+MkVtvdD
EUCp8eCPHrpUZAcCPODOIyzbmGNvHMU9Z887EBR6UtaKf5eaCLeubPip72VvLuU01hgRRmkdeg+L
yS3yYxTZag3gxsjgsVi/tcNjTywAD/V7an8tCXmKvC9iJL2B49JOoSYulDGPDJCfxvxyyLC9XtD0
peDhVd35LOzlDyTUBP3ahvvJmMexH8UetK6qYSqc4uE8gOhyJMaiK9QgxSIQDYjPQIV6IjJ5mWHU
Y8Zdrxrn8AbA+5KuUcO7e0NIkxANf64vlrE6sijHPqPUC4j9KaNy48mqkb9QW0sMr+APxl9AODsb
rPnkMb96lcr03klmX7bdAAQm6+pxjUARcaBtbAzThm+QXkMr8bP7U+pOr2BaBSuxpqfqI1k3paXp
/f/Qz1NQctuza0tIXjqUMLhwVRyKdQILHhYoYZohKmKg1P3W3b/2I7VxhREckbph22J/OstYte+q
bA+CZn07sjm/ppNeQHTkzQblK1G+Yr6KTu0dgm3/eHqUSlvuaYzx5/gCbHCw3ZXPWEa2rD+jdyJX
A9IIAdRpdn8fxdeKP388ab86DRYgI9JZmv8UnHnZIXyd3KddIYX05L37H7OP1mByrvtMg5u4CDXi
E9+jvMuYPAHLhvjqpy6v4U+itkYJ6OKrBjHiAwzXIm3jG8SvTql732+hMQ3RTntoliZ1yfqZNG27
mvy1mXwcbC2aKPHIMKDo3gYMmN1G4kzXuXXxZUFVultQIddKXfOXjwI10hHlPdlHO0kUyyG9/Ftr
4f7jMk/S56jEFckjumGIPlf29/rIAzuqfTAt8aUEUgckBFrWSTVG85vkZTIE8P/KBVBvyOamIXnX
7+FssgvC2s5Jv3CNFQ9L913dUX3JRHFSnicYJxfytbKAopBxr71oXW1NHCteHkAvdE/nqf6CfFKI
Y40O1UzOIbasExEQ+c7Ptber6rYHbhdayeJ9Uck577sNY7cq5DwCgsB+Fp03J2pCg2+CbMFeMobi
3gHNXihq0YsS/mdUCfNDr/fHn6nFIRvauvl2vvpTPUnSQugFRcyCVadGWRh0zgCL2xEddksJryFj
MJpz2qkuTOGlO2tGzVhnv56rrlXcrkvrosF2nfMi6dMho2ts9i4LXwlQr7MrYUr0FZH+UANvOMbW
YnOuG4ua7pF0anaxMvjgYQPVOyPqJVpMayKxdfgpxc3E3xBMiv4jleTQT2n6XpLXJEMlmMu5Mo3h
jXEwdX4gOdPqKZLa0YNVSr9oLkmANp6IJlKfu8PlVyjwtOZ2DFs9EsLPtCl7tWwXz7C0frukWSF9
r0FRBV4z8rUbV4reUjDfzps12h8y3LZ1vC8lKuB0WDlOx2Lf4t7WQpcDdwfkpbIc3nTD8xo6lvlk
EyOxBDYxkTKsqkCXm44DZzvNVIO0ZlbcxjPhL41+mNJEDLc60RwB0y6IZ3y66baggsZLw7vsp+y9
nHt7MHTOMu/ZzxmB8yl9vfYGuNZPbv6ZxqMVOePkvpgeds2ObDq/C1nXZycZCGH22QHwLYkKa6yg
FYtzYSINvp2h3/BtcW7Tt1al+/tXzcJXWTttem9HoMQuzttCYqWSHlhyB8ns7w44k2VP75nsB6ik
VS7aheydNkYN1x4xC3ycvBRSdpzg8RKKoUSUGHitDKKUqIgD1ZePBAqGZkOBZyoty1Xicn8ltsvw
Bpmp0a3ERqLx8Jh1zK77/ntsEnxI6FJ6hPeJSLHWBciY0P2UWqL3w1NT53Twd6yiq4SmhHdxzQSM
/REIr2z4nCUwlTDcLy5xCB8bo4tl+YKUWosqDAhMPgZsp45QMksU54YS6juJccCK7itrBKMzqj8e
WlGQngs6Dg+n6mbMBEVuZxBBEDci+uqcoOZFJKVtzyZEEUbnLLR7euUBm+iAvtTiNj35U6qqrYkq
pw6DZaYl+8CdLnTqUs8UtkDf0l7BsXquLqToU0aHdNaut6n3Ad2M24KELbTdWZJ0hGrX+RbUqlHs
LwFO+kpPyNio2GHcEmbHlfY09Z/4jvRXH0hAPeeZK/ufywrPFrg1nGfpqOjHwWSBhDzP3xJCxV02
g2McZqZGECzNvDRcyDKDL0cz2/17TEROK0M73FOA5Z0MUNYpxwpAqo1FG5zrxA16OooxGq3E1ZZW
8+ivOdDXxbtVgi4YYclK3ESgjWjgJrIfYNHZPFSKfyB31fv13P1SlgCw2fG28d9mNeUok0e9F5SZ
9OtUrMW1C32vLeEQSgE6vJIkeRTCxxZAXue6FDSbwN+IGQM0aeIk7goZ2lLsRoYpwWCm5xQvux7n
1tWXtlWkogkm9ksHs/UcNvJE/wEhH8g6uv1udaMLBvDm5FnCA4OwowLs+8FZLsMQOp48IZ/VEES0
NxVnli12F75nS6nGH5TF3FoWFW/JxE7HmOEuHaYPE9AIZErsjuhPmh3APWSlH0tkbdX2KHGFp9PR
DfYkq5+n7iIDisRRzE4P78T3rlIPu/4A6K1eh6aAIU3A+BcJeKvqDgaDEWOjqGsTW7jsa5XMi57y
NiQss1RZPXlaZjZRCx3e7knXE//pcEHgHz5Yr7h9xvNuWeecK3bjonEpg+zXOTy2dxs0Li+HVeea
2JQ/B1J1sa+oCR8RJ5m8w4MpBD/OZ6gMbP/HdYzLwifaFYvZo1i4rijx3GfWfUk7qXLKme0Dc/BJ
WVpUYqmAmWcodEFCqdz+1W3jcmRYdOZcW2JT8Lp5GQsBgJ9ZjjIGxdvA4nvX4ANH79bxvioCQPcW
E9ISbZW5Rh12+jWpRdGz5Vg+KBOc8eMwfObzhuoX4K311fpIhdjkglrjyFL2YoiZPsqd/Xc/BoNJ
37yJ6cp9sF1YwckKPhkrAyNAsaVPE8NfB9ZjpoFiAGl7emRqOdgENk/nBsLq1WSzwpY8iN1CvXDT
3GYRNMXRGd7+Is6Gpf9mt8MDNT0NCouglCA5RJJckB6el3R8fGacoBHouzPZcKOLc89kFJHuqm0W
ifmJEZdcfufqmw8kPid2cVZM+hc7vYHQTDbIeAl9xckQQahkhw4rSCABJeMG4MP3vojjmqgkEh62
WHzW3P7Grp4Q4zxr60vgi+1J9GrmPhqw7fkw4cW43+SOcFw0coDsO5eQ5xOHzv7Rmgs7u8H/r2vQ
zzR9askVKM5z/9q6jy452iNyRZ1b4NreYom3pzN3SiclN88r+MwtZq0hbfP1//EzbXmt5Tab1tUW
xt2OTwFoALXdM16np16ScqTUZ6kgm4WuijsF/nKJQ/9tIeWCbQ6UxEigQyScDI2vGl0/3qgFd8Pv
kIe9Z/CNG/zd0WBv5ZNvoLgV8h7VBMHivPrOThJhTxMlnICAhm5LR0EPOUP6SJ/pkvv5bPoOGTXo
ezZpVjGoZWTTsHwiEhI4Ip2F3LfCtpTrGSjxPv0/A1mespprxbCYM3he22XbkEWtmvt3RdHGEiKf
Jrh27+FR5UDI1893oiJdExkoQSoW00PCpv3MxIUhUduj8gi8WIpCAq08seVxKsArZixgnKrvspux
eg26IAxSTtzjfUGjfY57nIlu72bCUpxU9zvbJa4Cxuh3B6oRSPOfqHthEdet+T15NoPrNNQojYug
5T222yh246nEQxt1fpwYbIwMTLKPWt9Y33qXktXDrhZOhd9sXXjlg096bmYtaFegIBXlepV191u7
/O4f/Y0OC3k10ioXD5LTZlnq7ELWNMmJCGx5mlxLaUSj5oZlRpOGgQfQmUaJr8mfn0suQYO2uXea
S3j8fzg3+LYqVXoSaSE30ODisCm9Ovl++mjvBjMUwKIPliT1w2vnp406GbzDo3sufYqzRoxCRmw/
tH+6vmfm3DBcFCkDVgd6pCcAI+X+q+JwseLcnjt99waZKOE9AQ3hoO+DRjlFYIbcrrSaMW5SuKJn
2JqPAuw398vwII6VfBEND4plgm7RbtRoEWLsox8JAEwF2pKfCj3WDIRzdq50N3ckJ9Bm5xk4+RU1
HSkJe+CY6tbRv8SQ1upVBQsVeO2Kp4HGN6iVL1sgb2QRc+vBFxxgkuju0QNVLpWycg5ZzGK3fzlJ
D/uZBtU+i0kwR26CYD9FzQiGnkWuFaE1NY5CbQm2wgwRiXM5MQ1oJ3cZBykTHeglcSjzPUGVwoNn
UixS70ShGOf+mk4XLlt5CUKukIBF/SlygESSat3T+XylOz3MExESWPyUwtmI9aDU0GLkQ7XjI5vx
7kkAb6zU6IBqErUhLmKdY5lmBkKxhfk7JzdQsyvFmW/dowte1hr3KGvxQatL8dGMH6BREnlNSbqU
qO6DArh+LG3nilx9Ev6vlHI0oauK9LKCIIBZ0SnPqpPY/LGaP6B0+ShCB1FnWdsJDtBPNln3a/h+
NtmTXPSZDU8P6uQ99K9t6n7/P3uCdrGJ4XDBhzxyiym90LoX3y1DVxSP9IFpd04yCWmjej6wTm3z
SWVpmOLweWH+MeTM1AuoO5ODoEJ3xkeARXOqzbEy8xNQ3l1uPbaLzfjc4zjuNffNzxJbLI1f8pc2
ueiHvryforyvgt8i4GU61DQ+FOTU9ADv3Hz/18gRsu+rEuvoo5312b5+Jbam9YugaZl2PxNF8Yku
REzFWW08cXgfxnLI6a3vNXf9PgRz7eBFOPVYKlugGdgA4cTMS4a4i/KwrxjRK/HvyvTdIeZjXB9G
M4RVdTXAQhso5rbe3x70t2WbiXyqdSu5wz/7pMff6jBHJexa18uC77S7ELgSfEOr8SmnW19RCmAH
ul3u+ufoDIyd471DTDnHF7xgK3H/hIw/nVsPytjlKuNZwpl+uAgBvCuLbxOtZTpzTbbm6GeXv3WW
vaztW6cvb7xx9JAQRdn0an21pVK47xBjK+H57jtiHORXl2vuLHFxYSeGOilcwFAw9EBYsq+wkFFA
gvIZEO/MDOMriWB+AIIB2Pb4AYgm3aM5KuqGlRcf16hO+elQBuA/IG49sE7meduGrCmGcZFm7gjB
x3TL/BMDn7MQjzIURwuiu3FB1WfMDSVa0ZmC94BSVpF4DdisYAs/LuWYL9CTg4y4cpODL/I1da7J
3ZDMYPbr2a5WKCibpkG+zE1mHAPJIP+Zg2xDvxZxuMCN2sDY1kQDhKO9Y7nPdSI9g3GUn7K4HKGy
gr41VcPQwVjVDNFfbvrS61vPTA8ar05DsE4+glNpVHeyvWzAyfgK9+47OL18GHJmh0RNT/W5wvrs
vpUNBDS47oLCNbS0DbRVz4+l9DyYHeRDVR1yP4qbjTE0V4iERZ9cdWGAQ6LKB9fW9MVnFG4gNcMI
AIV9HiuRnNg+J7nPgGVZpJAS/m0B3Re6u56ZXhTbV64gkAmWATlOsZ4nKN7RwG9mzeT7E1g5C4W4
5VdB+8W9FbMUIh9N+Nh4S9a0YlAtaSQXxGEBU+ZrQ9P6Hr6P3VNNHiUWg0IgcBvOpr4tfmE3p8ek
eoqoNdXvDmXUr3JCjI01H0Aefgmmso1lztnIJFAAxV0rojRYxTTGv+DRJYzu8VIYq2hbomkY88nL
asd9dO1mgQ5SJQRodAecYs9auO5ep0ZekvUH1DplAEAfTPqt4AgVUTFscQ1PHuNmlFMUwV18Ph6m
QJQqZ8GXqsqMzpMCawfz7ntX9iizW2Qr1SOODViWJ0GY5aIyhMm3Iz55bz5uf4dX9+zk/0oenu2y
MFjvIpKoTZ9YWzzuDGCtPZ+wtaThCyNakMS/NphfPLms8lhrgdORkrwvxPQ/PtIwxDUk+puUp1dB
dbjeOdSQNJcEo6VgXg0jh8Y1kNNbr7Mtahs48zYGNyRF5dpgULn8f5wo5ZvO9syBV092Zf2bcwIC
OXSKje9w8nWsGngJPPpieplF4HB56esgRgGSCHKsa9eQdzUnz1+LF/olwFamvI35E+YWgtj4ijy2
o/9kTlXTpGHs5RbSSoYKSD6fUg4bQZzQcr11m83LRRH9AxnQdesFkkjjJO6NaowyEYpa3A016ioP
uFL754SlyyOKWag+0AruAOiEBR/vWM3vIlxg6SB9AastFkeQQgcuZmq5LMPzr9aONqray/rSE3sO
6x7ijlSjBe1tbzVAzskHkkxVpuw9NhlpyTcvLuL3DLgQIVjLLYxW1HfnZRrUT7DCekCRYraHE5NH
0brZQNLfK3cN8HElQOqnDwB0gLfYyTaFawxcHTMs6nqeRyp/NJ+GTVsVH4Jq+/Vw4YAhBb0B6cTV
Kj7PnWQ3Cy1b+oxQ4luwT82vpoc9rR6RW5m/X1EEhX7IxPy6bH5TRnSPNMsYrW//X53+JifDwAjI
kfYxdrS98hNdKcczPyHQygA6cnYDtcHmOVmsxdZdqgtQUqcvUTyJeujd3PIHzyRFL2T5TVAfnWAX
s3YrC7BA3fnlNHzZSJFxCzQ+muLEV5oArrPt47s1ZWaXtS2csLn0ObhWTBelSEdpR+PsSsYzwlpl
UYiAb3b2W6DoXQ07rWLwUACs76Psxj0TT543MW9ZBk1PG1wgdHCZo8cPMp2MALtOuyLUdXVA0A59
H2YlqRTIku1iz65qYA8UlrLHLzbp9yVVHE2aw7CWq1yJJ2Wr+8/xc85GNEk+29/ra+vcDP59rYbg
9ZIekRiONpUNg+7pLmZO1AhGVRn1I6sQrrZ8RNyDQ1STnzmP35Eqwuz9Qcb/iVRVh9DstNWj+e9M
uX6BLqULQ7MdDNBsFe63nDLSWXmYN/IN7oNaugz6eWTAPJsiKfRhg0z4t8/6NLeUKzQAvVa1r3lW
TnEKgcnVZkC4T1SWFKPtZFs1QZTXkM+4GVkgxEAmpBoEPuUL2gpB+tbJipNvYQRN5GiMDCboWQSd
KjjM1Qr8XXqCBtBKdE46T2aB5nQFQpjEadro4cKOOuwjGICe/anPbxUg15LLo3cHNdre1FZ6E16j
1GPrHWUrhFHgOWe7CxAlJMatml2XP3fU6/Yc6T3sNlut6ZGGf9FisAkuiHQWb8p1TAs6HAz1k0dJ
SMzDEhwnuN7kgIG/ibIn+KRtD8fRzJxXubZJjiISLUADmdTeqx2T7PevcuwccB8mdjaHy+JLEkoH
u11zO6Iqeghl1lA2s0St227WzoT9P1zWGJvPWgV24mb2MPwPhZeaNI6xQdKERRqBtppKb8m9JNqG
qqe4ga5Arn0cjQG9j8SLoAw9ZX5pe6hUq68+wCQmyNue6typtDH7MLRVxQ5DCeysZlLCPWQgbEqb
I14bBu2bscdg/gubtWwVx4iWNAsDO30OqpDA23VGzgyILko3SUC2yLdi04xR1u5wKXL7pDM59JaC
sabzlFXbm/nZyvrkMVd6i2d3s3XYcZtqra/jvn1saNvcPDXKFqlgn4pyhZt4nfJK4/BgSxsQBONC
pjVkI+34xGgy8b6xN1ze2mlhdikCnX3crFaVYyVQpoUps6EzEAi7fcgr8GPLommd9bYHZpAVBi4b
wcoiIq6kuqSewtouOlEP79xzST3/Rsqlo1PVdXTcSh3z8c2TwOds7V2r+0kzFbImx3certu6ItMU
gsUQD3bA+YOII4tqG5n4tEKTYnNU9RXvfY5pPppNfJLIVY5q+51INfHpgrYitQvLFF1mvrXiKEIA
kAKOKh9+nXz2UegzgCJeCzIyBkVY8Vtkt3UEvaeRTyeobNBPd/mWDD9RAimfe8NyBA87OpC2P/F1
NIJ7bIiofyhhWHmzttn8IW59yQathLM7DCMx4MljwCkO6YyGUWqm2bWq0yx19ZtgDxpFjbb4Qw6K
4lPaKIx1YdBXBwMBIC1CSSnEZe4VpEYGh0E0LWSkK1G/RM9tdKTP9u2rwdnJkIbUvaBriBGT8EDK
OrDa76iLHM8O0+rfkDSM4+FdD1LJo4RYq7BhiA++NQzYgFqRn9UmhKUiNkHUN1LDzrDedV9uVX0K
ZSXMtroQCl4Rt/KbDLqz8PJlJi9VwqXxc2iSg5U9FjAKe3fgeTb0eKep8yhbY7fapY5Ftdkluo+3
TF/md7qTVk/7TvMeTWagPoweO+U83MKMTW37it+UTbebnTrKd5UiYIuHidmscOcDIFNWbIqMaNGB
Tmi4WDGWOk5WlYKP2Hgtwfhq7p2ODwMkoNfKjUkZ/FVEdi2y1nPsNhXZIrgfT8WjiYmk95eQ0sqq
yiz9rZo8siYywu1k/AkexGNzex+XQa9D9mXtbX8ZprXhXcViKpV4PTvXOxR2+PUveQY2OWk1F+Ua
7evUoeTDpRHen42XQvhnuN0wCehJwpQ2+pq8LUZPluypHgcmWxwScyU9CfQ7dzQm9jdJVSUryBWT
RhIEG+VmAyqJ61y+lc+ypxLyVgUwaCXJcNW/L7Mi2DtJCSYjTsezqbZ7LnLYMrM8g6DiRg4RL8bB
7/l2ssnUppJc5ECV41vePYAZLb8j/ZhRL5XRjd+BU/s3L9vOwwiGfARN79gbkJhyZY6a5RkX/JuS
mzXN+1YLP2LNQR+sJIwJ4hhyuL7l5p99ypd2MhDeVKVC/yGkB0W0gOJ2/UIiJoC2Z+xRW57I7huW
CDeLRorbsMr8WES5cgv/ZzGuA2IaS1bY231nb1ojPxeUS/Q1w7R0Arfro24meo4XRdLcMk4dpsxh
jF++yEB5wZj0MDE+eoqB4je1LAfeuF9iGNxdao7AonMuk1Z+63NjjsBOkLGYVO663zlxnUS6Gofy
zwyXKAr4GTuow9a6isQfoSI2wzZ4OEHgODH3gdwwTNKBPm77sk0USz3DYsyDE1dd8pF5GmnXNWAv
i60RbQiZf8FVoPYBHskSZ7DeKhb19lcHg4410maYRwZKavxHqtK1+JpdXOPqxx5oCk/+jpoYGD6C
LBc+zsG4/ycOBzsivKNgomFNXUqASbItSfMHLYcE1Nr/tkqR5wkF+rx29gj5vOo8TNYzmZgGUf6V
VMmon1QK+uudmDmKpsvJ3nEZpSCc4S7WHXmwG/kkxM9TEzYuX8MylYepmJmM6+OmGvv4fR6/PT6y
QE6dQZvM4LzMgqbMA2TM7b6GTXvtbgVfgl9Kll9XejRjwD24Rh9vJENVDBGq9+zmVlIfh3OkH3by
phS9NUQwjaGSJmb8N7f6hHjh8QbB/utvc0xYswTbYs216++VdCM3QBFLFTmInam84M09/vIKPeNI
u8pYsARFJCXfzyRQ6WVZp5b4Fr7XGqQ3JGAVK1SSwsc7Mxmmrmvpeu9XSdeqwO3ay/QClyWf1C/K
zaWzB664RFwvpbugUE+Qop27ffPfO7yUpKuGUbfrgUIRcXN2w5Y4bJF32114kQMtY6vtPV2lu0im
LAeJPilPo8c2BHSYnjv+3BKR1LhcKJQBV+Vdg2N3J/Z7ZTnlMDL5zdO8bqQj5mbCSXuimey6BdfL
cPNGEBJqHFDvoI86wz0qoEGKMtEjEMmInhvBRbggRbmWYe4TpZAJ8t3GGsbsCZwRfDgJtK0HfDrm
Pv3fnqLJ1X0GLvFZm4YAoZ4IKYGDMspMrBxGYFgBJmOdhIFwP4dG4+qaFgFCw1nNtRQfEdWan91O
9ixsnnDZWmubchCfQdEgd9/0dENbd8qBofDnW3vPsFlg0dEYCxSSsE01lePtSWmEO+SzztIqSqgx
xPd5a/eIfgywSWsbFpUea3YIBhoNGG2Yqok8HsuuxktriW/e4HajJdVQdCAEOT4v1nkXBE+fHFRJ
byFeHAlqANsfl9wOTG87I7gycnMOIpKgGyYAmzd6hUlbLPlUuxbsL2d8Ld5VD2uYWoloruTf/9tI
dCuBD6AQVdK7u6pvAyXEASnpTtE6l9c6tvSgvXPzgq8wycSxOYAfFjVFJY2yMC0t1SphD38NlfNx
mq0orjdiTu/iV0LXBxV18BgsQ4PwzTqWAIdF0GkwfI/HJ3r/fLUsdrq1a4qwlYaYswxPRjEuICY7
zpiP96n4+sJATEhD3n2UQ53TQCx7+7slswhr2hkkgUQZG1+ajtigSr9WrfEiUjuTANsR+11+mfiG
D9jLwyZju+zZiLoZ0g7OTT+WFhLp8uIQ3Cnu8CJdqdOpOZjvQFaqBhhpBtlbwsxdIaD8DtlcI3Ye
tuKVMk6AxI/xAqb1oFvKX/i8KvyAlta6FRVRJNeiy23H6v+67LOut//vNjTnxDVJMDQ6YaZwy91q
dmGNltosJUI4vazE/VtkAg5mvUCb+0XgvAIOCT00xGi9CcLy4eIN99f8lYMwg8WqQp0vmeRMfB+5
gbpRry4bGeSjzpLhQjA0u0Iz5LsA5s1fRMSq6Z+S4MKVDjSYMidU4TbyYlmIPo4rxAR4+YnytWQE
lIAWLdLnQW9aMwDIblxgfFmZeM0qLy7IJY3mvlhJYWQUKxq3XqTxSdvtRunEmYcqE0sjJZxzG5wv
clONRFLGVNLjQ/3GuHqk1jejs7o5bH5mAL3kKOCSWZLQdEZ7Mm5v2+tcn57agDYuufJOBdYy33Rl
P1wH/qEjkdllGFYEjrPChWy+VZa/PxBoljWvA4oSih6biJmOmuX578Gnx4eiMcya5y8XrI+GdBGc
FY9cHZMKFgLNU68zZq7d6CDgdVgqD/IJ9VD6YqFD34/+iIZSxa8jsYEKPhgqZZMYTSJWPGOXuL4R
Kw8OQtHBWCvVEUMsn2aOCWFkd79sTVweggg9C0crpQq2AvOVdS4g/0bpMt9+xfH0oYgDLqEcC9Ta
cGu3thf0dJKgMAftreyb5wgjUnULjFCY7p4rN4E7Xw2hck/cYGQppw/Uy7mM1HFNwimVLWX4vP2E
xRp7UMEsmUX3w7rEdio8AiKviuholcPv+3aca455Lg2UM95glmN+LCvXUMqjBt08SQG7N4p/sNiY
h8wdapAiASdZUrbMRpN9/USCvq5b6t8NTpeFgDEw67813LmeC1M0Ktq8D6MErVvnJ/7A8+dGSLvm
XrVyCZkklo8gBgxOPosARKqxYbBtZu9bt729jlvDxcewxNm5PMeHpWjNOGpp3x+C5OodH1kKGMlt
zNOWYANaH4HFD6g8+ORVsOj2BBmYTqlcefmaXmLCbvDsLhTnZ5SycziRYxWKee+DvOYIxFSANpB+
4bibiENKW0K3TmB9pyBmK8tNMcfgOy2tGbruwVjQ6NW2pnArb46hEIUM6hnmo7CJg15p2KTWGvmx
oPlPpIcBu1vd7lqRUemo2s5Qnn8m/oVmdXKlwMSUK7RdKXMu513YPsrizd2pxavtHtwfelxEm6zK
qwgMrXE8srU6RMEikmbDe6vAoFgasUr90sgxzIZCE/7KTj8tn1rW+On7k3ajz/jXBN1nTXdUDe8p
Di9i9dzjSPwqU0tKIba2ztjOELMWpmK9GhGRHj3BVEo6Svtcqn+jc/M8dOvKkRAPqhC6URkmaiQJ
sBs6pTZhyqpS6GRvRY7RCUi+whJVOOhR8qDIGL9vdK8IETBQJrUeOTa7WtOQOxburJ0DDVb4VvPh
dX/vYwqDJZGuPUfRd79XDKPnrAgLDwt+aOeRKVw+1U+bWpyiEJASK064Q1FCiBOYiJ1Nup9jHLhR
kXteckb80QtpbHptZw6SnIayIrLNCEOwgZgjxrpvtG0Q44gvKj26cqvNyDUxfBm9CbLLu51zLAaJ
tD8Jdll5RxhWkOqtZtlfMKCpX/4u6ygbNYDv04sU9Tpbd2JQZa/gW3eX3sd8UlgWIVQRXNUO/0pJ
4jOPo1niCcN+CDhBiX5Q0k2Op8hQJYvj2sYXSZyg/UIFjsDKqAzNl+bBy1QL/1IaHK2M02RAPDmQ
JzKJijDVrXPLkmX4KRvlYvksfqfzKQuBIFXDzTtCs646QnzPOwNuzlItHHYTeyPcPa1G1K3wlcbo
TqNgg8ICD/lNs9Scb/Ubh8Tfz+yFD2yuQ9nRo5cBu0+iAL3npIC+nCeggx1FAKw/3IpLlNpgQpgm
H/rFhIwLkdVttTSo2tv/6WxKujf02yY1Kj8pS+fg3Ugkr9VSwy2XfxxdVyTIObws/b6/0f0YDHIs
MESiIHvoqiv6HtinbH3Aha7t1cdG95Wf7rXdN4ToL5AjWPXf78RPwTJann0nenY7VFY86tR56eUp
J6qZQI5w54KbHNRNaecR/p8scD5dtoQ/k3DLmkTFJrqeo0p3fpPFTROTWqKKzhTIvZCgrUz5bPnY
Q4IVCMnNep0tDt5ymKA3XlfzGfU1QbAY28SV7Z5Zyyhl587NgSILRuFjPO2MWyB/b4yMcodAwfqz
+W47YEPhShhZG7AYHdwkM3R0Mcl/GztDmX2gvy7ulUoGrWFIKmMZPJ31TT5MzmdlkiU4xa9X7JmF
y6kp8g2IKOPOdYIeYbt5KgMv8XoSyj7jKLw9JlQpCUk8WRsj5NEW9AwJe0tVaIWNewMKNU81vz8E
cuzmXOwLxOMr4NjvlHeYha4BGxnEXAgc/F/uBxSd+uzqx+TQOlYXmYlWOKSbVR2vIDwyPCX+W18L
dLTQSxMe/FQi9eaLyKTmFryK2eCaSR/sdKYpDSb0n6G7QRguQ5HzKuZdEmjGONyftwXPjUFQlv7J
3LEGOlFm4VOe2OaQGKrYKhmUxRC9pFzww44xYUq3QMNuL7zNVRtV3/Za4aPuuLWfydJaodqH3BsS
m85EBnwCij+iaLE8OQ7M91AQ7640yQT8tWGvVi1z05quNiDZOqnm3QJn2ETmXLsQlyBnZOcqZ5tF
8Tdq1av2ZTduxqoRnTovdCcH7HScmp98ec45lfQpqMyn4f8YnYHad86abd4FTJLLIHhhkTguJtIf
SZt2xv9rSLoQjiXkecDZQdKYuxltElcxKBomkJwyKriCWdIcHKWM60H15M625ne1TeeA5mC5i7iG
BN1mqcgwcDux6l0AJyybboapR2yPbF2h/CZLCN/ELEO9LDbiB1bjcgLHeSwogz/zs/oT0BuiEzcm
yYE6BjzpAhFxcNHt4uvfBZAu/zg1Qe46+gYl80Qsozi42fRxOIRokml25f66YWeGCGz3P8AcqCX0
avUptn9eDInDVijkSNi5j2t/3Euv64Asp71t8LZO30NhL8o4sxYsVromy5FyBQ3j1HOcDS30hVdB
1Mgd6k7/SK9zZmcW8T75lg6OFnSlk8zbXl1HWlgnDO9uQAo8lwML/JHXt2qmevG4kWi7YhHIVySC
SJFzAA5HSw6TDokiHT1omPBynloDU1DqIsvIJnOorHGrfC0L+BP+oQGZdnxVCzQ8Tc6VPFXyy0Gg
+xuiZhXqqsQkRnnOSO4KLHBMCcHlAckDMUlc5F6Zg/A4+BDINeRxlgs57J6DD5y3X1KE5eHg3IhB
a/OJUVwb1X7/g0EED1NmvDKW4CO0nytoR6iN1m0k/eAquLEqnHOm7CMSjVgeHWvihb7MiGZtScqo
mbxcAf1z/V2/HnCfHoqE/dsmykg/O+b1gxuTell4FpuvF7G0K2jnNilnUdoA1B8iIqOCVotFeu5A
CZiPYKJcyABMSQxVkS/7eDryFhhZ81w3QrIpoZWgUc0r0aRti102y/ubxqIl5wC4ne+L48HeCZTZ
2bmNM5gRBI26tKgDGusa+a46sTWM4CPifLSkkUgU1Ya4V8Ep0Q4TAP+aML9JB1hb0jx2J5xbh5mZ
uRJtohJLsF1zpiXcvWHO/Q/gNEBwBHHpW99eotEasbaElTVyfCprz3pqtVkPxkKb9mEyqRPF/Qkz
Ob0Co4gOBKOJu9GePw6UjwiMdvmFfDp3vmwh3lZktkKBZ8K71ZCdQ6icgEbSl9DffHk5n9enTRPA
ieUdZSEGhZ/wtKStp4o62FLpVwmoifZw3RynBTol1AEIeDpb5uTi+dPMRNFfGJDu6VxeENsVqaPr
3sj9mTJEK1Ot+Gy/KzTG7htxoG4Ve2lcuTzl4dunva2QYih0aQ80+BftDzeZF+hLWU1/ShVdXW5P
2B4xKTXETpy4AYUSHTQVVg6Ci6EybrKZbe406bn1NImf95IPhDaAx2K7upq3U6Giv1wR6XvQsOUO
XiRpuVedJnwviN/d/kL9WFSTKQBMwrNipXE/+uukKPDuU4Zbm1MncW14hWncjWVZGzCtwQ6/K/ik
1KpMd1SstQrm0JVsbOyCFQGA8zk84Rpz96Y7E/yz56+d1dcw7IpNBrjujETQ17D6k4akIIZ/QWTV
sz052sS7gDlyb4ZxNNN9ZyVD0n6/QJr2+qwZW7cEpjvilSU9t+W/qFq0T/50wZkSm4xgLuyVSymz
oRSp7Bpa3t5QLaD3oS1V+ddxYXuwxi8A97w4TWvhpVYvY7lkodLap/GEkHqddDuEZPxx5R3KwWZI
lSxPyNbMmE7V8/S8Lx+vqKNh/xBtku97L359afhLnVd+9ldpYzq1MXVZsVja8Ukk1mzHMMr9M+EP
QKJqOozK/AkHA9fxbh8uzaRhIo9xzD3SCP4OBiWSb2cCIT/YRWgmg2+lmdVdVnYepCwrnAo1jhok
alrxwEmaF5hoZ2aPdx6DBWN8e4xQHEbEoaqKK3JkYhJpWyBp2BcXJH5VRlpAF/4H278vu9pL2ICa
EKxsHlgXr0r1M0OLVPOcMDyL/gS7cTAPLjATRiZ7CxYsdxd4slNB4oJK9zv0HWwXxg2KtjlODORp
U7XCL1dSClfa8xnORhMzEpzTKUIu17MmspQuqzSyOToQAUs63now04aDfvWw8iMFOOkIiuw4ibAY
AOyyN2oMcC5BLY6DMVAkdUedWaS/mP96um80U+kGcKJtXumg8gdgauzHlkd0FaZK5riCxmbg6t4Y
MvHFjvMgzrflm1/XAhxFi6hzrUbVadmOvgQHyzExefnmyAKlR51wP+rNytpF6Ocr+/PBkJDryxH3
9rKvN45IoAD2ca500N9VQ+zb/fzebeKHUZ2llKuTgSvXais/SS6CTIhqks++aWmU5SFSx6I012nx
MqJWEqcjD2lb64D8eWVZNWHA7JOmWvRzBoVodrLqFfB6Dst0uaNnXPTD8t3E8TjjABx6Fv8NJxrz
0dMQ+dENHGxnCDxRzWZlQDj4zchmkT6Yi6612V2e72PCe3+KUDkjjwtmIzIJSuqc9jMx0djgt3kY
ITLxgSu6KGwho5ZVNEM41jDNBAQd6xPKwXP72QMwLFD4bpyGnzxANRWd2NPnI9vM+6o6NE9y0YpY
d22lqHILOFno/c186GKaeOUqP3OebZWPUWUfgF69/t1OoU6LVGXk2CdloqAkVwGNiKiJh5laJJRK
ZMEAzC/bFPNRFVKuqUsvvFlHMT/RqY8bqf9/AgfKScML6UkJwzyWUB/s6pV5PlI+r5rQvx9N8Zf9
3r7EbLvUYNktO8t8PMruqODgZIv8R8Fey3PN9fdoMoIo9o3nQ/kLfKnIplDy5I0XvxdqEMN53yA1
jqBmdqo0IrY=
`protect end_protected
