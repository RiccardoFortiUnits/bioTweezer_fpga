// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
XIzsYBxd602HCqgrNhzNlk04k/u/JqPRQpWjzIniYbDs/MUy82XJ3kqsrZHKnwL04BQJ8ppCo3/9
jrIPvcxypckDu9PjQFmy80zi9Kcr5SRxQbXRxG1q215vl5PVMfeOqdHdQcmQwlAvBXblvms1JQQm
AqdUdJ0c7VymCSKEfjCq9yJpmx4V9AipLo+JJ0Os4a6vpxcxe9Z50uDG7QoQdsxCqLxLeif1Z4sJ
JxYDOD08b1SAXGq68okNB+p1jXSv7vw1z2VKF7DpcfLy45JLKlqDyVZiJYB51p3iWasHG0f15Q3/
9vtNMK2LF4L2bgtN7JBq11hGLFGAe1WU4JqPyA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10944)
EoDiLUCqAuDBQJyoeqGhJnYB9YFiyw8cxQJ+HBzn9X6Y2q4iU+n1f8sXOaKkYBGJ1tRMegxUbzyr
6je73wNj/ajC4wj4It8yWWSRYbHmUR4nxALmngVb2+dcVHgGwKELfV/qghRwAn8xa0wN4B7C43wH
pq1+rhyaPdnT+kbqLkNZO1z5RQfvCAP7JRW6TKy3f002IkGnIytKjo0sHMFF7j6FavxewKQzTG2o
QbKPan/Np1NVT0FAIhY3lwslkLvgqfxfmyKhsW8thbYiuT3IJxWXUAaEUAh8jHRZRwwwkmubQ86K
BbVay8KUfjXyCYHDpTteWXHuGalkp4+fIOIOs1Lt8KCroQtcDJxFxDxejuYzpPdMxZVdEkDRBIpE
twVQ/5q0It6KipAprvOjlh3lkMzNm4HU20TwGw4Qdln8VOdQqgMvdx7oqkEHUiIuS41om04ooO/9
insmO8a6X6dm4Wyup9Xd5TBD2Gig+rYPX73CWoA6oyJkEkm0gffYcqBiOzXRidO2DORThxskh4pC
AERk+BOMmo6SU30oC7CtoksOpN6I0xeS+4J3CUmQYWpfGAU8OLUKFtQCzkizzzwXAMJa78aHeza9
FTIhJ8/DxMKSQ/FFfKaj9lTD2XzVHwGhXWQ6hmf6XZugvEPlk5Q9dEjgxkIGQkvBY8SF3Nx6fWxc
te9oxLejb8+Wd+PctuN5iH724i2D50VMup521Z2Hd/D1dPs2W1Mr5VQHvurSeQ7pMPnPCoSmqPu4
ShyS3e8Dv0C7NyheYRfPHwz8zfmtm07Sf6SZ0lMHh1wjFgqhuBH1+9tmlnWCMXuT2coM1TMd8BtB
NpIQXqlj+H+BlV8MjJhozQ3NY4ZE0hJEnRjGg814oqpHLN2/EN9KqT79OImIt9hP9lR87wndvkjd
Rd418A1uZ/L2L/GaTHX3pN5WZYauhpt5iCy7JN39QpniXagnPqvE9o6PXdIsxluVi6/Rhx14Sfd9
cw5QGKQ2UiinU44j7t416yrgyYHOPXJfiN/f+vTWxilxzLtxhbCTHHk9GL9BppFLN1r365IfZxg7
A4jlUXqMMeSj9O9t3rDZah5oytyW8ZI5BZdyiKU/kavgdng8FiLLlL4rv6Eix3DzWIDzuZlgUZ3M
c4kXr4vgEvWZl0RGqMzAZQTDmQaaHS3CR5Vd6vjeljb1UvjAMitwtjrJY0yZshWmHpo1AdL3mKQB
fCVSG8fTnUnyUiDP0HyoVaqEeEqM4mm7LwIpBrWPDXox2g3SVTzLcBkXhttlXIiH8YsWk1iLw1jE
THQdXMbJj1DVJGuKb4/eGi45ouiLjCtYRwQBF3bV9Vq0tvD80h8gvLsGi2O+8Q0sTS5TA5n4O0E5
hk7WwXtrid1uQVAxYnNQ49O1ZB15sPQBQa58NwoI75N3MDutusNwEny81eAscnz6pe0LcqbRdGba
ArGD5nb0fDWyqpEfeX1dmbsqpYbjzDRImYyxzYD/bUBCqxDwKcxkNMBE35MBaY8g09X1pCpfWnel
sDoxWr26kx8J56Gjb1xqdU4wTytVnNIF8PvdmpfbVdpn9OUd+QMbVJgcjwsYn2fpJUM0qnNp8tnF
8Q8bYYDXhRDTTaAW3tEund7r3r30gfAfGoJk4kyG6B2x/z3nW81CLrxtVjlvdXu1AVMyWDElaqkA
ajepgCUg6iSJH7FyI8gk4/V1B86j+ZJLNmedojUlEPB9lKbeiTtmEbjCQAD3Pya/HkZuw4nErpQr
RvoA9Znnkf17JapocOWT8idYrpqHm9/jKfGbcyrQuU6UDmf8IU04KBqddjLv6XbUBNpal0dFbk4f
8pg3IF+RcrgaSlw9RusEcyzGhNU7l1ViriF5vUT9W1EtaQaaBFTNN4VsEi/AMRDc5julLsgO3c+B
t6vr7mM2lmns5n6opUJ1xhH8OBSSN7ByTZv7b0UTw5rKM4zAp8LTC1OEP/eVbQQQwRcL4UhhIji8
RaXEID6fFqiinaCRmn7CqMrYTgqRmL9OQs2JPLI0yW1Z0SOPZG/lapq2/nFTl8DXiZ/e+Ia7JYbX
x7Fzr9t4HAAqA2nIRepRJ26c/w4J4XKJd0KCufmpvvvZI7jI7/MGd6yNFFG733O+XVLri8f623hQ
d28GZ5zqe2aKurWHjxZ1oeJyV30ReTLp1pdtlccuJ8uxHT4wNdiy9Dx+mfJtsDTOBtc415gDLyaY
Hgzob3slHkROkNlrUk5Kry5hQ9wOdKwScMlKPKAOvztdVtQ9VMYUwLKVV6wSFRYeRhagnIU2PswK
ytBUb/L48GmvQXn5w+3VEl9DJj6UnhtOwQoYjq1a9ov4j8UF3NvY2f6cMzOqFMXtC+BtGcRtEcwT
vvtig3OeTg6GiK6LefOmy9SNaWSMVEkjyb0BTJM1RCzkNXisCcLBCowEAcdBSmFJtePeUf8+RzE7
Nc1c7h8zkSPdBigOOXCorBiEmGlUoRklWK6D3coTaaIkL69RNpL90Lehk9PIl25sKYdZzKUrcpQ8
bXftFedINxI8bDSC55403y7ENjD7jJFZlkNtEPWhtlNI6evmhtznmgAZChQAeos1HnM+uVQao8/W
wg9v+3YE8a9S21yhd3ViySPleUXUhZclZyzdii+T21zoM+DZn1Taz0A1iKqmnZx6srglk96fgL9q
YmNGQUXdpzkMD6AfS6YMgxYUprg0Ugt/p9ZGOLtMMIlOHpj+joH3yrpR1i0wIvwhRYRhwFH9v17M
+cNP3bM7C1oZs1FzOfGbb2n1ReVD3azhFOm8FwAym2xZa4KLajZ56SUje/OAtWu6xpLsycGrsWd2
mhfMryXMu8XJ05LzLCK1jx8E0IoG+7WLf5V6EfyY/mSXRZnEfRJrIFNJQZvOh4iYmAWeTPWa4O9k
25si/L0K01PnuM6Cjmgicov2l0frrrdRYRE8SH5UusFaSUw8YMtJFR+Hzma7hQbtLYE830p/yeFv
hgxxhvb9zmRFyPJidQYqD36+kWMnLigusIyT8NnspvT3DG5exq1wwewSEqyodmF/gv0TeWyrg4Q3
mTKCTMnhjx73LnvBjf4BFkQtFuO3+zrNow3ZYIvFUaMcVx+C4iEvX6P2hR5zckN8kngaihWrEqiO
2q26oGWliFAHOmjBlLjeO84BpPcmGts6Jstlq46C/TPzhJHhrqZogVSdpAFmF2ag7R+LkKy9QDZ6
mifJ6YFbJPgag8biSJb+56P4jqXi35tC1gIbmjrzk1+CH2LB7B9qkZ7X7Wok/eTRt4q6ilr1ndO1
0ayM+s9Evh6MzUVGNyj5tHEzQyM1H5qiR3lhZQMu/PinL5cJBJzQgDaoex3T7dxncjyiVKalUoBp
3XeVyPxkPa83xjjiVPPwQStCyQFEHmLORwkVMBaPQn+YJpocatLijMjNiCKyXrzSdcnwU6y1WpLE
25HEGYC/+qe6gP6sRFu1ScZN+6HqHUHC+bWO/bG6Jb2TV78KWc3h9lnTXEh6FHlQo9U2qGEoRq2K
SHD7obvrQQInLGc63Ta3tq/bP66RCTK9E00F7RqDLqthAi0pFf9Hl/RhGWC0VGTDJmcNj2uTCUK/
iTHQO8/6gLXjaei5/BfmUWeNo2GwJJRVuAbRHR7xhw2cfD05fpPU44P+BHtFhJqLzVgFEFd3i3x7
suJhWLohOaxFEJGlahRH9iMrKgBOznFejRNErsKg4VoVT7AduqO9DFEpTZ74TGZpkymwVu5Ma4C1
16HVyW/Mheh9Az0Ph+rz0u6Rc9+HfBn+zyCIaRWO9GbfafVi/v9SyDpA8WQY1EpdTEKyjczkdIkn
9XeyPsnlzKn9w2uOesUccJ8kSO6PBRuLIrQ6p4EvRYcIthqF5KvQ+evVAh1hibjKHclUz6vVEPMc
5++jNcbz3gNQcnwWgYylTIg2ZlHkY9zYMND0YSdrpxP5J0eFcNCQLeqKnu8heR3oj9HBC6pDWXFr
adZzI5AEiKuP9D9bDnnYYTHwkriLNEw4Ye3DIZTDqZVJ5GGfLpHOiWFV+1n5DHWAOiFlqF+Rc4vH
XTginpjl8Qx7p6qzrOaU3hCfr1Q4nRadGbcJnZQxo7244+mKJ3OBM1ht4wnGd5wOEGgAX9Mwfwah
8fE216FbquBrTd93t73g+bH7Spw325QErKBvnoj5UI3GNcGxwgzuGESAI4eaKoE8/24LAxe0U3Gr
O8ZqFlbmuHnQox4aLuMKfF297Uu1YjE8Oyc/IqGd7rdfiRHkvCWn1Tsor26nXaHV/rSQtymzIfEJ
xZkKkxTzzW9vSIZktJTGJlalzxAqmclXG7jYL0S19ZuoNnPVYqIncCpwhZf4F1JaRncsZj6DZYNc
w+UVu5vI1c75PxDQXYxXrqCffgy8FBpuuMVyOc7l2TaEhAg5PchBP+5C78r33vL1gjhj2cUg9AzE
0Itj5D6bCkvy/ajHrg2EqKQrbBs2GRPjvYSBU/GT7xlYlbKivGMmXOsQVev8tVizYXFjkhm5u3yv
2F6PUhVHTKAgs8NacipfjOtN9visDo0DbhpWiF0vXhouBBHZVKcEuJrqqY/OYIEhdlKp0pV1sy55
jIvaScaStn/uvlIxxBZhhlWg0CLKSkoWS1WS+iEf2li7Y+glP7cOc8pH3aioIXnS15SDScxLncma
H1XptgLtqyWkYWOtdJaxQa4pQrBY26d5CVTezW7gmmXXsssrWYQ7r6Sm0BCVXRdQs4wKAR5CcmI2
hOY+Fe3nNnKtJbiKjjnCBx4jCoIWWXwCfbwjj9T7TMQ5A5QbE5I1nfJ7NrmkHt0mrZ+lKiKoF7kF
HH5DkkyKg9e4za2G1DZBYV5KRolzBXCyhpy77/xrrQXWWZf/Yrb0DfXKRdCEr5Qmi9nvEVOZDn8i
V2Wz47sfuHT2ll6xCok1KfTJZjXjiQWvFgKb3BpZDT8hSnfHdirUWJhy792V2wl5UErMv/ilAcnX
8LdBUEBrUPoloFdKqPJrptVB/88cHBxjDYztR8MAr4rHPbfe4g3tSR0m0bttMF96Rf5F09C79b6m
MGbKGIG5M/MNyLlJgK22EYlcBYafwK5i3gTmAToQpPe6tCO2hmdt3q2a4QRkpRpJcQca96mL7tdR
4vhT5N7qrBYPWm6I2PapMiozxUqDBbWn6NGnyGVhngwT7vgj8V1XKaDHK/ltYmUiNLoRrvKRC1ax
h9oyQ+VmKMCm9VXPkrT9U3kxGg9FaO9toBtYWuTBxjJtLkLttuPH5gm4WrKMVXCHwFzV5+duyI8g
QObyMH6Kk0v6hhi9o6D7pTlAtAQPZccJI6ljBBjH3z0GPMg8mzMSJhKw5ECdn/bUoqtezFKUHuS9
BlaOUOktt/MfIRIBfVG6VrvdV1rZ4Z/2F/0VkeEnaaAP0gTU8vFdG3PryYYK/6IIjZaXbtfhhIPz
zzkF3C1Bo73CeG5tVT6pPYS0EAVReDYx+lPWFiF8csfI34F1aybmZgYfDmR3qm5GeEdk6ZCfGGpX
dcyM6OpFajhZJy1cxoJ9hVexpWPxzYmZdcmpzeBJr4unUN14mQf7Gcfuma2XoBBt52htA40OdGro
rDWnXWRp5bInukqEXUGoQZBVY6qA7cYB8Bw2kHr2/kdvqUEqs9A1S6eY83fI4v6tpDxYw0vqMR2R
qtszJ5x/wAyXk/z74nvfvIU+sOVZyZJvBanEMgOHW95pRaFzhfpg1227b/jCs0KI9MCf+TVksVSB
UdskDXa0L4frXe+EZ103LXPnfxwVPUvPacynrHAnYbmNSM5/Y7xeKhEedNz3Exn7kKtsDRdF0PAe
Zk/b0QasE6QKu3ts0gLzEWyXDA7TzmPmPani96M0/qWIhFuGWFwrrSjFgs9hOwy68JZgD6Zm8A24
4puA094WfmZW3pxc+1gO/unr3AommsI3/H6kmjpw6DM/YujdqgrJOpjWsn6lQdAZyGfGu6OrhsJx
6XrwxiMlfhC4MQw2jr/5svulh+KadcIc2rv3lu2P+l21RKVWqX7MLYkfiZULT95HkohgaRIjFyoI
eRkU1mNdwauvYsytHMttQVchqjpYhXcnGwtSXEisOpUqPsvRKL601aCCmyh1ueGbSmAg5oHjnpNz
VAxmtV/eoWj5NHc5Y99AO4+CTLyBi556teyQXOg6ET3OwJ3uXYk69YoVnkFkughahs+4TrMUxDMQ
2B9PFQbT2IhVPkw1rOpzO5q8BWtkwIAPHazruGJj4LA/3OnEMJlS+FW4MLjq4ZXigCFqiLonox+C
YkEE39wfCs8cYpBHS7HhP852kF1O/h0mupqvfdQHckgcWo6NwDo0RvYgEny+TQFhPhZcfl/2+MSS
2ZX+IfuB3OWV5yyXnu/PdwRuQlcloztHRJ0FTs2qmdxsC+tuXSPKFOO8A0+x3LJkKfdQ2wD31p3P
CGL9j46OU+0mg0KHVwkLgekujgtRq0XeZLrG38acITV9hTi9d2EBwy3gukkDhn6pX4XDxamH/R0S
iiOST34X9gc0FSsVYAXze4uJzM3WSM5k84s6f8JXdnOjYhqgyq922vUUWlBR7oqpnObgPLMG0/Nw
7xKzRw8qp+TTmIQSBn2OAg8YM0qMUrJuiHlRkNyn+Q0WG8xcH20us9hXux54bicOtz1JQ8sFf4wE
5FIKLjiFZ3iqf0LWe5Ow1q7eO4ZAeW8JvVq364bEuq/oU5gaQ6879dvvjrTeKGX/Ku7jyV3a4FR9
yQdaBBVPcEprxMAKT/V0U5RDvdREYWYuy/3jALb4vPI9jtcrim/XC9cG+58vIi8IHW5gWP0SGJDM
KMNvIYyC90YoKYzFPj6MeUIUsl9G4L6ss1BJpQA0ZhqnrL3OGlT+vq+B43eX63vqwy0iWlE92Bgh
jCrwutWT/S57PycMXPbNna2IyOyJn4O1d9lyQjhRf8AdfAxpqo7r4MHns5Fi+1+Rt+e/9WdT65vv
I1+HWboIGMeq0JLDZzTvMeG1PiGEGbq0IytNx5+YGM1z/H98LKSvwDdBauXq6DecLQuBcojuEywh
lWXRhefrC4DhKd7V+uLtA2GvZ6LOqbxtNWljHD5R4RlCUez1PbOmnA59cEuBpDvcuCWszrfy0Bjz
zcr24NVYB2bY8L0BDUVUZLYeHFmX3ThR8KkNaPD5SUsdiXq2Ap0nI0+YiGmuwI/J2exoGe49kJik
RGAMoBTlM6cPBT5bZzCmSZwGGfl9LTlnSCaWw3A+56WkqlGHw1rMcsWuiqiC3TAcqjZI6/ruqPyG
MsNYVVOFOlSDNErmgl2BgLGn5Y1IqqneqbINoYZ/HSG+3ev1qb9E1yYICYr97nUvrEfvIgmZJmAx
wJbtnhpkO5qFn8Cc3MFpVCJ6mfc33mq+npqvnnfhaqJivnnwUAYU3DmwjS0MGTCbJvplw9L5EhE0
fKr8a9YGIF399YXn47mYgG9miGzis1m85j++t6dD8pqaXanSx3ncHZF0TxaYIMjNG4AX7NOPLmoK
ZORFE90EEyRcIb73WtU6gqIeQ10W2zkrkhYv99Fsvj01gmdCGyNVybawz4Y3kIYlx+gZWe2YEU83
pHAbFgzA1bdYApvJe9fTSu52//+6xrsxocILDkz3ER2/06WDPDySBsmebzWf6Izqb/vlh0Fk+oDU
3vYgvMhQt0qVOvMamHO/mPT4TyoLB6WouawbaqdczZizHvb29txxBb4JTpokzw1RlTVSUM9EN8oB
D5HURrRmiIZNnglo/Fxn0UUq0iaDbrC4BIYel1Nziy6FhupWM+IKrMHpyTkC3zzlFXprTNS0E3mZ
eU5IrHjRTdsHHMRUAWvkz1sMqCZl4fbPUGJqqO6v1bkTT0e7ZN+LxgBQ50XMztyogAZ55xr7Wwch
BTvQwcMQCESAcQPQd6AmhUhu/0f5OT2URxUWy1DNcOE2KmkGnXTOnXzFwHS24MVP1USvvxRimShE
bhsMuUcOJs2QhkSv/nd9U2M6xfJyC9sYMOxVFnWv3x3faO0oD9CPG7xaDHGH4ZR9zqH/rClcF7PR
CZPvRtyugz5MFKKipJ/ex7NUYN5vB9bzHTVszhZ9qszmukF6odx+H2dlAz94i06W5uwyBQVQCSzC
1DIIyhWQONwmb0BlBH3xo9fhYctPor/R2QPrWbYtWEDhL3kTnCzl7crWmNPhnbdGaXjVSRkoxx+d
9+HPN6bk8TF/pCU+f+7Wte8L5SAsySuBTbfcs+zv1GVZpLQeZGa5m5Bl9vmQKBYE+f53muY9ZqIq
gDmJzzoXLITePqducoG8k3cP00oh5oLvJyp9YHlHwRT06cTaiBCocN4vUHPFgT/rf0dU6rH2RsbS
ajPPRNSYp/rc+Zg0g1g8oXebj/uQpqDg/2L3qCVNYtNn2Yz6VVXcr/Mb9rjmuxpV/ggtxZ/Bu20t
t1YofQuj/pT0/XBf0vb7KPaeXq3WWQPev3m0abm8lJFQrJNN/JfadUj3P9+BkvY/Z5yGUOUsRGrT
ajamc8TS09wgovum+qlVTZpNKmRsZBBuxLDYhZeVxoDLPJpjV573/GcmqUSveSNb6Fx1GtFUloot
k7xqIL8AxpLAspmxjWEWeeC3CaVDwR9EfccI+0g3IOyQnVbzBm5AgeLBz4zh1li9cV6MnEctqmM7
f092CrNqItvqazJhoF3ComGMmShfIoCrvKzl3NLmraMK7iddwYkweHtQzTnRw/t3LmsgziXQRXXT
2Z81V5o1I7rajmc3gTxcPFGPj00mec3NSWA69fYvohXB3/ppB6vCyjt0uR0bhrAP3RR/l/gVRiVQ
2Q9CFp2c0QmaSUIieZZCJ/QVrVZ69GNepNTEoplh1x8oR2wLgt+zYHP3NuYN/N6PZcVYqF9kXKN0
fwCLD8VS9WPJ+96wcutWLTCZYwjnbYtjFp+lqN6/zrdb5jAkR3Qv1MiPCCNTUt27R2IuL37GjpDN
kcpvAm/tml/jwSg+W+Xcy9/LP8tr8nqRpAX3oy9jHVCT5WUs0TnKekubEobcN9BAuatrlJA+fvae
JKj62ekYMmBu860V1WQRAXgJCfz7mJNAv8cth3kG3bLYHrf+fs3Dkf8tzfQu6P+hnG2eJtFmROGv
R2gdnJa8k22eVdP6ZiA5jj0XWkOM9fBUcFfrnUfTBkcVsbaM+SsoFydgVN4p5Z13CTA1oqS/bxjV
37gM0wYVsREMIjzuDYleabUfVrokcvkG0cc5PaaZ489LcHcXZuxc1vtv70R2IyIVzNa5hHO3CH7T
Do9qtiRP7QyEh7j6vIqnTkbr9C5fxI4+v08yGmn6pmAEbczwiQ2amh1HjTZ9GiXplJkgdww/PUIS
REPBMb6baHIfv7FLhdPsEokK1YeS3lZmgWxd51nnYqknw++sHtFZpm79GCBKYmqpIIsJV5l/p5OJ
ZaRjFGaQ6qryCAr+rB60hPd+/HzRxGTMBXBLlbcsLHeRNXQ/tT6Oa99zfDmJsEGTKYws1U3i05to
Vilo+oYDN5qfJFSsqSxDiR0DTwiCoEd3ZOBpLZbHkPKs8m1n88TAt32UAwqTG2ql6usMezpo5I3M
QSXfteoaQ3Giz52qPBYZTWe8LUBWGUxwUTsCdZkKaQRN5GzfBbAsQenYJ+xFdmHlAXvSIpSMLN5+
xlbVzTjXMh26zPN6zvQ6XnKIdvtNM0xteVLqY4Ev7Qt48Svmnjwernk0OnRQSF1UX6bu4QRYSbhB
FLeNvA5Y/5+dFVbl687kaxpC0JryR7qfRi8dAJhEM4DU2mQQctfFn6AKP2y9RAX+Wm5S5/Osco5S
tkJE1ZcXa+N/HhjOIHSyjya4V6PziEtSM2cMKoK+lywulcdsspZhjbwkLXItT4JNNvaLu8YU5xqX
P1wmOohpZb6k8UpW8IqHHZKE4JzTim8MHDrmItanTvEEYZDnIIPkb32jIun+Hib28qtc2LGlebGh
4oCLasICMyb4l11j93HORUTiFk6h084Gz0Nx+wCQVxqjsGSK1OV2sHCcTN68YKqMSQzZEmG3fvFI
CkIblNzhCCbSrh+0gVE/GesS33jvdhBlCF8wbV+oTyJxBOSZcovbDKOUZFyycJkbyHeKyj8bjM28
ree576mJ9D2cBaPVmP8V+iYuJo+pmeTH8dWDVIgue4JDGaNpt3aHmY1GldAIonFxNLRK8E2/5XYT
7M7y2XKa2k5MO81tqYK8aXc3pv8VjSqKR9H27BgjT36KUN3R87knvbSj8KsS8VdevZU3kbq7Zn9y
GX4isMIpxEbyh3xIeUSarGKoFpi20pAZUgZH/QKqBJqAJl6ZOLVzCCmodG1AKFJ0uaxrFbvcVZYO
fgwWw4HINdh942E2CSNOV468AExHbsXvPjpn2yRzOX31gDemNoBo08OfFOwRjc5geXAfW3/muAVP
GXyYTWAZqqzQPZyGlwmHxnZ45BgiOfsujWBXFqHxsV3PK7O20mRpbX/P6znZXt7ox6h45D+8HrpW
+vS9MVXQmfBS++9wYmbn9+ce9xFy5dp7sDoMR2BvMbdb6+bbOosJGTcsSWZPZmb7gphtZvIe1l9m
DolGlDuvOsq4ReTvnZZqM38nLgP80vHmh7VHuk1iOMB3fmVCWrDeHwXgrH9Es2Rt3B+VxPsLBCIZ
Xg+eSFMVP4YoEp9sOKmTLIvP6OSwJ4BgGXUVnJEphEEV/nKhFvcRH3Hm5lSwdcbbmpV+X2IeV4Ph
l3RgGI7TqYBDrMVZ4DHBI+nP4InNPy2x3+4Y5aBgzNvrMxIwHSAalC/0zMHnK76cMEldo6hQ76UE
R0iisXUJ5tQNaWKS5UyF+xDaMZydXykmL0ezj3zdHheYMJvMJud7j7aPQsxmslceJN7HW6VksUE9
rCcHtasTNwkYJjVI2VbFQJ8ZYVo2v4wH8vVpDTNuTLnRzDek6D97RwZPduOsw8TVRbopCUCJFI08
fGvtfGlbLlyqtN3wSRSw5MDQAhuoTBcYgOamKRgyBedYIqayS1v3BqD1632LZrGx3+FvSd2xmVrG
QPLi/Y7yTDBv9sxCXedQmPG4gFoDfyY+WfhN3UUrOa/jYiaCfHItqN2WLeKK07i7merR8Qo0XLqW
sPj/enjKYvrmy+1jPzM7dnN77ceUWtOEk8fIAqp9wAZK/MwqLtroQiy5zLu4XWV21SrdvUtu2yqS
BsNxa7x+4QAwFExVVzObCwotn+Ol5vDyGTD4e62EO4HBwgz1NGMxeREeuE8Hk/2VTgKvMhGSrQFc
WgBnLBcWL5SD18QfVTtycWGgX2gUxnas+eSZeBoIpkDLfKN2b1STlMWl85D8sS3vbS+1Z4s+YWyu
OQ8p7oCbce4f0JbwxYOGQNCR2d5Dgc56OwYP8UqkLprGZE3sgpseEO1DOxxN7KVm8CPCo4IeUROq
1bb2VUg9IsPJRxNrjMsdJVs0Ar9IAvz+EFsLKkmf/QVCGZ6PqRIim8AgXmarjMbdLqIZo//oZAZn
bC5RaGeZt/tXS1HlIJYUtsE+Re1LYG1OuWR+V8sZ1Y2b9+wYRUYSAIBO3MGLYy7ZzAn8yxYSvPQi
BYpiWV1HrSGl0z6VzyVLtKp6HHU9vZPsu4ZUbxNJRnRqQsEYeZKvKIqGcswM2WXO9tT4o1kLh12W
4V6PSeFSqdsgsIHm0gmX9eNlVBy75y5AlJD7TTSA1HSqI6LAW7U9gK5OgReTX9EsumK6FViYmJoq
bY57SuAy527//rL1vLfCHn7yIPOHBP3IpIcb87nkXD167s5+XNQrxjwSq2Rz93e852kZVEivq/vG
/c7lETdB6YQxFD84lfOJFt2YSRJs3Wkdp8q+kVhxQBa9uKPR+kpN1/C/LOgB3qgz22Pjfr5DCZhH
n0OB+l188c7zAdFgYqCtV8Z1dRTNHPRe75/Ffs6+AG0blaZlwTeiC81zX2vUmxdX1NdUpWNoypz0
EUkNjaT0uMzA6tud+G2y+K9YYm66criPtqG7Iv3P10MesCdRukRCgEnXQRE8LNIFMv5HK7pqLoKr
EWW+s7Vdzdnb+aaP4JkeHSJxK6WpY7LjXLOyyXzaaq+ona19pnMnIEMu12TkaoFH7WEAtMU4PQ+i
OYWY3zuM6bFwG08Cyi4vKLqSXcdNutl/j+Scxd4jsHWiFIqv3PrxmXGOkSC2PP740NbUc5DLEDHK
7z/ntyBUniCRSr8emkZTpS6GMbfZbmjAVcTJxlyDLdsNRlT1gm/ZQxd5tmJqAb00XkcBgw31NR25
xd3xsKXQ5ZCcnelYNh7b4qIDkuGqbfLB7eId2HAOiET6zBdYOokE/YHkwAKKMGiZo6XXX2I9BiU8
veLyRsQGER3Ed45wgBq7vEbntV8L4HXhvBbxV6QFX7k+2MzpzuJ7cbi0R8ZTYPn2d+5qABhvv7Cj
Nh74m/9Gqeu8jgSk/4Nsf/dkIXjyGIMpriMO/dgq51TLsN7J0dZ6QwBeiT9C/7KDwGVi/LOHgp+J
atE8ZCY5pSTKaoxQoCNLo6AMmYF3W/f6H+Hr6VUlRwVZGgFAlcjgM0MEqGBuyBkaT/y06Ym7ONSZ
aKevJhcsoS/wbPo7bqM3budupu4iBL/LGIMg5I9iVT8KCyBEQasbZeFF3Y//nppJWdMNe5J4dUPN
2Cw54HszHAgXpuT0GBMrI0m8Fy2TxhFdYc/4EtmHDLR33k1UGdwDU0DPni5ObKC/m+XsdZIBX7wV
nbVixkxqNUOgLHC+MT2Vnv4ED/zpHXZAOvkZbxCS11/mcdalcCwV/nIwql5HfFnR9zACPPJI83wM
jyhPlMyGRaOM+uRYTJz+A8Gss1/xNqxtec1nUUhpqzcoVZpAJ1AG958bBpqYlX0lyEQEZLyUN4os
/LEFm5wsEiIOcniE0DLxsFyfv6rm4vpoLsa1RDU7Jegotg8L5F4s0lwMh8g9TGV96JFK2tMfelZQ
KGgK9BKXpgdO/iTfQEROcuYb1DawSaPHk3z2c3isI1sVVxVY96BnotObI3+qE0Cv4X02uilatTNY
oNSTTLwXgVKVZ4i8296vbNiepmVT0mP3J+c5w0JLHN5GZfvK0Nl3xg07gBJ29ErnMeMDKAuOVeLM
w85zkfaGxr/iRT//X3VH93fY7Qmv1/NKwdg+lB1nNMN2jQBSbhsC2+TSrGanPR/jSjvjrZxPigeA
H++OPNmFDGLxQ1NdQwUWzkFtRr7HT0JjW/lKMDUl56GKnZQue94EaRp5RXw+W+Xq9+36rLs6AS16
a/U0fUeQ6SIUYj8GkWd51yfqogx8N9VKFCnQ5MgNgrc2ZvV7A0o/OdDr8t6WiPsy6T3zv5t/LM+j
8/HPOqBcdfIEjPqDsHQnzP8P5SSxucLwYc2eTx6/9peVUBpsdGGwLZqhze2neG+dzxW6wUIC5kWv
3E3k19/ntf1rEDbiOSVTS1lPQDY9HnvdtNM9z1U6Hnp1zEhQJ9z3xIyUPYCulnswbs7wHd2Nxint
dcXo7VZFEWyp0aRQMvrzdui4tTSVQbUD5SA1H7xXNp4mPrRalLQHWdBpeCFSvnOp4k2VUDcM8MNr
DpIYQVp+G9/FY1S5mU7/nWRJaqfGDdpGrNlAWLpf89ouJfuZtWP2RjJE5fS8OTloM9vDpSJyYk8B
pEjUF2pD7rDihDmeBdS7o08CTAgma44FMQ3bX70tnPe5WHeTGPNqkdlvgdYdkNem45qMsRcnpZ8D
wSovZCk/RhO71mYSN+vmdFgl03hRmp4sORaUx537aoYevOIKdov1h0tciQh5qnqIZtHiZqjf6mEg
jy6kFN6IwWVM/S6LuST3Z93KxBaGrgGGkD5fKhZ3ZSNlgKleYqqE1YPUbNmpN0LdluekQdUyBVJc
eIaDw6aLfmafT1wWLxfj28ExtKQ1H6VNUJHgeGkb5Y7sU6bOcy5PtaINKoPIntoL2jMdTDKQk/cd
SSNRN7MK/tK7F2MNWXZnAsksbA5FOeM6rXENmUH4vm/UcaRzn1YG+xf1QcKopJIZJHrGzNzgH2uu
V17p9nNKb6JBk4Mor+P+h5hVIUPndsTQAzUKwQ55AyK0rYtExN7IpJ2gOp0NPvJ0R9vb64nIJ+iZ
qAZsrCpZxGobU3RwInme5jbd1get6f5UG4YKjzk2grR9yPkvPsWwY4tOmMhKJuJaYtxAxe8JR1V0
98E61kMAyOS/xKfnWAdQqy/FzXB6UnFxUYvb1K57wVkuLMLr2j6qV8oK5moEB9KIKY32b6tde69e
nnPBKDf4Ve16mhS/RAgp21kPlJTZHoIugeC96+eZ0vR+8tEKTrRb306NU9yl8pdJutf+q3uLFRmc
Iqf75nFuuGS39n6q/gPaD5axjqEcceBBfcVgKCiX77+baYj2UOboKf+sQ1It8ISjPDOWS4VxS4OO
FuL4F1EXd1bVdTYJezdTGPCA7LlDXBXZkzug6TNK6U7SpYAWtVdpCR3iEZauFut3XpVM8PBLb3uU
SKyNDIYnDh8dVJ5qMFZyjZEq7dvBitwUWCulWaN9YxQKnrv3deVu1TGqfPypnp7o3T1lWD/Is2Jf
6mD4LSOk28OZ87MaQHY5oeyBhW7BcRio+jJGxfQ54OFfFrmHeMNAo99P3g+2OhYqZjcvej4fqWgl
Wol/wvhtd3VSwPj1Jh18Me9g6JsMwZmN22/hX4aTkXfHPJfqvQp0HNvEdIt5USv842DsAUwPxQTK
`pragma protect end_protected
