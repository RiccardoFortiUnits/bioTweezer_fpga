-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pLByJy+2ac0CxqBbRv0cPPRTQG7AhIENVKqObP17STqJ4vygZiu8NcH3JMNAxchYp2wxeCVmRrGu
mnOWdyJk2+LdrwQIO63hiPDgqt/qubGZRfo/HIIKVKqvtJX4lKoAPQS7QQ+xjoUi7o1F0lAiDekr
gWeS53eVY5I2S9oFGrlZHbEgLjhpiR6ZG7w7qVg6B6n+mG9G/bAs8laUKDvVubfaaMLbK4Drt2MA
XPJ2jTfPiF6vrV6ods191WyYi8AKQGFA25rrem0tFznPVvj4jMKxtGaXzggGBKncTxg5QxD+bJIe
42HrGY9CJokD1Yr/aTFebk/9Po1uYnxVgNesnQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9712)
`protect data_block
umYB16BS7sSCYdZXoazmHkDmlT+IhGakBQ6Zye4viN2rSYS6chj7wxRpwmvOPLYHLTFkt3bjDkHx
8yQ6G2C9Ttkhsjtl/JeLZMybguvL/X8F9HM64YPQXa2iX5fuSSr2YQBC+0tH5KwSw14ZswOy7vJN
SeNKig30lg11miYECXWwt/Wgbd0zME7ofx+TuYjHrofW6K4Szq94fMPetNHzhXfaQzXkw+a9tdG8
lySBX3UuEBZnBatH/ZPN3bb9bhJg3XGyScaBoUXK++3DJmwCQjtcPwLuHEsXsdcnnQhOovQApVrp
nAnYyEetKw8tApjShq31GdAoukx9GTagkQbE+0tBJPW7q5BobagdytKPbQ1PZaMR1zAGqoDtQyCH
zA6REF1+aiXBnmQcnofnmE2hTePozWHD85fWKLRNQPIJtSD58SNAYskcPQiVjhUACRFMxnc7A5MN
E7Z/9YJUutkC+n1SzXrArtxF0msc1lXcNEM6HKt7qmoXn+W0fZEE82RKcTf9p7hFnp7Zhbdwq3hc
zmRecSvz+jcjxg10jIjkJzmVSsTxPSURSgp/aybzDfrg0zx7P8hin5notMKiO/Z6B6oDT28Wq711
RUqFhFNJTn1dRJT2IgtHm8DUwOtrupVOSPKhEh+EYufaW/F0BAgFW5+vAIFzi7WOHFjOxsVT1tgf
lFQKiigogDRmb6eB+Y1C9drA+/TiBClaHIEW+8JkOLsGG6sfUxpbZpDCw6xZhRhPyJULmbNBYS1c
HKkzrQgXBl1WW2x90wcXnGJquGkwzG32+J+Hv4r1nrGo5ODJTs6LoHwMIKuboFiGy95ELoyioa9g
lNpTnW0XluTq2L4fvlZZ6HKDNO0sHFEk26UwZgy8YSrGKVs5sK2ZQMXgJBmZI8LcHfAOyho2V0SU
k+fo4MuCxQqOFWNV1qAhhX/WOPLAPAlMiGLL7pTlljWhyihcvYCqSsJmzbue5q6Ty/sPDD/y8rzi
klA3sWEWUS475KKiU/BJzqrWWKNGzr+6NQulZqJiJZBb7b0qwTt4Hl6R4qSIVh91/NBzBxfphqgm
oo61KmbETj1iJe3rWBNTsB95tbfT4Q+mnzMWsIMxIRTtsfgzV/C2C7bdovgmGndC+P+hm/uPckpq
YiTqrNopPKTNe6c5TVewrrENAW7+weOc2MBW2Ba5TY9DutbePitzv0VziPV2TzCGiLZxTHbMPN6q
ii8NHKOok4fj2QcHtKkzp4bodrrICfIxraukpw6fQ8uy8tZhqmA4OBQkeOjUuBuSAR3tGK4nNKAv
245o4++MUeh/WlrB93mszyHWkHb+6nCSL9FMf8uSwpeOHaJ52ak/v3N7fJKfdUB6+e9o6i4Rmz4j
g7STFCI2oiCzm/B5ukJtMkILuE+fjcPynhOVja2tFrswLBYiOVkjlDMjuThaOlAS6I0jlDsh7fme
m21lNdEFDg+AEjEhsigxWKCXCw1iEyxYWC6iurizn4HitTaaXa1gig6vntjyGmNmKwbqqYbad1iL
Q35hJM769CzYgs+tRtkepL1sNLkF6Q67yJiY7rsvcoPGNadnHY5r1dU4VIenxWlvg4Gc37DSywMz
8qcNUW9RRN3ctt68mWS7DHLQccBjO2rK0Hyhzjl/yfSMd2ePrD0pwXfrRmVRBQkuVBiHkjCmheJw
SXkWWOHyA6+YN3nABHVzXMpFajCxdbB+22rhClKDgzBU6yJbqxh4DfJrJG5kqPea0DvxelMj0SPT
J8r+OlKdXRPgLV964QaQByqxv2BbRVKeLivDtTy0KRfppqloPLqyMfOY6ag0Kjl/RfFjvMPuAuLe
izsG4WW+/kXj5Fq2KUWIYsbwn1ky5y+tkj0L3z/R86FQOFIzPzIWPoB0uoyW8oR2Dn8zJA0xWmY9
NIjLNOVUen3GB6f7ILfp8hShI7Ktu/0nFTSSz+8E4ioycT1y4FCOdm+VvUEOsKlXRgcVvz7CB5r7
Lfj7REObpHMAh+/B+37i6Jqoy/EyqNQVqifncyx+/XrbxsFlrnLGJVYh8HJvhFuKpzG5u/jF5IaH
uPRupVFG+/zk55MJjTKRIorEwLIipktDqnKWFRliY17D4M6zwuun9yELvI+894TXEcvX/zxD4HCa
FAR+4Np07qp1Jgehx+Tzk7xzqhUgNBch9CTfICCIlb6DyuQZOvD/BwWCWnXgUK39k6WyNElncx1m
m5Pny3Py2aR/kGNXSOEWmmQOueEWp40n2QwUiaJaNDpD/uChlH5nYPfpd4/qopc6zBTXXijwGEdZ
GKD5gMk7Nnl1SR9iRqpcQmAgh8kfO7oRq/PwGEDYc/K6ixsdByAmMor7iMiXmMTjofk+NRPUiRqf
SmL2XpGr34gD3LNX5T0Cic1oDiPInymtoldT/o/b6uTcV+ogpYb2g/fxfMPQvgP3rJ7AEDGtBPds
tck1afWRnhJ6GKQcNGmL5mbw+zgY/DtoCP83bT/v8eb/LWMEVjqjVcz/XRrdx6FsLdcBJXcakOmZ
kjLt96LvumgHqL75Q6CAgyPj939go/u21rRJ77lrYrOtkhV7w54fFJraZGpDWXUXulxps8qBwBoN
lwBfwSViKwVjCkckUpqXoitXT5LUj+2wlxXSWb6ksX6/fwZm3j/zkqV1kDrSXjyhVhNF6/3QrQju
qqgoY/HlTOd0WCyrFEf5LtdYkIXg/wQMSBsr8EcZiOuHmwd5dSfZd8lxf9niiEo3mx610JdkKqj4
fnIbMX88cwOOCpd+QWFWRkmhF+h5tGi0P64Lup+9ka3hwp18/rUwjKL9LtfGk99WGjSaAprT+xaX
xccfz+1mCy4YyjmIC7MxWD0ysZJgf+u0EYaQEBGYG2xFzx2Dg++BTFkN15teGve5u0K7kaxVGVBl
Bp2fxL9Qgw7z+9mS5GkB6mgRq6mZk0JQERibRDpTHeVlIspIUckiulWztr2EaMAnK5wVuxNKoov+
YyvJk+KyK4Jy/IW2+fvITAteNmlUVnV93PIO43c/jU/N/GE6rZpN5tfU1Ae1xRCa1BADRVN/pzpg
pvBJ5IAc9DFj8D7CBw7/Q0zTZPXdIJN9OWtO/KYl+b5QNyYRGl7xWMjV9l8ys6O0fkXd5Or6ptTG
2hjjmYLIimD28vqLxc5jQQpWEXjIIWN2YDl5qs7nR7mTS22IqtvH/1ZBccX9b8kMG450kuj49wKv
UK+mW2gDtHcJMEV6xNhVbQQ8f6KioQH8dLysM6pi3zzGnPUQgCcyvoctBe92afQTpIODv+5SC8l/
VIeEbC5Zv9RrikTyqItMt4U8yI1laMhc6LRnEHBdYBYz/C2UMwC7UwoqENh9vu2K05SnGpnfRxfK
H32Rwdo6/HWM3oxWpBUtpm/s7+5PjARklVyKr0VINPdwbIqQjRSm6rwV7Q3n/9V9SjrQuTEokGay
5MgeNVUjhZMj1aohb7daeoqg9gi+j0czcteZdfiBk1L5K5XScMke/iodeeySJQsmD1c9m9/KxUH7
zKbHQvTcYAkLA39f5N7aPI5cz0ut3PdijblxHOFMAp+wuDx73EiZVgQX6H1Njl8poOIjXxgh09Aj
8b+++7iVfHotoe5inwiu934yOFoQqUZrVtFhN2H1ZNje8aTGB+/xwqHEPA1oJYik3YMygfBRiTQU
6jrTTbv57FocQQR5E7LSBoux/3Mi7qpsAUN+r5GMfysIkdqUAIemLANO4XUOuVxWt8hoPCCxZ5H0
8OoeTINj33BneeZ82Ne+M3GvLkrJGT16TFMBRenbsFoubJU5ERXlSZMWYhmdzVQhThvJ9LVdqm3p
dn2elHDPuREPgjrvuKfMzVe0RQqI/ZqMwwoLcdob2G76dnrBL5qSIY2H2GKjcxE4wCuOvswJqaza
jQKXnPCR6iodSAMUz9yEVOXUn7Bl3L/MUicI8zUldM6JrTgYzhr7CXGQV7rP+ZLH9EIEFwPyCyvm
Euec1+G+cXroU5X8gewyfaVnpOttb/WaIYKB3P/KRmljgYiE8XYtVFWbk6ckS1sYFp8hMjhebuux
yjpux0TGz3+RjoHuuErs+fsGrnMgajQyTP7aFvvkVm+3D/Jrr5Warcs8nSTQyi/25h5P4MO+TF0O
MhO7+HLvgGNmNib4MxCbz3stOpIY8oPeEmLNlrwID53aWv2f2UUuZ4rgZZv1Zb0C15VI1W96rOnZ
zwoEvZqkc5IH7YdNSxUrIQ03o35+H9dd/HZ2fR+feDfHLOujvIWYwgubYmKMyvaYfvz/mvCtbCma
Ok4sGTX6ez+49tHTlOqEAG5oc+Et/bvobxusmZXP+Wn0YnIpJv5q58MxnvOvw2Chgg8Hn0tcgt9S
1WGauV3A/sh+l3c2/BhL1EZSIIucmo+g7hpUxeU28yr251Rj+c8xXeM1+EQV9hkOIkhSbGd0rUT7
HeJ47o8VnON+WDBYpoTMJqTDdZ7v+5T+VSnz5rGEvioUJvPVryJvePFnFohu4Wh1vW/GAygpRxO1
Js1AfncStQSljSmqzd3gHnuihjxET4DjqCss+cOr8JTxhDejuz8p8yPBUjHxxbI5VFjxnzAFb4ev
6J7UoIwdjtbZwcm3FPup8TmFjWT2Nmi0rphb+t75WYpr7QgCJyumBCcB7SFgrfm1SuUEvbvxczP1
JNS6khbCfJ3UCYBIQ5jsry0ajC36gzkbKOLhpAjF5xvTi9DA7k8A2nQvvHTN990k+/cFsa327XD+
tKXRyqvCugOnBzNBBJwgk8VbZ4kpQwV4CrKeBak9pWwXnXSEbexssEsVsfRCJSBlsITQ8/OMuqPM
J5k6HTxADvJI6QuNvu/CtEz6wWVbi/D+eS8+m4rpHgVb0zZE5GFkpxkOlofm3+66pCM2cK5YTUGG
coRxeDThALI4IkRGIRSxHsBCPBIgnLwYGhae/VXDNkAql0MAj+Id7xu5d4rfNEv8rvOo02XD4zmQ
UCE1djOrWYlmKAEumhf/2GrIr9lfsAYkZmqM+Mfp2SkbK8F9X8yCV9UtUYOJNZ+6CrsMGwLu8RSh
bb561W/MKKDZCQLu65N4aWyyNG1BJfH8EOA7D+4m5qVQbV3MY7kVoUwtYWlooInONZfNilTFjJlz
ocY9Uv2DjNJW2mzm2FzPX9PTpd9ShApfavf83paydH1R1PH23sy4iEm0JiWbdV/ZihGQgpAC07Lm
QrD5bGF+QrHs19CY2yZD8SfTZFCWfvodUeDKrQWxjgg9ygxs8yjnzwjhOlKXIfo7HFjSc9xx7BYS
sopDfVQXMmN8PKsyDk7vvuKbYGxNwhEQJCX/BcAY26wxwFnEPRSGkj5e1i1WPss2yua/62mXyuxK
sGtl9I8MMYWOpMOMsG5ob29+o1fQLvyJQxQjYdGT/mM5UKis1pqDIGKaoCL0ZaCyyuNQls2TkJW/
q1YB4mJ8qe/alYTAivsGdVuLd0lRg9thPS0S1MqOTaO74H8SPcf/t5PJnKWGXMvEKSVPNRLwhghi
0yR8e2Di9Jr+01nTpPTBNlYEEQ8Dkpdi5WOLiuCkqJxly0nnY2IAnthHRTnD/QJ9wXfMtszPMCX/
jMnKNAffkl5jyKXaCZdW7XBp/gLrzzgRysqBS50zMqtS49Ds2sq6Isq0BT0jl9FWRpzYO2Any2l4
YgVOnWfdcYwmEbyvxbjZu8BwLS+CVrdxHpRhl/GMxrMYpE5k0KN0fSmZdV1TIczCxYWlmph9v9vs
QqUnWRbJ12VEVOAtpQY4uotQk0eD7OIozddkECLQn8VPaH87lzMCbEjodtbKRVLpNG8c4RK+G+Tl
UP5xwG4TuPt4Z2ZZrB3/fTRPhvrOjMji0bRwSgc2jJMdSYBUJrAbPlluOGQehdxI0MeV6TqVDbsQ
ZozX57EGQFiUhc3YPmxgVRU5QEfJOT3l23Gb9oONJ7kQm5GwSaEzSK879jxDnBUunp42q807FkoO
2j0zqeFjb5IWzUhjScdObDkfKcRvypm+36IMYbEgVCDGvCH2V+mfkeqfoBiVgosI1htUlG0iN+Jj
E+i5DNZ7Vx+1IdPNUeW96iY3I+BINwBq4AzxOyS+mrOI4Z9VrC/CllnOX3FBAjKD44JqPH/K4r3r
lf4EGi+lxgqCmSSPfoohGPg8VEpaK1pqqSqNzdyaga/eX0uq6RJUJjIk/L67aKVj0tl1Lxfc5ukq
J5bUEPEJ5wnjfUJe9ndiSrD1MdpyNhQwQqsnBKGam15C3th42X9CXlgsWZPj8ElKst0CnjOPlkE0
c2gNSu3tUKyCRoXxKnYushbcwNuodHS60MMxSqD3kUzHV5t/IvyfM4qRDhwo01jyd+eABMw8mvj9
oL6yn2HKeNtrc8QckNSfBG1O0fS1dwd6D7mWHbRlRz9fYmaG7VTRis+W7ZKNcMAB+u8ymmFEAK7/
Cd0S/J9hiij+F7x9L6FITnf8W+/7Ay9T9ysKxD03W15gLNy9w9Y5nbUROcc7cArz9Zl6FQ/BcqXe
ONkhbLf/7ZhmjoYSW3EXF5B+kJzPBxEuod88PDYbsnWzttQqgMhopepSjZt++qAyJYHIAH5GYR0M
UuIikQGUtAaCqTECjswGqBKo7eJiQTPdg5gHqaflX1joqz4mH5IWIg+t/3FIbk7uVrph6pooph4z
xGW1laJWHARCGZum+Qn4niiyzz+91W7H1gksIZemADalql1bmPtQ1dpTkJYCDXq1osMz+ufzU0dV
i8L6/s418QOOD2tHOrHv8uEfw4/kBthte+iSoPJVz+U65R7ZsfYhqJmYTG+HmTugnw0IWJHh6oTG
OrGhl2ugO8FNvxMTfNiYhjQYGsO1OfRihv4IP7AWYuMuGBdDCgy7ozHAN9jDVAVK8HL/SuZXGsKe
KpwTXP8vlPC1QYqYBdHAYCz6H+0UOU9R6PwT+nT5uioSPV70GCBeSthIGpupZcsLP7oAjUFENH4P
SSpoKWum8uJm7Fz2s/wxg0o7+lCnq5TMqZwrSM6AiIO/02vucENCuGzdQax46RCHQkCI6M23l0+b
x6sBYB5OE3C40X9naAq0axyNgdyvwcDBLygU/3DDLsA8rT0WgfEJ89gIEA2OCaS/vs/yqN7whtRh
pzUMRumIFv9bZwkkXXw8AlGUjegBEOOzc1QI2UuD/F6gtwxpS9o0TdyWrpAlpzcvOFfXRbEhJA72
QpM9w8NWVww+qfbbacf7RLHfr+zJeVnWYYj3HzEPfuzCiC5ddCSEi11EVJTFbacp/EgcC0SUHm+g
8QlcDos315EQEdtdABM87Xie0+yK/3Mv8L/zZh+fNCMPsgHv68IyqgQoSnjrLOFYJmh8KsvXnKVY
BKICPrIbft4avBjiNaz0eMgQwXQPZcJdCyrt4g4W3fHhmHTZs0QBZS+zhFcGn/ce9JQYoKWwm5J6
t1ULj4PwaELbjdsLbI2NiJshtrObwcVN2MthzWzS56OwiBzbf78qy1Ey4civnpS00f0LfZADCY8l
WP/78ZYMEFHM+WRQnztJ18CGZ7AM/tk46HiXtp1lEWRu8n0PnZvM6e961E1SXbB19tn1z9XwtAQR
PcadwpD4GjCdcNfqDJe9JBiz3aRuOYQk+SUb3AQx0ezst4zJDzMwNuwziH28QvYn+0ozZOzeQwHu
5y5G29dmPo5KgGR8Z0Y6eR3gKT6T1RN9WolbrDEwNaqjORwCa+5EMTGpdMOLBLYMHvlX+TYdgSMp
3qr5F/Tk8O3POsvgYGRM8WMsPJO+sgiuGDOeaevLHdk9z6hp/hzDjCiJwpAwjeFcW0SWJaeZ4O6f
+vm5UsdVtHsBe0E1EVxV6DRukc/Y53TMCtT/EgjkVN0I8hoW/RGFrhpS9t2bpvUxMdLQqaY3Ce9B
67ZNdKRE49KhSde79oI+VPbNTxNNNuNisl7n/yjwm5QUBwTpZqy6p3LAjC3j74cZmXkDfLd+H+dq
MBB0i9ClH+I/LokIofS1n5Zd4AXwuXDsvZWz0/FTeZwH4+RykjexBGrzakA5sUJYiDEnOIXGhqeP
cIdZvap3sDFlxRkyWOYg+VCHG2Zjhg3hBJNvurHR3pAMbp4qjWxetH4/w+Mqm7ayq1aMjZR0vTBF
cWo2ztEz9nvr9aHZmb4pgHRzvhcc1eV5C9T+TzP5oKO0gMx328405K+kywz1euvfR+Uq3YD/WIrS
ffJ4F8tP+YUiaxaUixoRm7XH6hC+66t2uTeAxHYj31EU2N5iQECNQ1qW/i80E9GFNOOKOCMbvN+M
vnLz689EYcqm1uAnRLjR9M9P6+W0+1Y/diWEOhVQOGHanPrDQMsEY6TdJJFx9Os4DSaF+XL1BG2S
JVsc3Hd0zST1Hz+7cMdRRZJ7ORGfjiqIb3A+Aaj31t/qOzGal6Vw+oxUxmC9GDJ9G8Oxp/20oi2G
gqRdXlSP+kPuBd3ckURW20Q1kWxNmjKv6g5/O7tWfpAbAHKKcYo5Nq/3oHewlI44I99ch8ZKTSPW
Xn+tkFpD1jr5HW/3FS1G75CFGW13wIqLD/cdRBvHTVyOT10z5H9NC0jlqDk+NWagvL2ihkXfRDrB
pyE57bBQdDmcJ3IqDSflTsN3uP/3lHUIQ9dN1YKojjMG8hkbRySn2ivdnaSzgRCOaNkS3ilJ14r7
GdyzW9b96hctg8BpkjQET3HpAVjCsgPvOI2MV3pvQYi3wO4WNZR0dt/4WRL0vK87yAEH1Zw/9FgI
jRVVfmMMRvdB7zauYaW+hMxOboOSWQUWqMJnvZytBKutqEUZrShgCd1PeYF+0cOo9RjKSa+Kv+Zx
CKyY8p503Cqqpyh++yYITkjCHQ/QnB/TxtmHT00684Tk6JWDXzLKg5bDgm7N2Wrp5WMpFr8revDM
0ZKmjowDeUB++QX268lzLfGYHrhwtoG3vje7xnrjdNUSSymZ401XOjruBmMtZXuYCd/bpZzAU7Kp
cT/MmGXFaipynnkLbmrsbcXfsNPnXD81x9RNPnLcFqtSaZWGXYkEaVSrdRapfL02FINn7Huc4rED
b4XGazXgnk54UzAv7/QeHfqAdx2FLs9Jbc0WPUoWEy7r1XcNVLSDXQ6H0s+PwJseVqlRbDK395YD
btMGarP4pcXA6hYesikT1YnceRLVhctr2N0wYxCZgUkYrqDcwqrNUrmJhKdOXiy2T27O4UVbepPS
lA0p1TMcdew+F44v8RjPe2U96eYBRpBZLpE60CK2O7exRetfEgnzbh6ZGglv61KcwRDBtHu99l5o
AhPhgqZGmehMvah7iPqVq7kkSBoS2bHcDGU3+4JiE8SfVAH3c2J3mFGJDIsVQGH+0FG5URDzi1D0
AcIxARbMLlnShSPbkfRqW7DRHI2PfptckcCXIrSY/DXIywev5oQdUnS2leyPwvnTsbesaOeKCexe
jDFTqRxSb7bBKavA4JAoMHVQABCnNxLIaE3afoK3UkjTd9VtqBXRqyNB+P0ayQr41FtvP7fVYYPn
LfW9ycmAbQw8GkrojJWvNXVefvV4EVxhGU1GdSs/cUBAacv1eo+D0f4XrNMy0X8pp4v8RXcMSi1G
W36iizTCch2NYgt7TWeVbag1Q18ZJB4KU0T3W42UsD2D0ieiqhrZmIm8xEoD0Unl+Exxa6/9QH2B
12tQBpEWdDI4bsHJQ5BxmgpsEIMeU+aRL4Zo3ADjaYeLDm7hV4ta1pREPoZCNf/IlJgZzBDIcV5q
qqvh2G0mgp7SJtUM0w5rlP24J5r6VYh+cWqVq4Z5sZtqd+M4eZd+AmHWYjj1pvmAzEauB3njAXGN
qGsxuMMpJ5ztvtMICXipo6jf59aw+MjadMYgSWC0EMmq7foW4LbczdscxYQZ1jJJPkbqC7vdAj+R
grXdb7pmBhpLjyHm7Vz/InT7WyLSTNU+L042FkYQDQXrV1x+BWTjsQ65RSH3vgGyfMlTS1Jq3BGd
x6mxzJyk700GFKpgfmVVuSYmfsbnZUaVJ10NKIi5DOqEfaJGTvnG5dZ5ShGWPwo8iAozoo2tglnD
UhaD3l2nW/HV4QtWnIIGuOL7d/1btrvVfp6fuL9hbVQq5m5BBDU1fHXRDcR4UCsu8fggtMiJTwMW
CG0RnrrUzL7Bnb6G2IsftE7c8tHTSLt2cMLnozTBc8yD+7yKb4MV18nnt5qymNxrNCNscBVgohDd
0AXzBi/+uHeJKByMrcCiuVUhxCReXipd0rmv34gQqBTH7kRknHzOxtJAW2kZSOOrgf6bsA5DMX1k
bxriVOlzEu+LATK8htY0OEhZhHqbCQdkivvXiPUYWxnnRLYtiRAQTHhqsbktPlvvvaoX5ix9VHnB
E7OhuhP0Ro+3821mg431ymIv7woHC7hFFJG0USd3GXGl41go1henUSPXR0faxOIqQD8jSArk1Ukk
DGrAJP+t+4a3bwvtCJXNCHx8ZtEptWvQ8l1JHngUellI12Bfw8BjY12yQ02WwwLGR7KMdXhD7yPT
HFUvk2Q7FLhiLOM4VBCxIjN4HibPCf0Oh/oB+tNG+DSG0acWo4icMD/7xKq8XZU5n6F9IJLwsSZb
tZfMDNHE3FTmEFpaNrKOTfw2vdQ6D9S8cqhi6J/h1Z6UdPGLTK6vOJQBgDWHqBSob4z9g4QGww4Z
IBM99hguEXb11bcYyux8AkPY9EDrro1mGgh6dtP02zMmUstXj3BjtcQrYkOJENK6qsfTEHFUCVq4
TvpTMkWfhFHyiKJ8HBKemcuf0yoQMInpSWdOrzpuUeHbt///lSmKk0eNXU83kkk3WlWnAC92larz
uI6KL0bYvJh7vw+7tA59Eo5qI8R+Lt+m2y4byO/7mYTHFKknLKHR7cf6t5ml4kfg6W8VK32EMFB6
LipkXZ3sXW5Vlv955tcpBL/ZrFOpydEj9MancGxUZvCn63FObvXU549Vnb5k/Ae4Q2GavM3i0iHt
tp49F01038IzBmZGdNVKxJwFDprYaTRIKTjSSxK3KsZGvYc/QbkWElDu9HrIF1KFqW5uHWGz9/p/
pOf1EiGcoKxfxsAjEPuvZtNFDuOeMyZ5q916TqQrPzGxTKZx/aA1Wa5hQzfqYRuznt7qkpUXORbU
RpgwwiJWqWcw5ByEioYTHx9glKM0Q5m43tp1koh7ueryQzI1tiXeJPEsZlJhzf3cMz1qR1iFfpu7
OQtCcrl+RM/JcDZ/OCHujHy9cX1ADel/wh9SoBOollEnfdqKB2lqz8yvY3bT6PX4iezRdAFdxCSH
vGAygNG39iAg9+5QvZ0AuBjuhKkaSdoOfHahcxu23tCFTms9l8npV+hYsEc4a5XmkGlL1KbfgpdB
pEHnjvugXw41QL6ILeIp0dz6sIH3+fX5nL7fBFHulRWQ/7QStHoCLeCkpp46jcxKiB13HrGQHysP
cNmtsrP4531BrDdLPJEInhfGLWSAS0/rX6oFQFnCGws+mpl/rc6Osahqw4Ob0TL+Gmgs1ukn/eo7
dur2ZK15FyKRadLUplwjF4iE8Z3rJIMd2HHYUVVrY3QnnMNm5o7GYwxz54J4YYzNBMSPLAPZFt0E
1RB4CLCtb85VwiR21loi3j+6DcO9cN/KJ3lwviJzASL8bN9UviV2EMsjgWZ56Dls9A9GT+wzzs+c
YLtuQGx6MynCWAYKhmknjXIARlJBMnUsvRduvwTNk1JAvyhPheIkMzXR1NvsS2SOunqi/paCiTFH
6yu0qFrHdNyjEreoclWGMH4Zm7yOowPxM8xvnzyYTSO2xwYphyJWOqC6DVctfVI8d9emCwqlKwVa
n3bRdbsD7gVIsBnJp53DR59U2Xa+cX95uC2dioo+stDgphkMg5Uj/ec6hIvkD6iYCaEEpvG31UO+
558sPz8p99/SPJFhYRMqCx7bZAqIaOEynDnOl8EomYDuo4i381fVoIubM5KQujMz+KGzrtl0SrBM
ER2MQpgvwKNm4mfQ48Zz7ERG9vfezHxb037LCtDa0LHJdA0gTesZYbr8oIQC3+AbRW1baVvDb1+c
5xQQitYALdTHGfUXh39YwOIgtr46eyGhb2UkuM03i12t6OjjLSSLg9cCQC7qBEkhJRQIT0KTnE7u
poQgBlRs54NJgRjLnScByLtDPftiCaKKbMgfG+NDeIvLPjjZUcuWHrSrYZ++bdpPFj5KWxluhufG
r6lHsqLd17NsRHxNkofIwh/LrBYaRFixOvNVHbFppOebwtzoq578g4tE8kGgzdpdg99fP8vHFf5g
v6SUqlQ55TPjsZzAwD2xJ+DFRtbHe0U0qMnN+cCgi8R/1zsviQt+b2Nphud/UKwhE5Qq7XiJj914
I7cCIqQUBc8R9/DcMe1OcUIROpE+m30GFYUES8jHVOxj7/TtZ5X9sBAvnHtMM4nAp1RusgZv5/tN
L4XfGQ8qP04A131O9ZwhkCfxyXBZEQt8H1A6X4mIfdhcf81k7cDkHA8TT5Pk25qcb7oC0gE4xFZd
2SpNxn6vUgzEmnkZkaa9a8SB0iZKo4oT4LqOr4dBg6E78juumkmugKFTbFzEyAudvQ5s+CGSTJUg
4MChF4tTAmrH02LgoQ2VUdrZIPw+xQ/E1ZdJJzQ4cOhAZtY8/D6FCg2Ta5xbMCtcaYDYFVyxzAn5
87GmL1AjaIfpEB8oe7RFhfRFIuyk/V5I/KNkxukLvS1N37D7SsPwYXkOkrVEEeFUf+YRPWrNtMIB
TLrGx6r0DU12nziQyloxH9byH2jUx76xKy0/Bx86Njivif6+C10LdkTtfLKu+0H3NH0IuMLFDvan
9fKGTFwKIgT6SOsIJxzMdQrmR0yivLss4xvTc7CS9UUUP1DyWoFKDxfWpm6YcXWJ+yCixCj0ogup
r/3RHOULXFGzyb9vUhSwdB6IpXnP7FDp/p3L1kN7Cz8rC+2UAmeAAbqvfpGA3AgAS6kgGGyzpqdE
hwRaSL7Mi49uOgLRNigIOVuJ1Cin9Z98b9Li1wdIZIKgewsFIEQ8yLmKaLq8822cGc/2bU3kpovK
ZaRsNjBciiOVgtbqvLwkCbbMWpRujQ==
`protect end_protected
