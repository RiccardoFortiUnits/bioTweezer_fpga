`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tKU8nfnd9mrFbxCAa8Od3i4qqOUEF5xLeHBJXa4Q++rPuen0BhpwzCftLq8il2GY
iYFR/wgeKFZkOj8Sz77NsnpNZLZ45+yWReqmoYmd2g3qnncH21jDIwiRD/zlfPAU
xpQoCo0256fXjFr5OBycBAcb/bncDnjwQfg1PgPr4uk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4192)
qEJLZPQJvlAwoM7XG+x8f/23unF+JKGWUImUUGbgLwb1MOJlTPlB9lfajqvFiT6K
ucuinjLpFZWmjcCXQvjctgq18CpK47BoyAIGf3VXrWbrRid/hfCJwSa/oGHqrQ+q
yQZB3NWso7bOqKN5owOftdEno8m95tXxLoXbE4KIUw+JWgCEez5SqnEXKQP789uT
dqP1/XfvrJcQaFlkWh2DXGJUlxe6jQF/YDPnXzU6qjmOnwzv2FKdcrZSlO5Gk8fD
wa9KYnu0VKT1rk23vpImO4wrUDsBTfNCW6J+3xFbsf85sPFoOnBonM47goqL8fYX
pKglfxzwi324yv2uju6KxDo4p30OtsmFcX69YVohFYRIWRY/gfjqQO/kNRy9qgTg
qfvoLZPZ15fDliEVMDp5VpguNvu/+AZY1ZHVTajluzYxLtEjBpwm2WotURxjiYzB
fvgM9ET+RJK0mNZedkYQnLWEPfa+UCdpVAvklSR+W/wW8uTwSBeGyhTUHPxd4Z3J
Mq3BmDZ0CHtBkC5wv7xBksTcDwZlfI73RTeo3MJhqX2xLEXmEHQ2puhTi87mqY8F
uLKMutKZoTdZO1dOHwdGa6iayDTKAiUWFrVAqY5FCUUPxLKfcxnSZhNcasc1AnVK
UXXJWQ7RqtAjCEIayp6RsepTGHFVk245av9/C8bfybZUANX8uL4NPfwPL6f90BBD
Gb+wcMB5MADwLDSkm3nEyhpS/gIhaC549i6DD25YuQPwzgRQist6KmNPwemZhQsi
uzDGvwE3Uv/XWvlZ0F67gQpW6taos3ovetPD5+L6ux/pWtllF6kQBJfKJitnQxrI
PQc7wXca+2J00tY5JZ2Y5ewuypHtS6DyyLshobED2BpAQRMp+8lIKWtrNhU667LF
/OkQHxlMmH+W2RP44lz75602dhJlcNo4JO/ajBNfG6MAfOif+IIBFWA5my+q+Dud
72PysTCQ8iBvl8ATLJOOYJ0x4YA9R3I1MyMTPeGV+aeXriw31UB3AA0r0MyVq/27
yjEuyzsEpvE76EcpuJ7zY9P/yQDkRqutdhpP6wmqgNJrOJhtadRuao/yE/2Cq7xg
FBbdj+k0go1uKhN1/jDujy9hKILLIU6hL0U7Z/tcL4XKo4hX45MrXTagd98n8BZt
Z5xcr+c6QTtdHIFPq1ufZG1AsRi+ttSldf5fMU3P/VEMaaEEfB3R0HwTOvhyyCks
dat32CjaAi8E3l31q4qiBrUVe4z+1sccGHMpEENcKiu7UiWUUxvh7RamjsCgsA8t
f4MULmgIlmJ4EFig/DrvEQI8oI0fkmTwGM2ABHsJhmjyMBdxvX1BmuLfarNGjAO0
DG57YE/YGIvWnhqRMVTdBzbj9igwbe1PhPwnxtjelAOStiQvGsV5yODyQqoMIrvX
F8EBMpWmHSi4ZlfzqcCOZUp2cZx7UVzrXGfBDEjLNNwUuQ+At98yEDM6AXiu/bcP
84ddTHlTQDP74BMR9N+2FnzKFV0LYk1S3vSr/aAxX4cH9+PI6mzVLjFCx4ctlIdh
i3VwkCDWTSCndQRUaz4ZjiFgYrJ/p2s3IV+PValcq46U7YHFfFGDSmE62oX/Wxo/
w2FfbQIGd2XYLRc6DDd2lojuk9rTrJ6nABEFEmJU/uXGBY+uLfbYURaF5QfayEeM
1+JvbVXuDXvdwsfrl0RYqY9wcR/3PxOH29bzynEzgkFCeo1rh1XTxkgg/ocBRVF5
cwKf13hANkWwK4QzF1DKk+ZOi6qCq5ci2OCf/WEaTAxTDK/gHUi5IRXUjEo/jDa+
inWI8toy64j1ikWD+N2mvoAYQUEwaHaoi+QY0q77ZUZKT0fV0IBNyLi86sjYsmtd
ikJ0qyTuVjaGxuPcwE2X3yWil4W2WfqBJDtST4ENiVDVzUW+xkqsXHkKw04gSI6B
45D0Qml0AKvDtzSGs+lz2fMN33fACWWuxHOdi+HxVjLbVwhg+GZVimjC7UPC5J2/
Z5ll+du4b5yKMrBIBnwJ2So7Lkvl6Zw5lBOfAP/hUjcl4jHccVCJv8v/U+LQnQ2a
Y0mj6BcPV4CP8BM/JdifMgRgrnIuf/pjT+GS+wYoCSg/VRx8KMRJOhz5FAjYQen4
NqWM4a2WFbvkC0TXVkJbwqroWtV96wJR7X2EJ86nXV38cnr7Sb1Oz8plt0DWE0aj
UG44hcykWCY7fdPB9ZSUXRenEn3Abke8flez/3m2Cfp3pP4/w+lrWuUaM/46ouTd
vHD/B/O2v7KbJ5NpWYpCcbpWr+SZIH64RVbIqrxanRoghPqjvGDCNMBf7qb/1x0b
S1pBejMlowqJxyMMEALnwomwnLUBL36PEOu3saZmdH7+wwl4xpjPb1ixMaTiqn2z
3B60wJpsCOk1MQR+7Pu6jTKvqXDj0zBW5cidtFauSLpfPKLqiJKJ5MdEP6beoZI6
xsm8YsLM2Upn+fTLeWH2j25iZcYTIzG6ibKlIRU2eCCYwCl+WDIlYB+cefXKptxG
F6lxp+JxuxYnOTmhDkGFq5GaNEGycojYStFwacrTiB1wqXuhjBYbvIBOqPXQo3m+
FahaB8xj3wwSnYUNnnnEe7yLQnuxq64+skyP0fvqt0MTjWa22IoSkGfBwuYo5Dt8
axzD6OLqTGX27ddT0lXrea7usKvnwihHWhVXgyN5JZefXT/eQ9LRC+WZERXf04Nm
3Vvptxmmnkl2ZoJ6oEufwzyC3zfPZRLH1MpiSPieTmdm4LUjJPiNX/6QxqSWMSCR
a6Cy/2AOV9AcXOePFjW45r8PTJXgEqIx0wZ8Ylt5n+DUU9UfdARSIe2E4OgAa0GI
W0Ai6gffhfG7QuubNsFRE29Swcy04XDU+aCaSD35UnPIWC4+QEXCf7ZrVfFgYQvD
8rWXAaf9KFr2tEP73+JXB0nSIPhfdvECcztk4eRF9dZjK2/dhVNswoVP1tS5YOYB
8n2NsZNG+vpjPwAHPgwJP9PoiNGr8b4XydlosRaYOeeMjJlkXi9iOiUv2OI+IvDp
3oGxkX9RD67YH0RDAkJZsH4tICwGinhkrleh43Ir1fk6XNtkOThA37BM34O6qyEM
eFwUunAYBKah4+GcrrLFzEfNGXqLwGjEGa1PoYPosTZcRP930BJD+0MLDHyetij8
XMDOo/B1BWrch7wLK7OiitYo0gj3Sm9NAbE3WOgHR1+ygOIDNJuVBAxBqUc9fAJu
AfO6Lg/4MiTEbudTRaCRJY9a15nMNldpduh+BAT6N0G+9CwdWhuI4KlnT2FEwtrj
ZNrfZ/hY3Gy95R0pxLV2r5eF6BVBf153AwT4SF6bXzATJkfNJwtugxXVArQHTIxi
hpCy5xJBRgBl1E4gz3hU3ulpwTiFlY6iy17v6VMPK4PMFhYANsltFDCkNXmEgjWy
2D/Sjlug11eymQmdBiKIFLXCQRmb5MEgF2d7vhllMNmy+xfIH5DsE5m2niZK0Rj1
2dKN2S7JfYVsHNZs077LFnjjxaoT7e3NbfV7Fakkn/SJbIRZKiczkD3SaZ2NuDNO
+rwPiC6OOi28ni3JDAsbob7SHZwmYBpGis6i2bNlKvxGVK2g5WxvBXunbICj5bO1
pbTr7klWzUX3yw7oTqfBgWr4PDegDX8sC5vuFLMOHe6T9bOCDoLvZti9V2pZr01Z
xTXdOqdGzAOiaCiGMQdokvm/dRS77GpWzBmjsNbOA3sU2tyErDGe14+XruH89+U8
BXB0KGj/KWGoz8b995eg47wvvKLVXharmi93n22piGsR4d70eN4hBIfmLKBSQIPx
8fAS/ShQIQJLj+ie7kAhiRhcPCUmMlH59QairOdmNH2ly46lQY4t4FOHE/sc8Epu
IeylzuQ3Q5bmlbV15UUKtX9Q4VpnFJmeofBvXqDyt3qp45jMmpdqvVE4OtRAGVBc
sG0PLfEWpaQc495ixP4/K//s53il7WZ+mqa7BrOr0EOAcIJXn59Nu4EVP2LO4a82
ZqPNYez18RYLi5LMgOmwCz5VL4lD9S8fEWGCqCEltYh/e/DPLeWNacVBtfdaJOcQ
chtB4YBahxA9LO1obFt1vfQJEenwfVk0HljGrOSIFl2HW0DcdsXtf4NQB+w2rM1F
hRheFtWqFUdTrRsYExGmsDp4f4x6EcN0EdhdyrkG44GsOp8i2iVeH9SV+B1cgbs2
DETyeJzhklNYFIaLEJv3ieejXc2IJ8CaRBIkOYLUj7rMXUPkY02vrmwXxf86DBnr
d2tqwLmknhK81zrZnt1mAdCjLODlky47D3sv8KH/RhJZb3NR99hrD+G9ity2BDMn
qToS/oYtuI+v7+z/5MPzOBEXBgfEac+spGsA2MbDoYmuChhz3UqHKbqrKezoh6BG
G0mXzGimMXNGjWmT27SMl1WNuAV/OH6F/mUJ5HElgOEd+yNzt6Q4qEDWbNwFzpdJ
8JovgOr44vZRDXCEP0mt5+sh4gJGIeC6O+GliozCUs5UkBBKpKwaPJI0U6AHx0Wt
vXnT41x/Y+r71or7vZ0TG5w5ITzEsnZpniJVQ1oZhOpzquTtk9W2DDEmPLSvVD0t
41DtlHerMluJ2tt6XKqP8noCzI8nla7ikyaPRnf1kJg0Ndms6HaILIIgzyAw7GY7
HPGXyiZkMlNsz5faEkQS1QkeLhbYXLIqHPyKhdymyWRCtVpeGgynq1RI2Z+uj4RK
KCtUDy3hs4Eq6MtGBD/mvWWB8t5RN+WOfn7POH0C3EYmR9lv03SZBHxo12i23K9B
OSKj4wbFBG/QHI6be0gj98YuJqiH2UqaAM9E21PQDr2rMDoZj6q1j2c7O3gTvds3
hudqpK1iHAEs1xFXWn0j3mFao76Qr0MacrvE6ykf7BDdsv029vRCG7gsd1src5Bj
KEi3GkUXdsCuDj4efUKB89A2OlHVUDOEOT4CTcSXIVw1RBMOyhgd50HXeK72jAw6
CsQf31LvNILcSBERlsx7xMuZeNz97Qy7x7/vQQ8Q9chkrUaMcuMOCWhyD/9bPTXz
TjTv19ZdYUAmIHum9xQ2faUE1y43JWbfgKG3xmebFInfIpmNg4wCGSF1buY/jeyk
ItTanMZC135RbImh6kKItmey/U+rDT3g+i15xDTl0nqXGIExt2VERXcgZGve288T
RwZBAfzvknWryCMX5vu2L9UaLDmESBoW9KHddORZSKOn9zpUZAu9Oqsi97lbP6ae
b/zeLAyoF9m8IVF6g5m4HilB5Tw4ReYYwVqZQdwjJoXEmwV1awcJX9NTBc2nJNfQ
/UnHIsXAcSegyLlE8NfzaLb2vcbEdAn3Kd7zPsmb6FYtvqA3g6izMYr1v/AdhDB+
Wkss6ymDQkuOgVGb/T/JvFJqgY6TsP1RUVfpC5DnMTkrg9UoZ6rrk8O/bct9K97U
ljFjNr8vGN/UgaNqnZs7mMTef2Rc+s9C/mVNxfjpiLf8aQHAYqeFlUaNdNRAXuU4
OSY/H5Pq0w8Cmr9nvRCJlqzhA6LP/bCJz8F6+uR72IEafTeoXE0GUM1gn1hbEz6/
DFE722FDu4SXc/I2LtcAxOcMhcZ65U8b73vOj2Z2/Y8UoUiwM0sKxYT7OCZDN9q2
WPV5+hJeg9sRakQyyJaJfA==
`pragma protect end_protected
