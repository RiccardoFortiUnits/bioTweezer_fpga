`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AJf7a3+ZuuFxTRUX6UvYPvzBQphu88gi086KOGtgoaHX4JNZ9em6LU7MI80tCmaj
S6JDVzlKraZi0wJ/wT7bkDh8RQgYeAMuq0sauvXS5THsE9SjOeLo98BzR7qjurhU
yIaCfU4l4lznDIFbLJoM2gAi/4EIVupVAtpzYMd/Hzs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12336)
V2HkoxR1JJBtpNbp87yf4LdFIt9yZjzh9DfeEIfxapGnwYIbDBgqk9dvZXxjzWO7
cWVhKYgFTxzCKf4fujuJ/pAX5vS5h7Wy1nW+5/86n7ULGnQsGXNx6mM/iwbhWFqA
xqGUrvxlXiaJDPD/scWlVp8N7J2fEm/6DiqiH2jtYRUqbE6QqGqagyKD24CtfTdB
NK5pqzD6oGMAKLpXePqPFBZhXLEuIetGILugMUgWadriMH3eRmUNLsWGXofsE/iM
g4mPxp5FD+yN5y9jm/wIoxWfzRfumPJf3k3UsroUMu5P0wosBlBLo337oKFIpmaY
g/xwjM5d1hlpNm9/MRecCcp/EOA5Ah5Ykj1ebzbSZm39tmfWUyCElMAG/oY2pFM7
4fyc49Q1EtgBNmSvIzSFTqDHJvs/I5Pa6V/OCcFkbMnhnlimmqa/xnbHkeNwfOdc
6HFEu9JhxfeqnU8mQ4i3KPq2yhGxJmSt1gU2/jDuCGlSmPv5NtXh5dw9TTW3kzEE
oOzmB/xmYTx81qgHNIp99/b6s0yj/Ky7JZEnEOx8CwnRX3KwhfI1OvnPWBGeau87
ixabVnsifCtnt0zB18DgJW+MYSftAcyztQ0WPeE/FLkKppwNBMyXc0Q5bThFhxzz
cL7ytab2Vj9hHmmAXuv9q4ujPYBa8bTDA6ZNDXU5f4h/DfrYiGiDlAFhOkdDcdLI
jajn0GtCMrdgr8MdJTvGllosE0XjFCFyM34VFPOKXNSkmmLeTAKRa63ziVyndYy9
zwtXeJz4hwqbaUGnmx32WxnoG4gbhSrEDHV49wEpOH7H34yYI9HZ3TFZDy1T9N72
WbJVHXGJwWkSg9uY7B9TuFYa4Ge31E+AJxkLfeY8UDUI66Q2iMIjs7nFM6v7fO+n
pgxEg3m3a3ePJ4WmZjgsS43RyVFPQWSwdOpTlHfSj/4dE94QY8JewDTxnCRNEAft
y0cZVT/9mkK4tTW63DK94sIG8XzqM84lv0nTqmEmFb4yqy9mAHCYcWTsOX88O0jF
+n9u/GLGZbNqnUiQ4B5VauHiB8MAhG8KzEa7f6JjWPJ/SSywu2ypbTm/oTZNSri2
iwqg/4gVYUxUXVM8I/jFWZtJywGHj5YGrs+1Z4dg1bSnai6Tg0y4jSRm3o7MFDr7
bVB5RhRF+XVyofIgEmDd+a1PZWLMRwWScxM0J+lpsRtGwLKDroyA+QSPlYG1ZJgM
9JGfCFR5mNSnVPCh+SykvmRepekqcLf1nvEJaUVul7TtR7FAfjcAo+NJtnxhUdwp
enAd7ZI8Oz8hipT6AC7r9i/zYFhjNMOQRu24oNMTftfiOgWiIkBBFS7TRg9f5i/S
reLxWizHLThRNZYkH7IhUjKryJ7PIbh9fWiCep4gtWLuxQdoEeqm5pOh7nw1VXKe
f24Ao5nuDKFvxZTrncEtey8FomKKDsJtzn8EwpqJP4SpWM9yW1cBFipZ+5cjroVO
6wJ+ScygE0yWAYsgd8YnqR8RxV8OvTjMdiZl7AQDG06we2mkG7CvtqjvaeR0327B
+fqa/Zm7ZvgyAyhQ/fULwp5EvuJ52pkCPoai2kF9y3yHdXEGgxxjCf0Z5/l6RccM
Bk3IBvLnIGx6U9en59aZKPsg86OTSZiYmgoJNdXILUvaV98bs28vXisM17BDxnqY
T1Zbj2IReMKrHIxedchux9Kd7RFGqD/glrksFvr1IBkobK4d+VhNTZvaozlbfkGa
P5eWOI4W3I/gGUmjPQ62GNv4L0QOl2/0HtHeRSupaj3ucIsaTrcYrOkdyN1I4ZXN
GsxfAw1G7uDhzx9Tmc+/YEL1rB0UY64yuAM+PqvxuXbnOs0ElIcfsHuXaWoNPRW6
3AaLbdCWzIBIn4Az07GTo4f+HQLEmJ6/PNakCPYk+h9SXW3lqy/7JLX3gWXNS4i8
iHGqXJCsT/XXSySrZ4XUXGJKeKuWkRS0ywkOOkjIsvp89BhGcmZJvoAEyowkma+R
Zg76X1GeiDbh9X0DzLSDCFE0parrHvASHoZqvrA5m7lpMuuTvfr9hojEYZqUf5KQ
M/LLLFvwVW6XstVSa0oSlN7hR2uMDbfH8Q0OqXu3x1G9GPFSaZ02GYnZX8/i0wVq
kEce9KwTe+7SLRF0mpoeI/FqzFSDpmdthsj+UmxIpJYStxN22su7PVXGUJ7LJUp8
zlDImPF19kh2YYco4lz1Y8WIcR/MpOptOS5UiLz5INaCR4EzjBjc20GKjhNUr4wx
vwHUl0P97BjalfYaqaU2c5PGGvsUWGTY2Ox9ZPbgWCaUWyNBx943QowKSI8ejHKW
zN09QINrYIk2MJ1V8G99jtZW8p8pQBewEsu6GEEXVVThgUNiNOI8cYVz0fUV0Zk+
BeCHWKX3ktwygqZLwT1aAZw9FgEHRt4saaHXT6PbJPvEukEh0Fds5eeMOHYaYh0C
RjPKKBRDiCVIFqB9AJGnQ9ZS8XsdTSwZnvEsJhJoDENbZP4FczAWWWK/WZSUcvmZ
Swt53kw/amf5k7l5zyqon9YPGfwALyiZs068fSn8x0WBi++2RG1ThhpVsVorvSmf
vYsdg6nPQvqEhb9ifRsJAeaNq4LVyqzbAD2cfh5lg1CgsQmaVHIkReh2d5RiG1Aa
bNcRgUpioE6JiHQZvjQh23nxupYq9eywpsL203djnuWLe2CGu/oo40oyK7ZjIsyu
gbu7m11LJiRCue79fuba+lo3qUuWToc+roi5KnPgYLmcKjfhWNAKonqj74QipfbH
iiegPfHlRujCnQBDTnhhxsLfd8wRGZiO5gRPWvvmOfIzd7k+3/KZMxMYZqoLta50
UgtDQ1We+2c6Y/AWxKEADGFWfYLT0XsOl4owRfWfsH0Q3GP5NhMB2bW853TbA3mt
lNPg+7Vlo7qDA2vp85RxWKxGJ3Mt2CxNGrandZD4oxkvJpkkaxTyCqSuyWM5CZzY
vBaVqysIeL9V7XjFQqnNvnYOht2CEcnuogteQfZNWy4mVzVdHK+AW0y3pyHo+sVF
yV9952XEzxcvGQk9B7l6qAzODMbaUNgwV4M77sXrYIIPY7JeXrKb0UKpG5wVhzz7
+D9z/2yGnzgnkkk+oekiHjtYFOx9Hzc2LSwtkuRA5Zz/sCjz71EVQhJ2dgKGHkr1
bESiYTE3XBVInpdU2puiPW910/xg6OxdPyppDQwKNy6E/18+dss/G7S2AYeETjJo
5Di+1X1wWRQsS3IJHbTKw7x+rGdkVy86GK3VEUKqOztwFDg1OIEQGYPHA8Qqc+mM
9EoH0zrSsvAqVB8wa3jGaidLuLiIE2cD2msidgi3cYwnphJM0+efQQ3LljE5tPHK
3tUa4uNw/1vXHtR6F0WCgO502qmYOmIx+4TW7pu5TDOkWDTFAB4A9HeXpbFzbn9X
IX5gvUzZ51BH00R0cKBhgwf+Fme3CUZQsT+WcMwj7SDTgYTTEf8bHKjxlvCnbmab
ntXoQTRe2TgqrEv6wLs2vZYs3PfQE+8OW08VOXEWmuitg4cJQodN+6K56uMQJ5oP
ZK86qWfPKXNY0m6QaZwnmoGgTC0HsdzIABJ9P545uw165EoOtkoLU5GMuCQ289vN
yfPM1U7XzIn1zV1Z/m6C/uCZH1bGeHw8kkFZcLXO6yO1UVSbUu0g9b9flyvr9dGQ
6Zj9vqXntMkmXSNWJEoQGRlg6cgoXfoNPwWJOQUnLCFmcfkhtHjV7wOFBGeZuKak
ArpTlBQZvXtml65CYg4r3xSX0DAKs8u2YYk+Qx2frVF+Ozj3GddxjQ8RszgMSPun
+1o3S/pumgSns/rsAyx6Vvm+nUk/TTok1Z9uZ0CGPfrTp8utl4A+zzIIBkPFKO33
xfMnPGpbwfEjhEoms+lJ3uY+Ooo9OF9PCwNI/Ao459vMRPMx0W55VKAu++YKVjgB
WfMEuJj0C8PWJqced6SJaGnDflRfCsVCkjHYbrHD+d/+cTS+MrysCKknNhccqdlq
tX3x0jveFv5+KljlW0odNIMsEplYEBVGGuBeeZJtyKYyZNtea039lgldwRakaYru
xUViEj7ZB7QwcjK+wk07SeMhzWFP5F32eJBU/WuMqCFtLScqrZCGSL1ILN5jLFpj
+ZW2Usp8+M6X4SrcPQaS7K/ZXaKZxoPiug3EJJ5zA0g6gATWUA2c6C8Y4PEZEc0T
AzwdWqiBYKF4gwNzGYkb/hqp7IkgtebO4ytKMt/tVFGeChFxzr+QPjcvZcWZu8h+
aq7cq4uQVCsmJ0c5AxKEP24YnYOuf/V+N2Ttlav1efGQckafN/bHqv+YKQHC/dbx
Lr0LVe6nwi9qJ8+UkRh7QYZS5+bhcrGKgt5SC+FqwJIna5YGDETySjH3No3mfLFY
eneuizZ+BQQ9sE+b2H38hhTXf9fAkx2xyykk9L0dyBZWraa0onTw8NqUAjdEm7lJ
C7h9uAF2e0Xe+t2yZ2EUIRXFf67l3XdT5Nd1n5PbU/MY3UEN+7MfaFrmpCBiV6J6
lrwC3OzFWhaedL8EhQ0yRd614vX8ssxX9KGJWRpTr/JaHEt9esX+T6FQ+Ph1k1sp
+jjOl/RccPe3WNFwl3u9NfzxDPjobtFD5NLWFKwJrhw9c29QA3merxzF6IXqthNZ
r9DQCbKpqJSZVwE+v6xD0PQ6tysNKQJNCwWmQYm9cSGGEyBEHqmQI7lXd5KxzhUs
5vsfxzichO65OBex0eSGowYihUXK48sSQRUkScdI+lyggt8C7nrM6yKAURsfZC7M
Q/nNiByDBf2znYebIVJPgAjl6ki0LKcNzoQ7l9G1RYlwMT+n1lKPP7+GcfkyWayM
FrQmjqHIhCN39r+V0LkEZFhXiBM800sue3M5Kg3k6zugLajLV+kn+AhuWfQDv2rJ
BQKdhYIlKXKQ5sJFK/ocItSG8eQk0dEMmT9gsVzTuaS3hLMRSgZblCO4yVeCOjIy
LdtR0TosDfjS8nr2jUZAvsOGuCnSeiOSpk4lvj+etCR2mtH3C7lASacc5afUS5uH
2X30HGW96IDu9ZNIdHHSZP0gO+1gBRvbLXO9oCs36AlwKtzBLzRzJxNrZ8xlq++K
dqdr679TVqJ25oiu0b7daxLoYB6eJy5rfPyPy7PnNnzD/t3V+02EHOaPHh0SWDnU
nvm0Aog5sxuwr6hTmzfHfBQCR2I3laOXUfVMgTiSEoT3rq/3aEA3FA0xXCaYajxX
R3qP5bVKcf2kt2edsrn6rwnukFUrXVM9qySSAmv+z6iJ9UiIaepKGbUcgjLlPzHH
iVtk6Bj0csvM6K8+JihDt5jjgLG/VRxIAZR8VxjAuIbXZVP42gfQcrZruBpWSWTx
FOKPbFEaZ6hHwklarBfo3GeMPdeiUeMcdyNjweVxISSBW5Y/mH4Ep3tSFeaXcQVR
fA38PhD2D05OovtalXXfSA8EeNdH6crKSBb2841bJpjCITAaVZRaCL4gMZ+IfjYq
uOF9mpd1+r64QH652z8lpYYXr+IHLL189qmiymoq3DCvwCzeGHu3jMDFHxaccZKZ
n8jypOBfWxq3uaRqaIGyHekwkvaC+jv6vNEU5bdTflrIzU9353S6cdXQa5TkbXlV
wb8I/mGBrJs3/XeVppCdp+CdZyfMvju+DJz2wfBW0qF86qfPwfLF88tEHdjdPSNW
LZnb+/pnWqolH/HyRa/lFk6g8iMX9YEz7PRNmqm7wT7uKqV6bnTpgCg3BYNupoXi
w/lC7FvOZbkuxok+VcdlwUd0O12Yi5VBduSxgXJlzrnMTXI8x0+LDfiATqg7snNO
h9z4J/6EnGGHEvHr60qpRRkjm45kkoxJj3hruTdj1bcSuqk/CT6YCZhdm2Vu8uJ1
xS5tzuFdSKwv9ayEtPMRi5TkyuY26Z4pflY7YwyIlpum1VOuJCQ09mHnEzt0q3Wh
gTeGsp/g0bJI+BSiuml4WBqxYzPLCdO7/28riwNIYXyRIohTePr3PLBZV2aUifdK
CStoBT5FceXCXWWncNgNeTnstimfQDOCSUEmOsH+K/ZYPxpa3UE3evsGr/Do6XFa
Xgvy/f7v14/6Ma6RbQKi+Sl9oynZYaXLAmab9hUgBcceoy3xQ+UFrqOU3xxMP3nb
b4gNCaSQt0yIpdUWHK9B2tFd5+M0E/BgHo+MehpUtbAQxfa1w6jdlhGPnNO+hsKO
eIRwI+8Ch0R1uPmpOXIIP9DoJkVyVEYhDY4tMB2mdKhCpa9GFngAiR8EP1sv0Qn0
3uIbBOq4VR+oo9JF0BwtQYDtMGzfVgYKGT9H+ePCVlJZ5JeeWEx4pvDjJuI55j/S
Dk3Pm0udtAXG8O2kY9bqD47H2A8uga59iL13PvJ/giirC0+bpVuFNhFuCEmxt9wx
94nYEwVBxmZbdV1LJg2SdUzAeiDt092ZFmfz/AlNz/Pv5otbbosmnx+BKd7A4Qs6
i43NfnEoYirGB7YuGOcXvwxL1XfNFJ0aLlnwmu4UBGb9WkcIA1NTuTx9k4WUPWXe
81WXEYRcsglV2828dB4j2rlfItAsGUoVldumxCjBbg6i16x+FqKG4NxDI0yPvrEY
s/51mgUmtQzkHyNtnSB1Unb7evllPATStS1NvVZ7GimDgzg4Mff+Jy4M6wi8d50h
9EE27DGhSuKPt9rfWasNuRPDiX3iFRUeXPHJONnzts8JGydHyrXzHV3AlWlaLX/K
4//lo8fVp8/hEdSeTN4U542GXIkkFHwq3p8WGBSJjzrKQt8O3rIntpmG6Mqy618J
bEtcC5uyc+Z4GICM8OBN2MbkdT/H2Zcp44p4/qkpEuXPgUMBkVFWRFZOIzqJ1vG+
c9Uo3xbRJ+KEptxPgNPpm6kW3HNC3oYf9ceyjAAMee8nm9D6YShTWLMqx6fjJZr9
1xfUIGOsoclbLE4srrETCfHpdZ1aESl0/Z2Vum6+vVgUnNPImW87zhsJJjQd0dHO
bQgEIPNNvkG43GZb4FQJ1u+S95enmMWP3Vk1Ew731ZQjnBHAIDTbZxkQ1YM0KXdR
/4e1EYRq8tyicNRgcUhWRW7VMJHT2bKCwNcCWiR3lAUcMyTVLRkn5lfyEaJwUqfd
uQznlljgUTjgVUattOqzxt6qqzzohIpTziyGroqaiWQiUauL7Jj0Xoo+SMIgM2wf
XeDi66l2+AuGSBtR314gV+iCAVX7ZVDu2DveVowxCe2lujloOlPoAktzzZGOOXee
nDP5MFui3Avk7ptdi5/u+zQk61brch6xsE+a5+TX5Br7+lGCkEBuUO+nrKgahNv1
JQKEPktibHfKT1LL7y635QArNh6VYUYINzQQzCykSxY5mrMDovDl9e60GbFLg//0
Qigj5obGFNbTyifvyKdOHdixDG013NDGA07pMMXEEu6wxv73oHClMQhrdIgNppnT
4Esjm3sdyiTsz+ze2PLxqma1Aw0V6437GVmF5VYUG+YZ6nj9XmYArKJ/rBeI1x2Z
hdicvD3AoqHtw/3CrfZgS18ILsYTdRXdllbdoM1mYc2hU3lpjWjiE9dqwOuIS99U
KBUGkja4QEGbyPHW7Xmn9atrg02JO4cW7qhejX2qOMVUbFrSiOtQHVkxB+VNW/U1
iS+TMuaJZ9citHLJOBASWnLTzdU/oKiNDibMrZuAJnUnoVpRUcN6vVRZUo7ud6+0
dt4dK//I3OB8xsOgjYnOvALYU6HEg4T2heDNqgpYY6AYpjAz8SHagSrYxsshNRAC
l4HQiG9B1b+smQWx2XIgBlVAbT6cPPevjSJR1srv9hv7IKvyKzmXLuu4BSGaSlxt
AKTky6whirnelfkNlNfzDIoCHu9M/6A/rbXCq3Edz0va6YIHo0sSBUFvjlzF2iDG
C3MtgPbLAGo+ofLNnHLuvS7uLcDBc8g+5XOYDuspukPsgSaiDFl0OP0La5+fXiyl
aZ4JyqXmKa2/7gu9TiA5iY7ZPoWbaUwzbqzsccUfTFvqG6asHb8asN34mZNYzoWo
icVaTHZsQ4iUxgkWN50l7slC137vx3FhxbcHXkwJONlFFi9XW6kAiwpdl0WC/Exz
S3YFj4lyZOjQygapXIokfYELV2F5LuAdwTFTrQyaxvJrm0izNtneIn2BQ9JamITN
09n+wnl1qzz6pEqWnF96HXuetH99qfBZPP23PIT/larCp/oeF7R+nWdMdJ5ZFKyk
zqYqxrwQRYW+z9ntaNpX3o4q7VvZbxYgcz3ofLSv3cCVlo+xYrH4ire+FPtehZOO
FO79rn9C0wj+ieR4TjKXoFjCC4gbxMXUhtQsuJw5CTFDrth5GS4E0UcFeDiBhntA
9kaNUHvn74hNkbozKxy1gAOYuAGQphGjKnGNNO4Z7La3tCKKmqZk7H43k3diG/E2
iCo74iPxqp0dk3U+nFhG/sDP0G85UwnM0AQJY4gfLPam93G2Urb2vr9JK54Ohnpd
wkDQw3Wpewd7Z9Sy/wrGTwgfsxeUKsSAVH518Z3Fini3bDbPgxGD32xCFczu9Ow/
3XeoZ8u9BIG/GtTtNeP3+jKYG7fXA8loEpvmPx5bex8aBUqITQB3rZ7raTxqDVWZ
ZW9CnOeSApQqE+iJ4ytg/cHT+bRc3VcYKv0OLiokKNcReX9cQ08MCYg/t/ahDvBm
rVcpC74pBh/+hQ7o+K6RCdJMGrM+0vGuYRuMA13CAkg6CY5x9eJjWfvZBm16Qd6z
c/SKjl5XsWnPegsQMc7Fol54QoZjzFIbPVnL8HUD4yvpMkpazbKlXY/hl+koayP8
P0tLNEHKtoDTeo6J9zEAGy3Yhk6yO/DlMB8v236cFqlLK+afd8b/ajL8AONAvyP9
X+dofamhmyGPn+j1pkUKcEGyQYVKpvaIc9CLQunccjMxple6/k4T62WRRef8PJPh
GGHXeCqdhcpjfbyT7Zd1xHOigTIj+0rHeNyncclLJs2lHePpuFUqmCxDZCKhPpbb
sNF53b3O99ik622hQwJp8cGa1ha00QH2WmVQfXvCpi2zCORjy8Owg2cKwNMgMYfY
HcggGEZIpazdSefudjHAT0KyoVbQtXfpx19Pr1TFzP5x8DFDxvAABKjwD2BjR49p
Mb64viCptszWNhP0uWYiO2KlYM+wiMr4Gil8En851/0HOFT+m425VC9Fz0r9mGtD
0UV7uz+heqO3HnkNskZeMYkiE9A6qta7OJGwUzVo8169j5wh6+NrVyK265uOZoPZ
Zb//jKt8PO3bEoifRd4BXGmX5zdrcDu69sD4Yohk5Uqkg3pZ/nb4yWcx17jD2/XZ
OYrND0h2Hhr4jAS+ZM+ALKkECYhmsw6nHJfziE9EyITh+l1NSePeASrUfIYcCKCn
m7PdCxvdNi6txOubNhhpkjvaqWHC0deRFWNpWyhveeLsA3hZ/rUxKqmowxVKg/3s
wwkxILdYrwnEvijvMcfkN0JstbjlZ54kZXW9Jk4GA7V6py09SPeZe7K5od83vcxN
lYQmaGQgE+pUmMgTFF8F1VlPv6WSpl6sTmwF7H+oKWja7TQPhpR2w9azgSx3q9gT
wc+MWmYidKSMhZQJE9v/FoI+7mCU02cz6dR7c02+gnrWWQaM/HBB1pXAN485SJtz
vENPCQhK285Acn+wjLlpSUHa10f6i/At25/PiAUNWuVBtUAx1o3fyRlXkNsCjicD
RI4XokZz4QypL7YEVcR6m0Vt3uE7SacqQxJsNfs7qqLKHguMZSnSOXpG1ig22pQg
Wzl1IoUyHh2SwIL3WVsHPuuKGVU5x/8fmTcbRwbhJlczIjG7qY4SgW+t7tvfN+zN
nXIebufeptJPVbpY9EK4Oem6fTE4ifmjHKxKj97fmovjRbi30MVIIk7fJZ/aF0WF
AGjBSzEUq6J/YDNsbsXYt8AE4wMRzvp6QziUh67vS7kur1WVk4yk+C9ASkWwbsv6
6ptjmx2As0O8dgL5MmcKSrRW0pui3fDaEE8YvjUm/4Q2zBct5JYdWYbWwxmP62UR
Kb3R4g+EIHaqWiHo6QadLuBkbnQON1Yq4NaaNSL/VGHAkueMy9Tbs4M+VsUCt+Tc
5xi6PSkF2+gJ06fPCaaXsp6pwCuErGIGtUPnlTpWKdQC7gJQRotl+ynXb+etANN8
kioHtMef4+QUhtR9V0WpFu7tc/FwedGo3uI+CIOFqcWa3yVndyZcTkaRZdeyChuo
FgsFo9bv6iQTsV13GLd+ebfBoXRvxxwIBlYeIwYC9jlJgTL8I5sS25iGLkTjqn1l
DJegx0mXYLCRVpyJZr9iZGFBZDJ+FLeYGpweI61NDATkxLaiX/FeGII4gW4Hnoih
PL74EchIo4l/jdZwFKJHpLo6LlxmF2squGzIVjyinhxM/2d8KexvUXwTiDzz6rw0
/e5t8dp3onZid/wOPZ+MSb/aX7Ue3aNQGx+yfvcQbW6NsRSU+OTYg4rJNA7zbhBw
5MW20ltHDa5M2jQlKhxAslr+a3dQ/LITE2DIfzC35mXqqrEO2og25r7AlTEuBoT5
+3aMouhzzBEPegOFXCZGjRvDKDb/uJGviWe5vPmI+oY6ujuyt8h+wm7JRbvbEAor
dfcmY1GGt5m8RBIXHmaojEIHTmkilA3IP/LYfVgPOoLGqyfTOpT7bF6DX+n9fhgl
8zQBpcKV18RPMG4ejInQMWvPQL0C9z/ZGmWlfqNjbL4cTVwv76jw68t3XorgbPy9
IuSPfOze1qeVyzGganm5hoqGQIO8EKkCki4VAmzIFCQnczh9WtBfG1ZbKZFUkQAK
y+NCi6Bi1BMd3o4hAQeKBh6X9gluPXubaTvUnyQXARccBj4UVSfG+JloGPxgUn4l
KPvORZJdgVRGswpLDhvdaS+CJss+pNS1gaw0WIZ4WIRVbr4+tCoIx4sQwz/uhuHn
4xiskFEO9I+V/wOITzg7eF5faCiDu9uxRj/vndKOecT+v7LHOSqsMyFu4kglE2Yd
fVqmyo/4UEidE7LNk9Mt/wiurPbFnEO3UIWbzniWLXq5N3jz+57GmJYnpE6C4xbC
CDKuqm+4Oq1Fx0ClDgKM6M+ikD//JfGxEGPWqpvFDFQ++EA5QWvDGXRbwgzisGey
icu70S+wGaUF0CTWn6VKkaNVaRp3+GCXPd7BnM5tp7o2HRZBDnxMMjF9jiyCxi8z
EKuIYLmwYTkTTQ2ZwPjAiq/ZWCrsBUC0CR+2efuFFTGnxjzMZkV7PGMiHWIbhGfF
yZDz1CeAdanUoBbuvHbSqIzDeczDv7HNcPNSmf0JgNfsM5438AA6iODEheYSyPYq
TAZ5A8V5/eQrfHVQiH96oWg26oeIU4BlidpECOu1zIVOVUdWTGjHp8h7Mep6VdB0
e4kczQJakC4KBKlH7DkU2n4NPU1NqHVsGmlrhYRpD/nPbw8lsQIsGwkaDA21hh9w
p3HpvpU4K7luOgvgNrYa90OmYS1RVljzDEVPQu1NNFYcZp4dOHmE2XjqsVW66FeR
8Ur2DSjSn5+RVhrSdPwAvuX/pXR9vGFDzPIBrsZZrOQivFBturzl0e/kmkfiZ60t
WgceVyieBy2wukO/FR50X0Iyhz0SnOt7AFFEi8G8MaK6nsun1VUoI6jpJG+166DE
77XGsHdQt6G73O+R/+874sJiC5ypOnABptk8pOWd2NIa4vlbSWrJ4G45Ie4kfqHV
1fZLLb2cTybnajnwjsdCF3tzaH2LKYp18nNwgYwkUwG6fzNGE20qAIksAvEcfGkF
RVPc5aq4+/+l2uhxMi4kaeFzp7Em4lhJk3IrZlrxSDY6CNGGOaoDEIYXLL6V0DSX
3wRgCCoC8XSNAanTy3a6kScq0izN2ZSOfTi4X0dZgGiqa/hnS3p/LuhixzUX6p2/
vIqcJQund5FL1so51XTtdubXof1CDD78EeBlek4P59z1U4t7Q7c+73Z0A9tb2+8u
ZGOj7iB6fLiiU5iUfHm0Al2KWK44TV+a5j1BgSd90WKbtHoM8xnp7S5VCOkirvbB
65GByYQ5eoXiEubJE1O7B2So0qOpcc0DUDgcQMahPOuMtOCEK6Iy0ua2//vGgJTI
KPhMv94t84UK75L9dlqWxQEqWmwHdIoHy6jO0NfM2MUlYBMj7kBvchhwEbKLJXFJ
nNYHWdFPZHX1P83D0iRr7k52QYHipknBtkC1fbHNlD157GP4KdbncjsYILUXreVH
KdNGMRGNw1Lb5ZXP4uUram6Q/4HlK1J2wGP5rfeL0zAQUF/jFi6y1SIPFbp3v7X1
nGrEQWYq+85bYmQ+ipClEx6CS9odnE+R/t/qxLIAHwJWAOu1HTz0yx4o0nv/SlXD
fad2lVisQrur2WODFlGmP96tgsqp1bsyCwAQrOhstdnwebYTOhshvUFqPKkqWSRF
4WuO6OY7WSoWOpauiJR4boNJ8dn2KyFCi5tAQ8R6XSUL8ODX7vE1KENPua3peAkn
FUHIVdVxJTa9D+rt7Jwci76Ml4cYYXxvvvYLQQQI0Satu2HregPVYb5L1HQzHqZ4
e4EVyp1/nXOVlsbisW3Cd92/lDaLpV1NvuRovMbjUwxtvgTubp6ToaCDtbjP/dlt
HtrlQZxrp46zUWV9Yruoc43YzAHMMSSZLdVb7Anw9G73QcFtgQtuVkvQpJiRnDmM
74nOEIJ9xXa5NBiz6fkGzRGIcKgj/EO8TGSDXm3EIFCsPb6too9obROFWulSDJoF
m5x60cHqb+tQf2EehEhhwhRzy3Ew1OF0T/8XvwkKsmai+y/DS/Jku6e+tGm5XjSl
JIOXrvFxrmWnKZ4D8YzWYmqwF1cVa1WMS6KXfyuLuFevopQF8ji0mLT6cZ9qD8QY
0FOyuqQGN17FHLFejxY8ZXbb9SCuizrMOSuEHS+kZMWfLo6w4IrI9UxT+xd1x24r
WaB1w4QK7wusgXIrcny3Of89WtY915i0LHU2D34Oy2N9QIDnL5qVz2f52Vl+UBDB
LYGRmRhNGkiLTZUnjC8Bo+rQD36tSl1ZBXLqKJ6XCWWPXQq+EVxqDTXh4uq0SaWr
O6UtbJnpwtAeagDSBA61Rc9BBPvMTExQwH3OfqzU47YwTfGMqWk30bIRX4wfehTv
13mu3pQnU3UkV69vfWYOEf4BbXs2ynorsv+SoayAYCKkpURXsg8gMNnvqq7eMvRN
o0mA1UC1L3kRH8yetbILocBNgTjVsSnnVycZrMLzTFHgHGA8HIoO0/QQn/aM4qgN
0EkBgHjs7avKv6upUF8AAU2zMBfmII58TKhota7O1eyFcrUqpX0yMyFWPsLJudSL
QlCwpWFpTcdjCBOg0Y46+nibPjLHAuCIWWhQ6tG8TmwliGoZHmjuL0yz/N24oDm7
F8PwJsyKz+gW4RcRKxJU2S+CiDA5zOPZSdUljBAq5vAeawnIwPpcEAFOu3OnJCeQ
I4vhaRk62gloPZGDukk+aKaVgHmR/aNNYy8lrhwKqnxOd3hBTC2G1UYByZAhPSog
aAGF7El6l1I4CuGzXStVGXObtd6hmTA2znoWcj1JiiW2KxWnsx0/trjThtTcVoK+
4G0IQPzgbZtrn9Z7IxLhQgcLIm1HvOT7ryGvm+Rdb8kD0uCqsA7wkPQ8LRGoYvPt
LT3tAgWQ58IdkbeCQBW6mn2OK4B9oS1PntbTwAC8f4aDYdAr73liIIDZ1vLZ3PbA
BQxiboW80oHt03/vs/1jH635A3Gfy1yRUxWC5jDTANb5AhYBqc6yLez3CVuBuNAH
5JJ2DExHwTJEUip7ebTknPv3lU4WYXOUU9aR8WaR66gFYC2xSJcGOo1eqfI5G+QB
7VY+n/V/aWmDQEL4P+9dPSF6iKcDJ7p2FBhqbVXVzBLqw2aHZ71mxjS5ahgZRbX4
fKm+Poue3wtveujpmrUKakPOu1DqiXIChl5QkswMa/G0LEaNHY73iC6v+tOc/jpS
JWInDXj9tgErjKHaeNErbUZaILZDTn/7vd55KJLwtdmLMCsqIQKbeYTH67uVIrm1
EdFte4Pq0oCYkW7oJsDTdVq15I+iRjS3Wz4VF08wB1Q1XZdofvYwXe0kge1udJyL
9jYkmhFg5FNmnN8RkAWuSORt/VRB7f98I3nGv+gExCFnYtsmKRExNIN1X5Un/c+9
YzzU1SUrBKbl3nc23OAWChgU0p8MRAacCqnE9/5g6E00BlYQ02tA/rchVGytM/U4
bhVXmtStBlO1X1hsSCw+n3HoX/NqZvVRUlW72fMjPb/GcRHf77bxPahS49ibx8/K
gtN7yGxH9XQeD1DUxIWjGIJ8BQWIezxomU5ZjOb/vUGk7Db+3KlGYlpcf1vbMirr
rricG3e/Lx+4vsefRN3XuccDkiR9j/0k9wewqUhRyLFlhoasipWhiIwML47FJhRi
1pjOhiDu4GeTIp+mUN29QBmSjTQXVk9IgjK9JIX+fV2W9wUds9wzo8oTyTkNuYdd
iCFNKjCuR3EXhAux5ooU3ag68NGZ2doKRCzgT4i5y1j14Th2QuvFSbYbnmAwPbw3
pjdqxxdDYQs4USANnQE2sBFaE3VtpAv9VfTeg0qpukrC4lKIQqNgFw0Z78y7W+im
v62xN1JUGpyP+Otn33BKh8jhajEiZgdZYy0AcGEotSBGdjUst/DfG20T4nEohlIc
cQTS6N1rZqQkteOj7e+3Zts0s8wuCi2mmLFoGnhiFS18SS1xdQ9DRgwMPMqs8r8v
wRhimMdA6J5Ttp3L6LyXSNbEmlTxq9W5KWwUKpHmoxcjFiAwBcXqPh3JxYsshREZ
NRl5jM54HLjpliwT0+frfUJu6vMqnLRwHG9mEnaSDgwe0BhTVed5o62+UtGKO//T
FghcjPfplN4dVnvyCT4uouDzAM80YzDDUAMJN8WdaqofmUrv4DKcubmK/4KQIqib
iMBjWSZ/1XQ/fiC0a/F9TdOZR42sSrQDWikAuy5qHCYiJlQ5ZtSQe5m9piKuKvMs
JfWaWxzxBLRR5YYDTkQ6yiloiJWGJeXJgNyD2Ho1XgevJDamNi/GiLi685AP1mUj
lzeAEioFg5ZaDBzkEoQvxIJ9cVPtIoCZmkAfYxXANhmkEV8mE6cbnGzPBL+j5qpd
bOPtAQ40PMjM8EnIoBHCuUBEqOlvtGZVxfycqs99tllooNFXzwTnJ57vAEPoDXr4
mA3+wpRoc6YQOsmSYkNkgRA28oqBexPV61ZCUqMBjbxzYojB9Qx6x9QKWLR0oIhD
QyhOeqi19S/11SVFMk0eFw4yTwpO3PeUDz6vtep9mJRUM1JqeWo9/tx8mj9bDNCi
BnCC4ZpY6s2FPo03dzW8ZHMNKHy2CJVeEthPZL1Gi+8BKZuT+Ztr2ARCFYawUQOI
vuEOwFhGIQTPCsGxghWGv/cqGA1wAwpsco0rxgp9TM6kcFCZ49ddDbGLU/2WmYW+
qHEXaa+LKjym3755CN7SrtG4wgCv1+d63HxGg6ilT8vQsdRPvrzj/Ws3+CuMkTJ4
i8VKmgViH2ccievOZaZ+okmYTFVjU1ekIlfvKieZDFqzWE4lVHbFXsK7DbTaTahG
EQPEo+FzPo135lK9wo4OtvT+0VDlWnfOlOujJdYiOzijkK+igaNR9090Opt0CREU
O1PPGvhbJJxrpQNWtHSJh2dv1yiMQZ5MO2EQjJmMd/gtXYkp9RRyNRYk7qO/5VEf
HgBPRHePz7JtmqYBZVC/zl+WWE9Pro7SVSMHoKY1h/A/jRHW5CPkM1hSVeIWgoI0
Y3ciiHcjIpoDFlLx+5vGZzfALjJ7iCzF7ktr2970wcVZiY6WC7h8RCu90w0YcS4x
uYT7OfwKs+mWiov7mBJMPgPxH5/pnjAOa/AGDvLwXabUqCljNyPSDH9FnTlaLmWA
8k/YFQteiSvMTMrEjoazblqVr35S8ZrQhsl+xs0vCS8xGjAQXKM7j6XNU0V9Jxep
wPaWbcGa3j8n7YWR0hj4dXMcGhEsLW1/GLWiXEeHILvMVsWnjGG4b1bH92Eu+KJe
2uAgFpeqgVTGmFvV4Qw8z+5m11pwTjYXJKH0tvdtUjKxEaKHOnkqA7bvSrd5YWjd
j8NivBFbdbHZl+nR4kaAIoOTPsPdE5hlxJy65IasTm6GQCkeBYlwSOC2LtrsFogQ
cl9pkWjtrksKuA49NCBgUzxweXChZ9LARuLcgwU9INLzUyTrqz/XKW1gC01FzsKl
W9LE0DqOUIFHnZm9XLwSLvTr3UB1e438b7UJX1l8ln90mABohoZYZbW4OtNtMX+s
JwuJc7g5TDk7IDxmTnN1JVeJDpEL7VDaLjfaPYjAB4Dy7oJfdzoxTIfZvcQzo/3S
ymtU11nve+9NqwW8JwqZtBw52wLxaphmxEZpqaFxr9eNxUdASVi21ORL9RxzjFBe
6tsP37qhzwCUiUmN1jt3XkAmgurIeLzliaT26gFg29PXOa64A7J1TqiDNvCRy3GL
7KcNTZSWC3irOX9W9HKuSMRSuFMTwhnXAqXOndmHGVBj+sBHvCiFi2UUFLeMyB2V
skQymfJb5n/yEEeWs83bzFqJq1lRAVlqU2Ap4CVKP4b0iWk3nm7OUjquIYgd+vTs
`pragma protect end_protected
