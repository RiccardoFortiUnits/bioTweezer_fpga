`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Kp1SOmTXoT7STnQDEH9VUXR1M4Uq36yUCCcebBBiB2JZI9DE3VMrHfSUWsqvTNTF
P9tjrPr7VXBcxzrS8CilHmn7W4j3Hr4ElwdeBjL0IuxKzhP3RxVsL6muP+uVI9rq
IBm3fgsCzqjUSF3UweDreGuc1jfsDFKsWUgxGcOzzqE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22080)
XtVATCy0fjqYwAiMK3Z1LfmvB6wTZ/FA+5/HriijjH8OPmdqCLmTJxPgfW6w/3gD
EDA4+os0IHMHIcHnI+d6GPOdmSy3NGefDqXe4JZ8Ca7T2+uY6RT1SwVYkT05KbDa
0z6yxbS6TJTDGbjOxB6OI8vMHEgiMgSx89wRlSYpGybTbq7GczvQHf9YsaOMKUdv
EiEgDnlyRtMNVZrNVy+rlunWa/cC0B6NtdbVfpdZWPgHjMhEnvLKRmLjmXA8mWEC
rqmF4rTyVXd1jv2Tlg1ZkFPCUWDqKVYiadyFbu03NtC4S812A+Ju+IGQDKx3f3G7
m5Yhb12TWTMFbA6X+WBD41h9bRo19thb2LR6dPzEYEiiB9g29kkl4nk944ZaN0cW
1GYjP3Y7FzOgoKiOi87g2TI4w3E2ipLUibZjL1TY9dMs3m6exPwJYknem2QXpHhL
7pa2YhU40e+68d3oRGdzJDZI7hxmzAHndZnkrziAurWwQTygJqgRmPj/8o67rE7e
m352m9JGIvBSGnCPBEJmtt4CeRZUhjS9gp4IsDkMLoJV9RRIYNIHEm7ZgkHIC0OI
YvjABOLsyO676ys+jN/AUPldpMfcDZ6xMiR7wpDIEVoEO4I5uImrmrduPSbNYoCi
BQls/zneEt6QoZGA8yWSn7galO4ze1D7v+s8AgvMM801lBmaDvlqq7f7FiasMxzJ
TaEfusXVtJnwS962AU8CvvhA7di0LMZlwxI4lwX89fmljxqOTrxtUIUq1Cn9rLei
x8ust0qluFzOeuQr/S5BDoRDfMYnNxGgvp7wGDD1uu2m2Ftc5vCmV+gT0uWC6gTP
ZVcmp3Uhm9ZCMh77ktZI8zACcFHTH4V7T6lONN3ooeaR5CHX5KMJNajn12clpbv4
O+GL/TGw//RPrauNLx+4SIhsGe8goGW+ENEffSINrRuYLlRXfhz1AOOS8X3a1z3J
bOVpPHHcmKV3qcIl51sES7zWnRn3/pW4j+dmn2TtiwekpoEydaO+rS7iv6uZqVXo
lOfnDle/o94TdUBz4wDKfBC+BS2C/q+mHwyzwD4qZ81gVI+5RMgc23UD5mbrNjew
YoxfCTGVemHyffLOzt2B7bwNZGKWlEl/kNXW/Khq9Ul+B+lOgZosWRQQ7+lSzIjE
h/N9BbtFvcAV4BhkWxCI3wISjm/qKcJTH0woPsBODPqXyS1ZgwSAXqPWtlIAURel
FbsDz1DqxuEMJ6fuazoFHKOiFqcpgAIlW8Oi3YQ3o/z4srq2UcWBBfftgAjthMh7
7z83TwKNR/P2a5xPe+ma55ZBSRVT5P89BfdHrt24aao3/O63Ne6BnWBrb7vp2nc9
B7U+OjJcenqVVEYT2kHoik7ba4dVsRwZ+tQqMs0VtmnkMeJeIcPTqdhz6flvejVS
foYiEtxVzPx9ZvqAqgNsTg2xqscSdIz1NBXk/UF9Rf8UsTpl7dl2iqVXHbiVxJMo
3wBG2i7TeIuQ/lY+8kkdUtC+ViPWnq0plkQRdswZcKApuYN9eSa3Hf7Tdk3GU1ZF
c/0PgxWeiPs/hoEvymVMsHG1rxqsZTHEyC820NXT5Z/bqIEr1eCr9CWwgsyWnT7Z
XGIGywqvhShqtsreOc1ME62p2exhGbJZ4qrwKVi9D6MS4uGOw+XFT/Oy6b3BCVKd
9oa5cbwgto7gBexi9gOr3kO3pT0LZe4WeDQcAMp6Pxak0cA9pmiuDQ9pcll6Ru/+
jnWoK89pC3XJrqPseTg7TmkE4X+Q1ho93VUuOsAHqD06qH5yhPko6L2+l1oTtHAk
ZKfNElRsSv+zge8ObxIp78CYnKLNOLVWsMvypBFE7sdnb3Px/aDZF2oy6RVuu9bQ
pgnRIDodIYD6jAwOKn5SplWhSWSNAb5KbSqIy9yvoM2EZnVTG7N4DT9I9pRVHO68
bqMgtKiWI3oqHacwRV4Iycd7az7i9YxXiOxlKmpbemXcMj28YXDlvi+oUyJ8Gqc0
rEHRdfSodYMW6cX9vVd+Adh6r8P0zqT+bUtg58GsCiO8nv+enrqICkmp02lp3hNB
GhUwRtEXPZag2T+U941Plw2cTXSooaTTyRlyoTk42inlywK/4LPMkuWGu/pynzKG
xWjJZx80yqIMPimFkgfa7CPyaFw2qm9XNiPSuUYRIO1c85Aw+K6r4vPNlHJTxD2D
vOEZuDjIOI6zYgexRQOabxRyI4tYnFFadeZ9mQ3kpab8XmCf/493knFJoHsl6O09
Jxapuk7EsAlzeu+XjSjld+xSPTubZb66dC47Z2sOBY1wqwKxh0x9BtrTsvQ9A0jI
Rz05HAMKe843gX6uJ6r49bvIm1xeADDCtCAxePuUJMsWlg/g6S3BnwXzBcTzs50R
MCMg6Raydcisz4kiQwIWSYWMg8IIzwp5Zt5qkAeBCW7ZaKk4hZtg19Kx8hSbj6Ol
zgs2l+xVvlMpsLAdIQbooUVAIClgmKQTz789ks/YXDAecA+f7DXyv3oGYZzP/DXO
bdCqnl0ZByAvGjxNSDoHaUEOK+B/BXrQnTlWbaWbMAzxa1iNgOj1fe6lHYXfcVTb
l5Lzs8gCJA2JygJh5xBNMPjzlpkEqMfOOTtrJrpvMJj5A3xatPwcaXPvj2y0MDiC
/9q5QXedq/fmQI2AsnAhKYm8fgIybnXNuAE3Z8zA8EhigJa10vXdyrJD7ovRk95h
dDTno3GGHwLHVrt8iU5xjhL34aHq4BNar7z2Lus1/y+kDmbKfDvJdXbGNRRl5GLQ
MkLcKoq0bCcERftDbGCp93WQxlA6GUkmKimUJ8PBbFdWbpQKLOt1hcO5JFrBp6Jz
/d+nNwl+5OWqUV1aHv4NhyvVlwBgdJDrSQfEvDaq8OwezbI+oJq5lAwgNwY5rBB4
YyRbmLxHY9S5p38yWqa0JMQERCSJa8klulQD3bYeQppIGaGX2rqbOcOzbKAJbwMC
FBrrrigvbqRPaGjz+kxUNvQ3hiF1SvicJpGTQZWNtmjMf0AkOHfWH1iEkgLoACkE
H08GpskeK9+G8dzwONlb9pNZBibCe5v/nHGfo9ty4fW3kj78yetxk7FsNXBQsCAX
1p90EaNpGG6WD0wfhxgbOZG9+xWSWSCY8fekyO2Llxr0OmVBdVP56g/HhBxtHFiR
1vrAu1gDYT4jVmjv75w7Ug8TtCmtGa/GiCyzojdJ0gicFCbFjI92eN8qDP5WA+1D
DIVH+3+0qPxZL0GaXCZki/AXnWUh99I9IOgQxjfPZGGusBot2a6Dq1dJAh3xO3yE
w/OUK4VQnDPfS/iTxZvL9yudTvEUJpzv/Ksoa84nuXK5gfOHy8EAiSm3f2nQk3Fe
Apkv9qsHTpxU7GBKCnO/hiUFSA34y7q81o95XvnGD3/1HTQ2FAWCAHeDKemkb3cf
8rWDkqZcpJuyCLXXHbvG9ZTs/nene2cqg6E40pGTSwGgJGpQKqrfc42AXrGPiTca
00f+2TioE9Bc23r23hyNZsX0EkBvvCZboJQO6lCJeC6dU1/QTab78HePv5tsoGfA
0eqFGwxkOgcnFJRhnEy0NwXyyVe1H4mHXJDrwDW5MdIKvNPpGBu7nrKaqKzOT5Xu
S1cmodgChhNGpl7G0VoM2J80ogqFhtSwnwjkn0LzHCDqqU432fqsi3yObIPUOtiL
xJtvBNAkRgrOKxGQkKNsdZEGJstfbca2HBcPX2R+8DKGSpuQ2Vm7ACvhe00cAXUG
3Gm2xu5FyZqlGSpnMEzTTd0/yStsQ6zLD1urT786njXL1Sni+s+ANWkyNvmE/3Zp
AnZHcAvXs24yl77q0+MGiak89k3wWIzWwZsnzZgxCAN/czEFPP8EdW+pCGrz4lTM
VxxeXC+sEqUme8PNYazIVSahWt36HsoKss8SXS410PWXk18u8kw92GOXk/J2cOMj
gI0asd91q/0uHPM8r5AgO0s2wF6eGIj3eR7aKK8sBtT7cWmXKKtTwca3/TtCYkzB
cac8x3Bgmxc5GVAE3w47xUhy6wGDYVuctFLa4yJLchiiUonhjHQFMuW/KUa1Uj9S
EGwvprqWswpt8T0XDdR/grCegKrMBTyvPyJnGtHVnKYHUJKBbaz3j3iqAO2D4agR
dSxsMyjxw2cDJAJQmQ0gDLoFBokPFBymAn/oRLXhmlxQuNICAkVyJ3EN9Psq+CDw
JcnM8Y+ZcdsNORMmC0DxcNDgB1g4nrzMvA6CzHd0HJuXtOW/FLJ+s9iph9RF0vyN
pjLwiQUdrkvjqIHyKGGpdueHBEGhqMmPycJMzwp2K0FOvBJEPhyltqkWRFJI767J
pg0Shuly9+CUDl3vQuuAa2ri5uCXNVfNxRozV+f0lesNytDNeJnEoWMTmtGC1HAy
scF8GLwv9QaaXd2YDM82wVqiYHlg7x2JYcsjUfrO9Sh2d2TVEGGwnqAdPvGOCzmJ
Yh3F6n+2MRd61wZlL4XdOCsWVo8mSebMj1MZiQH0yltL5hS3MlfyY8xFbhyXj1nf
57H9eaWlxfhZnmGkV2+aZmrXc4n8+hhR2vNfwEO/d+uIQ4fpuVGI3F08luB2S3Zn
PFPHQuvM8erpUsUj5ncWq5cbBqEhl8xZwJO2De0XdDUSfkkXbMXk29oDhYitMzKT
XbNzJwlBiUElsHa11aNqfsW6ADQyNo25LRcIIGA3WAraMIjrce5+/ORHH5vizj6o
PFWdHfN2ynPH5cPaCdZVNJvxY5SrywxqDRV30F0C0xVa6H1iMsZAp9NAZgKWaWuD
20W3IC7fXcx9+fn0mlqDITKFKyzvOEVVYciWyR3qP9Px+XtB14+hK3NQ6DjfhjKC
Jm1SQO3G9hByRSRVvtsvs2gGcxU0fjDQj1hTn+Dc6rx01MquUu64p/1etRbHZLZL
jjxWH06djmsSWGKKvwLDI3EOR005uSXx+fUcm+c40aT5gQ/RaO7ryYyrit3Xpb6x
CKBheobvVGeOPYDgRQ7WO0kFBOu+CTSSOYNWlzGQl8o/BwJh3srhz9cQHkUr5L/6
hxJd2zeCroQvM9Ecamj25WSFvOO9zR9SoKDiF0vWvFRudB3sjh0aSnbsb+Z7PUYp
2GPwi29dSY1iO9ouXwt9yStpI7t+nW3Pog6B3lTuKAv+cNU5BU/pObR9wPrXAEME
kmrWKAACYukPdmiT2GRjc4pMd2K6fyyUX4eqxKX/B/KRDL+D5Lw+VZi7LGSyvWgD
HgdwbDHPhpLUe+HJKMXJqLk/cDy7Bj4s4rDmVzv+YdJtgU3W3b1qMBq3H8vlk21g
D2FdaDgZtl9kcQM4Febjo91P1Gu8aCfn5JUypx1LNhfhpKtisnDAm3RupYOy06Gj
hEdETd6Fna5N1ypM6rFpV7Ak7etuwNUeDA81+l9r8wtQuN+UoNQJWtF2cZ7R+vpB
UXCdMTVqCI1x7rtgInOVo6iqAbmFjgyYoummTIAIjGgOyLA+iIiyVHm5XSh5k7T4
0mH95tt+tPQOZyAu7cjcLSom4JcM+CO0pP9UHF9ySeD9DE8YKSo2lDgM13eJcIIx
dP9gBDXzw2vqaIruyW6HLqGhNNlmdM6pPmD12ZEPlOE7gIYh357H5ABkDQlQ6iIC
SkLj3615DqUp6+DSQpoQQQowb4jhdppxuqnw4xkG+pPG+2B+zXqQIj9+EfLYaF02
MxiK8dsaAQs+Av6Loz9KjDVFRZvVlkhhG+5j8ONvmLeDnR9nVTx9vSBolw+pptOu
sMyJJ88y6RUgUlVl9LC4oKJ/JHGmIALOu2qrY77Qj56wwZGrLpCCYKbBcwNBklCO
Su29Lui7wFz/2p4lT2Yf7kcuWWrNfmbLD3AQOfbn5SUTM5G57h4YHiina/aRKz/Z
DSS5/OQoS6CPZIHc5XHG9WdG0eezTne0YXTLLdQzwcs7fo7rrZiX39Kw+YValOMJ
ucqFuU6VToWGLMumjj5nNYElvEeXaTn8L9cRYVW1dmOFdoC2luCzQiPcBLrBRyBM
4yOwIa/8rrxgWFaqZw0eId7aHBzl1Jq5ZaqlvCW6/8FZVH5XaVcJyYjzHOuj+RHJ
h+LP91zwqyO4D9wd6jG4xlqwLAFvVcxOnSieRh4x/v+CmRyraQhBI190JRva5PtA
4B0akDQg7hsPq3LUtMU+HlggtkJBWJZy+SJ/HDaJajjt7W2bY4ElvV+4kZhwbU7P
VJS9UmoGtp+ntkwaPTukDPNmWSxjxCabdOd5xZAIKsVb7RDpy3DglMDQYeQIM8IA
LptDjUWiAaK9nTtDNtj5Tbq962kdycicfTCGKAkJyT6sOFy4sJCT4+0JDleNRxom
ppIp8XpMl4Nk4vDMm/bVBzKfyo472cKvFRO59sso2mJluZ8GLxZvuAuPWutAkR/o
NonNirnzVnFuPAcyXmepfiJEKj3Cs1/ym/Is5XgEA0mQ7ZU5tXprN//GlrOmmMTn
vMcbbhldGThcv8Su7291eKz9rMiNhuVENbdDBpIPRdS+0ze/IPzZRnA8RRTf+Tyy
3fEbDpmTuA9bKN88BhRK41M3d1ruB4LuZqE17IVDQVEZjYaNQ+8wMDJxcqwNiUeq
BSa9A2TuwGYxWDdfSTgsNwiAf+JFzZsNc0A2LQVIzZzgY2F8qoWDQL839ybr9MCG
+2oG3h0KMofiQdccxI7UiGni66Q3OJtSnqkTLdw0MndfI8AD8FfUMkz+HnYVM5v+
UV56Fu8W/7553PF9XowA6eGr6JpmusWRZ2SaAFkS7Fql37xAVWiWlSI/tgFy/O3p
5uIvB8dbtJbh3dr9gHQEeBexL/UmoSs1E5n9AKEQTFZREro6GjtWzMsg+B3l55aP
gbChMo+Q2Q1mUZ4HqYL67b3sGUoYWv6D/JuAuyHMLOtr5HeZd71Ulz6Apq+7UIi8
D3mi1wyaGamCJ621F5CRBwyFpLZN/MLJlz4atzuTGhyD2Qs2rCQjNJvvAaCwRCkb
IyRbu5vxoFQmzHar08bQXRnjfQXVtD63kB5Z0Xrz8s2oBtnrCkNv57qPER9Q3DYg
Eb7IvHyvPIv3bCHrir0cyX2YZZTu7eLhfxaT0SOnp52u4XgFfgmL1R6YwCPA1yeC
nnAg2R+u+2fYiz8ZVcxZED8yhkD3cN8o33m6uLeVUTqZ1NfSfSCasMqo9j2ybv2k
29Go2qM5/DKdn3R6i3MhymN3fRz/1SPga/8rB3svqQ2moJt2yu2hHHeHPllStyCN
W6PWRs8puJ5PIK/qr96/KaDhgpjEeU8lsJSi0IbfX38irR1G8P3NsIIeQUfk5wxm
I1JrbxzAG3sMH9Qaef5OeG3Q3Z6mJfev3xiJC2XFFYXZuXVnDkuLIDzNHX17m6Ql
mMX8Uao6VmkKigTdBfRbktTwWJsBomakCVns9pd6CEPWLSxTjDTCMNUK7C/f/a7V
NprQzvBq3mCQUcUkmJpdU8N/2a5TRMvhkze+FGEyT4zwdejXQVR7Kem2cU9J/6YT
8xmuvCxK86W3KI2PZdyNsqzyFrMrXEgnDNsQ3PXZp56NvoL6MckvkZunFejR9o1t
19uXuNlYqLvpthS0urGpd9AUBo4XyrE/qaWPIv/qk7IogFXxxx8m80IUsTOCVZpv
efDcOytSHm/MGmoBZVt5Ds6bqtHovax5L8TaYyNq7HNB6le/rpphFxD608/YMEL3
HrP1lu5/Y0iqjBwOlI9WT3R9VEKB64RF8RkSJZiclJx2YYUwzZhEbhh/sOlIHZam
OwJ/FWkXiud+FmSoqXS4NvnZ6hEmhNrelwhQDwL4cIt07+ARF3XBNxemseAA5pQO
wiataRgpFshlXQQaDv+ybvF35V3X99RzjmBwcMbQ5A1pqhwD2rIrR5T8zvT4muw3
qyTNkEIpgQbNDqrQabQ7g+vp2hTr1mxtimH7lfWDYq1PJyuR8DHgwiRYQXtOYIxx
0WMbPpuncaId+0ohOkV0YYESR+KE98vS64/NBhMR418pspAqUqm72qwdCJzQeEOa
owpGP9BtBa2EwZOZzBiYHb4S4A9JDoPiZbZHi9wfbWH2plYMRdE9e4iznGbysql2
fOUE29pp4benfd3UtDbG1JE+Fnq9d1x0zYE1OyYxrmfgNm4IBGZnlFvg1j7rEMsE
5jnp4NNJGsKNxg+VAOTrNkZfUXC9FqWaVTfiBsY72enzHRrdrBwOpH5Cg5K359j9
aO4U6xT2dg8BrtMytUUm1dLHo0liswqDDVnJlkloFJ4OzjNmHo5/vkZxuSYTivFn
YQDVATEb51Pa2ucv66uLtrcHqjkMxC5qbpq2jpFTBISo2HxKprp7j+Z4VgDjQr8L
sevHfTKa0Ft0fNoH51AIK05m+Na4/HgpYLAdYeHESJVI17h5aPG9NHyJ6O0alUDL
OeSLfK3Em5PXADRZVGiGS6KyIPnBbXbXqbgFAwLf1G+G7U2EgE7NGSrjpJja3J/+
Cw4dXXkdMlReHx2dmUYa7BDGtlLerXfX2fmWTevz8okroNyOqozPt/deQtf7c5Wc
snx/A1cwSZ7EBY6EnuCIqYNrPO74c3J/yQdKFVYvRNdW/ejCAoRjY8eLwT4PUONr
k04UW2jTK7H3cp3G39jiIGV9u/ODhPbVPeePJ0Ci2dxV3WrKJvzYGx9Xm7S5Uz7p
GSTr5x4Xg49FMjlfTC+Wzs1YdPg/pDc6vC4kb8jXhhFps9t8Ui3ZADGwqSNE95KH
+CTxHFf1K7QpbTaaqbAx0kzVbZxYUkURwgSf9fU6Xk+xePLf8R2qRjkw4Lg5Uema
yWi3VpoqDHFAoXUJbkFbr199EQrx38wtz/gkpA5+p1L51Ysq4GvhoPkvLXnB0pqy
pxjkb+QDOGwHNAJYAfnnH9aX5lGSu3QPJJZP9lBOGlYe+rtVFw7XA1k+DrfWzwK+
cXzWNR5tNxmy6al2J+0mHWyx7wU8m7SYBrRl8EPzSgQD8/7Ro5nn+wcBdThUCCL7
bOlCr1TvU7cKXhgSFgh0oRsNq927cG85BatTa70GK2e9UZm0ssIwbnTcQLmEGrm/
ubuVMbhIu/bXmuDs1qHIxOa5UUkeAKHSA1zHF9m0MR+0dw7Ou9Bh2xo1JeVNJwp5
ROXc2mFCHjs4UyCvuToeGzbs2PjhlO49B3cstlljquq3xOICO0QyYSa5kDomekwW
XtFZejPQW3WyzlpD9l1/TiJavK/RmwRaKYnEIwMCm9u2Ws4whSh37TkURWnSs+aW
YQJ6DhcMivtYnOtle1HQ0WNg2Mw5kvUbqvn+ToHr1/E+RjqFfGntFgTjSh6D9MQz
sNhrRLmbGOEtnZxcNZwoLvfosMHW+y9xwR+J0o0hVR5kcCDF2U+Yq/KtjaSa+WxQ
FLtcdhS+aF7crXgAFqkTW/60OXghIJbERZHCgk3PG1tHasgHCgaKLTsnRYaNmIKk
XOGymYeZH5wUKm/AIwag1qJ6hTox7rGFSbjiVJDvWLnMgPn7rItgKmpckZwJ805h
zSLBJy9NURfZOFTMPpYbS1PwkTXf/hLpTxwPFLEBjEI1xFObLIJMZrIGnNxUsYHg
QWKT4+jsSzSDjdzuLR3Jz+TXr6lHszSHZx0e4YdFwMBJIoEBlWA8wMJ2/MOzVYi9
wuAXM8wavXSTovl4xAgU58ALGO2gdTW5ckRlX+RkTUgRKLA7r/2170DTp2ioe8aj
pHfwa55whHsbW+rcH+N1K2JSm/ZPiijIvWiQ6pZr611mld+PnOs6DmWF2Pt1pDEA
7kKJnErylMrNHLBMipbxucBnyVTUGJ2xy26NFXCTFc6/RCbRijvWcu9gWWyf3wgP
NAmZtf2jWP3rei9geqm1vNCcmVXEzDUNUA6K1i/Zf/KO9ZA+GxtegzzEr1TZvr28
uEpLsLXs1Y9Qc+3z+EoZCJ+UHWE47a9AVleCDE1yDG1oBjNKf2v7MBjwdN6xXUm+
POYARLfhVNqNuBvh7JGHDpurZMf42QIhGbL/LQFDaD84n08A/CZiNva/5VNEpnPR
n1Bi8hcAlL3s/c+5ubK4z8SIczvHZdD5q9q11p8Mtwdeg5fAPKcOQU2LI/m3p5yf
lefveIRq9s3CLDmRnqXGlerjsAQyL0mUiEOEUgKwFK0GXykO2jQgFOw4kD9gTTsI
lWyIR5dSWJTPoL+q1f5ioIztWRrguR2yUej9I/HVP2ew1sreV0AdsHc9ozlme6wP
MbBJSOJAYEcXLVOYolquPjUaMdRI1Pzv+wL6oJfdZwHluwXxzmW3a3S1wyG9mx4/
Dpvg09OVRIeXKUy9JKR0zAWKpeOpWCgiuST7yFUubq1abzXyFSD6kjPGpMRnuRY6
jtUNCDoFoYMTIfYPJObno7nHDAC1/h2IH73dgl7l0NBzIqUmQUPfMlqVtO7zfpoQ
7424XiPGhn8n5Ll/qvdpBv4iTxBMu9Tyyz5BEI7z7srKYozSA6LTndVsPyPOQl5S
Ube/rZMDul/qqLwXeKWK10zOHZNFQJwhfXCg0RMJD0xRf9Hk/v0D5l1KCSZ5p8Cd
ao+Gm/ODmn6oGO/4MjVs2u/YjMD/2Lxv7rjXAxDd4ECOmvzMwYn9/RRTZ4BmevEG
tv/YhaGOrttieW8EPpxpwuS697smXwcK+cWdq9BOi7fbi+QnPzrLpoAGnq3RBwsK
YL455aD4dqSnkNwGvChcfOAxP0obAo8YJIRYRStQnz4grpQHdLqOPxZk0NPtNp3b
NFV+Dcql+3YnamDnMETiq8jWRNXTDGC4wQ9Fd1nc5vPwvixnMlaFtCwGBDvg/sjI
cSC7CPYegaXyANHMszdkJE1WpZUw3Te8DFUjpw5NmEu/+EDWc9R86tqYAPZoQgKe
za0X/roupWSTqDttSIj7wtwWaKu2UJOfBUEXMjPiS3KlczVuzqLnno38ndJ4k97F
+eUl6B++AmcNeSnuf6FmwfLEsqpRR0ynrISbZSX5xb24wbknJvhIhMKkj+5KpleN
XLv4BLVdYML6ZKBQ98mzkVS6+04530xCmOJLS0e1XUQaeP+FSdT+2XD9Rmwd0QhK
hKjO/6lGZ2KArJFvXBmf9b7FZ8szgDeh8IjbO7JoaG7804X4yr0D7hJB3AZrvVf7
jilV4V387hZ8O9wzkMzu0L3ABwP1aKRfqfCj2xpLnBv8f8+lJAm3CXeYWbpKAK9h
IB7Mlz0qEimIYYsFU03HqNnm4Lrp5z1u5lewXrB9jXT0FbY8Ze3qeVtj9kNc6Pak
OYc+G15EhvK+0BOQCA+LwZtD1vB8ZWn8VfriqYZHairQf/wC0/pHmm3tNSy01Wq/
h3SgUvubuMMNd/0RaTKPxyPYd5y90pMn965g4vOlB4hUd7l5G1OLeZiGuG4VzCAU
SymPrUYJnMAwvIDJvFdCMx1ELEQiB2KjjGwhHYoj6JYhymYNiGZGkgcwSVOwYO82
IwsZ5ZpMwocNZGVlCi+1fvZ1YnJwRXIyW6lAl8dod8gH0GdgM7if85N4owgvmE0q
Wr27zDDhl4jwtqyJI+jnY6WwZg0x+Yb4ahr6jva2RYjhJcaW995M0nUV06M11X1K
rU+zFG4gS625W7wd+f4xvstAqS1fnmDQeDs84KvtyAMxkcO/HRvRjvZ1ODPITVik
FIuCCewRUAFSNj8jBTCaow4ZYNy7jL6YEsTVE2ZNabqnkvsiTLaoj1ojpTkfZO+e
LygsJ/jijDZcjCSmkuzDkOomqMSSH1cqbnlzS3eVZHqpq+Fm1Q4EXCg7PjEhmyfi
ME1f0xs2Fd/c6frmXH4oQemSYWuT2aU4V4cXhR6sfcRbO+AO953o1GRTYwWoA5kL
FovTu9oNhmvMjru5yiggqdxc43tOytPrVlo4rMJ2kRap4py6S94/yR4qWw1sBe97
vTIt1P08l6nymR3XL8o5tmK/igcw7Fn2Sq7p/cznB2gcwPgD7erjR1yxJWSRfQIE
HKJ3/CFzxqVGVcCHtw94SNcCmG+BHd/sSSLkxTpYEsqx/06LJwHi/LcjDUW/hmwb
nv/E5DtRgE+GH4yQawtjj7dAbo7P0Pf8cgQaIvgZ9c34RfOTdV+/Ev5s//cBjjQQ
ssCxBkO2DZ6vqpsdwTCoWe36Xig05TrKIF/k5jPYqO3VlP+QeXV9P86+9ECAAOn+
0ZdCrTHINQsdavg2zdBg+zVgG+9fAHYBRyKU2HRz/qJTcK24HU0OuazfFfdKXckJ
0Yf/VN2UPOwX/qmPah+TN2b4y6tkLNNdB+3E1siszPnN7pj0cg1KZQVM+mKhNJ7b
ve8ZafNOk3HusqNYGkGEB2JXXuC9TMWTjRWLGmTlL8XG8MtgM1zxe5SZ/N05IGZF
I70l2UyA3NnHv1okKFlqNj2N5rRu/h+MXIRI6uHhJWkiUQGGYe07V+MNHajHaG3N
RD2p/Ujsua8mtTweKm5udTqdoNFNmpcZjlBtS9GHJDrnb8khu4tyywxvJOezah+U
BATdCBxtCr3hQV9y3W3frWlnY2uzOLlGeYaG7TtvZ4LsRenC0kGPcOtlFCNQlGD+
GyC8les5izLC7h4Ns4HmQKri9LzrgqivFF/eMynMxiByMG04RTi6Y480hzZnwV64
4Kt+12DwxwUaCqkPrHQXMWm/lGtFn6btk/YSkYZmlEAvsfNJG8p4rWjvSQv6e2S4
2meOIvUrDEoEAUBrbgPgDqzibo+6eggT8dFbBG3vQ3KtD6pw0RbIsVWGOvcJUKbS
mhqSJKCm+TkbYUb6p9/PaU4OQDnPdYEOrPlEiswS70Z0fzPv5P68tZyrrEIBRips
UrtGUJyv0ies5X/VLHTYQeW7aXJcv6PeU/1rEZE2UGNl6bgQGeenxA4TOBnpCtiX
/rgaOOc1TY4r/3f1lER5ROtwsqsjMWfB8fOXNMmfzI8ciixlFvEPMZv2kN++Zc3b
UNmVv1fE6hxQ7+SiWZUsZLVKzLFF/g+gofFDA2oK8z28qCmDdoJy9rwZnaegcB5q
irpsnRc+hs5OVA0B/RdNmxpnSnuTFzyhYnh25NCWl5RrMgC+QcV3TwPL+0qQkZIa
jxNUa0tPfiUJ1B40480Mr7yPXsumJ51PjML/kdZrQ93DJ1hmCmgckWb3hK+AYXga
58Waqd/VClVripoiNSeTRDgJYaOkl6iNyzcUwMcOBTCBEDYTEGzcTsGUWkvLM8jl
F1HK32JoU8z+s6sWcmTBmnLvuSmV1rZBnj1401uJ9jgAVB8YucBpXhhEfY4CnryO
d+8n/oyXW6RWnG82pgqSOdheV7v9vkTmsIG1twJxiuwM0wWDfc7/u7jsLYPe03lO
6jQwsHis9bLmIwK8XO3VMUq2s8o4/DKh52GuWaQov3yoxXLWh7l9gSikOx/jMNrn
06gJTybB/T5wpKICBJaj7UxUX/joGN1NN/mzpZ5kjjIFiOWwYMdzMutgCUwD9tG4
NW9y7q5XON6r0T38LyEWieZA3LMDpxX5ge4ZH84U67cvGvNOYEj8dIPaZR3SeNk1
sXueg4obMAdIpEZFrrFF5LPBISGxlOnXC0LYi3YA/wVe9G2bCSLNuo/ULVHBAXpM
ypvk/QSRWv4KiVj35/hl4rtrlDAm4UL6vB8+E9fIVcLoGa8bwUSzwE/eAdPfhVM7
uFyWZhIwd84Z3O37oz+8x85wtmF3HnxHkemHguLvj7Hd/UVH2pkUQ7WrSITU8ZJG
Qn0oegYmKVFQfKyyN4A4U6taFLotUcZ5GD8IdRocA8qSnnFKyRZAXIqdpLTjXYhi
K5ME+ryZk8v/OyaMPUSuU35D6VYiYI9EpbuVJkC/FQfiHvINsZqTHVThi2EH3TJp
aEDVQgIYowZ5ZkAn0yjzewPgL5cfO5auqrwlu45ynW9GKZg7NiY0Fl4KUvmGdpku
tKEemylVNxaJoN4fSN6AdWOqY8oMc5hvqd52SLRT3X5aI8gCKfbJAZzsPoOQnC4e
5DK/C9S6a7rgeWgy3eCYN8bjSziDIltuawjTHbdnaNgPl9V74kYtMnKMx8xapGQW
cDbddI/ycE9IJErimo/GpPVfNZfDIjJXjEcPio/3StWXDpdKQsVw2Z4IW/kRsllb
vkVbaEidTNHctr6GbrcXVs8NGQbcoFVJgyZgHMb0PVtb/fwDm+LRhpNKtCB82xcy
qomd/25QdvCJKZ6BVCA8vpUdZ5jBrJZkMjhfse8925Gmrujw3N9PkLi/CTe0VAiU
XTH5CqCkyf4ZO9ZTSReVsbaYufpcRDgSCO3n+S9cUHcv2J3yu/zCe7m9+ErpvsJF
VHTG58kkaww4Zb6BKUS1nXoEZvs3M0MESLgxH4WOFyE5XVfcJlmj7ygsNRRC5KiC
AeW2eY79R8BABh4JzUVIhUYYPsdoKG6zR7qA53OFbgc015cgc0owGePJoFWsmDfC
oaHjq/2KP+dYVZkVKh35lKYYZ4JY23dP3ZtoisWHiYnguUlNQtQjtYh6SrcTa6GG
Xg50a/zjDeu/6GwggFdZ8CiIp333rgh7lxPFViDNjcUi+oTyc3HI/RKrefJPnGhK
BoBWCVeqb4H6o2d3DiE/K0Y/wCbkdf9r7fHgfwgiLXn+mVfD9JBM5PPYinjKu8IJ
ix6TPH3kFmY1p9DTQsXxm19m7kCWrd/QAwcb70A4mRHENW2JcQ4D+SgEwkthOkGq
mp8vUGUP5zgi/yPi0bKszzvCA0s3Yxi2U03E9PwRgdDPN5IKwkSwZ0dQouvh4cjS
UuxOvUKIjiSaA6GnbMelFg5Ov0IzhjaSIG/iPt9Egssx/CVpCq2RdvGCaSQMVTjz
jOytimCqmXZtkhDPcIjhLqm1ojVwmeTEwiTqN8EI2Y0ZuY0ti7TQ8cDWv3U+s/dX
mvozqlcPMZ+DKkQa2fdp1V21OSEVeCo3kT0ijeNF44crjuv1uxPGa4YNdNuyweC7
/ScOx9ZaJwf40Pr61zT5zwIOUwddfrnf8stnPP/w/YHgXWfdKJEifubkQazgxbHb
BQ72U4bfvUz+6eolNCPglvlSBQH/1WWIosdhtHIE1IEwU2IgBgMElZPaSYNQ/z1o
P7JXDN3ib0gOVxiAoxBksoSNmlB5Zlek29xxGyLBu0QTBlBJmgQgZWWkKgY6joTX
5cQtEOmpy+WHJ5a6nZVFVbZFoX5EYxaLMXLpbQ1d8Ilv98V8rQb3Tp7KosHw5pZN
H2sWN8EPoSg0/REH3wVwpuemdaUp7QWbSTkxujIE026k+DF4C+tfpuql1+F5a398
g8uUlZ3BoLi76ta2tzgLo1ZMvhfI1yM3PbMuvGNla8iSPaNTymaehRC/BoTuyC9E
wIAohXvxvFGsyTLMuI9rLyq6PGwYvlNgOJm3HdrBu1RZ++XdtUQ7Z+QePbsd2Omq
neWSYDrBcdIaalwA+K9yZD68RwpufmUNWtOJkaOtJqFQglLjVWlstoQuvIH16J+E
tJi3eVSYfAuos4ZlinwTqFwRWNj7BiRbalvu7ni8s55Ek9q4xqo1fDpBXUjBrHVC
78df2SD3G2TFnKkNWCNSq20ygGXE0cSNHPiNUnJuR1GWAbCQb3hQ9px2t7UCSIHz
OBgfhs8M28EoB5m9jwEZmIeyRoyBjo+8YIHXTe800rDkCOPy+iPLggkgbWFguzxK
oh3b7a8PKN5JEZkN80FnUKTCiZa1v1NVTBhdyiizDc226CXGkrlX7sow9QHwXlfO
rLOPCKyeK+C8MP6chV9IX+iuaPZmYJZECCSJLRhL0pNUGqzpnZFnhi/jCgkyvzfn
KLri4Eh5k6S2B9erieh9wy35FvIrZGDItlOg0nNRihLxj9CRkKpeUCu1Gw7jR6k/
a3V0Q8TqlPxLGptJTiyWdX1/7iEFesyRxXX++30iEkdNSozwnX3knWr7oVcdVVpO
lV74nrFAAoAZRLUwS17w2ej2oo7kOn8k5JJR1h+EVXV+xAtQJ9nK+3vmqK9n9Av5
oO501ifFiFnpNe219+8uGxRfP4Beoxjl7eb6N5E01IZFYJq0fU8H+NFZMe+eHdPe
AK9Z1l4SaZrjObDD6mm6IrXjnW7FkqjhLDUjjS3uFbqTnN5NKPD0mKSljF/vRb2N
towmsL0ddQsiJ5EzZpqM4LE0fXCpzTGXvteVQB7Rt2dNnV+KwdlImeUMOXhxfFgq
+Q4IDQrKew3UdNDqlf4wu/01SyTpOFYZPC1oixdQkT+gcmxJfPlMPEIm1FFtcrse
TFgNWw/u2+cMnkRbSDWc5bHAUU9HHTZBwhyVzzxWR2oaGpKHH8I1v/un59byd6dK
wD8hx9hZ+2sewZe00fHJKFQ9LuTKHi8mo8QmtgdzFNiFaGEoph4nyiGh2HRHUIAN
pLCktLAEtDID8Did2Sfms18hFwN7aqrhsqKJb8C/nIRFsBwUlb6NQxxv8jxKy7bO
Y6DakP7CePwrS5+kLTNVmk+ZQH5+h/bxp2gNKuSm08OaTpV0qLwuFWPfQscpCXDy
i3/kQc5XXIYFQjiYD6P9aSCPFTNKPbm0LScyv/aaipFMHkWJOMnQdAlRre97RDkS
x+bCwVKQANPl+N7fMOwyFjGaYKBGiUcnU41IalggmzAV9RCC9Q1GnwqAg2nj3E3b
zEf+E7kAsgrVoi4t93zJKMmt+F1ZnwgBC6YlPrJ4MUGRsPpOKI2Lbyu1SRbHTAWM
8iO8OxyjIFm3/UkJkLpLL928yNOE325WNjk0iptv6QBhX4EZ6f4yhFBjdiwMckgJ
ZIj6gCraZekXtUgEaxyEwpQdH2mXOX6JUDwywOtJC+US2t9L/fjZs2oHlYpQ6Zkl
mr3mC3p7hyguiyBQAD68ew0L/Z83uAnpnAslhW1nRtPomwZcUGIy78rIG9/7ODmx
6O5J5x7q8aJ/C1SeXidmdxgzrzd05vD9ftvpnveezRSM28g6Nh/zCkU97eo8bJvA
G9jjwrJkmH3AR9H4oVAT0E14t0WP326R1MokCsAHD+xfX8kNJ1BrnqYfbIl7UAMb
Cz3eYdFr2aDPcIjbJ5nAjWAYM9PJh8NCNVWBCB23bfjxoVpn5q9PiqUH0jmJBa+L
fTNKyAIzQ5ASjOpsbzf88TG1c0w3+zNIPAVvlQqmnNVt/4aJLxmt1HfgSGsQ05Xa
Ol3YryB4P49w/mVQycOFDeTngVUwH3kQc3Bj0cb0wLlr25CyKKMYWR+d6e38fEXH
NFDkqOa4CijcUUh2xaP5Ia4OTR2qCHj0+VQAC2OztBceeRzo+ReyLRRNgHuzLL6q
zZu6kGE+DE3VCSx0rtUdBQNUBnv3WwPesXfWZIui+yL0HFBB/qNm+2q5Tqwts8xX
Jmsc1On6CItZSorT3ra0ZMiHfmhb+Pe/jDoka7z+xbkuYrakxHtJ7u/5r6o2rhMX
BPXcShGnJkqASJij6X8Ki6JBI+GC4zgKZzgIMSDy2n6cgqsg3E4YwHxO/4al0WDH
2JsYVH2f52HW0penVbZMvQAhQ3j/jV0gvJEXdUP95neRbm4CcvOtJxKBrRBzGaYJ
EFEISAbZQl4BlOz25QI9Fj6GvUteHviGbjBK85Z4RY7eaq0M/7iyz7onybUt0oC7
3fmLF40HPN+srKQaRanej7bwowpGiEy1snTHUju/2lUR8K8c+6AS9xrwJOwRYd04
2G904BQdfmWsNwrBIkcx86wxFMzRR4LxIhKKeCpu4rv2MLUAEmTsvuMK2kZRUgLT
tZVHQjAbgLid1f0pRJJ1UB3n/T2S3KEJC1qJj4/aMY3TuYiCVq2FS8gvyf+9t08a
1U5Uq5dfGlOTH07Tzy3qhRjP1jTIhgr6sazpBUdpwSnfyAZMOqMcrUPsVA3QzRsD
WPmWDnWlt8GXYEwItoh74hKPKG7SyBBgFsgmr7jCDBWEJ5qH0Sjm5UcyIY3s1GvM
NVRooiWDryzVsBnFfoXhE1Ahy9e5p96lOA2ZpD0rF9pgYL5Cdeb3UVyw9hs1mVOl
mTd9HhS0oyvIgP/UOGdxlcBOmMLCw7bWEFiBwUEhjbSg0nKnzwsF+e6T56I8s+BB
9arHzjyrgt/+q+qzTJ6hcCpy5wq6KwneF7fCv2ahhuEZ8afCbeqXFj6LGsZTN2bW
WMW2kgnwfaE7Qtr0WmEXo8AFM5JM6P+vOAhXV90Eo8qHaVbQQ3MOEA+kJBPoEaBl
5vpEEhdV0wA4STijGOI8uEmlugs2yprFptCqwwbk01LxUh2Qm0iHYyTZOZi+oAyB
DiX9BVoyOxPkyGg/wqLOXBe6B+vQuyh2rjnPOFUtXc3u9FWsNzTdIKC8q5HgzcFP
3xwjzoY/fEPfa4ofZ8XAubPy6Ul9FhlcUQb2TFAnF03SKBHxa0hHpNjiDpkHQGy5
+GRuwoUamac9bR0PjzW8kdplgJER2upbBmjL6FQff0kKUiLjCZg601xn9YAtrE8l
m7w4JjhZ1GXVqCwao33lxWS5uGpABaDRuCNEm9idR3PMkaAkJVzvN/yQnFKSyXTj
ZaWTYayzRp+uZpfm7dZ7vkHHG3zBqQd1HZ+aaY4YKWkFJP+lC2pp7xgNxTypENwe
QdKKcPIx6QNTHnRJo1q9b7MOI4qUpQf5kV/Za94uPMJdLtDzwVVAIRUAYeTCcSlM
lfnhMCef3X+r6hnj7QQj7b2RFpWclg8waIG6zTMNXDZGoufPdQlVz+t+FCheQZ6D
uzP3CzweibsZqp/9gBHCQYB4aVP77B7Qx+MvATbk/naW5MAd9/sVopDoexq1fzRp
cXZEcvVeLbgn0R4fD35RATFf4+rV0nsWk+i8gILG3PhnElqHcT9vmWy1dr6yltE4
joTtA/sHga+SJ2adum+9H+wRpAG7VsP1aohRb/YPVBR0sfyEEOwrSPmTpNXZLX01
bB5qrzai2ahuWSLT1qjtyKz/NJH7jV5YmbrsJqCH8uB1SSsSpqYA12SLsJTrgOI6
r0DypLo6nllAwkSt3/qFq/mZxfivvnRPE4vz0u8vkNE84p4gMgm/1gA1LAZlb09d
13EHhLPbGeGInKmhCOJeVrj2iT5aR+F1pJXD/G+Sv0PmwnfA7uHCOGzslWsEPdg/
7+IzqLPb+gMKdsHc24pXL+WJF+sUQBFudQj5+5RJ6zu1pAfOhn/ktjIYMYJV+Kow
Kpr60+wUqzvECHSUXSIav9VgglUIJYVwHBPI1XQ/mxNR9SLFrDkOPH19k2P39mtp
HdS8BMoHjgcKON6HQYHn3301dRzXGJLKjUl/JUYNRFQleMQMwk/xb349kpeuAChH
ogQXii+t7Z2zM6DxPww525DV7vG+yAopFn7HJn/CNXTwaI+6ev9xN8A9pjC+ph96
ODnM5TvLTTb1bHheDcD5t8wzLAfbBLUYfvWTk90SsEABel66seAMnASBsBdeAeDW
GOAI6eWO1qau8uzOaZIlmVJGUHrH3pzEh60PrqW0xtd8+Jc/McO7J0LTrijFl02C
CE6cznCYTybw654mY1HM+6IZ2MoIEVhDIOgC1rKTHp4p+ZuI0lADBrj+suIuIe4M
yz1KeXm6uYlDAyELJd5tBOuwCPHeCTgidJM1Fio0pdTulX05rjm9SDIYbrZFh4yD
8D32d+BVOhOIf88/U1ZmNCg0lZT3kk0ahMI/USiLjBQAIJMjeu+G5kxiOfgFGdrN
zbzDhYzXrPjFRzy6UaB+MF4xZ3cF/QeGoUHYrwLIllXDwxohWhARd1kmCdY8gQPR
073s4vvNkAmTuKo9V/qyyNqjN+iGDiXYMyP9+8uXQRCjO2bNHeRdcgC4I8Jk1elu
VlRbPhTsCTlO58fuGRTqecL+lWuOWV3hrXwt5oV66X5uzzH7rFgNsnztnpP2ShCA
kaqrbyJ+9Y3i35YRfQoo1X2a751mGPDTJwYJVU3GpoR+Iapo6PIP0haO7THe3YNp
u+SK13WTKkMulAqqyXW2gd21B4K4qbrw3kPGj+g3WdGw6+TEDadGMrIgx5ncEwWy
Tl9HNtoOhoN+bKYPbaXgolKGnBQIZJCEQOyAQ3WuKQKJM8ovIPqh9pjcNFKs9PP2
elqP2SyEJE363jA7Nqwe6x9Mm/0E42M3aWeUkNHkoNXqcXmARZkOtVSFghwIi9nU
FdDkmwIRfYkO5VWjpojfFOh+4GKnGfwKGjMM6pH2JccUp1ZShXEOcs9mjaa9UVMR
KFkatB/yROSDLRLjLty0Ya/Kt5vraUaiasSBMSNjRX+XSHquNEOXkWd4U7PDT5FM
bqGQMqfSMN7IU89I733KPyTlNkhREpCSoI8s/P8y46CdX1zi8+VWBJ+UerjUJT9Q
ls2z7hHJe1s56N113f6cYiMx8sUr+TPQJ9ObyAOkn4YTk1zREx2jgq7V3MJ5CoXY
h2CQRvizwMtRovgXizs+1cpy+eVZOiGUksCT4z984L+sLnNbE74MGV5eGxe1b4pQ
mCMU1H31BcsqD6hB9A40iMaKyBwwHvJw+6e8DxmTiS3sdKHndV2xI6v8fPVLp1E9
a4lel+i+XNLLNqKLg32yWfpkjpZ4h0MnVaTKTs0M7WP6qm1nq8akZ604aygqUA/9
JEslMftfV1qjnjOxg/mH4dKeiX26zZSzpW4MLwVYSNB+tnq2itK5G3HA1T29OVbc
a/zKRbOGOSrpJlg2XOHGBKGrqf8aEIBHDOtYL6QpubjiwB8AD1ORcW6ZFBHDGBeh
IYYIrWllguOvvzbgIEGXcojQEvYZSkEkvZkGmly4Fo3HVV8FVs4bkgv8a1P51fCx
uKCL2m75zK565soXtBRcG77LpoHnmklFs045w8ue+/yW+VghTEAC0E3e2LAKX19b
vYliRDKqTy1CEiiIJ6FUk6xlwx/2QJV2zocl6Rj432yPfzmuuHqGrT3zjQqefVcT
Y/v/9NfCfDs7kJK/JxSFJ3OsJ54lx5k0w/Guk1DZ3/dAQ55wxxX8JDla5klzkeoG
PQjOnGa++UblXf7x9hNtFrN3hkT7ggkoPfrJ3V1yyrdEPtTgGocyTQ2UNLpLq8ti
VF+opYzNjDYqoI9SfljxmZxBbUVW+o2H9eQvOItLBGoCHJ+NOQ4NGKyFrAE4M64z
MTh3kp4IBNiZbT/nsCAZW9I62zo//m+4LeteHzkTGbzgZjqmBOTOZBxCVGkaOCgx
51tqKeRqZkWktGmKehPnCFJi8NQHhNmFjHmpABiM6iQLMSQqX5BgSJWNFKwSNFSL
l9n5h8DiCWVOHrn++3dgfFWvNGO0yUm0uyBke1tDntM+kNd+vICKxTXgKr0rSNyN
TvVZgPyt5pQ0jtxE+iJCEISEI9dT3MgzpEg4KKQoUr2Tm+3p5xP6TKVLtwMVulmR
PwHkv3SU82qimVIiYjh4JZlFUEZ04aVUJKtyxqDtVMoFIN6yFgBJ5ZxHtY1Ohn9A
EUwafNMeMib1KK+ilx7bfhem+Ladv69Xej+mq5F7JmVZQlDgyCIf9slMq0SqIIa3
mdhVx7LhTyoOU6neeqeOv2pSf2+Tw148nnNfTSNWe40WC8YQyyNdGQly30RHYMwS
VB/7mbCJeRvj1n7M8hgibIdCjQJeoOrmHHUNlMyJ8Zio+8zEzSNFo2DHo2/Aqmsr
S1mvm10NaFbLN0aleNw1n8JTGeE+Yf/P/Ek82hV3CNlsozt73kHx19JT8Fm3bPLU
UIJ3WfAHSAyhxSndi5GMHOinhKq2KOLaOuYJRhFm0wshJD1foiiGx7eWkCOxZn+C
RDFbAohJJQYY+WIyj/M/FnnFirk6DWHZFo+pFP5oELOKdEksaJTVfIFYcy3MMBb6
iofz9jNY9jlZ/vcF8Jts7tUOkPqv4ydqoNPKo0ZFzym+ukovhNLfrMo6rIAyRRSy
nn3czRleQoGwOOKbiYuJpai7i60b9H47x6Fpyp4fJ8PH12+0dmyBTDptAtWNX99a
VNzSCkirHe3ZnTMmLO+mV+tVd1nC8YRqYPvB9skIyPeRPgxNcYZnT1pzNvM+86lP
Wx+WSsnsXsTXi/ljmGTKB946j00fWEafEzMA0rOmsql2G+/yv4RBdImsjsFdnN/N
E+Pv2hciPOnXSFzOuywZyJxTeAF1jpXJHgpysX+0p7N8GCOgz/4XHZQ1QhVEpMDT
Rddx0WVO4cuWaJNtyYNlLG+Ju7HIvFOyxymt6GmNFIZVlP9AoBsVKH00oGs3ZRog
M6GKzmpQI8/f19cr9T4NQO45XcTdUmE30M3LH5VsFsQ9dOu2gQWs+pgsuMv5RSZ3
QlHk82vX9nkPu+zjGq5bMBGIAslOiChXYJPGmsB3he+iWFb94QZPkNuRTcWk9fms
JyvAgSWzJyQvRJrq2y5bak0DDmbrQdoeh8Ppoq3yCi4FT8MPayigQ5fKQfl0Xuce
mfKo6OUESoB0PVEeUIa1il1WdG7+d/UmS0bqhjTI9vLioYs+ZJ+2i4UKRxDf5KfL
c29ZaR0KNjVJ+dOSz0erilTfE5G0CboDNBTOhYf2jI8pWv2HGLS6mBuPZBfbEHbo
isgw+rizyjOcmznpNCWz5g/l2ZpAh3WMW4AJotRbFtxb/gjaiFINoDPjmfenIMiv
d4XHi89s3Nr6PxWAOLk50+/5NtMIr/GzMaC8VboktBxHYx3UanyAYUlKAXn3o8YS
Cz4nfgS1yoDYnJrHPqdaKDZLZCbjqCeJUSpbUEuLH4GsIRxVwH2bMkKOg6Yd+uLV
RU7FsnhxO9uAnD+gcZNXG9HSRY5QBGYYzjc1+wu43yhyORqkWlU3EoZxo3uBkHHC
ORcGZmVGSpS9LnfaS7Fd3SrdIfm1ntEXZ8LerifV6ot2g3U7wTTLm4eGKAmMiJMC
lr+lCs79HAyktrFwpZF6PQk9wUieSdCWyaXys/a5cb0q5l8SPSpowOZJZHnpoy99
+Ef662PwO7oDyKvnimEeNVH35xbrZqd2D9AwZlqWAp2pCTORml7sDdtBZ+8JgoWS
YKTgpxPTkETdy/P5OVdNoV4BUMSuRljh/JDLuC/cE1yXc4xXocbS+84M52lAnFW0
E/i/pbUgMx2bDRkDmulzR8CVyXeR0rLYjWOTRuL8s4kiymj3Rc4Fn+94UhMVeYbs
KQkr59AWAVrAEG2Q71VxF8kBJz3es/b37UEDVR0AieozfShgAgA9uKG+QgpFWsZe
mV5g15pp6SCGMZvIHeQxTq26dLyZ5fbl2L0XQW5TKU/rm338sQv5ACQHWi3rxNwk
LAh8xB7uZFhnaT2hWbedqD9Fi5ZGsr0i7VnK50ODV941SHaKCi3rkPY0/pYFKYdS
JJHaCTU6wnbqlPRFoSJ+D1s511BIyWyIxL9o1dIx2mAAeSgoupNx56W20BUehigD
ahAKHu6hTdcMrCbVBaFg6NlVzXP/ZMoVcGQXyGNriLYPlHWSZKwxbLWqNm+pJN+z
S3UZWhnRKEpfwEtI+wzLOIA/pQGiV7+v5fZH4iEN/ElJCawGjBROL2GfAojpMg4S
2Vlw0zWNO8725MYl7LECXi+pekaShGBnT5Mfo2ebcOb7s/2KseYHOm3iHx7/ShoV
Zag9ZrNZOJzKNjL9hrIgm056Nc1Uahn8S8jJo5QqjBWbtckU5ENOuAnf6R/+w5le
UYIHO0DZlQlAsyX8y9mYy3YGtWsFaUgasRKVOvkFvD0ndqZq4IdvMhsOwyHH9P5G
9a8gLFG+aBGgK9YO6Y5CNJSH4by2QTSdpz4MxV091uqpwzJe8gyQJYRPpyP9oe38
JwzQbWGW1jGtYTXuTi13jSIoNpM9bzhg+E4ZahOSdmGQaM8OCedE5PIyXngTGfNe
JD+WYQOhtwI6TI8a3NIK5isDF5bG/reZntr7muUhbsFRhZEN5EiTYDv8dsZrdGpe
BlkiXGaQIQXqIdb97L+CGkTNQIfEW/bWVuHFXKqB5DyQQaLV8fplPH7dolsmwd0J
AZNJZVya4CvHZuzlS1AwPGyU2OMNpqxV1AHCpK8z54TGY62VZ7m4pyRQDY8A8zPO
Y3RDaZPLcmLoMjHns7xuYUhwsOCTuPMW3hN6gjLR0Uvr+0x8TD1F4r8K1bSeYtUD
yYzR07MPSXFXwag0sZf6k9VihE6g4XACkcOVVNC3s+hY5I6pCWgtj/sOnAhn7Hcy
Hgk6Km5wgjJF2plmSluy9wlRQVYjrz7jVqblWto7xvm19d7KkXorc7KOcFKstcH7
ibgWXM7YxiIbSplHzUnAMgS/C72x0C07fNNvgSBY2rPD3xqceW/3vq0vapDfSJCR
dQsgd6WVctBT9exvByiMxYivetjaFLL3qMcq6iSaOzKr+C6xVBKhzV/6CGYGwfCt
dXpytEkZyMYLvvemqOyBlMrF0+OVDrkQrPDNVYuvjqTNl7lnJbApgFds2tmXFq8F
XZ+99+Y4bNCkq0FWxh8ArAElPV/EHK51XUBX0MO9YxwoRrAyjpZoGi2Jw1e+Mawz
qPKYbBdqqjyrL+ed2uRRKwyohb89ltqqe72MoyVNc+vuxlEu459sBLaNAVLLu2n1
dGXTyiCDXuw8yO5RJMYBKkYH5SJcziitomFtOGbggwVGNXWIyfnNw1gxKX6GZ8DC
q+or9byanLlWdGCKapkxoojOS63oF1Of3CEaVBBaw5KEb9sZz7ZeLKFlRQBBcX+z
UrhIjdMY0fg2v6BsQL+vXjG0s7WaZx5GepEnytzpVAHwnFi6KEfwe0On55fhBuH5
7wWk++P7RBJA2UBKLuggPA+n5JFsnv78BQdyV7ObjaTOCtiL2v1BHvRkMGtypUe/
ygVWFRrYOGXurEs1rsQO8urWI0fRQKNuJnWZZ7h1PTRU0MOY32ELpsZ6bJTTiN9t
oENOA++6JkKxva6FElsudO1zJlJG9U+odxtVpPkkEjEhq1PH201ZoulCgD3h1n5T
M3ngWVsKfq3QFrEnyvkDsNRmCquu28zcDNKyMRRcqlGAFEufH3wvEjdLo6HiVcoz
Wi5BbIXZFXIcWcAU+qexRIpoVZg8oWeI6KsgabNWKhspAK1panI8W8YtMhHbSRjy
sMbccqi/Rd86qiBjHGshqb3Ud2ZQFE80buUnzAL0Z5yArWd/VTM+mMq5i0MU7WTy
K6mXhbPM9Kqsu2N9tDFfOmPGuSNuZ5tNsJj6keKvE/30OT6oDbVkDLnApvJPrTSm
99Xv7MvbvwhKu6GJ5r0vRaLkhzXORZkHzA+MT08P1uYSICLdbMr/WOPlA8FMv00u
HxavkgG33SFL8+EeFSmPY9fPCx+w4ftMC+qAEYqYGM7V/mP6g9IFup2kR+ScuEq7
YLtJWKfMpq7WCwLB24gFBaWuaY3XFHQO3Ssx8XSxNgg9LR5+69qtrlDa403+4JUc
ZCYTpdeadLDnOkvWzrf6YxWsWbfF92zF8T9k4ukiu9cCN4kzwpSzZ+JFn5yOJq7h
8b4WHjDJOBpFfyTxuKpZYjEg8jNaZirtXR2+v6eLdastVWmhxyuEl9dtnjiK7qYn
BQ6rW+xcDggYRP+RJw/SR9g1E4jcKbfhxsSURvGq/EmloVVs59odcFr8bYbwDCor
TePjqaAlOVsgXnIMhCqOvQFK8Num7ptjse1278hoqhDdTEk2OHD/e62NzSIXsao3
3YdrXGkYYTBpVOdcwaEaMtmi6cNdO8e0EP03ISt9BufueZVaH/blvQ5Z7zzXIKdF
NSfH505z6PslQbn0lOE6H0lkfKFD3b7NSwYZ1fa8855RQtetba9wyTanfVwoiePB
INMY0t93P/lmEZYg5NNbn5ise5JLhEl8jA8SDATwbMPPKOHLZYSmT3v01ZUX3ydw
bCH6bXWuGWN6TRq+CfW4EBriF/wtQ5aG8TLCdEAbSkcz4WDnOgSxw4j+Fl/iBi/n
ybncF9uToNzVG2frbB7SmC1DscGqzcYs+f+PYyT+Zrkt++hnaUSEsoiW+kxxGrxs
Af0JQ/OOEfmc8MbvagKUtiz+OrobOfwf3NIEqTSYD7zym1QnvyC1TYFf06inZBUo
NEQtu/m0L5tiOzU2OaSH5f7eZmPchrIHLvJT+qe8OLOJg9iqISLcG2g9SGp0R63J
Oe8AzGpa28tmq405yipbgSsNJqt4UrDixi/3BVszDm7pLb5S8n59huDVZw44EGeY
vxhKgzD9jxDF14WjXQpl0mvmAhtNw6wg1OTOeOcjg2CJWaVXUvHxldSTNd+upqdC
1OSxBbT/Ss/5cEBp8ghdoVe5eNGi2t5sRIAVL4xtMSyU3I3nhW4gNAX1nTnYyEM2
9Es39SEvwn/k4vC5ZLFF2UL8tR52jTJTa+D0xcZXe5R6QM4PSy1DUuwrgZgoyWWL
Zt8GXQAhGy9EoB3ufr0IQcPaTwxWO3djozzdKep37pOuXo/3QamMRnYtJbdSOISU
/3D/KbJozrQ2pMc2/2DBUoF0YJWBPlJ5lNEwSnxcXrZUslgAZ2Ahn2gTSJ8a77u7
Vsamiq2h0U+oV+68BZYjwiZtqTT0LKoMpaqB6xKIMoopP0K7i8yIT3j0dGDpfo+y
JlQJ4ZgCF3aCRXkeTjw2kfbe3nVxuUomS2pHrVoZ0dg7/8QNo0/PAqGvTLcqerEm
Ok4gmMzlj0pPBLMU/ceOjBu3xeuQ0CRi+44xacWRffRMJX6WGckNU7IVsMAwO2FH
DB2hFhwfrJsozkRvLIasOWy1eSMeFnLVoql7EQJjvNNmm4hwpr0t4w5mykP1xdmX
ui1Hketzj0YgNbb8xQRNDnRrj8Ipg330tIS2FK4r4ruZVmUyAPxuZYnnmzRuPKoc
a4HXemJoQMgVvRWyXR/f4cIxUEgFohGCtvTSUh2kejbEvNumDgbmo5C9Dv/FA6Lv
E00/u2Jgr33ze0Zu5Ms7LsNDoLOR5YFL5yMPaiINYbZ2rWrEkhxeywK7erp9Gzni
IVndTBBTNNq77WGtVcwr6D6z2htRDA6qeRhpK9ZTX3zMsMl7p5FiDS1ttngnoD+Q
j2zps5DZl8dufqY/J7YhXEQKQcgscML7O4tkIz8MUrOJNKIvZ2rmfaciWhuop1pR
61LI7p+6o0hpqxcqSLj3t0DnKgZqa/nlSx6FrzhOvI+UMM2VbF6e3W0vHfWnrd6F
KoqK79nei0zuDewAFPH054AabJZi0I7+h519V37pQAiLfeex4yATXMayMKPiu6kQ
cPf4Ecpk1ouonm5exSV0Rzn7P29DbIXw+rPeGGhufgIWk51yvTL7vb1Y6StN0UEC
beMP6qaI2+h9RCidLxab7zhF9hRvpnYpDqD0d9pcsQyoB7fszbxRenNJqN78MWfK
k1TjISA3EmsYH3Udbh1tCCWX3Kkwu+UtqxXTnGgDdh+PCsVzD2fQ22XyBfvXCgVz
L83GWSqKn5hvsuNPH1I1wNP8cscLX+Sk5dnUj+lxuO00HaGCIl9WEbow9xGzBFpo
I0Ae8WqlZPw9JYUVKiuz9q3hjzDFOz0bi4mMaohjQ4nBkuUE40aw2DdL4pMJLpvk
ak7b5JahtASw5m1uWpSG7dGHR2LKp8q/AJTcWS5p38FKSSn6FHMKnJSnJ4Zatx0A
c5bAClcw8hnmUbXOB+5FK8AXE/2BBXLuTGVHCFKUP/14ZNYcxLk+PMTPBgP440Qr
mMTrE7z9Fw8hgR3GguOwKtti8ns6DnhBinY2Bz9Lf7N6HMomFEMJ/IO6Uzt1/tUK
k5s3G4aJ9W5AuS2DRuzklnEwbIfxqyq67BqAFn6Ywe2IE+ZL0J+hi5KB1HZCv/ZM
nDRLz5K4Hmg7kE6yUa/Y7Xh9nGuT0blDugNFFz4O/hMi3B5zIMgN+xl7nxn4r2IM
QMr9w93AmkcCQCX5k2lmYgC1oLpTvsEPU+Bo+9HVrM45fNC1qRyL5VCmgGuNBCSA
r/LTSmv0qY/d0rLw5o64dwmOwa/XJksBwbUsENoGvVgFVTtzpN2OUGu/j0fn7H10
d936PCy9H/WrYMurkDC1+pgluagiEVbJC5TsmsO7X/kmf5M3xFH7TWVdfiGYC5MS
H3kv4jHDRCH7+iYEoCp8i7uBXf920LDVQFf2EE/9+83Lve2xTJ6Vy8dHgHhHXipR
nSeuI+ldeNahLdi1Z8NmZNwjXjVGMS7oQAxtPvQ5xTqmyoSfii2A60l4w5MfZ+pw
NlWHuXANgxuffsOcxMhOEIMm6+jYokYsKSWMx6u5fOVrzQjWI6tl4CCmMwRt7MFD
mQbcO8X+7Jg+f3UcaXapvkVQjb5sjyQk1o/HcZz7pTH27HY0VilZ5CcS+CskV8GJ
gyUVFaIyv88LZILlWv9P13VtLKpjTjcosDntU/eY30zybCepsjpUYJ3wHUBFV5U3
RFbFxZ/FNEbYLLekDuWYW5M3iReEXxj/riNUxu366Wezagw65cRCLxU4u/CCMT4I
H/6BsaC8VUq2rsE6afzlIJ74/iRXvpj1PKte7sFHPGRmthDOQx5+Y1jY73oSD3sX
pIAEwbCFuB00oh8W6UMTO6VpYKC/r4TkuHipVK4/NytqY0uRC+LQxoz+DYM9VF6q
sB6YmMKsUq4b/2fT50NzEIzwnRObxeP0KV1qPqva/PcxjKXWIPbGP05aET/ARw07
aK7BnrYiWsvCpYA13Z0Eq6Z51xzik8vUa239gDuOsdv/ZY6YBNKSSAa1WEtJlvx1
9vvsKgYVOJpzvGCxpszbYpf9z3NN84zyLFbivJOUM+c3kbyvLRAS8EqVDFfshDC+
BkQEgZK//90bB2v7O9sQNGsLGEe4dtMRoEcjLVDQ3SpypFAxEg5zETblKNH6N4qX
4QC9NZ/XRXb8Dof1eGFV00Yr/NufY/Y5FYzW0IlT/54k+HnklihGDsPdpaPjoaYX
PE//VlNy5e3bopURUzmsTIVNEDcRIFAGByhu8LOUoTuof+YoY0OAuyvZKBCRiATc
mf7NURriJoiAbMyVFLd9NGPw9DYvzaGrwd0lJ7esfbkKc1Vtr+zt3X79oHs8+xH6
LvARuCus+EO0OKeS+zVlaakSXQfgVYvjYsZEQnMZ2k8T/2ul38HmPwlSdoJX1D3P
gKEIrWPw5BTo5hv/skDKMB/vmp6vQ683rXhgAMxOoqa5VRXIx/trwS5QSSw6VJ7Y
cvqeVC0jAappRFzSSkf7i18p/GeZNC8IRTB3do3QHpvu49lnKWT9Rc6X9Op9HjLM
M7wHac31yNl0IFey44J9HU9t+DqiBB+laTEMeSKwVzvdIirTnJpYzmcEp2fDbyxM
4Xo5q7Tk6ZM5iPbiI+2pHLz5D3+Mhu7o62fupkUvc+kbeVVlKwpHqYy772PlBSaN
N/WnQsXVovbWE20SkbXnEPp2nwNo6A/v7nh52HlQmVWDfbTrNJXpgZTEC43Fxskk
lb7Ee8wVp06hBbV3eq6QgMy/7Qol0ghRBILpIyty8/tE00jzrKxVBvS7XdRSthwZ
X5XgVzuWJG92nheRdgLMqPtaSNnOJak4piELsRziany05OyNE8syw9s/oXgqfK5Y
nh9xFKZx1VrgDOQ9uHdwaPmQMZJZBhhvv3gh76LwEX6coVOe8dO0uBYw3ysMcoJI
t9kmxsLKi6HbGDPpioi2xR+7akDfbaU0IK4SuDzO5qeESzxA9fJXVCrmcoVLwdJQ
s7kqcsyWx1gb4OmgvdAy9mF3SfYfrVJceN2G25Y6gN+ZDC6yauQqfS3yQsFUYgL8
oTWKyMrxp+WrliyqSdUR9JG/0012XeADzSbuT9SeK+qdUrPMrCxbY/I8kxfo4MjW
`pragma protect end_protected
