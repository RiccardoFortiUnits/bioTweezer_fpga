`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JTJdT031TIpQLIVDZ380ajULyesY+E+18UmqvWYwiQNb1lfooFYmTesbR+LC7IYn
i9rL/g2QbqGe812gCL00QA9wW2DRaB1g84qwGGVaI5GyQV7aqi7cd2odJEEODr17
gA/swGZn7rMwdHVEa0o7jFfjv2Ooity4FyYcItolAaY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1760)
4MAeu8BtWA0nM3GCYAVg1utZVa/dpE5s+A42aiPCDFY0dXnkBnOBPlA9GYt2Bg4k
/xkggRh64UV/9F2QgVrcLtWkrY/pnRU1kzcOvf35yU7rWQf1o8kPKwjeU6KciISY
1LbIWkv520LNPJ11z+tuf6irCIJ5Z3CeKq6DwKwLf7x7rZ2QtS06jeztQyrWe0eV
TmKb0uHdyF2cuKkY4tosOtdUi9FK+DPLJ6Kj+nwglIFuG6fH8SQsOaZj8C8jDqCT
r7pGtCHNGBrANNbGlfPABl7hDfJ3yvYJZ6rLTOSvksWV8RI7u+sAobOtfJ73S8DZ
ygmjuj7UjJMmdL8RWhTO+DO21odP7qeLc8KLVJkN9oyOW8BvnXc9jJNFC7N7WArW
4Ok8AG/DFH3ioH+S/81hC47IMWvlGUp1w3c11beRHa9RAEGqu6zOJP8zJ6himATT
El3gfnOZYaT9haq3mBEenaABqpTo12cBRM7FMZAf6/XTPNzfbsrvesNMuHERfghs
yvEcKYfUvKVb85TDgHMvuH1EznBm9WgKwyzFCLq4wtmqbXqFSqBHnjNJm/AGyBp9
/9gvUdJTUkQqbG9NstB6GV2D3+TSPjoc1zs1vxqzBJ25Wz2eiu9OuFhxIldt0vgQ
m3GQs+uMZwW/oMZuBVXsq6Cx3LpIKmbH9LTy8YEjYor9GNLMDr1ovf1hirfVYlp1
mTW0SOWAtgtkxjwzmimsBLcIA4SYVX3XzEJGSHzmZaDMV4Fpp+/yC3LoG2/yVjpH
7AulYgR009+Yo2DYizxV2fkychc+0mecogkTKwfaaw0K9MXvhOeYP60qbQCX/u/X
eJvDzZWz2fQDaRWl179vMVGpYGWj03pr50TaYD4PDM+0/zC2mwcTsfoeDwCHGg/J
/OTGYl2n2HfjcX6+OcDSHllcvKuEXs7SUfmd9UtapQTD7hSZEAh/0WjmQIlHyAVr
a7JS2X0Nwq7jf6tHkakpyofp0aFmTa8wy2uTqF7dac7bEm2YJQFoSaoTQb9CFJDT
6Idmg0uKagnnETt7TIAmmvIIF+4csxApkya4umuYIiNyx7qQRFykXSrwG+/pyXuJ
XiODazNqU43A4Gvwu8AkHUEb+XeLxctsEkGQ0Er9S+7zzDb9NGCn/Jjxyakv+IAr
vxyz3lzKqKWErOVDPWxtmMnsp0b8KtssfC8KGG9y1k1bXg60l4q9s4kUDJ5v158U
k7awSWjwrWtEyHibATAv6eo2Rh2ZUOasaN33G83J4sY+yEbTfiUDUxGlkVfJEbxz
dpJCc9CT4ieAK515iAxoMG67FvbaWyizwvZNz0MtemDWwg4AjmHuHCWGzOkQrVAM
KiKKOMYDfLuhI8080EzQfqnQNjv465MA2boBGKDT8obNxHpd7sg08YHjznp/D+rH
qFEuCrYrPDd66BN/W4o+p/9Lx3LrVc0rM711N+sE/cvXV+Ku8WjXwZuFMpOKgVJC
PonpwyOY2KRznj2IHGby4XCWZ69Q7WoiKi8dzmFXXUPKNGGRy0QSD8MXzCAywQQu
IoQsHqiigwrdq2tRTixpTVFdxEXeEHvW6f+1+mdG8qo7Uzd4rlHaMGWJMsDax8hR
uBYKFBvOmuFSIEkGGDejFPmybtDnL56zR1mMoievl66DlQBhBocrUQPiR10cqVHy
wTcUZebcsUuGq8bD6+3gga6THYNrTjbbk9Noq254+yY8WDtz3MuTD2XBeYR6Fg35
Ns51fL2pdjqeghHpzOIVHXKocfkUptnQLqq65nA1jPMizUlC4XK4DstUKs1eR/8e
0Um4ykFrpN5xSkVOeXxaWeHTt3RNgWPWUgyXhFc9iOCNh0dshKSqd5gbcNqOv7eW
EYso5MXgGLALbErhAzjDlezEK3u6hIJWWl2ZalxyPdLjUVaPnoZCY//PhP7X/VLP
h3wsS2zp2ucs23omzTUhV7LXE1NrkSvD/tkWPBE1nyzDNa+UAZIwFXOgm0ivRvAg
XGxWQgfxFSqKU5BSuxivTc0Ip4X4wrNMNeR0UWvYs5W10qfpA817xfTSwGjr2xcz
7ecDiB4/BKCmwIveDIhPWZt1ya5TmnaA1xbvozFITsOFM6yhRkdM8RdSNBQILmY+
L35Nx0P8dmPzLfjmNmzPz2UzsPqwnYug5NopF8gYUXMKQDsIA3Zvh2jifW+8cV6F
OMOX4WEQQkxCru91DHZJ9GPefT3nxHqbBLp6riHWDO2s14bhOfvEbmRwoXfiKxYX
sqXqNcsHcVidCzAkFVw7SW7RHEknPy/jmyFG0GknOajfKZL6ReM4YSnAMzmKMZ9c
oK583vt9HCPdMR/HqXA4qKRoUbqVRkeVq91Cnr8550Q=
`pragma protect end_protected
