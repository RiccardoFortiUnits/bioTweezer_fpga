`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RV21cy/bC/Qf0yLDezjJyUWHL1FcAog2DTUcu4/UaLsIAXLigi8fP1EdXl1p7/wb
EW/uLUH8ayN5qGxbq80JOGrXa9ob+u+YA09KOiHHjjR862x+N3OTytjtZGTHYy+A
GplQxkgngK2B+WBaKsc8/Bnf2zECyaQDjhFT/sYiY6o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
/bm7Dm9EzKCCClPwvQq/VNGNNSFeCgfYEa0mOg/aElhiiQMU5nwM4Zj5JycQHb/R
EUf5jsXU46VdofR+53A7swc8fOxj5vv5Mo/U8pI/aFZ9LhL7e4n3UsiS5OrnMiNf
cTGY1qiWBhN8g7P4CNxvFMIhtvv6dn1ZfnE7+4p8fpa7SVJmkQSX1f/0eBdhnvdx
NDYdCtKaaKGb6xXMyHh56jUGhGxcW+Wq4OG5S3SJaSJL3uF2dl3mEqasSM/SMLX+
Ae6X5DOXkSzkeCJErGOnMGvOxFmtlWqaxbCY8to3Ec5+utzuB5ECcsQD53/VmWVO
9OYiovBEts+QtdRUxPSKPYOd3+Ff5qfOU3xs5DDIIxZ6ICVgYi+T01waKmDqkmYI
ruHXC3TJ1VG+b6KIbZnzEBdX4hWVmCqMH3w1Sqes0V+i5CxMhsiqI1Tj8qnc0zSH
9EVUCk1q27rg0M4M3K0H90PBeY+rncmHGCK0EpywxIOXh8rDKmaM0OZejeU+Vdn6
kVx6II8sL73ARS/HYsnJhp2aD7axJPRmpkhPe7GGszwKuYTSZdzUzi+W99WFo39+
eHJLu0udA2ujaGCgJShPCtq+GnyGra38eIPTCnd7LgLYT4Bs/rFsCNYh4IlCoQ+6
k29LSmBk0XiEwcthXVXOahHofNGOeiFiHvOeDHbGVsbii4JnxLzdssGAM5hy7OLl
NDbzRZCX6QH0iGD/OOswb7x6h1SrF8Nv2I8FHDLRhNiCd6Wbz7dxKnzJbmxY0HH2
UrxVhACGICwBeM9fs3Obk//wsq2nHBrrweym/FkN6nzOEWHJGG9a8EE+MTYgTGpx
uXKG3nOy/H3aIqSDHmn6M1VUBwtvcJYWy3ZdqihW6GIsMb0Qu+jxhFd74h3a7mb3
G/09mHzflWj4uTduiuHCgp3t2bFwmdbv3qZYNeICNHGL0uSU4J5+NFxa+wF5QO2h
k45zrTdbRdC1F2H8EvNBXdwKWtrVkUaTThPKYfy+H7hGhLWB6rUbgkHAcnOC95LJ
hOrb8DiMko6K07zUGVVWDA/dNyvM3PGQa09VDaxOVpjvyvQRzrxgDiTHJXv3m/i9
KMxlptIezqz1BJ+hYeARUWinPf2OI+h1UIK/qwhK8LXDr3V6wQzgF3mCD/9N/Ny6
YwQAYDPrJWuQMoIj7OUIeRP+J6Qme4TWpq+585L+w7ynCWLR4ioIStvCoPmgCarV
DtYtQw/1kVBKMc1CYjwHu3BI+Qgmapi194deZUjT66DV+5tlnJNPenBQeOD0GckO
dVd02bn6mQB6P2Gu/vp2u4jIgKabl+CubSIyedOUKBqfOt9BPFzqNFs0ldmh4PNy
Q5SKBjAZZRkRK11RHvmxn/5V98T3ixdMzwyjCQ/h9E6Gqs9MJ/BbGB62QvitBIOA
nJANRi/58LExGvkaVnmB3oPbQ6fzpVHFEqdUvGiWbyUhJ9oUp6F4fFpiWHj1P4HR
GEDZxvR26LBmnw8SMXRoRhAoIdhmYnRFQvxCJuvJMpq+nwPHFSjX4F22irq819IM
AZPHjkwiIXAz8d9i6agpvdbQUwD68hL+dX46lG3W25Ef03dnAqvYlOxnYN2E9FHu
aOQ68kaNtnWoD2ir4GQDKvMlPvGpoXBa5xQlqSAUl/i3SvbRtKnK0yTROsKS11Bc
N1GfnvdForYUqOtRQTc2m86BBRAlOjcVCZCiWPrtESVk1VnQWmebjhAaYXHDnHWZ
QlRFwQU71RZRVClHC/cckzsSqmx4awrqKFZC8BtaEYTp8zpkZPe84dkW8jxCT2hB
9peRLwqA+Qe6FF5RPNp6Xpq740HF0IDtXeiyHPY+uEaaCb/JGGhtuX7WtjIFd7lt
r+dS1NKwWzO6r3BcOar/GeH/6A5jDwZehEfBLB+51YarqMhnLFQVpm++0I10O8uD
n+RtA+y+YdCBxL5/mRPZeeaaEg8OfG6zIS5aIKH3S4hu+j0rtOzFUtt9cJgT6ixL
rD9OPMxug0immqVGWTHDrdsd2BxuhjLm3N1BSdISrzxr6ah1/8KeG3zidO1ITdT4
gbp0my7QCeseSS4kuhvYRcMb+DdNp31BCQxYljnlANhgToFgcwECE37seXC55eCH
/XIt6hQIOgegsGB6NL8dyzjZncoydJslULy7dwRTPEMksRdi2hZwBMPRDCux4OfN
6KX4QqJ9uWtBbgEqQrkIis29TeMZvNioA81Lunx58WskvCNT9RmLZCGXFYBAsXqc
VFCL+wwf19vvUonmvmsmaE2SU11/IfWHt2BOlq38MbxpuD6r+FTEBYpgi3Wwf6A9
YeU98oIUXQyoIaHEvWRRwH2UGARb3IGXPoBzZkM0GBeLhrEm8kvvRmJD6UGxH0Yw
uAsxQzmgZcFd453Yk2T1rtOkT12y/vA8nAqz97eVplI9avt4WJfUpSDE8JU1OiEL
O+PPnXZi1KDx70vTp+aid8dKbIISK5Ftr3n7lQsVC9f54EFN2Ve+FeuEGewXFgXD
cffBw4/OetPa2o2LxMC+tfDSgpzxgmVTvZEgyOAmepY4Nga5E8qfOjcdofBhdD5X
wDNL6WHVCcaY819YZkzl42vmcZwDMFeHa8zvoT6RtbPu48FCXwlZP8JhWWNRqwLd
feyYn2shqIeccXDXN5v8HAawf8Ag9zEQyXs1sGJtmBmWP3Zjt2Y/Q3VY5x9NelgA
g5HjLLtOSqmh05TaRPBqkTsF5bmmhxwtXrrIKcLiS8OQO26m5t5N/bZSSkraE6Ot
SRiqQdJdU9yE+veUWP6d44MfiQdfeBaURFhiYLAkvTYV2IQx5KaQLCwUnDm8/bE7
GZsqaCefD/bhQG1FkaKuAm7Dnf5UvXFT8WBto9sSWGqjSbrdc/ZuSyCbPn4gg/2M
4KEcAPZdZ14ubte/4/APvGCg7t8qj0t3isch2/urkeXHh9GfNAiJHHN3OFzst8PT
YkxLjPdwKzjAANMKM1mXKd1X1UFi6mumgCjUjIqgPOd6q6uhGo7bqpbiU80fWL5W
MGEXlv3+UWsEijYBI4jjGOWO9exZ9c4JEPO6VZjWJh8DhtxO3CTCjtbxpg5p+sOH
XL4/zz6MBA11pv3HfFfcXIIg5XfnCsmW8fNxM3x5k0lpDGI/hdIrE+pD/3ZGPVDC
ZObAFogZEVax0SzHP2uGwkJ2Q1HCGtkB6XJ6v5eg7ZmiyY4xtAcz3kT7lcOGku2O
Cy/U+HWKTjvA0SRuJWVbq3ZwBXo8ZxYbQagSDTdLpUao5h1+tzQ0PsVZGiH/V9CU
S9jiD79U/Cn5WNnWSmHPV9g2M9cOsKB3+3b8q5IRS25cMtpYBANuEl4t+J/W3PIL
ygCTBxQI125ySowUa+aScF1W3K4IKQotXWV3t0aXz36Xzl7HwKipmr4+ZmbesDDO
68H4NQELpuCQeqwGzBmc5dj1uZNha5NZWb/R15jmgBKxq9VS4My5NQsxXnlt+MRU
2cqEcgl9KEAe6wIZbmyt8CP9BXxnammE82f/8PcEnmNLVeM0mDAK/knj3lpUIcRU
dg0xcMs0htrWBTroXXCP0sPKemsMatbAr3Y/gMX+QfQR9eOSVEq2Vem/4u+fTuM4
Hcy+boQ/eHczx88CGpXgc3H4LKfx6IexlI19mxt9vTrlOswfsb+TLhd3vkpSyF1H
DM43ILk6i/truj/mH1Iha4lC8JmHcnQ42lpa9AbTpApEjGHlkPnCQf92NXAQVGsa
ecnsmN/shsBBpsQMRISvzqKj2hd+Mi790VfHO8UxRA2y++v0iU3MJYf4HrZy3BOi
pAO+98+SoXhNSgdCejtOdJTwTKXUd7ZoMGiTwtYKec3JdqnfFW+4Io+Etc8N8hlt
kB56Y2BqzXoaVm4Rr8ZCvyyn1D9uO3uP0ECpLsU4aAkdK5yO3MWF60fPZTEoLNPj
X1nV9EzC0Aw0XXUmmExwzg+q/W52Z5xSKik5mIksUtYt7tUJVOTgEasoN4up8QC6
d9xBD20eNnnDz1/c9AxaiTaGS25X0Q+XFwRYPyT2lIo3Vo0BVwLjSlFWU46vqvz6
Z6JDaoUZxakOXnQOCwPZcw==
`pragma protect end_protected
