-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FXeGRePQVhYMfN71BGLNEEgGArh35Kuuntk9kZq+DeCt2RXXfy0wX8C+pEbqCplukCOMCFOyoG+o
mOmKd8obApt1rt+TvTdwfAhXKXnATAVHAjro1GsKOnk2zIMopS1m1DBdLJZ24qamSmywuweppgk4
lNcZAAMuy6/AmJX18gViPI0uNk2Zh3BQjBcE+gQl1TZOv+yD/APp+o0b5YIJ21RrgkT4QmPol9zX
i9Z5qRnawYVrCMvjFwlQa/Nk/JiOgGA/jCrqnAUmYhxKVGdYAPQxmiHuQXGhB3h88tZO4dzWkfd0
Wgns1hMUR+TedspEo3iKuQLDai7xaWKmpzEENg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23888)
`protect data_block
29EcIIRLYJmjqUzvMtkHk4EieykqhQzJJiOSTz8ikqU4R0ZAL0glcRpxfH2PiM1fTeqd0bM0QeSy
NIayKYkg6PKdWpL14fvNL7ZMY1Z76JX5imyXYW6Ts3zpYqV5zmdHlNbpoLgldFAAK+AvaK1/1jTD
TVvcqg1DF+5WDU/xtbF8rn1PQi8VWa2yfU/sZNN7IzkAYO6NCiZpYW3Hrh0afYCNYUv2qoZ0QetH
1WiIRysuANHNcgdfhYM2GkV332Vdi9lHZsax+2URzJ9jbHwFII28RARkhNO1Otx75GyFm75fiDYd
ib2b1yCZHbuM/cxXqj2EXhs1eRBeSr3PNKNzbpXX4Tw5qTeBGDOyAses4eo328Dg8fJjil1u9c7c
NORlXWGsm7Br11qt4oR6b25a6YQapYBGw2hqYjiz0Hfsi71afQiURpYnLuRjBpgT4a4Jv4h5KCD9
mPThvbPSV9+uGyPLipLDH+9zufCuB4Y+HnsAbxqNR4ryHevNs3rPtYhw3Tno6u3PQi038YL/zysF
xrkqeQ9kuHyxLX8RxwIOWC+E68H/snhwfWrZicVgs4Re187+F0CTOmm9d7i6P9RyCc8OiHgrNCIp
tQNu1pxOjw2peI10VqOlCJDXCMdyACLv3iIMXgrc71/dm1NUCWS6/q6ai7jsbBwR7fZWd1GHWv7l
jR6bGJsEC6yA93W2KCbLhNQoCla4xZUQNhbhOQnu8K1CjQ6zAZk17L3audiGCU1ZaWWSLzjZ0Ts/
tShpd2d5ExiNnovOJOwOmdMnZ8BnOqHmWQGFPpNcN2CEdSw/+WBFtjYFxV+rYGj4vC1EiN5ugBDD
edS32XEFjc0grYxZlTT7agXxst1xSbiLEQbWxJsnoE2/0HVnSmwimCxVWFAKd2mmMn6qZXGyOF4p
AakgPTf43KAheXAnO0f51sSF/iYvW+DHoj9oPcr4lAS3TmrKbgQjLbPb86t74DhJ+NAINpQTxjDB
llzuHzXsKv51EU81yV5I3dI8TSm84dgJW2usjqvz094P3s2RaDh3dSMuT7FAiP+oXi0UbYV4Or0H
BHaMhJfx21HVVlSK/rUNMZo8RllMMduGt8lqyLJcasHhtIk751xNfmehye6Aj/OTwR7LIGD0Nrsd
yQZM++gBGjsDnhEFnCNyecBcKdxzMf1ZXlD1s4h8XcxZiOvW33ntSXc9z7BgbnAUU/E1h/PaQWrQ
oqbPOOafJuh14cYcgEZ6cwaG7UNC8F7o3UAkcy6BkXsXNvB8txLxoZlLCP762oSxQMkUV6O2voaI
WfZfKGj/DxnNFHgN4ISrLI8G8C8cYWxMnifgfCT1dVblC/NlgJf201HU3cFl497MBXvDZBhVGJ3j
CjB5yP4+8KxBVYdaXywLB8s7o97eIZkzam1Xujv8ABxtCKAvkNRH66eYJchM6SpwKaeUfH8XvqJ4
5R36GgMCyvYihnruPxRz30oTRfZsROZewyjVbgCMacPoyzgP0Z6GXcw+MBu6DeLbn77c86jfbun6
g7Sm46qrcDpa1bLWknUc3eEV9yKxgX9EIlSX/i+ElF4RNBX1jFG+1FBK71BZniu9IKdU5JuJnacr
ssKvBDNqKYzF8TrnrjkMFl6jLlaM3ml1a0XTKr+oxmSFH5q116M3lcVTsoWOvd891SGz9NnQsmh0
VdrqUGaMyJOEpu+M1FDv27I7jS/+677cZO3XIE2dTRMPiO4TebIbh0oll2EgmZczzGln1Ytye3xe
lWREw+3xeZ5//ciaMO3u2stgqiSGIm3OGhqdcrtv10vcNitiDdZreMCvQBPg9rBcqRa8iECi105i
hSxGci4usLvlp6d5SlhjKVOVX+igPgQEhDfozxms1lHIiNOrVRHyUxcISaO1Tx6ZgPSUsXXdFthT
xqg4mIhmUyd5xCNAkh2FZZcQVNk0/L0jRJuBzjY2tT9fjfWvKdOI8hNvxN46WJeR7sZb2jZ8YRAX
gmB97NpJk2AJv3a2QMyTFiWLGktVHai5j52k7WwNkFwSWC4sqJGU9B9giuNG4a9CmJVuWzVcngSp
FhDsum+R+lzcXv7kMlCu50n/ASdpEMJIGgOadMbo/kHJVeG573lqrqpU6o6dMha6ss/L7f049yrS
2WpsTafRvLfuEiHjQ78cCjwtwQpO1QCg7VYYSHkFX3cruNpVu760j/1xUN2NIv4OmG7wZV7giOGI
RokwerGBdcoFsdkaUy4rTymH8imO7uv6orqhG+0Exy/ghR4YpPh08ZoXMds00bqQI5L53w0L8fac
uJu0xj5LTkj+YMQVswYCxhbeeYr6bnCEHqHtwP+5W2k3rMi+e4bcIGhuPqB6ucrs9QPi6l2EI/0p
n2cEwsFGiUu34Ei/VJcooDFv1UGqsiBZ1eVee1rvV1PjGnGczAJBGMhlaFFtkqpRwoofWDnTTEn+
FPjW6euMyznKQjGfJMDDfAHEuSx/+ucl5tHSa48/f3fAykhkn63wDrm25t548wDgcuWQJYLKaU8U
7yWftDQatcnfSJiOo0EP8W5AHUc22WcBnispfxOj5ik4DBvX919XUqw3cbHKx7z3EsSJTmzGWHZU
1oAzmMsIVJvlpyVltD3BX1sU+bCsbCqUabDudi0Pcj5e7RCnh6UI2uGqeJJY8SzICV5YX4xEIPY0
IPn6e9bNyly18Q4v8UpZXSFMj+wimkQZThJXFPlY/hWCLzB2cLb5dqT2BskYNnVztI4Hl/UbJOCN
TkViYG+fQzQLI8VmYDYKLR22EAyWxT1nBBL8TeLSoTVUr5AQrpUcx/DF9wr/6q8b1YrBLFtm1lYL
kf0gpcOX9NbQi8YOW0Jok1CrvHC0KW5GWSJ6ipLVLU0COrc12PzaDTv2sOljeWnlsQDaI5GMY+Ab
bLh446PN5md9l0y3B09nDStyXH+ayuqCmScGXOn6XAn1MMResfIOXUB/7vO2H9LaTpQkr264pH3c
4Ax1DP/t4FbXsfTsxUvSiKNpOY9Mc74GQ18KZOXGo/f7mJbXY9IxuhWsJeSwJTn1c/eB+lyRXot0
5A3Cr8jPejsnLOrabdhdXbgMRRB92uavTPFE9eM5wKzs5tf3X8/XEFQ+LcWt/6WZGSrUpucxOQOi
9+v7qA1jZ33vioddosdS2KFadpkrpH1qSlLWh4nRErAsuxN+ccFkAZlL75Eb/h8T/CY+dbKFcz9O
1e0826X00O9k9CHeS5GiuxNGYn45KcRavwOmMbwM5xrkzyuR27JhMWgZP+XF4GBhpfQDBlzqDvVH
dMVlzd/DnYetD6ZbS/L1WA+gCTI4tXhkXfnI0GAcszrgWbH98zDlH5te0Ep/zKpcSTrKD7BaASPE
V33bCNPzT+PRwg6G1YZL6Cp+y8csONqX3q8RJhOda8z2gm8LfL/voe2LCJ19vZvxBG1Ub1/NURfz
eOSqWNbL8WCdwubJ6pjF1L4aHbaVaWymtsDAYRnrOmVrUm+s9OAcHfhu+XKnWCb0oD4+LYaPwgNg
NMSResWugURIYcduYjrL+XrQY5BcmeyLOgdo696j3vOC1Jk33I46uYXLYsmQypsiT47fgH1UUnME
Eys6qQTxHtGxXqtSawwa7yz/wEVPxJvQ2q0R43DqYKx/gCUt+/Tu8lQU+19E/q0nkUqoHIIKTGCD
ZAdU/zOzSbNUYas5LrRjMesK6c4p3hlEdvp7+lKacS04u6AclK70jbFeD/OerXbd7S+Kj12V2WcQ
Pu0lThZWCzXnWwi+T7gJ4WFYuER/iD0+2Q3KPgkzqTUinBpXApRXllEFInqTuL2fBCfV+kFavnxy
d7DLi4G+IfuoCga5nlX2xw6hQV5/3Ld/aZhoAFBUENlxsZQpoEZadEUlk1C7e+sHbcsm0e6YLaoP
Z9WhfsWWFgltxumVuH9wPYumq7Uc+0hrRnZph+ei0eUljSZLhV9QyV+AqfBiPfNWE+XwX3jOujuH
pqs8ejn19MaBTqEQGnHwmT5DuNgCm+v+8xzAgUfyXDBoP3CZT681wIY03Cfd2jvwTJxjvSAcSQRM
vAzGr027RyKgHdBp8VBKnxHbFo7xfafWY6gzyy0Iifhe25kQ+BUH6TWyL9Q6nCRmGQli/xLsAg0Z
AqxaSA5PyI+HR6i3UpFyVgXI5C2ejtxI6C9ZH0jhAEeFKlObV5LnSsZL06mdS5MPFtz5E6H2TdGv
otpxzVez0I+u1/dtGPkjZEYL4TSlATC6Izk+JS2dC/jJpz75BK6BROKbqXYx6TS8wa2OpKu1kYjY
+zuVodXFguAAJgZbu0/rmTnanHzdNmrKeFux/PQo1Dak8+ZcVX0VQr4+N8kwbb5VUSP0/DinpIXd
zT5D4ZS97r5AxDWw2pNfqM64zrkxx/L9myWdFAGW1S89mBNws3DRuxUmbwPs+FI9pSPDTA08bw4J
zpYB2rHHdZ3SxHts19v+hVYsPZ1g4AcNsKmBWuPAoYnQwFMFIMsGr46Io3kr/cpB0kjueuLzet1r
ekaNAbmY9rll1mXceOAfGygIXPHSd/fp2NYu1V566Md9qvGHRJzi3+R6So6Wnm5QS58ZOCdGyZYk
C5VVfrg38qknKv1SqlqlA85wZ8pw+tN3UT1N+QZkgKAFzqRrdWVZsGVT5+8og+eASH3C2o9YRMCL
M9x5mQHQP/EjC+R/LpQj1JNKF5SHTXA7coT2X6tgLi0DNxthqANcrrB3an/oKdMcLngg09qeNP+j
tj9E0+75J1b5G6DB5jCUeKoFQPjlxgZHDMC4OxQjWF1xopqmp/hy5QuW3D9CeLv0dkPeHefNAIxw
u02JsamOFOOPqT0EEmgOXzGl+y0rz4J3/qHFggse8yEl1ovSXbNnYjchpj20ic3EdhDbo21WN8PZ
iu9s8rSgg0RGPZeNVAI8LOJQQSrPJkVbVt7k6YicSmxMa9eVG5jhlJ7qt003EwcuGCs9Pz1L9C6o
RAwm7pf9MX318BGeUaqar4G8cncSmaYTxAguIke2I3dG/WwmuhelxGX+kZvEZeMyaEfSOeF900Jx
ZQFxXGquCdriXTLQr8jWe4JmNpQtSWl5Z/BT8+Mxn2yBjB9B8QbWC4zN6EYTHs2fyHpoha4EGvr2
t3inQgtBmI7mms937Tkmgkkdv3u2f45h8PRt2hD2YuaMijKB6uO/5dnpbhlFs+tAnPy3WzdxUPCQ
9/wPKmF5ZWYk50tUOkVHHBDAmp++j9Gh+oq3zmBTWORC1TwYdSP1yAJCA41x18A6nf8eScNBjkcs
EJAB/BWHnGibSF1mlOBF76N3Iy9OMZL8o2uy5Qh/YcODx0IAi9/mcI7jbt/BWRpcX2lp4myu96zT
2Rxica6vL1bJPC4Y7ioAiclPCRCz5HAl88JXzMMByMViA8WD+vlmMNDliH+VHOpwaPAJSH6sO+e8
mSNF1Kjt9Kxfu5+8L2Iqh8/B7OsiglHuMug6CRg4FaKMdT/gIAUT7NqyekzJ1zSN1Nhj0BwB5Ama
57t2AN2FcLPG8KDIAbZyBa3Mc6SkPek7V4fGEwixWCEZ6CMNGgPJHFFnOVZT3YXkwPG/4p+UZOJs
Iz/ypnnMBdd/DyYrplxRU5kM0qiNEUoBvWfyJd73DZnwYuPzOynjDPyEWyUSFwnmmbLVJTAn+kSH
9RivbOWjRMHVSfLb/a1+2LPHdh0ARyOXWg7RAD6Y3w7sDxZ7wFq3P7CAnbSZZfJzwnzQjTnibxx1
nZ+3UeCztEh9Koi8hUJMB9tWi8Y28LJPOV8U0bIvTWDi2TF74/RJTqVZRvoDv+eCgNHgRc4/Mg9y
iRwNjc+zWMf87GPYRw2JfZ/Ix9oHH1bAisjBbUanNT7EoZtYjZ74pj7kO5DMr0gb7hYsQlaIqGlN
TzRFfhs7uPHNcH+Cb49+zpYzPB10o8RTI0GPTE5eRX9FZsttIOjoRzIyLcQijUOPniIXoSLPkLdW
j7j8NKbeEFmyPtJnTHlMWEYyjsLD+F/fYwHlmnDMROkE2LE73xh7WSxQmEvnVJ19weM/MtCs/TvU
hZAagddhxCCucta7lCTIKvDHUqPwF7svkgnVYWq2gt0cSQ62sw0COs+QWzxf2kEY29lSOj4m/Z7A
JmutADd0OMXqVElv07uWNjQZEmfSSDwmYtJ1GDeyKnQBvU6h4oH30Gu88nVy2ynf3nCLEieK0G6O
PIEIs4Pwxo0TPyMr6GmHp2BfXWRLiDSvsqemee+DNJl2BS3PymG9DpS2iJO9oh02VplK622amrt5
uuyHGVEeHeZkpJdRQFCrmhDFoEv46QvlIrJESJWsPYOY5Dor9mBqmtBawdWasrMSXoZ640k02JPb
/0KhTFR8Ir8AE/H8Kl8SabzMVJjAMWpR0qsq9S2jUIZu6h7mz8Idrrd6O86tGF61qMzkCDPKIMmQ
kzWJxL+Muswhj/qvvimJEuoLvQIDU9RZZa0IjxSZ2MAuJgWCXzfL1cffaLT8dt7Syg5LnW4Pj3b1
2+LNbh6oAsyV+pp3+o3P4ohltzUBWA3FFGPdD5+5c2Iy3Yib8XdnXtKjHW6JzQKn/9hFVGu7on2F
sWDfkrhna6yvTvZlrWjPszYAiNblvlar6g7swZw2rVhTWQJ4eTrj6G1SAei2850HDFHPu7aS5isK
U3h0JQL2xuvEU/JThoTMFA92EkeFxALTEHF/XVKB8myLlmqytfWJX5G7DyLGaBm0KApV2QEarqzW
rateMwEv3jk7iuWXqyfEMnEuBFgV+J2UE2iX4G1nEV4SUPv5Ycjb2t9kq2ljARPHthkV/+L34OdO
qLHav5xf3WWf7QqpYj7gRT7XbXrU3IF3yxOCtbzz0kRVfK9vhbNBU7Q6c8oWy/lFQumrCrunvmeb
VToOj9iSeM2ehcLyjHJjdflyuinrL2sKwEpX3ysFQ8v1NIqVvdTeWO2GUn1RHxeDidqTof5vX+Yi
Z/5wQlufyKaWD97ioeZcXfBBDfVUPyH1mTK+uUxTfz6N1ipigq+Kznl8M+2urBCtdSIKMnIP/H5Z
lhfnjHDyIKjDk+PRqALByLUXGSOkLrL7fCze5bil3vpLLLBnu7mz74UnvHZmY7GsesfDmF+/t/W2
1Wg4aJUmJ8yYn+eBRUi6ictk6syQy2Clc0bm+E5/rxQJvbXUp/ONIdJWK5FQBJwCDld4dVS6bY/w
zIRvryaRTRJXgp1wZwpGPpj8nzHyHS0izHzOQiJfIA+1e6ThMAV5dOr0BOHAWl/KWZW9Xp2cwnhb
jlPTY261H8ShBkl8LxCyN84l2SXEqYfXKm56OwZAO9sej5s33bs4bQwYO/4+7da4h6m/TQf9MrTh
ljV+2FFvQqoPdjTEMaOU2ZPY+GQH/9/wyBM10YVjyW50ThvzYP673HuvvxisG7pbpC89V4zowwXk
8yBynkvo+x9S2V5jGc6QN+GbzzxQtI7psdsbsZz1FOXfpFVz1fovCMzex8VB43EYuvkO69vNSILT
EiR0+pY8BwUiCixb5uC7sDGVgjaUtSrjxq3Y1h/Ry1LMJXmw9ja0oiUrt3hiYnEI5imnqJYX0uLY
yTHkms5HgPIaAGA06d6uc2kJeTuB4FvLsLZ0s18xcz9HYfeH8HDJ1uqaw8oKEPnc3z3qdEcPZh9U
CQCl53gW+mK1EBMOS9SwiRCFh5TS+rOafdLvFAUlt9vogzigusUVFPKvlZ7tMSHBtJ/aDbTnK9ij
q2RlhZqffrZgPsrWd+GkeAytBa7Cs1I0pLrz2J1YIZTBnyiKSjXvIt+TZtv5/YmyamAYK/bTqXbI
eO3o3MD5qBEbFfMQ1/n5V/9Vnw9lekxDiqS2SWnxT/ez4RyQb6kfL241ew6vq/FdZDhFhuoJRC9t
ICzMIbdzA5ntRocNJZXQ1ugv+0t/VuINMB9vaZf3/9f7GR/JSI8Fekq+BtCg9E1f8ZJsDzyVuQD+
Kk1Ds/JnMLkhf3gCVpecEapQ4seM484uLW92DXdejDglzdJzn3S4uZL70cGbfW8Oy3N5DbwXDh5h
3OVEppaQR5AprCk4AN98+PJ/EPhw9hioEY1NcvEC+9UvbhWcgiNNEI41BS1ODgb2csmfUrd2HaBa
IlLuKb/gckrAmzDB8vO0vQsYEANHntQ+qWhdtsn7slXMcz4cNxbtvim7WiyN/80Oloj6514ALc7p
lLwrLBZjK0V9pJpT6e/usLfPNTT4bi+i7bOXmwl96UIZULXBMJqjOltUhqCUFvp9WK/IgywJeh6t
hkCiFY4mMahDlO0BTOKj3dkRXcxYc7pVPPQa0MyVT9QFwhHN32/hIKpZD2tI1FO8Y0tietaxux+I
H903mK2TQ+4i9e2BXtDk3wQNXYSeesYYgilG/rA212GGMrBi0ZmbVIawR+vMsMCCPpfz/QiJdji7
7oB1JBr0fisDi3qyKN1tKUREJrMoY8ezqeMZ1Q5KladyVP37N6gv/xGiJ5m0oC0qG7LgG5nvDhc5
7+0i/J8ImiiLjvqJoR8ySwg2LBKesEnLeRswvcJ2KN4d9AR0w19Ocm3wkC25cWNR5+Kk72Pa/sbY
R44orqlc1B0k6InWqGoeMYjSBMiukt2rlS7t/94RdhGui4WQMj9zL8hyhxFMcmb3TLNd6Piu+Kow
f2+th7o1jbC/2rXGHVHjuIQnjtH7lOl/WefTbjI18fyfl7ofXXjlc4+Xm5bs+BAVSZAxBDfMLoKy
rR/3RhBylO1NzRFrJ/3Clqd7GGnfiqpU4QqighqMJGLmOz1jnG7PrNavn15aPBgG1XVDgHzqUFlC
w/71SiMN24XFte/Aqtf5nWAypOzXZ9rpNYg67FFKpWJGSJuCFOzGr7C+311yYRxigN67CbD/rAp1
kJDjyqhA/zC8G89vsXth/V2+VvCUzC0T6Gi0Ts/iiP/+DOZgoSR1r5O6efkh816papjOxS6zxp4t
hidR+bR5tV0thUEAweQq/KU4X0Dloxf5uD6bLlq8ylQoNGM7KjK1aQvmX7q9I9O0Mg4N7y8OdirL
9Mijn2tvDpGVLcgoPRDMx4mFBeasc9inofAQlDrnPVGNX/EIkf1sMbHbwntSUrGMbYreHksAkj7C
IzsvhyHYfredF6ctVFH4eN2vjv6I66dsXmF8eaRO4obQhngbFrcunjT1Et0UusOsCZwslm4jq/Rn
o0KoAPSLKxkFvWboYeAfyoPj9gZtJZaePzfKzdCMEdoJ6Hw1pNi8CZW4nQxPXYhGzy9F8kHN5tsv
Ar4lc7QDj/615uPgwYxMwfXCOP6pPP0Q3DF2YEHNDmxU3Lcsj/E6uKatg/8F63QS1YI9g8vuF84a
y7o4VwYnPgv+HEYilcFJ5nFXa64bTY/tIbe5s1YrBfjhgjGCqoznth6eJmptaF+99+1KQaTljXWv
jQMoo9qkEKVSD5YqZstdcRQs8j+wRkVJMGfni4R25GjyyPk9XRf5zefHcNHtF4RFJrR4pQ01V7Oc
WGo6xPMn6x8RcOTlL5ZiO1iTJt56zY14ddz88537VfhmfqeAiyv6HuQUpc73E22BOEW+zeF4MXzF
GJSOTsSN/ywsClp3ZbQnESbyh2RnknnoI3NeQKT770X6lyhURaFIx1E+EAfUSawlXPmbadxKkSW3
+KJbmTGs1mOP3gA5Tce1FYtpAORxG15nrYBn076rnoiQdIvuzgrHzvuadjQfX6n59cncd2l1OkAH
CdAfK2J636J9lytMcHfiPNWYXSr9Ju+MLlmLZ8NoyisGpzXI4zEltKDQw+1RV9FckRjpPe9X5p0N
7rbp+tsShkxcx+scUiVRnvV8A39r4aWU0yxEG32rkv1N86PE+ex6hxQy3LvdXk8V4k6OeE1a6qDU
w8kT+X2PZR84i874e9BmvJYFedsz2maslcYPSC3XCM835neJ0fr7t6L4vqfAGBFtaGdYymNArMrK
Qr+uyUcYZmIPFiRB0RTI0+LV8GL9817hbcAxzIkswAydHDyUEjou3wk65t2OYWfy2fJ/SCp/b9yQ
ZWGyz14C1TjFdBFMCgYYYabJGanz0bA1e/fhTMU7zRHYAL+pVMbBpm7Bq8MxFo5iUUF3jyokmF87
InwH6hAoFkXVH2CiMwHl5X6xZclDoM0Dw+iAezG1Nj5uw1G0Y9X3i6y16/WgicaB/EgToJk+HBYI
vZQCiViGGY8v/EJn6jx28DcxD6lJ1pxIlTvyK/ITrmEPlmdIjl/ROPeKkn4RC3I3x46xQpibNhRH
Tgee/4cS6ju5tTjtGxr7broXWZO4+6YUBddZ0SLny/33HQVj+bbQObsMRYWJSELm1IuRD9bihEhW
OGQsJU5dN+YebO//7Qx0DqTwSQfYl/aDVwO8L/WQ1xpiUsw86UY/4RvgJIlCo4slpc46bumwc3Rs
aUUYU2Epkwa+0jD7h2Z1ovV0s6mdG3LyQacGvqlccYtnMBZ+zS/UptENErFTfjJF++xsQV7u0lZI
2vLmNbFT5kbvWGtgPe/fgL4sTNrCiJ5GQVPlfv5aZtEPc4yAjD4RtW7TA8W3XPgUURtr3LHkEjlv
vKoLBzfwfmezIDVTn5/ylkspEy4RFt5zja29E1v9r0z+3mfWikw5+v2MVYiVToJ903vxN6HOfx/j
AY2FGM3FHcl1P78DfIrnlKmwp7JwSPc0iHA/LNPURiYNXL5rzfE9bzuhtktKRzPDRiYw6/9uhhBn
ZW7HTGa+HOqrue673eXQZVOVHWsN0EKKhjk15UDHCYRwR57JGN6JkclqgZj5EPfhDrLbUuz0Q16a
uuGsTq8JhI2g9IvVAPvBWzrtp9SMdSnHynJj3MsQSs30UXCL9+ueEKkL+MAy79+cVy0ifZnDuhar
PtZyeHbG9QT6Ws+ZJvpDNVJgxudn6yFFbPLjRkAmsEPexBmrDF86DMtiQxb9sT3G/4uqoNNmpiIM
kmhG0WMANaJA9j+dCu2i+VEy7dDSiE4zZ8YMybiA4wGcTuITl/I39A5Ot/nC4h9pujPhtjFQn0Wp
djqiCNMJmx+OTYCBohK3Rt/Xsh2YWvzm2l//JaVwrSXJh568UwbKsMOA+vH5yLqnbPcINJKMGwXV
EklO5Zp9hqHX5Q84RBWA1SgTecN30iP4E6JsuD8FIWG8NIfMQT/vUAm3e3IV45aL61n+31uDchtj
9qnrrRioCLVn8u80wjiYdH4LkM7CDRA0ydKj4d1/tJnvexQPpKuFPhNpieGt78E/T2KFsS8qySRk
FLRVGgYhxX3+82kNgOghnqNpWOt68M462dWm5BhKAecVeYlxWPxv5Jt6HzksZTEW5FmS2WnXVDcC
vbpG1MdqjBlKwf8GYRB4zZHHh8S6EGzWt+J4HBV1TcXOqjvAvh83Wi2SWtsxYX+5MRC/Z16Qga5i
BoMgW5OZHmE1gd83TsYxgV+UZypVIxj6eeCQmv+cRoTrANKHBZ5uBhdoqTEESXvW1xXb9qydlQ8S
4RRvGp8YaW2aVJucYeS87Om7jrTFqkFAsAkuEDEvSiD9sLUOLX+8x+pu4KSfVckxnCKZU1pCclEt
EcXQlxqte82saqEe83Mj+nRshWO+d78weFTigYLGNfBrcpBuTAWv9jk+7PQ3WreuV78YW8weh2VS
4lPTDkNiPoedm9h/iSu8kDIMYy/2iEpZmFM+VSyrSnlSog5TYrAcuxz9UwHqQitHKI+zdi+CPngU
CVrpeFObt3Ypu246PqvaRkSdCGniXv6zY5KTe5zm4uTy+OEQW6NdaToeUHfh6ga5bLbe0Jlr8L3/
HpvF16xvxaBA6jfpvhZqrlAxc/cG7twLsgo8VYpOW2Lvg4pqnHh7omv8Hjirrk8wBWCeTcdKQGsy
080QLfCRNJrGZamXG5QwKqaYg2PfAY3GohtnV8cg4i2PXLU3S1Q9mueVhwKWWT+t2CfCXE/125eG
7xKmEsYjkagpa/MaVg/6sDDrohPHw+9sAPz8MUK0pWDnWz6RwGVcsT+wjVffSCw5n6okiLfY1S0l
F6MGlOHLEKDOYKz5rwjSrGmZz5NqinH/owwcom7LSyYULuBHHWnaZjuLT8GbPZsmPE2lzk+LRk/v
lDI55wib6nXTO7Cp1q+0CzxWVh37IenDVAKI4MhuS/EpFziXlrE2W9n4/drs96guSlxxTrvQiDyR
1dlHH7ESh2onySjF+eYeJUzwPyV6BZtCjqvVz3v71pwkdrPudz4QQnyqNSxxZwZHg3uk86Oocn/0
/FiZ3X+IKna6zJRG6MEL1lRTCiUEm21QNATGSHQMliml9BQwAAS+4TbwnMYnHNCuiAnJ+S7V2KSF
OFXaiu2ldmRpwsijdrC4fQEIs3zaxxly6syKzMACoYiTsGyOJbUWW182izGV9MquTX046+gyKnEI
z+6Nh5aNHwLd6UTxoanL0P4lHzisHhFnqgHHY1YzYrpzGb3N5y5DjY4O1eOtAvxw8fm5h/7eKxsE
nLJnRngMQchi0KCjeF8z7p1fvuXd/lk6fdX5Kscex278PxG5c8h5z1js4u/MnIcRYE4Wxx9dSNcd
uIoLJpYbtGprggyQlpewSIUiuRwsWAsMjDbTMj1oFvMk7gIuFumRIq52GaeHCv36Qq/prepJVrM+
oqSaHz94DrozuCD8cWOekA7WPUEaqC6wC7U3Qk9V+vQ12lv70hwNTTFPyT743QD5R9lyLs47u6SW
FaQzzDm71141pLwNGn6ibgBiNZVIYALVqKBGIIpl9z4unTGYrLrr6xZFhLYaMQMeVBJl8KZePQbW
agTSAWV1TeGb9OXd19Fzq8DgP7IlYZSPYs4Y+84VjpgGXhN3wMhwsp6c0CSBeaC2nxyqmvXnAWsq
9ozMM9NRFr9fuzIBIq3sOb1KkI3l1ZZNjDrEndc/WQAlh6Lk9bF6psdX9Cx17Mpzbz9gRP3/gleS
pY1yRnJY8sasV/KidSMJ6eO+SQ0bZP0Bnw1wdXCmrw3roMlrHxNo7FezGvpZ2M+WItzFzzO5L9Ef
/eprI2/Xr4JAWOrU2jRP+Axat68SJdIlBg/4FKoH2d2hSWPTrZuxqmigRuNxuYPKfs4Cm58PrvkK
mC+OiWEjSSkJTm3FVRNNdTSwPTnEMn7VmkMStymLuYaoxrgzOJSBp3KrSnlUpUgupMY0A7gfhjbw
wUJHZM7DbyZLo1J8+8a9GGFrBNtbajrebH/7HFrZiKW95Z/N/XexQoqPktGFjNNdZ1K7rzAhi887
jpVVvgYV/ebLwg7GOaW6Ev5UIr1Ss+4Qg4ajglKl8okN26aU3gM7XTY3/I8bDkJ62Yma+VPZAkvf
cx79xrYNXfMDeH1LzMrvh6MR2aiGdgizqxAxy5svpDUdoOSCG9KjjdbmEsMKvJ4eCrCldZQy4eSD
swD7lmKv+awT9ZAy3VNz5G6iDwcBKyKykKir+RqIyd0JEB2PD6sK+Fuyis6Ue6hZRBhFrYP29v0m
++CarHZDQ0rwk278pgy3t6lO7RwYU7V4+2RxvugX04tlsknRm+e4jUv0ESlWwMH3ATiiWuAmQ/Up
Tghhhg0A+WtZ1/sJ6TEHIiQKlJlX519GxcL9uS42Y1EZxaDy+pWb3xVhDJQGD4pvsW2AVvRIJt7K
7IuGv3BCFKi1x8vOVEI6Ev+LhIfDRMLEnL/OvjhpJ/wiFeF397bDsqz09D0mkq8+G/79ryDxebSg
fHCwIfxfJiIyW1ovzhKpkz4MTXGEZBuFKSZvtD8/2AHMIREkadZ40Ozp+RPf7x2h6CjwgejxlYfi
1i4n6lA+GF0/jSYO6hi2SIzw6+K/VxRpPN9RL2gdmIT8tGOWW2owpByMIDLNirbarBlbFXmDRqxY
B/bI3Ju5TSmqlUuAJYN+PGXer5AvBTbFC0C7oTvQ3qOhDpoX4SE7lk44IgR5OaE9T2UOy9yeZv4W
F2y3SQbPZLdnY819cg8czMJVyZHprBsj2KJbCfe1Byg8umCDmUAgFWNzfco/kRWrAFSO8omGrEO+
J/260j4Y/91TJ4ueLFnFL8xWwbqqIeQYPZrERy60ZgePGKmBaC1BrASVq3kfiuJKBbMbrQj+c8Rt
GT51gAxkCl6LeoHCbgoAg8PUBbD0ZIj72aJlKskhUXY85LpJcBhimhqs/7wD8Uz/N3OnZL4IFF2p
1UevRJydbeyBvfUemgXh8KGn/HrYFsI3UWkgQaQ6dGaRgZuwBC9PetonOK5uXqerbmyCDipeJmbH
2CEMlwfYQeRYbwgEqvM0hSl5zZ7W47/Y094sVsf9F8pQdWJjfTJWHCIXfRJt88rj4BdQSJCg5YpP
eo2VpRqC3d7xGYdBTfKQ7PEo2cYf2upblUjI4LbaWRTgx8z5VlK8dmzc1YwYFP3el9kxfrn5jJWL
/809RMSj2yVMOjuePHhtbrJ7CVuR5KSTRblMvT1aPPBTa88yrlrYr6FLtpasgXDwsYN5vx5/XzU8
iRh4fN+woMWwJXxQah5JXCBP7Yz5WcuWC2m+6fqt3IXxvOX5jisxdCmDPY+eo/6fmIo2ojwqJjO7
N61rr6a7kpCReWU0TtGpXrwgOlTgBd2jfxQePTfJ6/BzL9yoAQz9xlkerw+SVcnsrQczuCzWz4Sc
gThFx25c+8ES212zrrjl2YjWY3hzwqzI9M+SPNtqwCIPcAgVjpLqW8WHTDDNfD04G7XTc3LNTGWc
WtZmxvC61gCj8vxxKPZksbjvgGz20rB5MyPPjYNZtLLc5gTbJUFhpSs+lWIV8feqjuSBQL+MIm7s
/elp70lRbImUQejyfadh6Re8Iz3am+1VZQd1V02dz28l/7eQpq04KpLcp4mhyEvbvJhBr5vcuCdF
+nRBa5e/Famhd4qgRrSCgwNp1epWrRjzz6W5jOoWU3mhKN8+F/YPOB6aMzMQJ4MNNYHYWxFOL9Hs
0qzT4hwjOojKE8pxdmMxC9hxR0Inr0ys6spjV2zTteYptfnIivnyvoMDwcsCucyUsRW/EliGCSuT
wJffhjPYpi5zyDuFrDqYc0ugEbntVFbn3vsNwTePV3IsHguRr6NZO6/qAMvwvIHmifxd0DfCx+1O
CvN4RHVxVTyd0xtRrP/sG2+zZbXXL6+aqiNpkq7kbgYguK7dxTltk+xPTO5U8p4stI8cSiUC3n0e
CR6yshITBGYIGDLViUvfK5kijZRY1SX/DlD3kWm464pvMCD36xAJFkNtQPIhdu1zfjffkP0H1GiZ
iZ1krC//4V1iv/wGWRb5AqIbHjshDggYdN2Q6dlFjFlg71uO73lReUm51tcgeHhs7xtl4Errg2JX
2bq7RrlBjHqgRaeigGrX4WXvegh1gKV2QY0pYtfPbV+YYQuXgEgMTH5IBGIUIZ6EePiOIjJwcwQi
XjQY/xKXBWH0t39BiQLA34T6MpwWnlK4POADOC6wSOxXXawMpQdQ5cauM//sGZG+aSHaPT15fySX
mFDopHzKJnVFPaiG4C1Fy76KdfOhy7mpkOInsb5XBBvD8w4CErWslVFrDM4fR3uKVDCNWurPXU7b
DbfDIvGMsugDLS7g6puxvSelHkH+WCMe2McmGuYRcYQPicE+MMkaHeGzyGRE7XPM9i3zF3p3L3h/
7xi0ymZm9MyF6f19WOzrRVzTem1qoXaRekb0dcQMXwFVv5LrUrEccawK7gtWgm3PqPivNgU6J7lf
Sk+j6wUoADIkWS0j2FmYBrGJrXxi4WmMXWlHO9KlL3U7AmMXEXelUjjdz2qApJM6tEHxZNepgD6n
17MDLLYoe9wFtp9BwEI2MyhaF9IZctOl5lonvI9wC9Rpqg8ap7znwThh8GBZWEU3AGXctVQHQayN
20r927rOQPKc5b+sgUwCI1QhYnsXzoQyusmpvJX9wtIxbtbFfrmzBxWRg0gSq9s4ljY39Xe6G0ew
V6IUWipJAccQceGNIz1SepCf/HOpF7PJvFetmzFiKQCdF3mMtGqOLB5Jx4JfKrHNd02eCxWXnFrz
v74YKoT2M71D2UzMnS/jlcSjyuBVPgVYDLhBDx1f9qv770EGXbbwIVVqJR5IN62Elj8M0jxdC/AC
cRg3HKZzgAoB4TVYZS+Kxo4oADYCC91RdCInviWfH7pVmlx9Td13OADJwV3LaNXVmPk0huT9YJ4d
qeVzrmY63Nkv6DEbtXFeMQUDrXQmfYiDlr3c3gycmKywY9VdDO1JfxF7FVZxgaE0K2+QU2beQzGg
z0fQPR5ol0OfQ6+dwy42okkoVdfVDLLl/6QQcPbHjwUej+G0rAgse67mim/EONyuCge0ocwgGh6S
iVQ6jrckpGlvf8VpI/HjyDTRjmVImLl/1bna1thnWPArwMHeFyEzT+uvUHEYcZeAK+uH9hui23o9
7AOYCmETPo5+VaVFR916HWLMkGjXoq1lq6kQn1lDnoiC4MgpDP9hJc96fOm02eyRz9anVjPMLGT6
u5Jul3HRusF5IYUBKMJPbx+lI+qfM5OdWyKQpxcHf9NVNDKP4qm6Gh+f6B4eFVVckV7HfhcceHJQ
gNwXJbmiRk0z/Rsx6igQ5gDacbCfsXb8TWGbcBcxxhaR+ZqSi5VJWDizdWDQB76Py6oKbMxxyeb5
zAxYE59TcotmWPmNh98/a0K1/F+ScKK9PSzorZEojs0b2iKYlDtft2O4pYDrj5Ap7EKlLANKAWGR
douklXzvLHpRdhzIElyViiUo44WsPG0LSeMkWTjOg8CJAJXVWiJgezksmHw/d1Y7r6DQaLjHX1EF
F3q6SuFVn/iyfip+owD7KQXzKlzmE/0axA++nO7rhX3XcTllltbh80WL6V2b/kCgdVKhTCinVsWn
v/J3GrJDczZXsV2On2hAOFTNrJStwmt8Rf+3YhbT8RH5iw44I1pGzZuAZtPphL5Z+Q4bxid9xy+U
lOL4DBTqmZMrEyX1ja5ipbpz8sbw7ktOVpiiI1bo6zGSDyy6V6faI7dh0UhC1KcxzihZm7/5jA/J
BV0FBG/LYss15bkK5lWxh2gTXZHHyxXQa7AAqDcberYNeaqlc4HTNHkrjmcFKvNFdSnXF6+R8uMn
1e3yiDHOlN2aXU2v1YJ7ub4bOp/WRxbJYkDSbKK0kdC8pCMeeFvF5uUqsve8wdtQUgBBMJgIOCFf
8e16NPOOqOuskBZRlKFCs34umQTZmUdNR0P0XJ45ZVPpaVa7oyqKvdjrQvnipZrk1DAHRQVV2ycj
+kzz77AQRMhnxGMIgI+93j2m5wM4yoYh9T77182z+IyssSPR5TzJAGUAIPhIrFrS5pFlzkmZ0xXO
dW6l38jbVYWtnAInzbts8C2O8mi2GYYgMf3djVlfHi51GwcN25YwvuiJUx7tXRQ2GamDkOs5J7EP
UbplAc1ZF8jmCTx+BXmbqid1H+4quFnbH3Vw/ouZzblQIaDAi40Ggok5agqOhW66jyalI46/BhwJ
sZXpXs8Nlcbq3JJFk3PbeKikF7BcjnC4nCs8AKlZPbzaYlTGQKX5sIjmrofcQ/dYDrmXdkjlYTLO
183DTm+l7l6d37pwJ5Pd7Au51mdpUl0KJB3Q+mce3ou8/2ZNvSEMMKS7wMzdP5wppl0muBuIFFPG
ShwCbgZxk7H6W+gYJ6U+XBKfkmN6N6P1BkFnH+FL9aE7ak8w6cW3NVJDxrYUVwCYWfulh9HgwUZ3
GHyXeThpgJlx/fIWQRvNnA8Ss6BITHj0Frx5egSCTVvDD/r6RT3VuI8az45AFk06FXyHsRS9+iMa
TKP7tKGz0wsSFc+zvB9coYoYNr5M0emZ7tquN6uSe4C8HBYKbj2EGPRq2QSto+wz9WoRaynkLyMx
HmE7PRBV6jpmXTzki8tKyUMjiHp/qBRghDL7ks1naZBaol1/BkJ2iArshqVQtx+ZZ98IHDE+YRzz
Ecg4mPoJtVDvNWxgcUR/vKAhwhWRiKK3eMGbZemqaQgVN4dSc+Dcdi60TJOO9rLSeRk/Y2gaZjbm
UTCCExTqvvdMpjFA0hTXy4R52fkAznf/QzRarpBoY2Hn0+yInV9rg2h6irJ706h06QJnzHYbfTzX
JIjqEMogQO/edBqb9HLsEvSF2uO82ndUD/xpYdAPSD3gGljeoKucmeUBUhZ27crp3Tc+dp0w1y4B
xPe0LX/1wyC8hbODlF26TGWlUDCjcnbd6cibKaLbdsfY8rJ6pT/YVrj9BZCvusHojTV19pjs67Ln
FuLpEwrLoCUBgc+wSYYJmyXvmuzymDtuNu8PVNE8Kd4PXrP+iTIn0t4QvjRrZZYvlZupLqXoQRkD
255A0NXlvTJc2iSTLjDyYygfTDYy2iRSUxsvpLmubgWc1vAAadkJmBwe8c+w4Aa66lJEuXdW3BBq
C8O1tL/FxYVZmlvR81nWXNzH5LL+wX3DaI2xLoBD3ZDFib3Jh3C5yoS5XsOIV/8IIfkTuyxImdjI
WCBFweKusxBmZn2hUvrQQrK3iuKUZ9Ts73gThLplvhZ9gDA8lQZURh0GklMmbYURbQABE87ItJDL
plOhewRE+bfwNHy5vpDn9fDjFu9DUj56pnpB+T95aTIYfLNyAxQEpnbiEvhh0dBHWZ7CjBIiyMFK
8P2AY2DpD5GtTpnTU6GQeaFrss/3thU9hvwDFGN0xPOb2TTEnuYS1pBoGHg2fhWFqBAzL1QsMIDx
fIdWiu3tLUwcrsnFg31SfiXkadryyWp0Lads0sfBi0zXQWxmXVlPxjNiMN3Y4PtZAO4aCqdOsNjf
+/keCqLXyvbsAcKEVMrfHBqh8mCw5gLlpfD7iisPjH9SwZc9VdDIbufsSpJuCnSMazW7rZTHgOdG
x8fV1tkmWlIOZurqE7VFdMozRJ7nc2OcWZX5cZ1sI1sjK4Gd9SH+oLCxGc1XhLAlMuLxSw3wia3p
uc90MHRI2gMTSR95vJKY3rL/mosvKRuD+ey1tdLD/rAUb45tG8xtcuQGO7oaTBDRE3G54tHTzTkN
PN61R4Uhql+W0d1VuLyF/pORpp/VO8hC2K4d2XQLq8xz+d04V2a5v1Jn+lgKI0f4AgKp/H79HdM1
mIVFULQgPduXm96P6BDlRNL/Y1wI15HE+fj/87/FBxIavP1mAv/1ucYJXx8iN1/EUM6jWPGS5yaf
uCsaN1jUgcmUBn9fa243L2eQQemev2C0S0KZ7CC/Xs3tV/aOhBBk2VdY4/T4cpwQkjKd/G4XkmAd
yzyNWTyTG7wfLcUZ4W6ZeWBg9jlEnPtyRd/jjBNsnc9Y6vYr33gZppXH+gMN/b1/zLQPmZik49fu
L3orlfDamvywCUnWDPY8EznUI6xvbKrKoiHQUpRNvhPyYe4WO2+AWGImfSLk3w9txG2fZAKMF3Py
HBpIHRqeHcjS8t3uBei9SWqy3xT3sTIDuB6Jh2vhm+97uTxlPp6GDoUqXng4FmotJkLnwK+9lS7v
LDLJcRpVBBo4vswZjJ4i9RF5T27s9h4wvDIGl/gGHoQCgPB86jTfysUJU1gXnAw43xlMwXHsPf1R
qnOCzo2AbKQdtP4gaqOGC+/4jhBzE0cXngB4N9goxN1K1LY310rWUbfOptpmw5clyEoZvHnnjoND
8xpvSBghJ3V2TAcqrLUt8WOdiyXW1X1YM7LB9gLVydYYVWoqARaZqrEDAAOv/EaYmaXPYaOP2yRb
gB4TndtpxJC7r7WW2uyoFCajxDGBFW+milCB1GMVFT7nkmwZbJaWoITK154zSm273PXw0bTQYNFX
n1AiKCKMroj0FZcJjumo8141pTJSdt+k4+8KucnxdoXbdlIYalfdtJDnNg4P8vnAThIvpwnpG8RC
dwUR6ZALwYZ6qFHYtf0pRyPXw24TdfxwrF5VFnk2Fk67YZGp5Z4AZWHv4LALEw7MfIeQVIwZE5r9
pi+yk7gb7j0Us+2PZGSmea9szRDbS/ZIUD7b8XVay8nU7Op1bUutHJ/PkWTMHWwCsgZ7Im6XyRuS
kGS1Y2owWTgtCkcwpeDp75JAd88WWMkjjzh+mzAKCn+5XtRh9rrW4va7R+W7BMV9kSVsfbcH9XBT
Wb+u4+oVfBCgmXES3+GLCrd3LFp4cMCrc0d/J28C5utZmyTwHXahHCYeulEGGST43+j2Sa52LfuN
sYWGTSSiX7zg9OoGkGtNHwD4LO9XXcnGGJdeRNUEJgskAms3am7Pkm0l3HmMSmr+9MjG4ATbWJmc
1tPJoai+5fivsheRY04KRbcfe7yNaaT35uYb2teX6bB1VmIF90HuCUS/y9Vz9MNtr2y/JXd8ppUV
DSH0Rm5ppn2nXkVQ0yccSfyUznFBXBzd50GggsTjBI/xrrW3iHEKiCIaTWyV3KYkCFoC4M7mPVp/
O+sPmeL+hJOIAXAg/vjgJV8zfFqN/PURr/tMbMOI28l/S8M+S/bTfycCWi1VmJRYl41Q6akWVF9v
4/ucoHWL5ng6et9pmTcff+hfYXQAPlJDS4YbJoaTnUYDWjGZpMHjgQVtU/Ph9Rvrslojk0UKnQ2A
c6az4XwlMvyPsEHnTRYokhEiUZmFg3Ieq0mroo/kc6xGkGA5p1ffesCtU7cw7Jsj9OhegSL7GckJ
k0K6QqlZsbjuqrZS0RYMitvs+TMQxUj5SZtXJP4z5ZQnbz4nj+fpLpuylGzghiddBqEut86CS9N0
Vgc7DzpPOfnhnHcw4lV/+R1JqAxftFAoej7SfPcPXm2GKRSRTPJN6/5fIizYhx0ZiZjuxX+NSOXY
XT/5odPJPk1AsNHrYmTDtCo0y4NvGZwazKqo6XAHrHKJ6A+THrhnx/uXNKLreGx3tTOSLMOJE6L5
sUQlzKqVR1dc2ZmrKvbObmej6rzY1cDMu6Wva7dnY8IiROvVZtdpJ194BZ6ZyvRj8Ehjz6aGvfle
24oXor/z+hhNxKC5QJyg2t/J1iNHUniLkVDUpgA3X32nsWluzLZwlTcAdBhwMrlK/uncFY2tiBl8
QKW8CFGEnQrL3ML/JiFz7GdtORtF1BPhfGk0Xa1g7E+jDgeSBCchiHDci+gcgdUZDYYfhpgA1M3s
jJd7/P7bML8K0D3YtcLJaCYuB7A+90vvC27v6Tr2Nyf1ZFChOVyKn7jSPb29RwcbK4UuHHuxM9ip
R+NjvTzvlT/R7ugBGNTvoQSlS5Me6CJ9VI4EI5ZN5jdlqK6pyCQU7ycFoNxePvWMkzBPBSJ8jXBv
+0eSIe08nA9uhvk6d1uYOa4eJVxEaVlFHWsuSIV4oJqLXHXwuB3oG1Wz281OQiq00WiCBmHKErb3
/AC0ZOOcc2Mvr+Mb0XfT6eVORimZZWWgAW6YHPzg/3zM36kuB9YzqL/Lay0dO0jPWipRpVPNvYOY
DtFx7WGPFliB6IIHi5XKlW09ET6kYBieuZkNVvQT8UBvoxkTqZ/svJ3ah2TkqP3SsSNs4Kxr4G5k
dMLkiNckNzZEXok/XR0GRsGoajrf162f69gw1jkJ87axR0eJDPCPUOZrxrITASxf6Z9jzsypN87B
hcVr95j9sS+VC2Vg/3qT0RFWQdj0RxI3rbEZpAh/XrJ6jzqy2t/XDwAVllq37+HyggC8D/igfqs3
h3N2pQR0ZbTYergpYXyHEQpRVC4C6pBLhXtWx9OHDj6SetDPqFU6wsAjgC3pgzmfXKUAaJUiKf89
W/GWqJ1Mgp062xrrgGntrNgtOV2bqapy4wJLhFMtIXnXwmrygDM7bicb/8t6u1no393S+xzVzujc
XAjY/F498Cmk/78E90glwGlPCWyoA+6aX9wEEhgjHCiG5KzAuAC0bpdons9JOowKDFrZGNicWWGc
hcGVI2redwm0emJTVehc2QmCnIEQNIS4vd7vskB46SrFvSTEz2svqJn6xjTNxQDOQLxSot9uUfhl
qlkezUsZZvVl1ksTbXkvJZkJigJYvlRxy+VSmin22XKYD2Gktc1qyZdBzGe/PJT5sU1bWvLAf5Ef
AzTWYrffKiUG6/nBZL4sf83oa2b5vg1oqWjjpvM5leV+C9RQ+rb+Xralrorr0MqxUtvBIysnV4fe
kzq0S39ezsAxlUOy69dhLolf/yJjpi6cZSqrcHcS9hJsVnLXQouWQ5pUL+RWBtJvS7H8E/qbLTlZ
RLfqt+PqMOYhwSmYYUPsBsh7LKbtVAWNfRycUxW3NPYbQCSjWXEXao66KZKgWqTahG6Yfiq84g35
Gv0e5ZV766YeK2LZLdg9vf6hlkYTMRYZPDuD20YH7qs5R/11EP1wX5e10/ynS4cVA7BTmMZA0u8y
RknJuK6hRcW6At8v/shGvZsOJ2SKhOgQ7Ghz4Fmft/KgZ9JSH5uf/AkO7d6Xn/Er+MYPRMD6W2Md
/ObUVxFo4KxfwBaSqXSPl3bt7Ii3Deea6edW4TLRzcQqPUoYgwHC/uDcYyNr8pPyVbkIyhRvnuHb
3ukMujqebxRPPQRqBZKOyZ0n+F2pdcoDOuRWFGQ2lVD9uM0eFSHEiM9oA6SUQBObjcIiP1rUlccb
7SJNp+IeAz0Y30udn1pqIDS1tvgzP62Mr+aon/7AhiiBvbZtURxFACUITZDwg09i0+xu4FN6mW5S
sAv9UNKaxO8BsWCO2dJjN1NyKv79zjqr8iRUlWOzBcUEUdlW4XTXFBG3rgcT5aHxOVGb53eO0wHN
Q3qyPhPxtfaYpPC6efriEcErosAyUrduLw/70wXIuOvLUDHiQdb/2Ip4damMA7XeNb5D6iepD4qp
ky4OzJzxgqk9PizLYu33ulpJtoFvBvrsCGFbPx9lilbLYqUr8MX8dRf1vcDvcBCLoYykY7SKCkfg
6brNtnSl2lI3Wu+8I1jtwxHpmr2Kgc2XQrJnVDT7JXVjNB9F85IIvCdGSzalypj+GCxShI7Y5dNA
4KXk9RRyYwOp1TSmLW2FJFaR+be9EFfSUWuiKCIgty/Q5Xll9XHIsE/UcTRiPndrHSFKDq5/4O3o
zpI+R4E8uiplL4Lz+TWh5MFAoqKlQKSFEA90aoZJdSMG65teQehzuuxMkzaP6XPy1IfaEH8pfb1A
qmeqHmUz0bmH4Udvpdve/KCV5Qadj7vQ6Pz4lqic5GJoO3qUVfN0luHOJfkps9ZiXJKphRCG/wY2
5yQY5JNYRavZ0Y7t1+6UQbNdzero9DRKLqr2Rmg6TJJzMZDBLTVwefuZyLPokIIL6dAJPlf6gdnS
zb8oifxy8OxFXgXomvq81xN6Bw+RH4ZRCcZjp/jOsH7ZSo3EEcM7Mwv2bP+7Hhj4MzPGqOsxKzKv
XnajJW91HYIFtOAi0kfj2+yNr7Fyz6xwkB5m9iE6J6wT1IvdfFaHmsoyIcpQPxAU3ATzwZXJFyjT
PzNwC78moO8kapz+wT4ZSDg5eT8sTmvf6dbRMdcmjoOO/97jI6GKTSB81/ApvnmYlvmOXBTSUdqr
TyaQf8QjF5Y0knfKQWIAQFU+NHMIYfzCFHBiwNoDcMHmxXFyeaK+QH3bv9z9VnP7LfAjs+sI0GP5
jrUP4qdRedV/1PKkFJcgKbWtxGExCj64NgElZtnsFcXZKvZgE6XVpKT7FRdba4XUr8XZhHtYOUdf
EPEsXbs3DG8ZH94a0BzhwdAjB4o2JSsbI0zh3tTma0n/K3+zreKFFLUDiRVedVF302cS+rNYWSFb
vQOI8ecLNkM14WPsGO4C5p1D2uVK4tPCoTNSj8a8UpHjEX2XCg/1+xvnBb4tBWst1HUSi54HBlX4
W6np1DSYU8WcSBrlTc2dgNo4KjpJPhbu/5lcqKBr0yeYAB5j6NUKybTZKYhhf06vORvRnve/NDLQ
/69AWlDf+MKLINVVXb1uMkSKdGUJXJ6iPs+H8K30ouersddFKYIP9538QgXOHdNQFik04X6pt0rS
hs1Hm7U/lvp2d4elcvw8V9h6iZP5EUVBWpcDEbbCWpEO97k2Wu5qpVgVrpxzTr0o+tojnmD4VMEZ
gB9NehwUdrnrieZwqyZy2fZ5RImQZjSEK9Jy3WA4bqtcGVc3e0ig3AlhEPjVseuzrIxhaDyRDeNM
uDEiWzfa1nNks2UpReQcYmhSYM0uEnTwqgRSyUfxxnOPPQGPpaj1Mk4BYGSerh37pZ9DfmNbEcRK
GATa4tHXCAp4p7RDe5vLWQgJLp5sViIsXzQwHdHucTLG6HBdmHS6D2X/zX7JWAS3lLSKPIQ0is8R
B5AQ3UqjkhdxTxMBtzBBAOZ1vItqLNr5G0pE1EOa4QCVOSY7CK/KMZjKmq4NrJ4x8tg1zgMSi79d
Tsev7LN8BdEdcuLlEV8u6KTxlda0boxt25bSsYV6RhhKGSOGe+jVzQhFouxJPZt7boRIhhZ7A4jl
cxVWUU0JcJl2BkcFoyqJCMSABqezTmqWFmjRGuMLqmVcTY4JSlzU9Z3WM3eSUAoNrwtKuWkebPph
NQRFYFsx/mKjIrZU250dYDANh5KI21G/jG5sTZGR0oYZe9Q1VDlUJjN8SV9gcxZ+5gzPyUnj9amT
cCZ9NXRgON1GJkBpUc8eX0O6UHtXr+9DHRQs6gFEEHMfo+eQRqrbb39nAeipHrd3xQOZOLl1dl7Q
e91KfmRhN0YDk0d7EGA/73VSI2l9KuSzv92byDA3yezkp9obeN3QLxZ23nq7qIySxmNpkHFr5lG7
o3UkzwhAgOwv/LkVkTOnq9ceMoLpqdZEct3+Tg3b5BceeOokWU7x7dAudaZh7z1xEalC6HYQeF40
E1KMTtdMnAzlhJL1wMREArhz13JIoeshCB4ZQ6UabhaA4quQ3w8V1F0DMHgEUOuBt563bROn5jBt
h3pJeqytZeVgwCwCMlsLEYaOU4ZysjmRV3/7iwoB0Ji7FC1suwomIBJt5ICaz5Y51dBk3rN8YNzE
XpwmZKcoi0bq24QjGQVl9zaiCuCtOvyeUzdTmZBgiC2S5jIB054/WQoILRQ0x4ffspuXtJClrCGz
OuCtxntE8y20kMryunwyMEd6Q+2CWDwG7JDhFajnqwM3MLNJVaWDAMB2EgqRPWZCQ17HTqYYX59P
6J32cqS03/wukrDxSrb8Wwdh1npGKEz014wkdM1+dUrGF9VkJ8QazoX7koPrESLSeOOCNIxrjL92
AonRa3wulvfa+bHXqlyohKEFh8/mGtE1PwtMc6rif2lE3wgYQiBiNGjYMNvGbKdwSsYGqhbyUfoI
rXniYTP4nHloB0xwDi4qWiCNCkroS8ytu+rRG0vA/ozWg2hFwiHRVZ7UID8qLA3+fY3klYR5zRTG
JCCrRQd2HR3lt7ILXipHm2Z0nDEQQq1feD6Mc4i7J3mDQhA+SMtPRYiQJfCErg8WmjM1vG78ItvF
rG/HInAIyheUEBtc93Hbzb+nWNZEtbBZ4W75tVbQH+iyrYgecN2iWUcI+w81UZ7fsXbB3625aDmG
MnQ6ElxZpxIPvwvxlC+39Yb1PxSs1ogo37lWkYtjZ5eMOLtyrVQKU/SWY1BrhOF9yBoD5dd968L4
yFNNkFe79W4oqhIqM2P5y4mI1hbsXYT7H+CYrK0+Fw8vZHCwUH2tsZlR3rDQYG5R8Mm+ycTxx7lc
7AN648QNoxDuYWH/i5nVVMsmyqR+4QQoydexZ4Atfm5sgaHGYwKxmhH/YTC/yDFlbwgdTCk4qobX
RlT7R08/C08z39Iqju0Ex4Evh8t636a4MYik2506FOeQ7f6J5fpZU51SgG3uLin14HbJLVghbiCZ
QA3d9Lqz2e+sopgwO1ghr/dKTCVU+8LAjtoyKMqP44LNlH+AHhxzktr265z8GSlTdBqo8gOv0ydT
Gwjn86DAq/y7T/17M8qw+1LpOeC7rFUq8e0H1gZfGaefReUq4U27y5psfFQrU3enAyE8JCyrmjEI
evIDhEJ2LJISiXYU9E2mmLznLFOXCW7o159HX7FK9vTX15UpHOjcQHKAXxKy0eqf1vFnOpkqYA2n
H4KAjIs45PjRlbFXT1bKX2lcLrw8It9FhHdXCE0UWoLcGd2wrxfj3plEjxMUlGT+mRQfctxyNTeg
YYlZxei641HqYJFfZTLbpx+1LwGAz0zI9fg0hKZOljZr0z4gE3PTRuq7R2NVY2YsLePxv0ctCare
GxNr+QNVJidqrYob6OGPmUQIgo5VQpbCj9dynsgb4IdO9kRf2XnarS5nwAIZ2QZlMRTIpTDYjsyu
LwH+ZIFegjUhivdzWMv5u+B5t9gvXFYbb72SI7YFER8eqUfXEdcds9ZVsbEYNvj7tfvLOZNmNcRU
++zEHah4OLpZcH12tAHjt1uyI0v9w0mqKXyQ4eyl1Zecef0uDBcsd+JJdmTjP2CFVcUZfZZMmpIn
bFJCvHTJdZuuHZOPhb8ZB9dhT0sZw+K+qsFsvF5Pqpzom6+E6sUwW1E5ogqhP2Nvv8m1H05ehXYE
ppa/sVwC7xMRQB784gcJyjgeD66lb6aV9Te0/D1zRJkcZEW4NmHrjq4TE1DD2jhkKdgb+lAfvicy
ZO6WffKslKzhDgddBjCi91/ImsJbUtpSJ01XyI0p6OhAVKh513gwC9zyU12M4CkrmuBAt1FcUPu7
uwIvDBK077lgZBqrpTMIJ53tVMLhDZ5o2iIW3VmwbdseJXNIpftMAWyAt5/QpKDhHSHzhvbFIYnx
gaRLHk2pCN53IHT9y60QMwOnoixi3X/A8lO+jb8HwFSmeA0SQznElEjxyRqPqt92JuAJaIJHr+9s
8O/7VRZw9DGMJHYdBGb2612Yjb+K2oTwprPC8VdkCfhSq1oInQVF6v9b1SmUG9INWKUCFfgXNMRq
pNkFhrDIx+z4fEGpICZsnz+NcZvjSksF5cBAgfMd12rWt46AbhMwo1vE4JFR+5499YYUxwM5ZesL
9mGYT0X616U7RX04q1D84qnDfaHx0jIC1f1162V4q8GJ2vqjTYne3Ztf+rHKq2W3RSFTHuDSS61L
jQrpkMswqCShlF2ialMSdMe+Rezn/z+oKvbxzNY9uDjGa8yM1lZrNZL7oyLWAZNcjLDTsvIFb53Y
7Bfpp3y/7lYhV7IQGAtFFzOvE93dkl+mj8RESU7jryLzYkgab9mRAeT31/eZBp0uo5mdzpmmcxZF
JBZB7OaHCAQ1D9JYsoCJ56KgxFjKBAWc1nWPAcbeT/7YI7YRXIdY1LY44UTfgTkqLTgaCgoNRKNP
jkkE6AoKAJvszLGlHYbgmJ99UO5WclrR0/QeY8hYRBBTlRx7Z/YTbu2Cy89EElTOlh7iQXBUtKBC
sJFdbSN4dsqYLuj7+J7fqOcufoZWih+pJA1jQ0iATmAP+hsGWfgsFsCHITWWBvUifLfnhfMmxtFy
UShoDYntFMjwbDRrWrcwfb5H97ATsFFidrO5p+cct1cz7KNQH4/uhdN41OuZ2663sEG25JBCI4Tj
DPDQtUqQDpkZ3apVIHzPQ2wrQGszkvFNvfLAp/GWe8AvzZm8dUahVqstvzPyzR7E9fL+h4rf4AJu
uq/YKS6wkZvVRhY4lka9nW2bCQCoqRvA4GMORllUvSIcJfGRRqeHassolKu822GDbjK7DRQC2X60
xKSj3CFQZhezZtfNcaBzuTfVlkMEyQLK6nDrnM2/py2lnlnus1tvZoIHkJohoJCzQFRn5+k0Os1C
i3g1R0TVwGf2iP9khMHWqfIroHzsblkmCNXQEqE85wFrDjBoYHF9WUx+Rinc94DYOuRvm76ZeKCt
0vxNu1KLSl5UIfKHIajE+ju7jbuu3lD45r+Ku9xEUmofnwragjvUBm/hP4HGw2fOU8ik46Uj+U7C
sq1QoYLvDRX32HWJxSUU4RhNYBXT2JFQGeruF8kgNzZ+Mc/q2idBw/JR+6LzxiP2AjyJxfA1lN3o
YkuUEs87LkJOOcDmOMpdmBz7VteSX3yUie2l5Abj0GaxND83SHLaVC2wY6fkg+92lZu77Y8Aiq71
JmqUOLx0AwQaxdShY8tDWnB+MbrShN/e5PPQ7bcdtIIwHI83ibeE41JiQOorfWPOr6+8xMFPK1wX
AnPogxMqby8bg+gkQlK9C8akHkKZcioxZF2Dgk4ZFK7z7mVzcMxWMaGbm7YmqvlccL9mSUrSdyVj
M8YP9Z3uW9zvKhacpL4m7URi7OIuojF3ejYdnvhHOAsQDsdyzSEKsuJz83yPt1Ima1nILuu4Fj8Q
4Mw5mZkw5uk3NrekklTbyU89NRgyY4Ig04SkXCkmSgfAjobG64eqqVu8DYWOPfmmzncWFRXugGku
jpWbR+VncWAabayKZiin5SrQMW5ZaMqQSd068t+13R5WAfyJNJER03i3b9gWlPx/cKsihabznpox
rFvy7QDubxnWF2T4HagLutE0yCzeh9IqwdO9OJeBQDL1mLYui8pmtD5H1TIGJxMErltv73lMSDaZ
SHwy3nOwxF1CxaRo5U3VRyghEjYAX2jTm7QufTZphbzBrEdA4qcifHeZSCEYJ1wlr5/Q7G1a8ayH
PSAQow3QThM5d/inn9LpJLAfkx8D73ip/ABEv+U3JyQeUWDTXF1/TSYJdgbmDmxwq7uYHxv0O1Ol
IRZCAfniecWJ1Q1U76KLxKKiqLwy1dwgFyLKI41RrMj4ggVmDvgzERxEgOAXXyDt8BBA3/YJVcw/
CNbQfv1NWZ9Zw1cMLxYeZM4PwEQp+0/PKaTM/ktRn56k7g0EgM5LO/a6i35NvMAOjo9Rfx5PXFEP
VUx7fKY8kAZ64iwsKZpuifKIoWRWfJwqlsOB2LArdtS0d3bfo2VxNV5BWaKHzKVCiqr+YUT5xNs7
E0jAfqkiuuVzbqnqu3RSqQRjengqF/We/xAc6x6z+pA/H1edv/DdqXY/01rJfBvd0pXq+L5RChTE
NzeIEHXbv4ImCTz7Aq/s6DDJLGXPSgaQ/MPl3V17M8Oslo03Loj7ZFy/d46t47SUOwscaPWvy7W6
/dN7GBZuvtvjkmNK5A/mN4GukVxLffAC7pWqJzpDok96rtTMDj3z9Nw0HRSE/j2PSTKuH4Lw2F2U
+xSBVfvAUx/qR/OCW3SQ23MIi+ov6gZtnizgVl8i/siHk9zH0pnWFD5N9n4ujczwkYKMDGlSI7TR
/PAfHjFbm4XkB06YXu8fST/tAbfNNeBg3Lp4BTnKi4PHFEHDG/7eA25z9cxJB5lrsEK4DoEZ1m7R
hek0I/gSbfug5cA33kgnUlG7u2I4G5YKE+YLG7yPCYphDcwaSRBPTbIQkIrotjgEpnoGmNDJq1gm
+CJ/yArZaqqqJWY6uvLD37LuZbmM0MsgmS9ThLbf7aJ4s4UeMk2zIetAkseEHFu/NL4T0VNYBUMZ
2xw9dp8TIP/ho7DQ2tTud4X2FI/UwlnvdBaxeGQc5POAyQWh+RFOJ0+vL8xLj5TOG809oU+dsuNH
j7dXQMWQtJlq1pWvMGJcxUlIhtWW2x4YAYOO1sfLnkJsVQk42cBzdZXn52ny6skR77267M4NfMbl
oHt3xFiA+UERi8IJPiZ7FpG1Tubh3BRLZib66PKL70VqAII1JTavb+YTJbqadwOib1X47ArBHbDC
NFPqVMh0J5h+ZTm58jOMj5OUMBQ5HQkoRlmUYQQLZwsFfDOKcR/WEN/eaUoqS/98Njwv1mis7T9A
AmzydIMsGfN2iNRPPZa9p/MatR0PVaTHPvT48nmmHuJCYfRqdeoP9nKxJbaH78F7J9osjGPRgGcu
VZ6OM1m9o1HX85Y7a9juaE81s/rSnmgkNvU9y9sHKtUWqcK3wGCFQ9FkigNhlKeYJy3UpAx9Ou4I
YpoXTGa1BVpxa0+H8rFZIDE5+qtg0Yda1qV+1neCU7txD0BM+BpL8s2UvtQTbdD2x7fmIoBIfuZr
fyAV0L0Fa41JrN5eLlWhBMQvMocwQoLWQVvmD6/RV63NvZ31wum0v/oXgSGAYzTvRq1IZUPkXt8c
v8wWeDt4kC79jxIYJ17FUYy5hx4vAsuxh4eYF3QIo0fqIM1aFfaO044NMp6TeXJa1HgORFkVkQup
wuWHGwkvLcJ53Rf+kKwKqMyk4zvABO61Yw3j1Bdy+C/da9RCfY0UWfWuezkdwNiAwWmeEc8YDmA4
tSCkYehMe27yUrpe1z/V3AOkM5LCXQHO52wjtBseu1k53ClyCaXxYsSbi9BLO6Y5PNeZuDOt2jWr
SYSMcEJVsMys3y7UYBEzNySsXKncNhiwteS6/+I7kZnxibtgyu+kUEw9DjxaI9Xsw2scjDZYQefA
L3Up0MG2HODVMkSgBcTc47we5AUIZfM2R4epnlh1eghIFN4b3P739lee848BjToBCKwd2J9MUiWm
2TOAntvs/aFMhTJ6yXxGjcWCBxR2eYvyZgpd5v6xLvr+1Tce5KPizLM2E3r3or6ogGs3XatW+yV9
uI16795tvF6JcSyHa1EMwVcAXHaSD6iNhKZrBVxISodyZYd5IdMPexr7o4qqLpz2IEvm0q46EFS7
/Tldl50NPIRZg0/FXxpg3S0JR/ofN0bKRyEFjBip372Jh4Dfx+hwiuk3K1HCxU+T1EWXwvNCelyv
T5yXXHre5PvycQ/ObTSBL3bNd/VelYdXQGKiNQMsRxhS08G23YyDBaKodT1lcciqEd1tovVhNE8G
wVoZ1bTcw/0qtCZ2FDOuqHLgvpR4ql6YtbSnTy6HNkNbI0oBhWDVD5+NDMimPAGvc5bpWkRJElKP
Uh3jaFX9DmMZrRqJYuF6L/Wg8pu9llR/nW67DE945V4ID9DALMS1Jj0sWbI7g+CKGjKKsmR6q77p
mYq3lT5NGr1ZXgAE+ppPQJgJaGPUBgGuIIIV6/xqzlsIXK+NnYpW+bgkVxH6OFJyk1xwswok6PVd
b9Gc7ifn4fGLGQpwr3l07yhykdS88lACFK8GoYig/h5U2qlpjneNd0/xZ0N63raFXRKjiGs2uzCE
6csuxLRXMx01QXXiOkptBetr2Leemv8Lcl1lU5qLz7YbyCGmGNPQgok0O6zwcJSdUCRLeQH5/Ttk
txzyebOrxYhH8akuIwWpVUxpSXGlkSGyTG5WNEqpniz8Swz7svCNZGOS8gXN7tM+1mB+pxjvDGaG
v3P6CBqBv4YpyA2JlwxhaWq7O+8DScQhVMoCvoJNXY7qG5sPpNj/I/+4kh8F5Y3my010QDecWZou
xa5AORDoipJJNovquG7Cy2mFYBFF3QSqdKXXBCek2i5BSyyhxXE10GOifk8HyqKnJYBPHNlPxFWm
5Affd/W6sWN46AwlsfCwXGmbiM//JB+nVuJ1jlq9qgNFPsp7S5ruhE18c/VCezUL24mldeHPqxxU
vhWrYFaVzq7F4EKL29CZ/s00D0vXQNwdeaOH2qZ+CAjsF0CwyF1LrPLwylEHM0xWqVPpp1cocI3V
I1xMblX+6YA/hwTHj85dIpOoTDry4frtyytyCCwZaiYP6eQXSvYtCk61Bd4+028PDpdzKJ6xbecb
SgU5ixAYi1dwGlH0kCIj1uAwhvfgwtfOsqV72Iiu1uCFIEXSJNgazvacY+cnQIfm/FUK3TVmIBaQ
LC0eIeHqtMt/5q7W0hRl0bEyQMwn+sRLmv28tM7vgMLeMw5mnh400CXW6mt/KIw5sY5KNNrpWGC+
4+POf2HweaHyevyXjz3x5VdchIeotDz72A1AzzetL5SY8JewgSogxwFohKYFCPv5PtLHF4IiQZH5
vSEbcUrkbQAYeKsNHM1sPYsr3mJHpQ253GOAbCq/N6grK4CllM2gRpWMDcnrI3jIEDx8yBaclstC
aSQePI7CwnDrCKjl4gU58aLLeZoPjZsSyjgn3BowoBxZXeMOiukABccx94qGqUCo652jGKJhuEVr
xF/PIidwJ6wthoODjMS2tCeKNKMHMQRfC/nZs4lEjkuL4+h267Ra9sVZMf5cHb4oe8U/7cUSDOa+
DYZwH9wPq9qwpB9CUUKe8r0nvRUqAyVpwB/f09cLcu07l4oYroNfIA15zUseE2GS/JQhc2HD/8KV
hAEBEuvxje4cl1Xd+bZDx+3xEScQ72oDtc0koTvTgCgk1M13p+hrHMvLzZcLb5Ux5PJguwIho2Gz
spSxBWc=
`protect end_protected
