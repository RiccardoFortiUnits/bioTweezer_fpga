`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wi06nFKC337Q0c4hgEtRoDvtnLZn89LiZEMk3V/jKNv5dOZjKvnq+AC70skwIlhl
8CrfyrdO3UTD0R4wOBbiZ4bUwL5c99WAQFvCM6CgdmGDDsP2aMS9tMG6mRAz6VQO
RzwcLQChcy0JFI96Rjn0URIbVfsLI/D9RN5NBjMBxfw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2272)
guZMAD7Tg0S/6Fuk1TzUqXvzzIVYGM1Zg+HuIZoqkpQ5URDRToNWVvdAUGfa0TD/
TDG2f/TlUvqhu7dgKLea87tE6RalKcSc3eZcRPqUHKZ0MdtQK5ZOJ0hGbE2jB6s7
ltziS0QJiiRYXYNI+nTFElECph0Y8QW8S+dsUJXsQwPfEZbJAxFCAC+1o5JhwnZk
2ZXRu1fVTeuVAyZPL02BBVv14o77gN5Qgr/EtOB6o6UKguw+TLLMlP8ayZj2/0Rm
3sbxUb/Rowx64Ryq/85nJxYFnKJnckm3B/gMzSqELR6tuhQKNqZJeixikGtidMY2
Q0DGA0TyaWEbhDuU4UV08JR2LNGyB7AomJ7zCH8wflJkBR22ktcU2ZkaO3+HsAZm
p2DdIxheqgsf0C/ki+tdQXE7VcFOE9xXq5Cd2A5oYQA5Aw18NRjpN+KVlNrNAkjz
qLafZxNsdnJCu2W7ECdllr603ER96sZOS0miIZi1PsNTsVMpV9D2XyAtuwHUXNA5
XsbR6hzdcNh5l5D1nM2yhsQBU/5VsCVlDrCngYetPhRIo49cfMakhgwgYMIokEqI
P6eK8SN0AhfXSJzvCpxzRxdHFIepkjnuYMQniJNa/oRUP8J+cojUpsTATzr3xiZ4
MAtF7l9czLmj/r55khJbw7i6v0CV4uku4j2yb/6upbEAHqSaLS3ydoIhZKA2vA3H
cNZFpSxIfidtqyPwURI6tN1AjftBjJC57r+Tmdf4nMVItk4z6IWSeAKInvV9aj6p
S5vAcA/6pTfUEzJVJhbKf50fUAWQ1pJXeVnszi/qFan5jB9XoWE9oFNWh4198KWI
3XNhDs4SzVOiJtpsEExke9zdElHl9UIrShH73lG8e+zItzKsyDjXiEzLilFEIFpz
TNGusV5mfvQRp5uLKL90FrkYElTAJVQhOLZr/qHSJDk70hBaCFiwdnP7T8kLacVe
b/sB7g1l7fRcntUAU3nW+yzBdnQVyU7S2f5a5y0pXSzng4MMPw84DXcf8QbOmo7C
NbTcVQOoQA3+I8JVSGdEiLojNJZOhonAgSN9JTwIuEd3AkX2xuxCXtSshzaSG1TF
kG3NyARn6I2Eevo7Ejhh2TkS0t6iyZpHAwHmhOFXzPHy1RBv9Ccl4JWxfE/6xEaG
5vqrg5nvM3lQS7Ew2ceV1hJ31SDVv4E8meStiYXDCyyGaYPhHikKALB0YYyOn1Vh
Hkq3dLtU0aUOg1WBn+bZIXEDbuJbvt/deuFWf+An02iSDJV4y+cZyvmK5ka6ykpi
oJX7V4/VU9O3TzWs64Y8lSi1ilp+3zlqxEB1bQoSbJWDM7+2tfGRn0K39HBC7o8z
R1XZ4BSbqQL4qqpoUqn5Or8KUfUkYWB4Fm5YQQgc1AmcXfStZ0JJErOoqCsidan5
66zNv/HtHO1Og+vRLn0rmfb8R8MQ0StpMFAu+04GefpjEcs9TQES0JBt2mF0NJy1
Z4jaYrKqEY08ICYWwPPULoV6BOfYT1wNC3+u7hnJBNAwDOOz2inxrVPGRZhfLNHz
uWekF/Fgoa9618A5W22ucqd8pM847dn3l689zyajYOEOIUTMbZUekXBjLXJugHev
oFPLx8/RbT7NRPLU/qJWAoysLhlFjo2ZOFYcTdtP6V6nbFintzrhOvQNND27U/5r
Hd9BBiJdC/x6wKpbMMRLMlPhG91nRg0oYzCZL3ysG5HjoYqQ/vgTZJWxlkXQB4KT
v0/4Vg19OFfNabJXPwd2M6NLhB1bvGkM206krDuVttDyYOnGIlooAB152xYMDc8t
0gw/Bvi3ycRd+lTgrZCutfoI5AKI6C6KzBQx2G8RdPcuuubwD+GkLQzHqb7e+3im
9FjPHrYiEiXRBmGOpm1mPD3HQJIAvB7cTuE3VuyH76scIUFriAWQsLkvw56XspIw
SvWJ1T/kzq3aZjVVL6ePn/kZZ2Epr/zTGe/JQZsFe+4dxEmcs0EQZO3vOVszGBcv
HtG/JyqlIrVVSNKNZRcnDy8PdS18vfVjbGPe+g+6sGrbGWBbOmp9CwSQcn/fzyrd
P77psLnsJNy9ZVv3+G6BmoySeeYtVqzMGtRAaiHfDJEmprSEGJSVgayAEfL6Vjdm
PtBCaDMJaGK049VWBwYFOHjw+k2BCFR96G3KMtYE3FMf7ne5tgFvv0a6k+BZivYD
IhXQiyK4fia/PrrlzpyioHTcyg4sM9dMJ+erylt+QK9ihvtAc+iOTfNMptrXFq5m
k7DjQBp2oX47C9j4ghurYIvlzuM2cL+v/z00qfK13MKZNRkEL3B1gq+CgzXNE2fa
X+wswD5OuycEJPiXABuaDlYUWZoJZKmW0llAkkYsfssnUnAY7LfYUSqSfEttTrXX
wUpbGWBVTj/WJObrmD8v3S9ngxlBtEViExTHGOnTsmdO6roHN2o4XRGIHxG/kNba
tMNwLNaaM9GbZVFHaAdSYneq2L6mZbW3fqcB6fMjvvN8fEgn4wAM0wEOpur58MAA
BFMkp+K5mbw/KIYRYTRS6Vl91QL6LdRd+FVtif/KRevA8aA1d8H12Hj1gIp94F7/
w2Pzdbj7DQxiU5YdnOGaa+pAIT34rhOneWzqj9+Z0vY2CNCRLSfX0vIX0t1MdZZ0
qhOj7QuBHTAVKrcN4+p6zQ8ldWQsf0RVpqJVrbqBFJyAE7qTu5UYuCuUs8XQHaYk
jA8a/xQfm8StFCcvApzM9n/NKS7EMG3DsZq08otCUK9kwE3lTnmKrBep4iVq8W5H
klEK5q8wQhjUYvzh5sJprBdZd+LWD+n5vMdsmLnufNLvjQX6jOE2r6vR6/YLJv9J
XvHQZcH2YSHtJmipi2WFs7C6AMlrsYMBDw68wm2iVEN5PZL3k1UWH50Ch7GjMw54
dsWPonErEMoTNn0/gWfLH0WdwYNkzZQO2iSp9ATSonW9ieN6kpLQ1Nb09OF3K12n
dpkR4/z7EiApLlX2P6UeJig4ZSS1iEY5pcwwVC6dsX+f2gsf0GIvmFHjfREMDdUs
GGXV9ulzxtCVFGJfl+t15g==
`pragma protect end_protected
