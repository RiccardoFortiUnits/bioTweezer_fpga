// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
K3jWxAur9dwK65w+MTl31zcOVuPvXybn1A9Lq1qNxHQ1y49IDakOrSbSfPSpo7hFJ4l0xDqUkWo/
Ibsq2XF6xyv41pcCY2fAmJyOWJEmM/ZR/1ofgbW5CBQd6EzVYWLz4NvIVAphDDYp3rc8FM7sXUTz
jSq6u5hYS4e6wV6yP6Tm2ZqdUmOjIpPcw3JiCPpCZSmcPcIXA2vJ3QVzwYC/rLCJhOBivka0l3JN
yzUwHfUp2ynv4wkdWXkt3yJCwRDLfI89glz6OCyOL20r1fpRMiDSUUCLImocN37p3AebxxY4+4CM
KZ8U1zY8ztJQiVlsJA0chRu/bYdKarg4Dd+sDg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 1984)
cIg5TBr5lvwVRsji0bO1HjcUN3+v0XV3kUV7ef6rCJKfRPczk9OEa+LR0RS3sBoUCKgAIVLKb3u5
w063JZ0E2sw6++u1PMvuRx4wwPLgqgkHHtH51Gr+LtX64YwqQAY4FqJaNZmsfgqZHPPDioRsm8Cu
rsGdQ9hONxVyEZrJgrOtr6p5Kl+fX0CG0d92wO6BTZCvcg2dBZcYzAJRNIJQTZK4zOcqre6cE61C
qeb5HUhv/gjeqRNl33pclUDpcDucvhzFMYbdpsaDGYVuERoi9RjnYNGtjf5eEay3I5PTCfkrdNGc
c1nCu9gU26l/P4yJ8SR5AsBRW5X7OycJGacciApunRT69cSPcPa47wkJ1oMpff1mUff8Nz8LEemS
ZeXt/ADlvgKGbFCjyTe2yXavlXcWIGA6/s7oFOFobtpSIrbvbPp+2qOzz1iLcg8OryKmZmtcFpPm
KgypHra2fQD+vulDH2Qlb2e6i0xH9Jcl4BTrU5wkYL8Hy4JrAlFDK55dVaiWTaxlo/HkFolxZ/Z+
cdA8jbDChTCqslfTMAjcJXbysrYtq6pEyMS9Sm7yMmtrrredA0YZZuhniLibkzcuUDSIk8aKBAI0
3Qkxp3ZsOkM+OaNAdZac4ZHoVawtMHq7Fd3h034YvZZ5Q9ECBNrD9WjJlJw8KAnTp3epX3RTV55g
pXlhCvBOshWG/BG+Zx1mru62Un7Yg1OR+Y1YclOu4aZ3DMASwSB0Xh4zWGWwlxO9jbZec9eDx206
e0gg6P/ObDpWvb8VkUmvLTu9f50bc4DNzIMGcII5+VGd3ioLFLy33JjWInY8a9ZDNuUuvTc9fUtJ
CIcUDFA6U2iW3knFUizeF7WGHwJBRrYT7Qf1PkRl3U9mDIASEcjz8tNuBJo0pLuc1GyPGNQl2B8E
3Jn+U89AOZZuW6QvWd0ULX2a1rH2OtQIabJJZbH7jinmZrYLqlVZ39csPDmYWDT9JvODvO3vSAA5
xVhWFFUcpWqhGrBFqw+ikTJ4K1cUO3IQa9LZaYXPwLnPbGN9IdLhIcThLWDdZ29RPkVGPMF0T09W
bbU6RaBPnsLOwiVydxXhR5lPCK2Cxrmukk33FIYkb6u2pJFXi4XZew4bKJPQYzVFlAJrFzSauafV
w41nF48HnerDZ6lNB8vOgxNOKSbH+8tSSCYV6WrIOUqEDjg3XUKsHnML+6K8fxvvUoffaOYbBRBL
X82chxCTbLBQvfaj3x94EK2VBZAmkM0jZYxGG4R/VXmBQG+GGmDO54flqoXQ3hecp6rLrVHxwH/Y
7WyiiJ7q5PmW17qRWBRK+W9y17XdMlK+QHX13y5AELwX+GKPozHCFMaspUK4/Pmh71Gm4oLGN94I
LD0Fo4dTWl5EJNoUzw9zW+7UCQ7swJcklBNV7IcM9CIx4tQ5VMvLx2PJAzm/G1w8wlU/P3RHTLGb
wxu/tsrHHKQmGOEAp19uXxA0fNmlOwgJhqQi0NooZHabL6kmCwaeRowjca5CHb5GqoMoNF9RrmwP
Ag3mezpN/SUXxpkLE8ZJFRQuJRxK6rmU3gTGsKLue7/HBg6hMZSTwa7n8IX6nbNeN92FQI9QOBS4
yKw/5V/og4SxdpX9wqTRvnx3cTE9l3eAZqR74B+rXiOwqxhrYVo71bNVo1OApm99/y7lufvXanAz
vw1dtBCITcpqeXHq9p43D3xCqDZ2+ayFwP6JTvhhkj8kSQzDkS2ZQmiXYqywCXReSRUI7GUTWj6E
KTvhjGbxBN2J8fWkLrvzfjOhm4uyIQ1RFMOLBq8zeSXERrMsoeZ07j4XfGjnUvgx17vhb01DDxwa
8Na6Yi5e9zkX/Ykrcjw2zvLA7gc4bkM7vG7ToSJNtYhyh4dWZIZNhg+sHp2RKij7NIlIdzgv6w1y
g7RrIO4oZwldF9iXhRk/m0yNzEE6a/0HOj3Y7BWt2bvOYxlX5nO4bW1qlWt9zrggOuaIZ79uE1Fm
GamiuM0eXL2VMB/W8/8bKplFqpUPdyLYf4MptOlUUCy/R1KIIHI4O5vEfD1Lu4tSD1Pmbr708ns1
iJdsrrjP3gNhia+XDbq62xupiPJzew4H7CMv3A+jhTXjXS3xix7mTYcf66cgzuD5e7Qt7l0zhfMx
/aqiReE6bh83IL91wU3lSiRcKFAYzIp5gzSDk2MDCRXlD81Fod41GVuGLImZIV4fn99JkaSAxN2N
laK2YWkRwhewy8QI6djg1UGLtASa9vDdN62muuNyucReTRxsbp/tE4hl4dOHdJm7YDa99F7pyj+M
BRt0IHIoblfOJeUhVtVFFaXO6dVkbCYS6st1E1tQ+0YKjYBmRrvqZ9uOSxndiZoxSCElnzBQHKvE
39fUpa4dUlsY/ilmzVVFZ+er41yOgyLrDQ7cX7ajGwEaxhg6sRxxBkb4Vq862UlfD1yNiOrKYscW
FvqUa2w/JqU1zEwC+y5IicezvvGLMDvsWYLqPHNuoA7uzTroeqBD2plqD4Pi6flhJuQI+H3KNgWo
HrJUN7GzdQk8L+D6vaDZJFHsC/ugPW120tzABxrRCdNpu4TLlQurrIN64HO237lX/PI0qbsk/QgD
UXi6tG28zGVQbqmFH1KfyLeKy19cugG8apGcrJHjs19rar3aWB/CWSyaKDlcpA==
`pragma protect end_protected
