`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ahFxujeSos5SlWAkomFvE/etRLAiBJAV71uqCWCf8JiLDM5yt7BvxWiZ0uqYGzEv
zTbzZueYqqiJv60kT+7y6wNR+1Y6xb3uZxIVEhQA2WAMAXa7w9x8CuF3ZaORV7/X
qPIFllk1ZP5T61EgOFkEdkOFQHA6GkdO0sSKdRR6zT4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9536)
plCdGZvn27K0alPCRIel1LuMejYr1V/cnclYlyY//APIyGJL0GPUTZ/vc2AQKU0A
lAwYrNIg4eLq6nxLwnNPIVK2WuzWYrEc+dwlo+BqknWV35F7OCr/p2ITXey+hwY4
xBmtlzIF5GivBWJsonMjHzvsmrw2p8gXgjVZ6+4D3nT/7MZ70/oAziV+u0dgoFPh
7T318FaihpMrOjMAPkzFn33ztOkm0hKPdaYpSN5q51l/O1n0cmSMY18iDASOCDkv
Yh5QqL0QwCJQrU8J6Colqj/4glAF2X/RIRPz5WEjQz4QVLLwjSV+r2h+nK10IDjF
uzMatPdKFowWmu6ImJKplgTpYmjskrGMPS1UOKq6waU9mYuHvMwexife5F7mQlXK
Mm7hT/jgOjE3NrkJ5IbElvFAHRFpTXiwruR0X57bQjpV0FH+84BN3k5fmvwmvqSR
yTDxJQzl/WvtpafL0Ma7jDH0bdQYJjE2Z0hkrTUZX1taTNtSpZpLptmP6LDOqk7k
Eh75B6nnFlbrnGnMujhtmM/vto+CfMHuPLoIQwnTUe3hkcpEjjdHhaD1G/VCi7Uv
kBEiLmde2jYmoezlBkQVwSsBfNwTiRIbNuuJIso2eufbwm1KP7uJRm4li0nRYIlR
VGMq/FKBARCo/sg8+t/fwtELjxRa7ZbRxtPcxAadzr86nTJ5ENpJ/yJRmeTNaT0O
YuF5XWiDfthm23ylW9QGz00DOeTaA6VcEbkN75NmAGkG02cTsqCP1WkqEOajwULr
6J+Y9mvsTz9oKdVA55zyl4s2ykuYhy90e9xiyvunnycyOqi1S60NAU/5TulzuN5n
yMxaxeAJQD5uJsqNNoEX06AxdrogWIvlIkydneFhvpDPu2v3SxuP0trdK/srnI8/
LqW9oz0EQNaHS1N6S2H7EOWaeKW4z4qN/YY54lTIysjQt+y6J8Ru0JHhJ9kiHk/O
RtyFyeatMMBZRLNXZk8AreLAUpsIcmQySURcx+LLpKSdWseymwdMH9/2LQhjQPii
xJGj2a+AYXRtVDtytHIWlm/el19RMIBPD5RUXpBWTYB3wMYvNGx0ptgn84sZzeZT
80IuyqcSTeAWhF/8wdpy1V+7PclzkCyoK0ojSWAq9rV8B3CS/5h9jMaMb9//6VjV
PQGp3gFjA0T/7h1Fikf76PT+TH9BS0QL6KjIxZKtUa2nS0JN2VcMxbXE8pfTjVVm
xAI3mLABL4EGgZYH6ZiX3uEVx1/jurb6Y54+kmfu35htmFZjdikLk9HNnr736JIS
EAS6y13kOohh6Wnv4ccV87uAHIzr3RZgmbj75L+8cbdAV+WkBRm6qznXQhfGCTbB
tX81LBt1HenlF6YUPu7kteW9Cd+qWeqOLSnPUGys0AXZGj7n2LHnHGvpClpOEUaF
cR5uJY5Q+96pZXIB0qOOIdijhgaK4kW4zdSzxP7FF/NaYl/pbpHfP19vzhHIx24d
b60mBiePqxRjjbmuOdbQgCNlgWxcJ1oFYmsfSGbbSSvWi9SC7ktegiTtoW13Z7Xx
XSEL4rbd/8ZSNpS3Nir12LrxKHOeL261kewdTVGpq3jhEvropS7qnw6BICeqncfU
6EN3eb55ZHRSsjwLeMDo7BfSBwr0HJqnRZawPyzz/apgMFx4cSNc4vp030Dh+o5y
kO715N0gbNX6Lv6FK6WLIiqlFNhdQuptaGj5KUcpwHZhlDr70oPcDAzKBHkM0tgv
JwEDXYh303IeKX/CIJ2919G8AX0Rob/ek6BX08oaklBPm5NCh//Frk/gob31907k
FM3E4ktJvM9Kc9iufJcwPWB1FsmjoMIavjway4+23VLNH9NZa4T7tRWfZ0LlLc9/
AX4lHNVIIjs3mNkm6mFXk48JKCtwoE+Qel5vMKoB5vurEfmDoYQryElMayCy3EqR
gJqQcJ0tsdIYsjFaQ+qJB0n4sxnVpX3pznE7WSZ/BC2aNQqTZZYXlBDIzIGHyIKJ
uK01ZV3Q8MpRChggfYZkZAoXS+6TWd1ErcAjMp76Yosqdl3xDqNrCqGsflNsohob
MyAfhYJFS4ULP7qjjpGpwTYYzecR2e7n4Hqr92vMeMtVu/QuVxy5ulbWHUjoEueV
3rnKUGukOrJwoK8dLdIbqPXz8i732pZrDlE/SzlVUePuqzPR427gId2gn0d/1ITQ
p74o2nWj3AWUrgk2bNegxJFMgdMrPYsNEn8bb4CciSgG2wSWPWIPh/t+U8uZYm1E
1vHremEH6/iNr0mE8Akp8C7ckIlf/0Z4IU8NVKJtsGw4CywMcplk7CYDrtDs5HPs
18uf3lH/D6wV70choxA8xmFgqtvnQb1CD7WhkvpKuS5PBA8HX9/BfKLbBBNVML39
Qr+q75oSBLRbdrsIqy8MywMIlCUzSFG8M2InCOTqV0KNm1WyOf0gjRvFNYvGNbNP
c8gJQuNoE4zDYr9KAH/21E+eeJ+6zhs/YtjGOlmZlY0a0kMNHtgmMZzawnnegCCJ
x5TwA/dGCSZHQqgMyKCrhxU1FDyBmpcMTuqFbmi7mjbJUs+4MLOiEg7HHvd/pZj7
e2RVuK7koNG2fxycQB+nlwUeapiYeLJD6PZ3gytOralDMSBW4UWDuUzTtmE/CPPP
Xexfh71GFGuy6eR3v5TFg5cJOHJ+Vo4aB1eTWacyJtRoQGP5rGPTCQev0mvd6ZX+
BKVBNNdBhhSFe4IkuL04nF2GnvyTeKi5ZJWeSPoFDHRdM5+iTgN65JciTZ+0J65A
c1o4D7AnB+cNcKsoT4PIhrA1FUznXZJFC+QTPJfOW1rfUoXXFLFc2mYc0ACEpoqH
S2Hwu0DUzZx0yhzhCG1s/7m4zSiFufVwQwXTGoR8L6KtYyMT4DwwCT7Fmyoy1+nj
T9w0R6zOzzJN+cRwRAeY76jNhJgqBdx4PGmJCEA2PHsveeW11BtLFw6ag57z7pi6
TzGX5No3g/vTqtl3ATL6cUg0njc/IHKasUk0zhSaVUgqIc9sirl74+67KzUSWZ+4
UGsj9pLmricLU9frJaC69yGEed2aJJKWhz2jXO4qFU2eo3E44gROChUSqZKxH0dZ
9V0kXHovFyeXxZJAXafN777n0XwOGdLwEr998lmcQ05BsKC7jIS6/TvsXlrNo6q4
o8ebfEhrWfSS+WkiuzXP17RKKmgsuoBDxf0TqjXnxaKiWJw7fp85Oc0F6gnzrNXl
nuYMxKmN1x1jsLFTFyfEYc/NDwMQYJswCYzNOv7UHG7eqVDvDhqDlchw7PFjFH5v
a1FVLmEyGmOjQmKPEZlBXjKh34moMxA5+xpCIyKx8kNX/OlRYkYz3INKD0TjMPGU
35uke9ZH7zYHkuv92/Bqg5pDtYKEO20Nu7CkoyjR4AjYwRaaP2HbS+Fr9j5crsft
BQW24E90IAO1/YKZq1xP2zBAzbqjdwx3lN/DK43RixLFdvaP41CpfxCqWMU5mqHn
d+SVANpYWSTgwL/eLcaO3goNGDwJi6djaPNLxFmgNIUzlYZFsfjReZKptahADKwm
x6Vtu5e/3dy1NalC69hIvRYNpKv3WKlrf1q/jlx7aWc0AKDkRXTrXHp8qYNUBG3N
ZGyIBuU1+vB3q/0GtE2ybNit8JDnDLcYTv5co/ITQIm/fJiU5XqEfJPpv2CeB8Nd
N7A6VAz/ltKTUiVH2fxsUbWOjVqTsIupCT51djNheb8E4/6+xinQqlxPFbzhoBlU
b4nevLUBjDLMoUidb4ezyJS5mBko2wjBvh9O5sz5J2I3bo3eFCS9VLum28Q4cusd
lRKji7rRn7xghgogNFV5pTqY4MKenqfhhtd3LIfeCCP+BEGY+mms5tgyEDV39lou
bmNzHynhoyQIOEqMn0cQyfnhu2pNp64chR7x3JkEmFYIkrF3jVoWEUAw7LSqIqQb
zk7BKjYpgfyVXe9XQfp3DGeQNdnGfIgQMX96aNqO4JDxxJFHW0PSsz3nTcS7p+po
j2yNJ1SkMiTHeVM4EzF7eWE4S0qcYNJ750Y5tGCy1paYQlGKDAooJwSu5xLGgBbp
380nKNRMT3y6iTQ3uTPolbubHLB/5DZ4ZiKDb0QWw6mkt0iH8w7SzepzwNlVw1FV
XtCrK3dpGawHvSC7Bd34VzNy7Jqr1JiW4/okCMKnwCY2FFE6x9A9G5Iuh+CBrfbR
kjR+2Zl3opuYmvmFXwMVQdGXU/5FOibPoA06Ed7SM4XQJU54+nINJXCma0CNMj85
kjfC00BfRDU0/fqeStwkaHaRAw0+3qjp9mbdmDj++WnxzfDqW2i9hPtNXl/LSWa2
ztwGyLsHrO//q0F5bqrzoEY/0rHkuzfQqEPrsC74t0CblBOYrT7/dsojhK3I4mlf
Tyvb4UgigeS0yI9E7ArVXknB85EbDUMTGys3Zg1fUbMHoeR+QMOx7BPGlMm+HuoJ
8BNZ+1ux7Lo/HlFOsj1bU3NTFOU9LPR/E3L/GTrJ8s9xg7q/OqEm4whJeA0eW6DR
wXC5RYLh/7am/ZCEapPZ1QzLOt0ZDOeKlmv3IqLrYOi8P/5FNlAFw7GZAhy7MO+M
UoZCbowOmKCqMfP4cduXDyxnu9Oo+i7jOXCV6ipulFoYnmUl/CefzwqQoZv/Kwza
fhFF/5FnCUwt80xtfwTj+TKsTsKeq9f9Z3r7MXekiPe0AJ+MrVcDtqWi/XjggxAC
RsxyHNokSxw1tOeiPcgWP7fxt6z1NfQHwNy2StsZlluAGbSVJVJBJ/7BBNVxA726
jiRd1ZnCadkd1ZVL1tz26atWIYRvUG8GAis33tEvOyTCEmdL07X3J4NE0+ezvJ4Q
ErDeHzhJ/WrZT2XCIPGLBFKolE1TcbZ55R3CicC06Xq7pV/Z8B0rU8SEKEJMvSi2
ahhkJmMEHbqDmnaxbtGm0jguVTbKafj4op+hJbN0+pJQ2A9ASUJ6m7vjOb5FknCa
qB+7eQDYb6Ml/3+Nn1ycRnW+LNIBF+g6PKwXC9J9Kw8Y7+07IPozk12fjSQxj0EP
bvxDkEYRoVdf3hLRTPXlqXITgQYKZVfFZqykyOJU5pxFt+2spycg6WpkSfhpZVFf
xfjXZp6CBFi8GcjK9B3sq9q3aFblPBq6r5qZhQuElhz3kkFUUo8s8MJJ4jkjhwoW
DbMnVU2OFDlm/apObmYGhok968viR9uZlng/3S6v5rzzmMdtLlSn3KzcWxIkjCmz
P7AQp3AA03UnrWv75/9z6zttyq+T2q53cGGGTWN3nFO7PVOyzhIbOmY3uHIKF2W+
1CWydiw9UW3yLOaTXOq/BZchGY6uFrSs3pxpvtKFHWmLlKbhV9YMMv8winzII/9C
ef1TkiVcUEXiMGoJsP1Y79cRP4ukjDMVl/kmWFPataScRoRA/q5+l9JmVvpla1PM
OwbX1D5I6IIqtTHDNwK/8DOfSdlhAbY5Ru8ctEbr4s3daqWS30YNxPkj8gVg4YBa
gVTWXY8YpeYzvgeLJRbWhRYewdaZsHZNQ5Rx8cJRQgAqa/aCCYetcL7caX81nuyr
L8euOVTfuOe7TSWSEworYSAEMRtydI4rTXlcNEQSpfzqW/2MmGb/NWXYvHIftX3L
vBufrJSRgal13jC9HpubuHkqLDxZkTaOV3tI6HpinF60fqdhonAoC82dKH6EAKkr
Fn3dKhmbdYJmwsBQiffdRfrl/o5djFBmKGg5mOpeID2Pthi4R0efffCp4dDJRqT8
cN7ed3TKRfRHCs4NNAYrS3jvs8kVBUcIYO93pPSMTaTRyiGzYoih1LZEaKWu/4DN
rLd+GPoFGfSalZ3484P+AtFppwPR3dP8OOpeBsirefhBSLZ6i7s/zjOl79Rw8LZ1
S8ZwNx26ktOaqceVCLm7YcqKJ3j6TYy3RNaXQlp5IidTc3Gkq3HwmaOCvv1432FD
6Zj8AbJ9pxV/a1ISJbmY2H/xGztb0tiA3o4U+ALZYSlNXXa8oWJEgPgT4mnFTXqT
dUKVDPjDY08YTwdB+zKhb1b43a18wjlU8rBWv9sK/w2wWDwEODE9qvrYyImRBexk
GH4ZL7tb4Yb+G6FqkQkyfhtisTy7jwC2QOhzLatcIZWDGrLHvm/PM90Yp3E2XUS3
dq6eTf06Ej+5WLPirWPO+jTB6yDxk2vW+48Eu1aXhh76osx0pt3HdpmCyiUstYEN
YH8t5S6CHA9n82D6WC+QIVbx40y87urI2kTbfq4CFNpWfC+Z2MQsmYGOWlchzg2O
wFIIiIZN6ka02bMOH/ziytLpaYUlowG10050vM3L/U7Tuc9ucCWJqvBB4fqenoZF
A5olsQ4mgtQ8nLFR6yFCxypnWt+ax+dep7i43JSTc9xtmUklqH5JJp4BsN1+Hv36
CxnvblCtamEfR7hOiI4SscK0RQMD+nZzv/6rsfo9zL8xSOsEs594GRfRlCDbuMi3
Z8vDeQSO6WbYzG91DCb6eFWO4yfp+YrkoZc5Wb2bTMR3mrrD5/AMjsszZlwG+AFH
XrH+ka4yzg+Nz6sHGS3vOV0tQBtps6yRnoIgIMcRmXJCUW26spwjm/YqB/V8Ad3j
HeAb/TxTRqEvnAieiv1JcmGpjxgbKulo592H7YNPMyDv5xRIrUPfvk6F00O1e34j
CJ3jvRDU4JZ5tfaxvzR3YILiHob7rdO0gEH/XPygCjtIkJgshuQ40ZT8yqXnG0nL
K0cbPgqWVOpXPqbYD32lgTsvaBqC/zFIxXpiwVe5TJeo2uIcZdhYGsd0UmynQWy6
Iki1AtSxneTKsrxk2pVj/SwVTkzvMNF19iYiOdKShqU7VPurhoq0kyYKVWW8q+Ys
Q07oPbIWkgzqA/Z9e7gg3MKNFwaIOXQPZzuiYGk/mN2VxrBzUuB7ZDa2GIUrhokl
n92DNI6ChOM2aNv2SyXqQVVzs/lLS059lcfn9DZs+U/hNgU3XCAd0HfBl2hN9fMJ
dxG9wGOBWRPid5Ohk4c5dLXA6rTDY7oHm3I/M0SRyNLL0eKu4+DUgf/5vK3vmZXJ
/TcKP0vlQyyjqkTBoHoCDBdmOSMIy56xcC+esgc6IMtDopXWugl9vmehenr0RUOY
M0S7DAbqA2tCfKEJmPMw0jcx5Fkr21k073z+G/3RumN8iEjTvDwLSg8lJeffxgdR
s87Wx9Yy0SOcqlOHINEgVbPdDgt5hi9bZRydxlATJz8V4rB/yduiwag0K9gB29s4
5Pd0Fmu0QNNSwyKpHxZ0wXOHQRl2x3bPhwktuaUAs8DhLIQQPoCEhwjG6YTXLOqb
vHs9wNqXcjKL4Hnx7QDujnNRNWguWQZ0m0pgP/rjPrwOM/eXtsp/2a1yUJf5z96a
mY6wKZ1rENRi/Zl1NAfMcF9lI0pW/3d+r4p7pEU6OyYKEq0iZZa/MBeRjnAPQ2ya
tHebI4yTSh3i29oZDqxfQ9H87tEtNo9UCiAB4vXf+fuM9lJQRr5SIiYvcpzeGt24
uL6hYl+pY040tSCWVSltlkygwmTpPZ7779HkkTE+iB02OkS+zMzggs+fdzCyzy5d
To1U9ifi4J3AUv/n6QS20FzDO3ZZcmZXxHbMwh6PXBVtqHP9v25q85Sf8JrxCnSy
o4GAFapztNLDbahrSThfF1Wo1BPlWBHknQF42chvh9KKpz3J49vTZflwwoKk2G5B
qCf7+lFm0e2XRE27HalhXV/n7CUNbLS8xcAAfdopFsCGDqq4HeBqrpNvStTuHnQZ
g+N1OYbcKRDUS00X0zmy+yfcpp0Y+3Ono7jrRNPl+SNSKk5jMAqOeJG1agbvZaQt
4KgPmb3nXPEX+2TWTuX7qhzNekoN+lzbSs/RFaAR8yzu2dY+NAPdK9ZqjMLtYGzQ
2yqtS9t20qsIG0y4CsiCmPuYjmT7sL4oaqB495zgNIZ13G5TXJZAx5DmDL1K6C3/
BQ3Cb6BBJd83YeeEYjo6Ga5JNLrsB95RMZsBQFn+zQBk5I7cyo+cBJzENugDN8cO
KX38O3w3KYhG2E6WJvEbImQ21YhCbsXSMOi95g7fQn3ScYagpYzrSTfzqG5lyreI
6nwLUC/Q69AD/HTYImjMTKHAuxCkkSfL7PBJ82k7aNoXEEXxUyTptnzWaqTMQ4+8
upflCSZVw3S/3YJqs5TEmWxMVSQu6mlB/ssrSFWxeGWT7grkxJ2KPDlOeZAarOoL
yt3c8mq56fxMm7Wb4PHc9y9lj7s2PkvcD7rIuv9MDQQor1iqj55RVzrPmy6ThmTr
ncbHatSbj9GywDWVn0H6rrNzVxKaqov15DS1CFHV4HerwrHpCHvfqDATqy/bXUfu
uJO7c4PYOu/0A4j/m178oYjTLT/WYQgU5zJnhrEFR/SC1Lode88qkgR/Nh3Akcw7
2DRkc9QISyi0WAsRvLO8+L/RM40p/Ogf5C0pAnugz4f15AIaJ4aWm7ELllQtshMR
3QXsUj1vd4KLz5GE/1btdnT8whYIfNkHELu1YBu+bOC1EvWX/AO4+3NwD0hdfXLM
5kcL/wtYovhKSEbeiycKELDSuCpT2BUDmhfP6wYlZtHsiS420lcJgBqJEupV+Iq6
7zKBbAA4a2HO6M9i/9q092RMpu622jb4Gx631zmrRrRloQN2EZlB0V5SZLitkhx5
R2vUB57Siz+/N7P/G9u0+c/e3qHvcub3xTP3x681DJwLrBUpKo6oLlu22VLDioBO
4oWt4PukWJA/R8X4FbZomhyN2m8rkXgSPHvhe6ir2qXP5ho9Btw08C/Ekq0/j/bu
PnoOgCqwhDdIO6oHcYpdd2qj7/8Vx+HG7NesJt+gQjIyfmk1nbCdc+twednq/R75
PcBIpjp91WnUrZ/BIz8pt59wj06dpkL/QoJyGtjYXk5YK0Hht+0bnHoadRlhfLbr
jiRma4fP0/DwInrp6RKYa16f+4FUsANlj2p95Qt7JdttiNyfdwIW/r4zi/XOfQIo
mdgGgL1AeHutvsUxjBFNx91SzlMBtpCLi1/2al6HqhmDF1/6OSOT4oEcaBREIAL8
C7kv+m5NPnRSEfCDaXm/wNTMpadUANEZDO6Blu5IcjAwBgwuJccRVMWAcTRu4ALM
E0j9MONHq9XRIengl1edQqxbKfGEHelBfXx2+KsECw/xsiucEXZCj9cRj0vjfUqD
K+ihPkNlSQ+gh3nf2m8ShGXPyRRsunAwNvPhxa0VXUzPY9wJjkbNbm8Jz452KNxY
BI2EmjFct9qS38Bstfu3AOXDr5Dm8o5B1voNVQwDvgsW8zry6GDU1T8GGBeRkP27
dSal0y96bE+qOiBBeaM+kJVGRZp6VTyz2q852EG4WNLl1ArdTHfxrkIoa/UYU4HQ
rCpXQH76NpicsU+tB/repOlZr1azNRKFIpsTYKIsHBWCYvuZBdWrwpG5yMh47oKb
gOpvEuxo5kt+onmHaCaez+c6f0P3RhgIHDZs6JvIextY0WNWdSekQJJDeGZGNMR9
umXp/I7TdiF8LSGFnG9hjPpoZT2LzUUzU05IGvKDJ3FMmvhg0QYo77GQabTd+7S1
EnK+L/ruhh9GDh3jKyICjJrVW/WXOs9MyJj+xPsIFNTZJSuGGjX3Ixdzv3VQ9aiv
8BsCIe1imXN0p/kljOA/3XzJ1lUA0oIEm6KRbEL57O/3VqxLhWA2ulFzTKZHKLbM
Lp8Axn/6R6Gvkc0IWklpW9DXGwvaV17gMkVwI2TqX8s+9E2LxdAFhlfDMvkF/jyQ
xb21pgzT/+C9Mx+bt7FnwrPndPAxjNuved5TSwjhK29/wGtFhnkvroA/7RM6NcVL
KEIHDcjj3Geu+GBOy37mT4jklHfcCq7MCh8SnOP/6mExBHErWVvRXkCNkVhJvVjW
mwAsa9wRaCjgR7ZeW0ewz1Sx4YOeZuNB8PziQmnZNE0xE6Tlzoxo2EHFzbqefkfI
qVIT7NcZfd6D1FAPavHmQytyqZrW+fAP+tAU5sTNE/sfEpg67iqZbQlXyxU8BaVq
pheyDmrlcT1jSohw6fTHHv6fNIDi52h9g30zObku9EJ4gnz4h3bkXkHnKi8uocX3
qOF1NnSQskFJWM7G/iUPgl7qzPdT+VoplY/ofGuMD1zhT5HAxpR7NmmLfE2jlX7F
v8k/Yb9abPSnRLg0W6wwMCnnjaccm23+GP0E95c02vjq77lMTbyLfx5iOi6IVlea
wgfH4B1RaFZSi9xLwiMqNS5h77JiqXfh2MP+WSiZKlTvvgp9rgHkErlZMr3ntVSQ
H6IY8icG2Mb+Rpglv7B9L1XcWRFlPz7u4L1//rRWKbrlp2Y/YUW5NHXCN1W8H6zJ
+JtZy2fx0mcKulxZ9hDezWTfRNk9ByDAFxFybqlrIMmfwh/JuFCqG+EmzWdf2+sM
dcusIRM2mZvI427KiaoK4A1CGFSxyQ5j7JGsdGLIJHh3yuk+/iY+R+PIfOtYu4e0
Mzlqo7LQFAf0uVZfp217bruBxTEnoqwb/oPHJrt+/1tKFl9knB4m1V1XbyPPukWA
8dhndh+XNLKmYE4CBl+RYrGVntf7qgFYXzyMTKby9cTpyz5kIbS22FQw2mBLvTh6
xMpHGmY0CSjsXqFpSEG0owZhCpz6TGdFpZ3nV2uWo/1/47caDc6Jke7SGBYQa5bd
QVwoevnOlkl5FmtnFrfM+j3kgz6zA9FTBBLNX8rFyv3PHNbmCBQ0eN6N6LR5Hu56
JuR5+f1SLCyxLkrJ0kA4Vc5xnSrc/LDZjA5DVNsxkQsZ1y04Hf/ja6d+BjRWIHAg
ngX2yhkJZ/iwRudMc1B8SwNiHSnTU71IxZq9pr60S7U3//5H4PTr2Dc9Yog9OvNG
DodawEq8ixyWWQOdlrZnD305EIZ4d4ptqDxD6NGoF8yH3l2r7peCdgS6hAstvrqi
WIHEVbNZy9xnJt+ouBCA2U9PL2TQCrg7haEBL/omOqJkqXATgjJ206M6UwzDhdHG
+X7NCLODxrkvmX22Wabz6nj72U0bcnWsU7FUj6mD7q3j2KYSL1hbATRrnooe4lTc
ittCek2TvMyqd2ER2WHH9hJI1UItB3K5mPnxqoKzgKTlVDHXjCMdyWbeVXX9oxBR
vw+ySo8khYF0zCS18D3dArwg3T9RJCzbJs+Gp3zsq21hSiIbiBpvBs3zmk8PF1Nr
1jbCkdg+nBMVQ88mCWi9m2RUslr5JIhGLEe8LYvwx5VIjz4E1zkhxNblNg84P9lL
epf8Ga5lmy2JXB2wYqY7RDOJCYx8dYWiIkvr/RYHk1OoyzztshuaWPHeHgn4dozj
ibQBYNn7czUFt8kaXkqafEK09Ur1ND34/0NoXZg9jWqM49TlLxKq2iKgXQbWfY+P
LTsm9pTsk58oBTJEGwAIz9By7tS1f+0vdRhKA7nCGEWZ+Qp0DfdnrxFH03e9ri9m
sxBZX0v/8tJgncu44PcsscW6pJY23YvTGRzKJl7ROpTo2ao6Cm8bHpc+XJNHHChv
ClHzdcQFWiUIBtPK/jCfFaL1jgUJoZcFyXcK1PTcwt4NWXfru5+ONi3GaSAxpKr8
6My6u3jkyCKyLnCsaoIUWoSgsoqFA3YJItZ/ADDcs8fF+VeQPHD/10hqyti3A7H+
8GLvUI6hMObZKYsfGbRjzzhr2OJinXtfaaCQkWYdAvXeX6r4zhArttAfF9t1k2+s
ZOYOfwic9T2ktUIFAPL3qWFQo5gEBVrAlM0xlcBY7o4faR9Kc57a3lPDe7tS2iWf
AKIU0rjGRxuKP4yLXgz7HgL/bj3Kn9tIiDSgBv8DOAJ7lsOo0QuNHHHqm+6eQ+WG
upmn24GuFOgsDOF9elkhMYRoMB8xOpz6KWDw8yYqRgjya6SKm46wILZKdSenlMTA
4lRbWyejs21SZ9yIy54pziyLfWejvuH8mMRkxqa7FIo0Ry1+G0rI4xtPUhJyspSN
prbWFgx125K3h6sBMEbcLpCa0L0+VY7VR0IwaUWrJc6v/dbzgdjmuIpWo4weJDlG
duR5h/44ii2vRCBSBS9Z2nKctZylqmXXNH5d48oDoKeEod6y6VYSU1Is3wZ4WaYW
VCzHBfaRsUwced+zYaNzCACeb0gZ71sis56uhx4RZtk7Djcm9K0lO0TUlw9I8gfZ
MPGSX0vqnJTGnlzAS4pdGNGhXCHVaOdXcuKmOLoWBjlVt7fWvRegikO5ox8TBU4t
JykpdC32E82qjhsUE9vKJOqGHe3YJI4SLlB5FymNaTfMLlsevpf5drwBSdko6awE
SFaDOslZGtAzQ9LgTekj556/sXWQ3IQfj0tgoCZdQP8iOke8M6F5GKv0kPsSyW+N
kZc6EQfoXJtZZ3HGNQzDDcENI4EfCl2mgL3+ENoqfUFv416X4NlYeg8h+eaiyZCY
qrWmHneXDbbo8LwXp7rC8ZtFpPekq2kguA/c3AlI2xxOucJy6vKvImQDjsMwk7/3
5a5k5+0nRXaoanZoxrAg1K0sc9HmEqfBlXQSwO+DyMPr0aQRHepEy5UcXLzYE9XQ
TAbvCpJ0gR9ffBRtblVFW9Pe5jje9HiQXoR+5KhFR+VNIX4d4jEuGmgOE/9p+pMm
refFrlZh7mYDl4dWb4yvz5tVJz6lvU7ObnQ6ID8cSapmbFlTkQsPh3wtmPMC5zwH
oPZmZFxy4cDsKTG66Sb1JNIouPgjnr7NDDIn3G4Qo33BIWjgadDwA7MHkxshoLSn
f2tEfKsqwXeW46Qz+o9Hfcuv2Hr2R4UahiKigB3HwzomoL5wEsACPLxy/zQexhDL
W5WynLJQjnnYLFmtTwr6yx06Ajr8SDrPOwSiIfvtLRM=
`pragma protect end_protected
