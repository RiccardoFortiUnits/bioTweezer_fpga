`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zt6/TI0d7ibXoSkDerM+plgTnAKlSuZp+bSzUAwe6/oFrekOH89xrcqTGvD0hVih
DWAaZ+CITYyq+NmHM5ZSeWJrSFlDsrfyGYvgaJrcgCz1rwJneC+lxdM/jvc6CMH7
ylHlxruBI2FgA1gIMETuqNqyxoAn5iZ1LspnYl5kMZk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12336)
jjOLqRe5L6RN67OODdX/TfheHRSEIIDOyAuO5YXu380OkptqxWCOLYmDYDda02ud
EkSYToNO9LmzyFH56TSMIKy0QlxNwJ8ekyHiTk2Px4LDyN8ApH6RM96USdnxjEK5
D8nEtZKmJAmoGUwgikr2t+bAv2oADWdHW3kORxRiVGm4MfMOJ59PSlsegF78nhk7
isZNaBhUOnKh07wKhMZzqKD5uVuSss1R81GBN2AsiT0E9uwTGCOwScw+xbjW0KTB
YA0jRb0EMj7RLfa3WhaMThFUxZQyh7zPinP9KQr+Tow4RU+vLnJpIQlrtv7dLSJ5
n7tr2Wr1xKjsD1tc2GbjgEIWOpGdF/QEBSOUY+Qn40dx1mQZmK/8A3ye0X2PbMhm
Hc9yy629Vw9X2hyKoNnovHAP0LflqEc1+XBzH3Bg4wz10tnSnkaovgcLy6W37Z6W
feaeQODCfnJ2CvEptv+mGox2720rClZmF53K53deMqtX+Qe1c8HkNMMh7v2Ypdb2
C6Gi1LVBI/9AgsLHY9WADjKrSDVN5+sE/Dw58NGydDoePtnhRgfai32sKGRidsFn
W3D6PMGbtqJu2wlc7FrpQANxkeydlsuZTsN/xjV+O3jO0aMVNoRk7/CexP+rh5ru
ELdbF30+tIv4Kw4DQu4sOOvUJNI9wE2Ythl5DH8bLriPqCHoc5A1YVvwLH5Ahwa+
v0CuAQ/BUyJzXek5RUF/0EVCuMkUxQZmbKJerE0cgcenWKeTAuD8ZcqZK/7HrNZ5
BKQdLXAXAesJv5Ak/QGxXk85ay6iXL9vPYoIvslyDMG8Sn+5mBgC72WvYw5n3yLZ
uHTC4hg6yW+XQnJI9S+HD3+xoA147DjfaMnk/q9FT8IUolNHpBqsRQWIOSAmhvfh
rdJUVjKx+sxilhjGWQbIe6CsKXInkDBZRfjbmyIJkr/kHfF/cyIaohdnyTStNScO
57vOhVkqg21bdylFk2NTjsFHoRbRuFqGDeUFGl2Dd0thC0JTfG0+AMJXBvFexfVJ
sIQhAObSCKj2Kvj8Zgd9nbre0rJe7fCecpqC9aqS1WDyQEy/a4I9MOzRIG/ftVp2
uK3ofBvNDHkTA69U6xxuikAPrA9R+tG7uJCXBDMSXfbQt/yKyNEgR6Ob02JVBuAr
Ihhig+jIpXiG/F4UJtgR7LB2M8eV7cAmMaNHOntkqKKa2UBcYqQmJ0v4gYalIcNq
OUwob5TpImDO80WfgF4Gw1HwasD163ih1/7AiIRZwonILvjj1MqZ6jzujop7DoX6
ZOso48ZkvkoZyPhQw8zI/vGO99ruOEvs/pCa4Wn7n/EDZ1/4ZzyfS0knq9IzI2yJ
Hca/aqib6nBUS+GlGhN7PUhPTdQf9A6PsbrYneH895Rip5dSIAOvXmrPzawLGH4j
0Zw1XPUprG65N3DA/ePYk0gCTHLT0YES96ySOlSFhm/rFjxg/QuwlTNjn1xrvYy8
YOn2jkO9TTTIdeD3sgsAnz/0RB5NmpwMXwHfnip5GxJ/ImbJheCoZfOhRQMXZgtx
p8Ko3FkzazXFFm2JtGEc4SsgIp/qkJKCNbNIHX8CxpHunR6QuLR7ObaVce/EmfzU
c4jlTtZw5f5s/cDJ4EEETspSYMUXYJtePHuIvA1bQnck1E/knZiOpUIEOs97I78F
wAIUxcjXnVHjFKt6YKz+pLRbNDCEVyrVv0qjCVKX9AfZv9tAy0eL2sqHEo0/wmuk
tZwdZbOC7/4QwYwyAeppftrVwMI3n5iYfTQRWn+t+p4WnUBv5qQ+B4Sbri61+9L4
hQEQUDaq8wdXj7fdiUlzGcsO/KgQxrlN34fUwfL2bbKyVB9J9zPBg2LrMN/wBcUq
VdVY4w50B2OMMoRBb2bdU5Lz/Tj3mglff+V1vvudvWohvurl1N4Xx+PlRF56v3T0
NW0vCboJK6sW57HaqvAyblSag2DCUobPLnHRL6vZXo2tuwVxqwJe+AAbZlDueS46
igpCvyCZtW2jZLVjfqiSv1s+/z8v1ZN+Sc4NZvjedBzd95syhCrc4K6yjxD5G7Ab
GKxo5aTFydQs3MYWPN49kkGP02ry0BOgK9Yc2TsDPrqylQACryU+nULtO4yenPf0
n7lkfWMWevyC+t8sNVaBp+izW3qTFs8sUkUgCYN84y77fOcVadfnsAhKmR+m7q8o
OhxAQH+57Vmf2bR+tNjU9oliBaE8L4UgihDwi+vbbO3O9ylQeqGzsjY1c9jClgxj
8OrMKbYerQz8dEu5DgAGJgamgimk8k4EYBmXFAazqvtb7bzxJnqGoM2fa7uI4TIo
ASwoqeb4LWkzRbtulVZ9y/KI7U2MDqYrzxAoJVkYSeKmt9+/HYLYnKJ0MzV1cZfK
4WWaTjw3b1ebV48pANu7Rorn5ma4QGpqC6qQxoqjxganEyURQg1rc/5Z8Mh1kxae
YZ4rvpU5pUSD5M6kiahW63Toho+J7AGHqGxDcl+rzi0RPF1oP9fu4oJ3kRq89cjI
ApY5PZhg930gqyzxSXJ0GLIDqUjEv1s15I7ESzTq94FADZoepACoTwwh+/WT9SLs
JlelNhJhi0KcIWIFwDEmySOZ21vTuM3DDJrm0ipKcAA3CuTLHfq6ReborbLGoCoH
PT+FQfQUhLrriK8MJRZS7Jy6UA7OkLQcPeOuSCBDaXaqQY94VbtDmnfKnEzYJAAM
qugvnqWo07jtDisxhNZ9O5HNyL6GH4VFjnSX+21FXrQLzuJmSVyZU59CWfDGePTN
1/UeoxJEOFiV0Rx5svpSFb5JoZN5Ajhz3RmZJrNYT0jQwiaRRQAqIwCEmW89lrGl
vio8q+dnSTlEkgDjllGTBPJF10XSocbVklm6ISTiftlJIvGwP8k3tPku/lWPfxWt
NtsJtXkDYPmQIXTkWP3HA9WPVHg/0tZo/Vt4RTPrcTA5nCm42LCzTelwzTVTMrjk
VMo1EbWawt0Z1XM6w3VCT4tS8DZoo3E+O1+rfQGnaalF+GOHJpAaTib/AcdfW22x
paU1xma4MN29wsV50NyETZ0mEh1VI/g7kVJJ7XPy3EkvP7mXD94ND5sbLuk0XsDV
R0sK8uabLp6/VKv20CVjtVw2iwa1Qn3/m7v/JButqP1zyfc4AbuwW+3w7SoRxI0B
qfbvVnU5+q9CbymyHK7sWDF7TnY7q+BtmGZNnEnKrmKerC+qYOZ54iTupTKBsqEr
XqMmsaoCssk7n5o/UMGUrD9cNW6OA3P/GkgLWMmbvTbzJpSy1Ox48Jah+k8YQpJl
qdg9Z1/rEEo9hEhvCGW/yjc5/9VkiCiIcnjbjbxUjiNkSRRKqHIqdQwZiP6hJ8C+
QcJ2ik53hTRhc8SZS5KpVDDPg9HNKDntA7ZKy7E5LjGVOykhhRc1UsOXz8uvbfQ8
5ic80yLBZiISA8DU0OUx005LBK7VRkAdR/uwVgzM8dr1kOLu72RE3EBbWgCXf/OT
sBl6Z7BL1JPcmFUTC7gNZ7WMzL8nMoqXrpnJVh8o/ILU3Q2IdW0toNQODtUy7rqc
DqmiX3h1USzwqQcH/P2y7asv+hgt8I1QIfE/WNFgFfX0+Dw95SIOx1WShLfEfxMW
655/Q2yktFQnVcY/+d3UCGXLqgoinSyLPIV+dprZqAMHHHSs4mfyquB5RT6h1PYK
LhyLHkX7OBsX7TmIFwlHviuB/LG+74tt6VdnXlp9u42qIJYPAwnsbqQwxOIFYdoq
cvgxeZ/Gv8Jyo+u9hHL70kXGqTesbMZ5xFF8mgPUEQgRt8DD1cRfLdgrucp2FlMH
7oBSxL+CCkHaxo4Vvf245CvPGrjj1PTiUM1NcQxUJcyXHCBdgZt/whV8xNezk+9X
S4PgGCf4ANUN851xBrC+XbCzLzZ5cPm+JMO1zoi1F5Av/vZPxETsB07XO5hc+lRe
AIJ4GdJABAq64C6Hj26MtwPaqKhGMGUJNcWKTWl1Xa7AHeAV7sMfCJ7x5Dn0Iset
drzXDm7wHPbTBiSZgk3FoJw0v5yfSQyS9eWQ2TEmSWV5OvrTKkX/LGAoFa2lqXPm
FpP+n8sjF7DZogUV1Ux0TucmeQ9P1p9pH/QIy5SLjfexfABq9z9ms92DNOEJxnOO
LJcrcE3ezQ4njaorweZgN3xqINyCrMdUgMRgk/9yyPFWovJXZVA1NDTkvqCzn3nP
ojaBecNguFUR+aO8tNgeryHlt4wDVZTloUIPqp5zpTnIxrwPY+O9jv/59L5Rcjse
vyGK+/Oow2x5PzRCU1VzNqGeRv+6ThwRpvS0gXZyt+TqJPEOpbd54QaWSV6Y4Uyr
Lukqy18MEd9vePB4l+952fn41f2gdMf14+2fbB28z3XgHojwfeK8LzAPZgYZGlDP
OIBU3AbgG0LckHw1pChnYVgSDi2swNvmUo2teypwH+8FvmCv+a4cGDUJQasbsHnc
+9omvu10MZhsKhpB3qjG396AfbhSw5TDzXCHXi7NDTDupNBmWclwn2LQLK265HA3
cKrUIH74nLm/YVgY6t5opdPjq7OP0B6CSfQWLA0i2e0MV5aqpLKjfBudygPR4AhV
ZVAVHxcJhtLMSWEB5cBmBb1C77tPvwptuUY9zi6JkfxzGfdrjvU+dZ44Gba7cXtw
7KyUKveTBfVAHzQ9uZqmedTfXm+OK5LvZcgzuXpAb1Rc/2FKHB6iy9GgQdLlL2rt
32LxUTcgWieGZeO53JsowLc7KjKVVzQ7wfYCdl4UOSbLoxb35kWY9jfYtyc2BPGF
+6TjmnZ/CLZukRvqBUZrHVkG5NfIEv8VHdhed8uIIFi4jPQ1RpVvuaLPSFYHTYQz
JZ2g9qjAVvm7rNi7F/vMxeU5KvxothColTl4JDzVwSiTz083CNBSMAU/M++oKUQC
8s2TbDammddnFYohAcxnGaDfR7gKZSOGg2OW8EQyfTOErNENGbIj1UoWyp4d0VnG
6Xe4xOwgpGVE9DMG5p8uw2ShWYPNVRN+OJTSwKQMNKk+hPfekVFDuGVLjQhwornr
zvxZovH+k2XabjxCTjbhGGLCUk9iiw3jV2rlA0+f5uSIqPXVC8mgIp8q0893vwbA
qnLLB+5HG4a2qZAkdSp4JzZmS2TNqIYACextSLBSw5k112BWcgIzeLcYCOSjbYcO
gWY/RfvO9K3Mp9pVuZaRVD/rlrcGCzU3vqB/NZGSxndN0rhMhdbQSDbZl9bGcDlk
ymtYOm8+2SH4WbDfc1tG8K6OWrypxIFhTem8Lc2H1pxQuuuOGGmxSNaDLod4qrqU
0PiI148miuf7OEA/v9yoXJfyqDvRvwE6/wAJReaYH58oYBwarOAjaSBb1DMFchDC
KmKelVrA7j3AVdutP11Q+XHu3tHgdKrlWwbH8Nn14l3Cafexh76wyGd+SkB/F1Lk
73qZybdl4I77/ktTTUaOrILG1rH2EfypoyyeWiD+Seo78OXuu75p4Pl4BlcREPkN
nBINpP62+8EAwjOrDPK0lRVcf3p0BK52r8whnjbelE0kLHg1Gvs06EeU+UAqxuuC
JsRKYHZ5oeUdRyCM+Ow4vA2UCKW3gLJZiU8tWDuWS7sCfDjrL6ZTpAs3CREykZ2c
Pi/hgaiYz96aYwykhI4M2eSGG0CHRNhE0V0esAuPUAXez/ZSDFZx897Q12e7P6SD
qQpDylvcNjUofSo5rVKI0YUSSPy6gthzDZgukdYH7d5sF6VP6raCpQ+aB0hDZygn
poVJcigfgwYwDK/t8Q66TB2aN+O5m1RxSKtWCh3DCBkG5LTlz2ZVyAueq01pf5eq
Dfa49TT89wY1TrkOmWQ2Ywzympp5to7r+qppwrb7bToq8TIQmSwtTJMWlnszMy56
4eSY6AIuA74MECIFZVmdRKeKA/1+oO09Sl5VMFXZf8/o2fEa7sdrnSV8q7DzLSOQ
W9h2ZG4Ga0d0z3f8NLEI68TUXHR81n0Cqlxl+7DhyrWabP4FrBa11hheFDtOytoF
6RSPimi4XpRd4dXKohgFaIs+V+YMqoAjOaWvKNHYz7q4Y9yCbAZZ+r+F4kYJxreL
KpJf7BYQRxM555Hvx/cqyNBExOtBejVQ4nLzWxenodW5a3Zad8Jb0j/uClkXutAs
FMRJ2fXWMRiUCo8eZHi3Jf3+6/2lM0IoyFNLcCtzCj5f5KDSJVWM6tqph7yFvo8O
UGVZDfjtQGCnC1h0sattgrfMJvIkXNPck3MWCkbAP8A/kmy3Lp6FB6uY4P2KHPeG
IjhLIxyToP1vXrkRTkSri4ESVlmOKx4L93r0r5Tz1Ov92hTEFulUdDw3gDhB4wem
w80zoee1Dz9373YydUmNUmYDYVRlns323DcARLcjvIjMkPlMl4YifQfmAS0TOZxy
7+I2GduMUDavZcPAz8GJ4P3fUjsIo5BnEhXMTGnZam55+aV/tl+wb/SsKfD1iwPb
St5HTZWB/k/OlSqLTpByCzwhIS57eMsTyQr48q4Mtf5JYp2E9hWwI6Pec/2PYpd9
s1z9yjRp9o/hL/Y0T1CoFhXjDQRXx2aSmaCP/Dlw5YoE48+SGLT3dUnVPJCKgLGf
Mh03qdTIiRNWJrLTNEuCVXdn8gXYWMXIsKD04DoBK/p1uHu6oHnu2yQNf1srrbxm
var1ikapaMpFsTUxKyUmcjPiJevbR4tOPdsaH4dvKvzQDnipnKlLxFwqw1MxpqNF
dK4a6/1nyASKUz+l/dvvzPL+2B1OwGIBjuk+33+ndaTckphrjKQuqA4QUxn7Ujqb
DQFlQdbmhAPDuOCk23aiNRC4JVnl1g4rf9OnzTAlq7IujkHcmOBd/yS0iOzl8ywB
Ad+/3DM36bk0Iu+7PyRtHta2QLk/EQFPwEf9OnRX2cor0lG02u+C6YukAln6/kyj
wgQmqtZ/QKGRDwrhJVwMESnXZJD+tkh2MFngq5AaHe+P21b9h//YEohoK3G8KT+5
TjOGbVObeo4YkgvyleU6dBKxIzu9yC24HF2ErXKFF7iJD/aCuuEx+OJxO3AmLDxH
+6aFQbCoiLkG54MpCaeEs1vn+VV2wDChZg96C4VC7y66+YiZSNcSsRS7lDC3HqKW
gLuVwXwml9tyGoud0npDC5bHaGZRGHia4gr7M6NotnR/Mqakd8fyJyieom1Cfqeg
oxI856xeTyp/ROCf1SwkouAgNWqDbIpHckLqo0z6QzEglQIyCahfNkjeopZm6i4U
RNc468XcWuW/Wx3UYQDVizHeiw75bEHLKyTtgHFjLNN71eM8x6GuUBF6VRPMTfBv
txOLLbMGo+s/gVFjU1GghCcA/cdvQ7G4FGMUPgk+NjHscNZa1y4KoXkEXS7Bgz/D
9ec0KON11MLUEaeI1ZPifXPfPnScPkqsp5K4/K5yFScRnkvyCM+y3HnQm9p0twGs
EOsVa8tqduJVIr4B98HSo4+wsp9D0fIRkSbYzZHYnHvmVn7rhz8fh8FPuoVyNuLe
ziMSJXK7GXkHCF4t4zqU6p1VxNTQxRDYVX+JZjsmtLE14wBtDCCjgzePGdw4Evn+
aS/wuquSWXj65KhqC8PLVrVtVlLaSPZu7z5eFXEsu9jgFxBfjvR59xVINbwMSSUY
07x9rswRW9iQfx3mQLXcvZBAzomoyRWTrvhItxDIq2cyNoIcc9wbe9kyNgVdl8D9
4uFj75ZfMSDMdSh7Q0cS3ibRTqMKV0WQ0B+t0x0CwAZxWwkZEcv4JA693Gwr2jFx
dKOGb/kTi0pZkvd2jW7kuFHtIEY8p18zFUcV0PuFFuheys0RaM29AgqJIx7dNmVj
CIXA6AOMYVnHiAW/kJxSBr5lU4EcsAvKVu5gHB32qhQ5qAdNfI8CKvG2OfxrNkVq
cbo5A4ZuGkYvz7QH+NJj/duzT9gGx7B800Jg5dhEZEktJWDdsrEam6CanZpcSsv0
GJB0BOlHE3tJas0HyTkhTLozMiaoXRLpc0D+nMdz3zERoHri8lMvJGZKf2Xl/g2s
Hrd5ucpKXz76OvIylvqJ2P1X1PzeAymoj5FklkmENQie+iCS8M1xtSQq2QrtGLvs
R3tEx/oT7RQncSVXu/EkGknhEVZjy2fqjGYQ3Gh19LcZCcqHgwZgdopG/PcjnBD9
p/tN5ya7PUbFRdxDUIXWGIyo55S+/v3bzZLGU0NWXj4ODKMHucrQg16Wxj1v3TwV
BIxs3DSVO7qd7F4OK63NCAt8XRHZXam8z9Dv1XkoR6g6sAvVNVA6KCzm+WWtwsg+
p9XvM4uh/RYwrXQdKTxsmNkHR/wJh6YwL7LQZhYUTlI7605gLV0fCDGaNbtAyTE3
GnXWxo7u/1EB2DCmK37wdViVoeGTwAzR0CCAyLsBtCyaVMEiHpHIWUfbNYyj7bPH
FUOuslPsobck76+QdwQTIIMqOzqrY0KsiJF5d826EQr6UAzVAHzyzqh1ZOUawv8E
Vqw+bt8frv+6vLum6YM+kiFwQ+6Q8E2gSB+jvXXIQw1LXlRvBiO4xoXtKqWN+WzO
KfH/pfpsYcu3PoU7UMiJsNbT7IMsMIIQEUlvcbSgkQ0bWBxW5mDgdBiF/ScN9nDA
PyEALwrKtdxzeX64+xylIu6xBxzhPO5+HM3XwzPWOsd/Tv5Vqu3pnryNr8tR1uPi
sgCuSGnsvPtTwhUm38sveXgV/u59BEOmMlm6sVdcddSMwuyWSsWF5AUfz2j5TROd
Aj+lyzpgLaSkrwXIn/WzRHsGhNALDgRSE9dWk76XuT492Bat1BOB/VYTCi91Bm/e
W1McmVY7RVo44UoiURtzNX0it0+32cdp+tnwdfVmYUcEUTZH+Uc6WRQ8vGGpOPHy
Zs1h/2qLww8mJsQ1VgXvUE4Rc/bbArhUGO5gsJYrzKmAj4rPFFKcpxNRsl4GUg8m
g3XkpaF/fgx1OPpBwbwWldDREfAfpAdnCCJq+lqsKgB3YLfdNxwxgZS3Hy2ZGXWx
f4Gf9bShvJn0ho/s4hs6Yvnff39ohOrwqnWaB/aNCHW0LTgNCuTTfsmFUd3vsEJN
o4iSZVl4KDgWlPLe4jMt4EooQMSyUGytZ0gpyKZI0Sne58Y2zmmOo/l44o55ImNF
kr/STkMhMDuzLU2zCM2/GbrNlTu/6/adVTRScJLvEvti9oCCxGKXigPqOg8HEabb
iCGoNejl4CAU2h6AUy7WEkEkkSrSyp0Qhfl3RKa0I1dqRE2bfFFc6kNBBYRA0bDY
L/JiVtcOsEVlRDjQb8DFONjmU5x+u1AfYSyAjvmYNnYLV+K1ua3lsPDi7zBt3G9R
em78wicz91VE65J3B/e8ui6NpVW8y14pQczBxWYR2bAgfHfDWIi0mQWiE0M+nixk
arQFg0loG400LcXuBmzvVO3G5kymCPRAGytT72fPY/XxcFhe2UVjL4Dd2Xc8TK2l
Nl7gKJJQl31JgZiD6ubtuJicdDlPYGzd8/mhc6gJX6MKdqjoUSvyypjSFxsz3nqQ
x2am87pPsbCy+pA5N4OIOMkM2uk577vxDI66+eqkoq1nvOloIUN3fc6HRqMmt/VD
itWIPki/Np88DNwIuP+eGUnwbdPFCN988GW2f9ZzS3Ce+m1nJuyxRZRCbUHSujzK
HzsYOnu4k7Jx1m+WvL2DrpzK3XJ3LJVpaHjkVsNQhAOZdtKwC9c/69UTflWJdP1d
GV7vz6g0pYkLPeNGtAYSdE688WNsu/aFU4lOTP2GW2NEkIEpg4223kCoAe03NEjl
DYtQpTrZdJtf+Eh4PE5kCZ2yemAIXxJCOgTRnk5GFcSyN2S1eRHSNqRyMxjnOKz6
aJAe8ML5SCDC0eNOemUWyrivXONjOOz3OIsOYwlwQOlx/fna72KblLx10Q5h1JHU
Ok221bZ+V6TdD4tZpZFfu8BuVUlF3g8/xWcPMmMq1W9xZdz+3B5S/MYiD/D7Pzqq
ygqT0eeItO+q7fdoJHyPkhPoq9FbyiAgVlJFynVPV/wSffWXkBweZ1FsGqAc9gXB
qj+hyYs1G6hGFBAZ9mfKcFB2NmU0eci++967pjF7lZ3Y//PmepJZ9c0mWjha69We
Jnwa3NuhkIiU3EIC/GgwL6nmaiCm7t7haASFrMzX5H68Mu2F2R+eSpHOaaxmhFvg
c0YLpllRsbcL9lmczl1w/P9TomYpK4v0mG7U+rxzKY1Fp7FImxhYmOuva/HhucuY
xh46ENy0Qizth5yh+FpYk/2yy3UgxVC7pz+bEV71mAbnOvmudcIX9rkHthgA+rJg
0CVxic/OKlg0ffVPVReHTKfwZYcu4d/ojluHShu8o8Vq9pOr6ozfb8geVgKGxa5J
4KnpI6JF1Yhhl5Z8FyXvLBax7Da5pnbsieo9I623QHONIgJVNTRlUOalyaHUn9Cn
l384PwfVMYrCV+Noq201MJau7J310yML6uWRst3AqiRFYQBMSss3683ho0r0qgI3
DfwSEnmlozPfp9rDaf4eAHwrvjKgkp0DGRbgQlbInhRqbqdCETqXBeP+5SKLvuho
d862BEn/WOZ2wtqEcu0656ceWP0GljAW8PQTPWrR7M42SMs5EWO0opBx0IoJUzPo
xzuPslHBj9zhUkX/+kD3KyTfZozOIe5p02fpk/VPXN1B4m4rruaiPPMUSDjwLF3P
EAs9JrTGjWYe8tHdp3BXRhIUv3VwcqeU0lk1UTnIoUhZ8ZOXU6Pudl6jTSlEr9P0
LsD1vwP1r0FNGEWcFoM6F8jQVZN5vVo039FGZJ3eHWqGOlK1a/d8kb3+aMmdaqMh
+ohucRs2GP0bukNoHz4X83o3Q/O2mwgmbtAdJzDo6Z3zD47HaxXb5YniidnO76NG
Uc4FNVf6H5yS3C4LVQ50RH+87i2XrLW76QyxW0vYt6MNJqb8o9RXrhDtoK+QN5xk
GrLsdKkxh06eQDBhPPMroD2DYWX8x/lRLwQx24tgQzxhaKAYhd1hoig2IYiXcPaw
VvL7BTezyUI0SelmmwqsWjYz3ufNlEekGhfnbq4gmHkOPrR+Nrp8YtGHIWHD1bUY
5mWIFWLJ+WinllslaK6BRlPUwEDUdN2XDoUMLmlX0MiR+3VFyeo8aNh908Q+DuHt
dFKRuUUTQ4qo8AVfuitzyzd+SoOtsRp3KufP+R1A00Zczp3q80Q3XAHnwp6x79pV
tghvLbEisuROY2nXarHkWrXZyLjGhy2G1J/AuRUVQhMoAoh3CRanXpxI/NV41Qnx
G+4aNRntOT+FsW8+vicI/4Yl6Z2IpUmLXklUIlrr57F6Lih9MqHrS02R4ooBwPOS
tB5RXFamk7ov8y8HFPBraUTejEPR2S4YqwunZPK5tsNhCcj14uLq/7C6y/0adZCL
GtBqHkzpFbKPDxcEcr8z1gmAkT089CSW2Qh7WnoOife7JZMXpCv/vjkpKQDawLMi
jnDyLL1IpcEjP9WpotGHmocLB8IQKrQOXwJLMg6FM8N3G3pdNoLPRwIwXwuo05SJ
7dUexQUWuSSQRopz81+0+DaXa1c3m41l78WrVFGfI2FkVhZtBPd2F/cMqO+TgXDH
rQrzgtcgvmcU73IgTVwzQeShFK85VelnNMpaHvL7z5szbhd0DnvGsJjcnuYpDC2v
P6MnTU5eT5OfN10UfopwPi7+leMbk2h4/+Z38QRFDyphfB+lX5SsgNbeiu7iUyzr
PQ3c/57mFjYHoKp1EAt7VmVmpIrYHPEZhMr2NzI8wmOqeMA3l1co82sV69xwnwJJ
L7UwePP4Y9J7DiFfsn9QQIt1Q/UoaNZCmFPLNT4/wu2/VC93xMPnDCU3+QLMKZLC
q9u1JGe7hXIrHk7l+mgzF9+FO5WuBe+UZ2DYtGI5/tAP7HrwDBzUlOMhatZj51hN
rXl8Fz8acfx4DSv7ClqnPtn/K4KZDycbxFoUdvTjlk7FVL1ZkhTcsYvkHWGP5tUt
XkQL21qfLKIRNRyAE1/ZDn5jiQqiJUQSMYaaKjFBr6+A82ZiBWyuyj7bRWfiDrDE
Sw+xvIp6S6PBqmtNaM/sfW8bbrrXXKh5ufGKWi02/QXBXGW/F/FEYmxPG0ID0asQ
BlkeRgAPMSgv4zZD+Ztj7GP+S/aoaC4YQGufo6WewXP1Qo0JBivdGRgazsYVv9pc
2VL+lQh6iVp+Wtl7NKd8Z9zKy6kxZfNjyvDHA6CHysBU8FwoBlgiKzfyfXqmcgvv
klSWonIjl4vqgWU9/BaDEuIYn6tCnbcTZ+WwJabBKX/gW/XZxFL3XQAFXsJp9bjE
bXn0JH3f7849VvwXYEqy3qNDG1or3ywcZolW78dhA/2UlV2CkRWmIagxlWmpg47P
7rkyj+7RyaME4/NzkhQbxM7gBDt7xyvQZKR0OI5Wp+yTxhBUONKlZ7S6AUHX151i
ezJQ3X10p+8bivpbpMngV9cVZCUveQSfb6ertwEK3aUF03Xbz0l3tVuqtadHWtJe
SgyGChO45v8DXsW9dHqyQKcJmiX5OBmj/IUCvEz1+6DXMNCGIjCA6pw7nYOAsSpd
emEV9IyJEsZvdDgpf4OlTl/J95DILbV7x+FTjUze/jAVt0uwjiw2hL8pq1hE8wXi
0mwKm5mLgmePte2J2b1Ndpwv2qkktqU+upbMTClacjS5MqHC0lbqfmFnGou3IXXr
yvTsSGd5njoYf39rXVZ1cR3Ab34O/PmpFgt9/nclyz9tpU1BpDUcqHV32C+7uvhO
wCTm2afrmpCgL+SbgkB9jgNwIJSmxDoMTr1KxlgSGLyGqeX2d4wDtoWwktbkAGks
9YC/Z3jrcth9bSDaBp72BjeBjck9nYZCpeZH507XePCtO2Vfcbx23WpU3zQP6QbJ
50kkBU9IodFl45FioL+LOBvL46n2Ft9gXcX88V/B/uLWuPJ6pNfPZWLN0F0rTuf3
3yepJrvjAh/OtKMcjvUSImQ57fOllf954tFXpV9fecLc9uSSFJHBiG3GP72tC2WV
Q+w0OzvK8DWjFracPlx2JHdMmtFDbyFqt2adGwcdepAecrdzzKXP5gs8hy3sLcav
mtS0Luu3Xn99zhE4c1qEnClfsVeMGbYEVmFB2vSiW7bLzcyYLdy3ChgrIKTEukjK
PFk8hy2mLITT45xkf2TLkc/NBGWwV9er43UdawWA0xGqv7rdgpcAKtpjGY5z3MvT
Ukyq7dT8cX3huub/ZR9NwwcyG5WNGi9qQX1/DjTD+6SjwktIAO8l9FzfmTmHaldd
ODCdv0Y89O6U3SbmvYzzXU15UdXmkt6NZ6kxgM7oj4la27Xvun35mUXN6tz9zAGy
aKOwZ+vdBH0ia2f/5pl8x815YU3XVspD6qrPDz4zkGNs/V3rmf9I78mhHyH+rnM5
61RGEFoVsCV//EgQIcExZre+pjifFZGy2L7Bev+C+UwyNpoDwmZTSlL6gqg34/G/
2/sD29K/O3chlhvwwj3vDeNwo6UO1QxfKcR+/vbJjDpdyipSTenxN+WbFSAROxrg
9nIKpzqRYyNjcDiau12IfVZgsPZYbSXaWOIvAqG+eSLfDQq6thIrOZDskKvDhoON
GooP7j3EiHKFHdzpVapqs1PDLxiVYvuPxdfy58TzrZNqOiWWavVDGM/0kXK83V/8
X+k4FSLB8sXnff2Vw9jHRqba4cU7oUHyOR5XOAqEyOSFwKQSM/zkmjMaZtyiAfuV
ru/Xc7bNXd5gtU7KGbY5qk0d+dq+Ct1XVYaZQpstYPQbdLbSk52ZenR6JEDC1pYE
j/BvumMUszIqmXMvIq2MswbroV4tmF1Rnb3pYNJBm92PZVdlIrfvgJgQL4Z4ioKA
zId7JmOq73MxYSCGTrzPtCo82Cc+Hbah5ZX1EVUcSW8Lshj4lg6MQ/BglwW0XTKL
AY9aKx+8WU6qUzJ07zMGiGpbyaIvb5WiP19UOoW3GbWM7uRDIyA4GKUji+mmodgt
+e3KQVlHSIjuSc7t4ry1Qc1TLVKX0QVSyZVUuqpd8+KIrbP+5ilhl+/RkbazvVcX
29tIv9MGzqdK/wf9ITZC9KL6b7g0PzfB09je/vfdB0AuemoqEbQHPhGthSPwhM63
I9ENi8kNAsZbh9Qc4EsgiCyEPZkr8gzBLHnOcS7c3m5VyhC8eYsuRKOxBVDf9Tjz
XAJk0s+BMDRxeebf5ieBfpPfBIpGRYUROdNg2uA2reFTG6yFfiISTH0YwbxAeB3m
II1/xL1KzQjb7xCZoCtj45d+JsTw6AqZgOTfsG0PvbiUmzV0HMWqeSHbALSPu13B
94849v1f9Wc6sDMrvk7rIAIfYsoYO9+oY6GWeBasJsBUOqJaEC3VEpi0PAQ7HXTx
/VNMvD8Yi7O7tfXbBlMsvssEEWqIAri0QIbFnenGOc+2ZiexYMrcIY5XHyXEW/bm
JE7Dd/VrfGk2CNNI1G1tubiBvkFbbqnyK5XBOw7hf7Jg+5TnMxH6lUfT/Xbu//Ds
Q9VbUhfd/adN0wA70U2fuNxDnuXFtOu5RWlcxgIDLl13J9rUxZI+jecVp18vVoHa
s8aS88tk2jvZdmLDrIHeyRZahC91WNLJbHDCrBUx62eXirPQeJ3xl/+9WKBWXkSK
FKO/JZ9/J/r4M7GdvevaUtnamG+1Zs28l6g/YbjIjCC2c8+7ia5aZyqw3IZ2c9i0
it+3ngJk89YwdUqrf3mBmnHY3TJlJPAaj6h4v6Yscn2WDa8JFLsIF88zIxFI4kDZ
wefnyoNckj6MOkpekoeM6xGFQMlw8hHBumkNy7uYFwG+3Gdyewf7qmHz5Uswf/tL
mKs0tIWTNm6tJURmJsUfStesMSsApMAvADrqfLLyOtSJUdgoFmkCue7ItOm7/LG0
SdIWqT/u6nFiPZzTQER4f7DEVvqxPFkchB5Vws1BpjDsYNG4Kc/HilGn4WMm2Nor
2tbl+cFbcJNRKMLZpEamM7mCewZYtU89Isb3CczvndaHhJ/XQFp+fzUwDFg+4gRz
587vSxqKes7jLwukv8YawwAE6/Cane+aqfefusBD1S3Ak76x4plP8frXitYHvjTS
yLRSWThYsk46oP1tbHBd8nFXG75vloLfSBEU0yWGaOOlijTt7+HYor6Sw9exTBsR
HHamjHsuPvNvmtNifqDG+kYlb4q1wwpdK8eR50ge2zmkK3R30MCDct0u17Hczn4Q
B0YqhH6hj/7FZ57JJiL3niz4miOLVLU7qMoV0S9Zx5tSELooHBcYPGZu7RbjttVi
ISaxzb7NtzDC6ga3JH2eMiPUCwCx1sj1I8E7liyNp28abs3FE3hACjIY8xRlKP0+
3YEdebENfiwx7kUDfJO7smfFgeIa804jjmJxEUqfJ6FAWc+s/FnLAw0+CsbUypqE
7kNUarcwJq81Y1u9UyrSDYYZ4gUoOAngnQyLEuJ3CWCHRGr3rHH1mJ4EtboTsEdt
c7hNHMLljKH4P/eqIM72+2iz9yTbS/qwyCoUdQJH1b5WciKcGKU8mO9RQaVNMg7n
0wgZ2enMsO4wwzr3LdId1jTnjWWbbOFfN0W+02Umj+0X15YmXlqAs+7uTzeOpBb4
WGTnvHUDkGYvVq6Iei3yJF7aDuCd4HrQQ2bpgUpdCtpC+cIgymOURHyx6SMaSA9c
vGEwetgZ5OankjPw7VUl3IkscQMjBI6OJNdI+XlAHZ0cNtASvfBPFseMerRV7cw/
epJw89I3ci5f0pyiL0M9GlUwO3sqCzJ4ebt/65/4MgOg4Wr3Kn48HvAxYUrNqjcH
ZUQQZjVmsfMz9qS1rFnOiMgj/rpaKPS2sh+C1ReIS8SO1RsUS7PxL/Bk55zDGdvb
mO/MxK3P7ysZi40hS5wTYPllvdbPBFRiKzyXKuehxDMqCSferQXotrOQV1+gTiXq
Vfv4R5XoxELoII5kJYRbmSio85/8rcusu9OiC3PvmAN7N4L1lFogFUIOZFLj9/pB
iW2X+xfyANWQ9JHcAA2yNozWdAbzlejBmNb17m1VqqgJ7HwfyBRvQaq9uU+Da0a3
umH0sQN3YjUL0ozHdmbaK77Yso31gxKAJovGur31nKTU+WeoWZMdO1F6YTyLh7IM
Ajx7m/7eDHT4fYYb7MeSWKlSxP8DjHMFYeldESlEBsyPs9Kz8ERx+98ujqgtOqo7
bVuc7EiCZTPpzXKfWg2enHweQm4o9wfktq3ws9Ys0yHnJsys+YRNTCHrcGfCFXIi
KO3jj2XvAoehL9LVTSCeEyoRV71efveivPuG6fRidZCXUrFj/46gwwKoF6btusmp
1VbSqNHSYLo70H+KdVU2x+39guhsKhDeTqqrHgCUtaWnnJki7y1Rhvah8BjA5trA
SLmOMHOPU8+HivzJTUR43t+TyAVPCu1eeECArYxkD7K1BEUzVMOKU5fvAsYHMOAP
UUcn6/uTikrI9ptXUDX6Aw545si1sszji2rMGizfgOjZg/oc0WdcHqu6kiyqBFY6
aMT/tjkNkKZXK9Yy8PXhwTA6OV7hWfzSQGRNMRq9FBzbZ0f+qJ+hAO0/ZHauIOy3
xSPkq1UlyvyK4PAeVzJGaCjLiPEBiO3t4AuB0AuV03WfzLZg13ZKC3Ytb7XXwUZo
`pragma protect end_protected
