// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
YFXKxxo3Ke0dFXQdf30NTFl1Dd5lvtVQtrU8H//SqG0NARzuNragovPS1rZ9lIiLKtU3X35OgBe7
rI/f0uQX2BCfM+I1sNQY5isMR7Amq2lhDfSZq3M9DMj11huFauaGYHE8qCBfRUpOzTKPEsj76PJu
Nu+ac3UagMnshGntCKwh6Re5mqqaofPBp3TvWXXkshwXXbbW64U3lRrpyEy0TeU90RjS8yYdwaF/
QfdnyXLVzXpx8Zv7INFg6dT8dr0oVju95RWV0s2xq3O8sHW1wOJyhxGluxx+DGJG6l2KiTVTXINf
m3Bzd8KYFeMcHiFdwfO3GPr2fXyVFlGmsvY16g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9440)
gNcY2IO8oKFRUir1+mb3sq8vwh77u3+ZS0DqcNj3XE+Lm64CJr9LF58C2OqJcAnBBEOA9Zd3L4du
ZpmEBm4FzY+aJ24BrGxWs67g5gFELJ9xhUgIgNT6UP8MY1QFmUxQpC1jc1EPucN8gUBopSnl8kgD
i975b1SgiscrWVvlMtWV6e6mJMP2qTa0pLWd+BSgiluWrEz1V4vvdpyCzO0omDtNagnHYQnZkxvI
h9TDddfYJsE+aTYbACXj6IjiEsmYZryxNWeRRUy4oNL3eP75O4OL19Krxj9Y2ZjJ2YuTTVjD5wGY
LLIkeC13O063zcDEjxYsuVPG5hLbjUr3414GZRZfKdGxLYd/HBgj2SqtCvhfrh3hkPTT7GlbkEjA
2778PKrOIQn7hPBTsA/NHSzjtm50YFRdvkyEa45rsntQknYKH7XVmZByApfuOLBnJeV1vK6wCbYI
1Ikc/bV/RNs0Qko2iAnf+0QTpCroiRWz5MxS2lfjIi703SENNNvRXriv3UMJabxiopZhXt7DNfl+
zLka2zZDXOtAVC4nLaamz+WboGQqSngDOJwTepuwgYU5VU4YvaEoELBXQX+4YGWdcl5Y3lipOGKG
taz0yhCsf1RIPGbohCBWrQWrfSGms+4QZIdFjE/CZtbc7SJ4aEwR+HCfuVPP8th1MspCaHMaxHQs
uxhCLbMLza8ZwHvoAj89hc84RDqR2sLJLFVT8jdUJeknvj+0zDQ1ApkzXGwVMkjnJiTfaTCi3XyB
eR6QnmQD0JNymCqszE1qWcjqCiQW50QNscsZjO4LVker45DU8hkuuHQ729LTguR0BSEqZYZil/xt
QEXTtovPRFp3hF5TzVFvQQrfb3lh6sHyShXg/lJyKcbE5q2WTKxAHTk3QjfeZ/sf8Ocav5b6HJZN
coRQ/89SkbjfiWE/20d4Y/VvqlQahVu/H7ykchhwEKG4/Kz0CrodtkXZGXOVzUtalEeOtv2cAOIw
wNZPJZ4mMtvva4sUL5x93fo2S+eNJngVkQ1PuCTwyyyBw2ein2MHyZ2CniKU3vc6lEImyOH+2j62
vIdhBs15zeG2CUgsyAzAgd5UESNiGqk3GwOTtkNdicXGf34Hc5KyS3AJl8KQCWrqmLuQzNOAchrD
AP+DJJnatYDjqpJMfjb+hTJ8oB96YpUmqlcbxFn5t2SVcawPDouPFIkkYzRaH8W7U2EKojOgkEEG
GFImg4EIvHtDhiVzJJq/gqR0C6Q94S+nnt43aMSWm/j42WiIG2DHnIf7exTPCNCBIpLUc+e8Vsgy
XUBp3f9jfPIujAcpC/OANdkyKAKt1lbodCW75VUrbf470Rie4piKGWfJUwlDMgqtTk1XAQi9BoT2
YPS2JowtEK7xKxLjdQpkFbarPaYhj/Gsw3O9di9Qh6Jq7RR3Dv8gNHxt5u13+Ir/5I58aQ31V7Jp
eVQF+tXDJ1KIdnoevv9u+035OisAT7VxCaqLMQYykNaGcdT9CH+tHp71FgmP8wRFWIjHG5nMs8ZU
gVxKtMtUngsUF8dJpWpUZiyaSabrVttL556gIVyTHWBTe9UcwU5qHl2NTyPArAoND4X6p5C0UGhl
bVLWP9zcRxXnlMxI0PbXKytD4RNnDuY7XqcyW8NPo64ZR0uf9vmL7SninYCxAR7BpU43hLnlqzis
u9Oir/WJO3JV+Aa1DKVg8eIaX2sX+VRj76e3F++5VmRv86H+PNPDax0dsHvcempgC7buqFPJ5wLg
tF2X6R+LNadHh6sil4dvqKfROpQ5Es9LQxWQZrtgJ8bfm3MQrGDUTt2entWuhSxwBNJp008hy9C4
RkfZs7H2H6UI6/cYkfHEyH0GHaA1ld8W/MB/F3tNy0QruHzQwj6h6vlt1p4WVf15sN0u7nuMhEP4
uAFxiM3MN4FshtpTTJRPVR94AsFpOWQ0oXl10TOIP/r37KhYj720eAl22C0p1eCb2pW2fvNaJez+
Ry5fhwuP2MYSh5C8oz1nvvv6V4gQOgAY5ufLRRY9K64VIC6lZplrsq4oGkp2EeD+yNleuVR09GtP
VIH06c6CGu7IlK4lN6WdynGwFb3vLn7hXLV8W3MF6iBKA6bJr3KhT/Y1Zufvoc99MKmR22J7bpqD
fgwTFv40I+w1C8HZ5gBt5bmrytC+3XWoipHD28msPwvNGIbgVnhitpdX/AiXk1Ks9cl1o/4aSV0/
M7tgAjz+tdM2L79h5nmf+hoe3PusjyrHFfLTVU1v6lKqNxm2N90C69LnRUkNCFq4FdG9h2stYZ1R
BiCq8HlZNEmRojaf5zTyu0YItghQb8+DzJSgJNLPJEfHJt3N7xiDkq81sgZ1Bkj4H4f8dRcpFNQ0
/PbZrk8VVzd2EIAbj5ZHoA+Sgm8M2Di+SHVCuPOLzmJvqe8cyu4qE8BkXhQzi2pcdDgPLg9dPB2Q
0J4UHm99bpOJnQKr1OgH2qisn/rocadDQBA+lzwsX5l1RXmtZajJc+S6fQoLccPapGbO/mOLM6sX
vnLRXdHROMhtUvOB9CDgf/+zKmvfDqUuKKEy6A9DAVK8F0jp9ECcxmzNuwLqOYGgTjyguoiHqP/E
DMBpGi1gLWJtCaadguZMV+Llzaiq4B8GsfCZcWl7/+Xl2D2osqOerKmFLq5mQLbOHJCp86xxHU9Z
DNf8sVo2EJTQespXZLxoC9h6BXPu6/hwN+9x/HYtWyj3Dkz8pxNHsmBafuV9wqEAChvUgpa/Og+d
oPGnEPQVB9rJcDDDbxoTzKW3v2KVRrQMQ65EorRKRcKupXtEyDsfcKgLgKFjntIlPu9JfYpkhuPg
KOqLPUASN42KiVEFGmH14fDxU7qbeBfZ1zmaMuL4lKcM1xJXm7uilpZQVkcDESvks7k32v71TwWu
NI1SUXQlbu0aLDtglU149xHVee6UQgcPawkr9X2uDdw1sV5dXxs/SMvfTRc/APjwBC4+utrbpVek
rkrUahWx6IQuuxEr6bPQQZZK8m1p4uqUr4f+dTUwxExkdw9PXXTnD9cGf2KcfG2WakLbzHAImCcr
BOINECaC6lCFkdfT1iikuw3KVUK8nusVygfyDKI1U7Qi7kmpX7cLA8eL1+04NoJr0ijedXWs2cba
a3C6OGbkqOiO5BHKw1zjS7DMit9SAzB8q7c1YJaZjhkErq8CJMSA7bMixryOOMk6gLOrS9PEDV87
5/wRh1fELcytp2gEFmW6EHy0ED3PvFQxVSTqQFKcAljMmG+1uRLJdeu25A73pMIajDshzAMzzeLX
NGhrA6DalW2cZNGnt6qpBTWBCTq/yyzwwK1u1nH9scbat5EhoYI7V5pHY0wy5oCMOLOagNftV/Y6
tkPjzYSmLVfR+Mi0/GAmFdXHRRVuLOrjsxXLhhfEgmGE98eHcamJJdUcVbIHgI6Oau2PaQI77jU+
d9f4CZk1m9sYsGk1KJSIao69gDUO2L5455W/nbkfse27I3m3ufdPSlnOGWqtkns/SY6KYXuWitt1
aYivUc9chO0jpwCqNHBccVqhL2cHzQrNCpv8gbfwCnOc/vjWndFTxAYMWUYtnZ3TGhErwCwCDwXr
MGOWf/En5W86Tqsq90RmdhbsM1z/pSIke8S6IqNL8LPQkh0x196dJxqK4EuVESyTLT1++5XBh5xd
DVwF3o2fNCXmgCYFC0TtPf9TEQnXUdjuwkmW3LAMQo/BDHH6UAX91lTWgWu2S8eyclt8hMlbAvnH
yQQ5ZS+sBGhEsgB5vKEiSlQ2+5WPsXnfHQxm+7YhrMF6R1rIk9Xw2odu/Ij1qSJqCMJUVQ93la5R
HxdShqV3KAfPfv2fhoiXb596rMQTuyevoM4fGRdgU/najxIZlrFT86ItAs8QfEffZjpxgDwc3/TX
uq400J7zO3tY2Vw2CSxaRtCtsMm8KbbKtt9MAfc0B11wpYyc2cXo6Yn5QPJ4nKF/zF4AbwZH/UzY
UDJ2p7BMxmxJgvw8t+wBoWU+VE9BHwWk00h8FKVX7QcX+35Tv6zMmxqamZhzTjRkKz6W6RnQw5O/
BnRlvCfe++Oc+DXEAbtGDZaqMIT9hNj3+gHVKvXTPOOIyQgrRICZj9nd9oCTcs7rIRyq8Z8K+vIt
uw0wUeOUlC55c3i7Zlux9Zfmw66OR98/9xhY2eGtLNKLpzudtHVqSU/vnsS/Ml0SR8vNN23bmksP
an5dcWoIufZNi54LCvQEefmYw1/m+rKZ6Rx2tgnnY6LaOXQevJvz3jE0itdRrLp1l2XUFiK9sP3g
HS57FD05momM1DE1EAN/slL/n7QmEYA9O4aB8ADYGRC2ig8MXTHEUeqv+eajPhJQ+pVrhLWzKBP8
Tv7hiY9VxgjJnsNSw6qREv+TDf1s1mnCAhVKQsgxuGqBD3vNfmTM1KlHo/4VL55/SdVIaBkOZSZl
Gci/WnnkP7OfOT91xE1PbadveWnHvUtsBq/22jJMDn/wMvldcRZJSOl7T6k1hsas1VsT5/8lNs6X
15UOSotd944GjAzIDQt8x6XA6ewAeUK6U2J9cGDq8Cn0FOzpcp8fzveeggx4NkRBZGM0CXtlNC3R
m6wqoreYE9FO3ukKwN67axqfGQzOAHJeDPuT+rUojzAuhyUb2S38cwxLwAJpkGzihH/Yfx0NDd/+
cETlXZLViXCkA7jVJBvNCPNJhoEY4NJ2+csiTE2iL6RERvqMvePcxeOcL3gmYTT0C+7lz7qRcv9W
3B4biWUAOmoxRtDx3fdbdHfLFmfzNC2Dy3qb08CxBzEisff7eSLvxPbL2vGmyjDY15rQ76cj5dH5
MqGnDRfQFXFW5c8wrj2kbmnXuFW25aDMFH413yF6+P1NW05lh3N3WhYRzK5haGgxXqiuGfVkYtj+
NF9yOZwCco3nksjd5LcOH3z5Z0xcezOQ4luRelUcJmwdjDcRI8Y5SEnFViffDhs6kqN6+ZD8x7O2
X//Xb/X5FJvgPKyIeYH9f+uqPL8xU9BxwKAbz0jJFB9N4DXE7r04iZM5jxWwtmCj3VuZU+Az1VrS
0VoeqcRJ2Z56aZ2Ca7RNvT5e8mo/pGHojH50MoZbx6ph6u21OgHnneq0XPeVsLLAMT+eqAysWcKY
PqkmeAi4v2j9FHsivfqdaciIYF2BUjQkQwsJ13MakgXzkhXH4URf9MuXSH+Te3YxhPt9YxqMuwC/
9qpSZpsdk+/GOSOilSbr4INBXAgGjxwVP0NUQlrKTL0LDFVm2v4lNrbBpvEnlTL0+SSt9oMiKJ9d
aN4iarEMQOxPprei696+5H8QyeA9whjOBc8OUjSXGHRp+H44VD96Iie8dZfVk+Y2Q3+Jl7HDxXk4
YSYPMm//y6LoKUsFiGmsGAfW/ukigLT7uQwIc1H0MzR22YRxFIIQzVfwviZHKcoWZYPQfG5MtYG5
QNQoy/gHQwZnOiQ280LFgsfPa0KEi3OZwXQtaAmsN9/wP4ZgPYucPZ7lwCiRcbHpkY8lLsut7geT
6Ug+WVa2iDzl3QKpOxLDRjHR8/ZsKZOs/5wF51kmrCO45EilQUt4gl/4x9kz1PfExvR2ihJ6TrsK
fsBRnWHnlRL4rEejMeCgPmhE3byj366H7NShfltDMDLkfAcdX2CLokJOCQS8k2THW2b6v3XC6hFk
l/UsbYjWoGfyES2QQPAIiMoZAKp4bSRPFjZOMlUoO1vJk5Tr2ghoVzkPqcAkms0QhPuiLJsfs3bx
gvag6RXUYBHgqZWmnZHDzgdIxZ9aK3yfEDHKv2j4qFzejVwWg6RdisMWNmIICyJ4acJnhx0eoVku
so7OvFyGor5q5idc2+2xhidtpPQaKg/BMHVXdgRYH3g+Faa975CWEFY2oIKQ724w3U7C1mqdJI32
AqTY/REdLurOiJPfW5GRugxO8JgQ4ZtKAMWOd8yb/L/UvVYPc4NqsFaZ1pvxcaz2hc/pSA9p6EaE
QT2lKLw/RhAo8cnYnWtp4pNR8l7EPrLvrtL5jG2SY1jQC1Ais61H7oWgdeGbiwupTPNMpKonCKT0
HAvQqwrcWm0qqfC3NF33HNSK6AB31rxsyErl5+zIkFP7N8kLDCocyjBmpf72TpT3e4KwFZ/khwta
R8SibHcmeT1IVi+aUib/FbZYmOADVcFPY1cRm2qSz/5V6bcHP8IXI88ZwGanUz0DpOZcIyMzFQ8r
4H67OF63BWmbnkH9ZtQXLuWltSUF5YAvF0wAMvPSY+B18sPl5GPcxh14g/JgKEua7UgH1dKBoekn
g47ioL3Tw4DECrOBnaP//nUfRQgA15peHZrmUSOL+/SpVcW95oCoR29yItLka+3Bj19l/za3+8O7
8emt5P/dzf0PfTMCYJsIbwUR8j3z7LL2ntSOHc8LYpGUWi8ID1KsnNpsqNLmaAR80yITaC68eqlC
9IKYhgSBwpeKLxsqWR3zDm7C8pkC6/n732SMh6O5Xq3qOP/RUM2YMgatSwLx4EQCHu5VxmZreupe
fSHVnIvH2zufxXZ9AXvBWUllus9Dd+R+8SLhkY3exkK6XOQGU2WifQeGZX6UELy+WsMfGY2ER4bq
46o8y90gaBtmJ9gdXdnvkhua5ZAgJtnNyzSfZWl/QmdihmKKP7VZcyYA/jhZoJAj3de6iTLooai9
p2A+P9F3L7lievBSBIjb0jRSvTfm3YHeil2YukVllmd4PJ3V7qiM1iScNTMROEsLpOVsiS/aFQNA
ozcmvaVShuHvJymjkB4bigEl3T302pTM6XtASYtrvRCSaIoKv9eKjI8ZYyFrf57SOrho7YCVaPRc
X2gE0DjPnosiu6tyig4hBd7prlYUZ53Li/R5qB3qSATdBt0diuZHfEv0KD9p3cyRCC3rkzcCerol
mzO1eRBkvexqEL55WgKFAy/j2byuoYj+VVqLAVYpDiSk3wNPUJNacOXHPziPspKfByd6nPaSthm9
//gnulXvPJUP+1luDQOSmyHTknhbW7c4ndPgDkZ0IRzGwAWiRW2/Nma7yBZtqrN5KrSACeKAbcla
TUTomK7g+3LgrNEBBZO+CS2JfxbQzkLrx2GWkb9Cw7PeGd5SrIZi2S9dHxcgwPh6k7BEZNt2LlDi
sIEyEZkq5t6M1PSvNaCdPzCy+cASbe3u5BlfqlhA7QDQHUyQqiRNtlInYqO9Gf3hAblGlpu3NEsA
u6ee4jAzrmQyv+k/UdErY7PVFGXEkX0JNG6zzRb2SLMXWagigraFg1YFCrW71L1vpkv9ukJzA7jI
rojxRjEXBYbYG+RmNBCeLgvv/LPI16OLfpp9zOHm6atuEIEFy+0+T2+1CVOmEpnbbOUz0kZCkGCY
cqGbAFcETC1v/cj7+m4DKq8CW1T+k1RU27sQya7NIypaACSKj+PKURH6s2/k+MCPakAHNxXsqqPL
wGqHXtKxw7QNoQZjUTS88H0Uy/Ch8dl43EyNHT6YWgZoeJNsRmwI/lKlVduxihP+eyapKLHxWpz9
FdsNWJKS05MvESoHYeVhX22xM63kLic1wKQ6gjiLY4qWqqQX2IR346zE1E6dOKn1o/PfRS+3QSh/
uGw7b0vFLMQqA7OtdpoSAXC0B2N/O83kJO1TezPtmOPiQGFnt04H3F2Dpri54euqHic5K+VzfzdA
2Ov01C3fOxvYlfLugJ74eeGwz24P3vaONkJseNLsYuaLY2XoGmddV6hwGllQkpMhOlkFIHq+nXUq
CjeGjenpDS4wS2vddZocx3dJJTTUqTDkQAr/S0BUDkgjrIl9a9ncZMsF+Nu5dVifrRdKVUkuQ4IS
SIRfzWxVt/hwrQQsUzmBIi7iztFkbbufWPOIqSqsryT4uhlDmhces0YG7a6CA9PVPriGhD/8b53i
F23h0b91Eg/xYrnlSpdmN69Z2PtdSw6i3W3vJGnZYWL/iYd0TAfE9QZ1+3Y7c+D4U2JnJav+JBub
JIvgrJM1hkI0kbtj33tEzjQVak3QFsxmAvCJKPIbGQyqxT/DHZKKckJYaovGa5xE5ilo4qTRNkuw
7sFXH5Vz6gKMxh8OL+MD10APaeORmp1uCCtI2RCT1z6Vw8x5lOSp8vu3P729ZXSdzojqx+ALz3BS
wjc0Z15d5FzkxhXd59EiiLiGK3lHY5FDE7wM+HMIkYSDpXdHUbqmJ+uxjJarweYRzHNJ96HssHHw
dGFt4VhCOtyX7vSb1NhaHWH1vg+aOzTanFAd4Co65YLxvwVSgKPM5bvLH1S25QuPqpu8bUo111zF
XvmAbYdN82OcEIWezuD1kMr1xV5jjqLjBkPDE9/jAdkrojfYD5oaN4EWhQP/HZGI1AIjOp0XUKRr
JUUwyPccoKteQ9gATI4X+J2X3j6kdyAqkbzO+Lv/NgXuK5fd7Gu4qwG6lIimsHeR3iTniTy0Jm7E
RGodQ8AEe0I3uPsJpopFnpTC+EA2pNb92GGH+DqDw7Dm9teHcNgCvaV2WaawZzsd1jN1bNMSsq55
OjQf+jP4plLo53mMmm1wWP1Wx4AGoeSlGI3L3dl+In6wIuLp6McrQzY6yPNl+SJrarqEcZuc2AtL
TnRopp0AAp756N5xr+wA0Z9brxXEhWz2AyG7HcCqeubTF2mimRgztZ/uowvRHiLnDq8VVrA0sXnZ
OdRd5KMH8Pq5/kIJIy0vuIuS7a5Y5G38+eG4dkzTEv74ZinLkomGakHWYyoZPX2p9Ox1R3o1uPEO
zIBab3VDu0Pb8IBj2vOh5jp0AT1iL2JCWugFIjIw18THikoDMmsYb++MOOad5PWQQIXEwoqk0x12
C4gW/TafcrNcoAobc0Qm12pqRZviDskKKiB28wr7kbuxtv3of/DSD36/g9h/qBdPKrBq0yLmpVZh
dIdOouJa8W6za8LR4OWiXkdtU6YBrTWl/sbTJR/OXsPCZLQKbGuuP330NkqDayBUAwObjxxNjNH2
lAl/oQFqqkDpAjb588KlxdLF0/oIcKpXkm2NOvT0IHrh8EcQU14ckRmF8hYrH8mya3S2oqUHegLU
2A2ADyabTK1sM6eS7oagYe825Ee6vj/XSNr5BXo9rW9h3jWaIH/ITVcWsBK9wwDKchEYIrAMfrFE
ZmuYumJZilhxFFt7sA5FXFFDCXJkxr/Vn9mk2iZ/hpLKBDF1YImHsZ8rIM8DHXodpzdtEELAT6G/
XLyRtgbZ5HHOqVb2wJHU0S5zGbwDqGFTK7Tz682GfZzBlVzZDfQwR8bzfKf2yUgFhOVbcc8xJM9u
vcyG5TT+UbXdRBtw/tQHEHBeks1/HIt0BdyXE/265xAj3XZu3P21T9rt1af40n01qwW7AX5MfiY7
LoCJ2H4bwvgEYFvjlEC88KqLgd1X63n1ALpt8okGtW15c62vAs7w98yuv1tU6En01TsC0RfG5+AH
9wksWIkyCTK6SoLM7h51yfiiBOj4OHPDY/dCYGKtXEASAYBh+19KsI8O/YuNqZLCCaJ4gYKEydve
gHYYSqu7FfJQj+m3a4ABfcV0iFx25HKgIdGbjXGh+4dBSAvWzbZ5EdpaSnbto19uOijLqnODGCmX
/FnFhyIC0MrTfQeWz2XAV0Y1vfmeGVJ1rrjpRfYPUT+3hUtmhBEEso2CZoMZ7/+46UOnZBufDMpp
hiABNRZStu8UGdUft2Vcz4gKi2RRMvEVyI4fXMoFXMUQ/qBhrYG6CJic8DkExNoBbXIE5Vy0uGJw
NAE5vSctUK95FeNsxJp4QH39QU1Mv/scKR97051ogFMEPIBxqM4nmXV9lkDRXtRw/+2mvmFYddIX
WQsQ1enAC4NbnoZ1jTaMubNkrEZmd0SpCWF4AqY+eKyF/qfArK7HDqb/2L+/NzQ0o5pzU3VqSl3J
KEfGXr9ymAa1H9ucHbJ9TRRYApPVkNXbfV8LQheeKzOQbb949ycDMZ5xVQEpHlgECgOUzX2+RyAd
Jp3B3EU/k2ajUnch7I7VCu+ReFHBiE84KSFJuAdrsmqD/OhizE8MYxThCAsunFymWd5MVdn9Zm1/
aKGuddC45Z3oNdF8dGjQw7RmTD9ggvXmAWDHeol2UxyIqudZcdbJ9BbObUyHxRFvCmRwhF/dj2tw
Oj9Sx0noTx7WDnzfYp7EXSHy+LhQfC/STZBJ70MeFrV4ue0cBtUVd9tRpINEkpbxGC2SIPE3csBe
lBU7hbjdGXpoxIdWjO5icBtLMiZ2rndQxjbhFzRvabmIQnfM0OQT5jaMezyXRkwFUOu9f4XpQkQu
BAvf2XkPSCZn9rYhNmZ31E2KxbMLq4vqMrfgxRuOFAaRoyhyCphqS7N9oME6lKzAnAsHLCh1mKHd
IQKpYig6EhXzOUPNXL7J9tsCUIxgPG4oXILFENbCP1oZJmmzTej56EzSXoe2TgXdv0o0h2Mg4Q4b
+gz9cOHJyGyr3+HUuJ0d3n0+JNcml9l/p+gCaDDby27WMOPkCN/6qPLGTHvdZTIEHJGQvjhkH5JS
CaV1rvgKIA3ognfDpX6U8SjoDuL5rEmUh8Vaxgbso0HZaWueslRoJe+DeOq/Vgjia+OTHJjGymr7
fCyFxgXflRuLGuxLL9ij2ZAF4qCdrb2GbyJGNdTy5EW4eBJPA3DCh3elTGMCReTUMhCcLwqsa2cX
+G+8nR0NCa9ew+6/pZon3xdflkAhbJGu8iGfS/8hFgV9RPLzeud41MOFpJnPzGMXLwp+MeT1wfIx
CsYbbIZ9F/I049OOXW62mpBv8p8Y5C3CJA388Qu0PPyU7ZNnbOFMOXIZ76SBaqxU7YwkY5egsxry
qZBcTlqScg39aOjodhsF8GZ8uj41IHPwcOibEgYnIPoMWNLLhaCQ9KV/sh1yhgUksBQSemYREjmP
TfZ+ICA9tnT5I3k3HDiq9EMA5i7ceZJvAbmxWx8uiQXycET5goK7YYPr0L9pvDL74WSSkpVgQ2Ju
53QuEQN617bi34GiW1oas+FW1YcreBMvuHvd9gImRHFCIQoTRf2+KXgE+rFlWUlZ4YHykTrSFAwP
fD0ObpRQM+YCw/R2Gl9+VG3mHX8COON22kys0XdfNWAwDL5DbPdQ9jf/fA1scERgDQPdkPOphE6m
be9WSDQBf2FeT3C5Y1xZB9kcigExqlwZtJqJEv8ruppVVnJ4uk5TA9IWUKKi47lSqZohnHeUkp/B
zBGrhmVKDPlFoSQzzdfYEgTtthe3b8ymp6LqfW8cCh9hH87KAP3K5ou/BzL/OUChRE4Zb6QBZosv
aAZkiAzzbOusvxUvA0w6RH3mDAFjwmB0hZMSG++fcHaY3Zimof3BJU7jrW5f+7+JYRi3Ol2P4IRE
c8fAc4hTyTE3SONkZlhaCicqc9Omm/e9fK8UqmYnbCYdyB3AHd6asaFTy9ZTSKQeIP3ayN903eOn
Z0z9vDSFmelOE12+jwtQ2xsFaj0EmWn1wiPpwDUT8eoXItkYLlS95TMw6z5lZ8oFALR6Lmsb+5qH
aY9S1LqlImYugVuIPGYSxN8U8xXcq3GPJaav+Lzg5kUPLPhkAHj+NSXb8iZZl+5JJ2LTsvMD/Ieu
do/oJx3y4nGsX1aGO7lTvhopp56sCwVSPOHfy1YVh7rUyvg18h0jbqohIpapvJlD2IknL4Q1wQb7
LCqiQMvWI58yVdlYRnKswxLAzWiWH4TxzlC7mZ9oR3IGaFFWFJODNeETv/VEIw4nqRG6Z3R8fxkZ
FhxT/T6ZlSVD+cS6lVdJcIeO0Ql23p+pLRTZGaCak5DgTmekMiH4cbLh8rTe42Ys4AuFieY6sqa9
UR13LxVDChQUzZd+eO9tnxSGtT9QVyV4HZR+NfJj5tXoz1swngtOZnuoJmNKnvs69TTeuxl688bp
ll0/bGnugsZ13oOAiGHshYXzb0EpK1n6zaUYLd8x+5bzgx2sTNwLITiVrenktqUc/bRXQj2Thbtt
rgTOkr5VH06yT0TKXc7w0Lcb/6zBZLMFvzqKbLFYKc9pq27AYod17qLSpssZJjXHxpfWEHcNO8Nc
SaqdXxqUTbFbSMyVLwYEDOc4obWAtrhGaUkx85H0N/OeC9escqHrzu5hDDZeLJ0Qe4qp2wX0tIaK
4dHE6fbgwm4P2kIdWW7QJCQulImE7WlHAel65O/hPF65v6YZWLUMs7b8yB1DOc6Snq7f32s8CWs1
QN9dlVWHXagmVqYH+POTtUasiTGcBfbzT8wh1gFfnSO1chg6nU5FbqeLrMMqKEEUn4y8rw73WT7c
gW/kvSrYC46pkOduhx83pLLubHI0366+nR9DZu7bZH7Zy3IGRQK8BnTHncJ4PRetu1SYoTmk5KWA
Z5jybRZIMUZ6pQmbGh/7VIb019bTMwJmyTYQMfhz5tMDepXZ0HOXX7eb0oej2mla6Id/g7KFemLt
avMleyTrjxKA/18nySPPjLi2zdRNDPTL85RBVMYWP88zf9KWQgNUMX6oEHt9nIJDre+n45tHMirh
7e2CuUv+T3ojP09MGFqiqYtYxFXuXg/4oeqck2y55M+GSZnYPYSIor2NI4E0psiHF9C+6crgFaHK
9AdBtYaa66DmMRrsp1FZAR7SWSjCOEwrfYSQ3sSCbWNsl4Nh/IK9w0K+t7nJG9IrF7zJv+z3MgpE
dClitvmSpc621zTED6C64K8w4qWHPQidcd+vhB3uvsss63o=
`pragma protect end_protected
