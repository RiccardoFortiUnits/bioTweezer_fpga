`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mNLnUyAXHStbogesq+azlNRYeIO2BrXSru9U2dGfjizY1OwBnzD8MhHS7Sd3UGm2
OcV+wO9hWSPO5H1czj1SxdFDwsakdELb22gCHmigRfOK1PhzCJtAQSSGJK3wIL/S
U7+6IyzyXTq5wGttDh26c+3ikSlL/pBDFEvxmJxAGv8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33696)
QwtdIUAS0cp7iF4OgZsSUAabMoxr/7WU18ousFul6u344GJ0tYI8u+1nusdjajZC
OWbwmUrswcq+ZjMtx5CQ1RJfDyPb/gAXkc1b1vjRrMXtsKYqE8a5FmrcTcvG+LPl
ZBjgudiXQ1uhf3zphf0a5oWIqIWF5556VZMBlj7T5oE3k5P06nzexl6ZKOinLDAh
3lWjijGHE+UEanoSFvNJLokcHfE4XGnZwGAqIZyD3syoglD5N+rk0mozaZviFwuY
rmjKIO4dZ6zHLesT7KqKnZkUwBINr0GqOETZHYDjQmdtn2xJbqEh0GzLEGmrsh4f
5oexIXo5jnd0zmsUIZyg6yDJZXbFxxifdPsenCxEnfonIDxVD5NYJ9cqtz5xKVTc
nwq+io3vRaiFFijZEP5mQUBRvNdhOT5SYxt72EmOSOsnucywVjIJ+jnC6Onsu8MO
cEQc88nKAdxyBehmDPEOM0ZYvWC8DWw7z6YTqwe6XyvaJMgYFiZjzqxMBCP9VcfU
kbDwIp+pdGUj/NE0UaujrnZp1TTsJwnUPznRQOTzp9jtaBGVJAgbZLltKEwJAMCJ
oF7sLN00y5C0bjWeAjKCmFyKomvneKPttZJ2qTFFJpDryyhwNwVXjSg8qi6/QkQP
R/VkDzbYdKLqF1zU4j67iSOeNQNzmyx6Om51hzL/HZRtJzp8Qyz5rHA9Pbk8QUns
V0ghbh3TpuDvZkmcZlll04D51csOi+aMvByxgFlUbesAIhWAI6apxeQqAEidiwXt
m2LE8F5mzYfbB0rcALYo1L/9+M9UZyQIGh/Yo/GN3BYvC40Z84TAVGo1+sR1zDX4
dOOYFZ+kLZGUFKacn9NeMAK1rpeKeo8OBaLTN72bN9rGzlLamuwFhGFE2ftw5uZm
yIot7O1VUxV/6ECPNS0nUDNdGKqAvSnCphrn4TG8AJiROHhcQS6zXIRYwL5wj5Be
xWVxvDj3ZIFoMPPbr9LAY3+WPI0Fy3I3tIiGdGNeONRCNv3hwaj0P69vih4RPAkr
SFmURFayrTAkDsmLLEUNNOyQ9C8P3xBotJn5QTi/vW8y2lpXnQ3f+Kl3etyrDCtv
XTUYB7n+kvVDOuIlirqApNNnlAhloGtdZpa2Ktmo+ZCIhBNzs0DWIT385TSIWgai
v3XJR2j2Nq1KDNOonw8UzNXG1eMTJ8tuh5qKvkkJGvsvN4WT4POhU+xAO+eDCski
+fg05xYBcQRHXpbEYenQbr5JgioeiuqSO9pDq086eYr9Nqc2Dv/4m91eu8gvdEV+
/wrTEqCcw33ymijX+VQx1qq1LV0tM2q/YZeWRcTzzdzT+kv7h0CwzEcRWfFxKKd8
8CtaUuZf4iCpQ5mjoj6P2w6v1wQxJ1VF6jSekxKsWJBLLF/4RlkMSKJJ25ht7VXp
duscPurL5SZvGmo0STvZ8jal5ntuhI7zrCqUyB60McbkX3tnqkXo41WkCwjyauOa
EdfeQBtfStfxAbyBQzSYN97LEvf1lRhtPGl+mdKokn9y7kcoHI1tMs4zuZjTFJ1R
46S9o/zv8If1br8BNd+3QT3FwQoTpEZw+2zLjuCc5suMfQYU8602OrpQdYWhHi34
CMfnox5GZZ5wAksG8rPDQXaH5QhaeI6syjKDXxH39Ar5GmX9Gc7A5OVnngtOWh6Z
BbhOydK8koUm4DrDtUNBoO9+GdGQCx/2CLk60GQvlfd+8avgXlgnd7bhb18no9sa
z7BSudZ5Tjgr3/diP/KUOG/vhixs9YR180mslC7o+xYdHk9LVXgYfpRH2EeOLdfg
7aYrsblqoHWTKxQV+Tgz1L01Uzc/z2ofYVIcGZZ/kaktvugcpzzs1Y1j4zdUmG56
xHi+RARxyndva5KaWYrndm2GWBx2F/484h+WhUmkQmcAA9sLLfuhhfkDORDSggvF
hedDQAXk3CW8QO76+IeWjMUqQS8RStkzgmiIXvcNcDmu/zNEfCpysFle6Sw+vw4L
z0qKBRZn1WoB1AhFCSeTMlSJ8u8iwm+ZZV+yXK8sFCsj8JezNI2GiDbw8MQCNRto
zO43zrnU1iR5Gcblm4OYnpnY/4sM4RGmUwz3TQSk424j/97uzNIqzdhD1drMbH59
sIqtRSzS8SwiixKleonQXzewfhJcXTaggm6+jyKeeACfi9S/AnwtpQbiJk73rga/
6F+fB5nF8z2ZoPZKmFQrtjnfSls0e6uuN0fpzAh0nZwA7ux0l/X8LtVIAj+BSast
bjFp4xMJXXK48F+2Lun/fRAy1KY00bl3csgFmu9Q/n0b5dRin3NXgrAUiirX1BzS
SoxtDR5IeDc0h8SIAiJd3Lgw6/kecyMiKnpeYPl+s+xjwvVpXlnauK0wey9BI9FI
8fqnHzqWPGMq0wNj9uyeJOVHClbFgUTVzIAUiyfbjyGHNIJwXTOkj+oL+xxt99Yv
Onxl2+Fw3lBYsUcVH7RdC+mBdmuPH1wdKe7718SsmQXGN8ZqU90vVPH4a2WEqvNp
/2YjjIu895c6HbAiJuYPxMK31iAEAw6VoNRqEuGKQeXYsdJd53quhkx7v3FUwSjT
+EGbWUHm4tI5NsLhdLMCNNiKaF8seeS07Enxw9EcCIOJbQBP3bg7hQ1p3If+2rHp
Q0lv20AvDYZ3zSPL1H3GNL9XRTSV2C3Cwut4r6hnWaeJaFaxu3gH0e2EYNklysKu
op/9BuTtxUse4cPQ1m5bo90+r+V8FL4qE9CE5R5HbR/vepYaRRdpwY8Awdfp8Avd
JnhJiXwF/OVEJiuqU2aBQXgHb9J3k/nTXKlvNekwU3/SBwMQCCtuMxdGD9f7AQq3
q2DcJXAKWnyD1dxMZkk0QVI9G67bpMrG8VPDCquoOU1gb/JQKhYWs7nkhUKJYvbq
EzO9i/waF38RpHCj1cKCHciBjVd3VyD7Uf1BuYrLIJ4QtkhvFRY0RV2hhgAJy6UE
Bvz0pLX4KZGbf2t2dpjLfhiysEXlfoIs0uNDiNs0zQ6zKyQeBwi9GgVntwqzuULH
r5QtQs9c1Svo8OOM5Gf6JVMr0wwPfklB7pW9Za8DYS/crV8MRaAUAncMVdk/xijd
rGcqPLWYUtlXdblXIaaEeQVdAilCf0w7S6k+FoyOei9jXydjx+RIvZVdrlwS/oG0
25wezloG3LJGhWg6g925BLN3NMk7YE6rrBLOtlmPzikBF6tqUKemECTsLJermdcD
soFtMYK04KLq3QUiwGJzkKw36qryg3g5TsgIj5EUOc0ciWsHfK9gXB9fF+rbb9fb
LtCysoJswnUCvxD6diyVyTioqChHA+55BFT5COYyG2CkyJC39jczWWfw4Ej6OYMP
IU2kfdD2exnPmcuVtfQwCwEE18vuyfR04KmUPrR40suS5bxZ/viX3W/5wy8C6EbQ
rr63zI7jJK1765esuMnpGR0VIrV6sOSi0fwis6ycsZA3ytERDu8CWNqYDlt8FBx4
WKhFXJVBkx3/idB5x94gKTtTuZY8bHimvlklVUJUBI1rRX+MbMr9XExzzGdltqXW
3okXbXJaId6vX6idABDcru2dpAVp9SwTA3Qpzlq17LDqjNmAsesKqeS0tDCxhOLL
ArTMXuQe4RX1DiVfJ3C+1xgRAtjNG65POS44RRaBZWXPzRBO53G1eDZ1v/8H53+8
8+r7s3Ji3ogHcvbYQLztcGX+XbB/Vqoh/dg+kw6epu75bj6d72fuZzocfODdsZg0
eml14HwsbEeK/7wRKfyRdHKNLUkmIqeX4WStwGXEGGDcRbZdLwZxH3e+RJtEqKP7
oI778hbpcGqCyGOtyj0/XcEN+XGd2WBC8nmTcYDRXz/bs7lcpnoKoTBLu9f/8iqM
UjPqrK+Z0H+ZQpTrgiwtqydBWSau4WKLOUpK6gjlnP/SbY/XPWxdZ07sCiRp22vS
55U6Y8kQxPyq2KYX2r7CJ1pxbaiu4mQSOAQEnASIGiJ8ERGdECSxC0eb6IS5hr8l
QBDbBMxP0VXrl9dkAeGiXAqi0Krvh9GGD5afSwAxzjDiS+OSgkTJEMonzbJScagi
/UDFgdXvKtEnC52i63quqIJPa1ZGq2xDca0XfdMvuVzW7rWUfdR5UFxPwQVFMOLt
vIMKeJJpZJmjJPXbR4qbz2jU1yJ6JfHrFqWtlNMbjk4ef8PXsc0/k6+oXmDfbyyq
3wU4GO0OUcpbzIQTmhtFgGIT0WmglM9fWWoGEcmZHZBHQesZFao3WPDOx83s6QD4
Ko2UWIwCSjz6Ta5TO9jcO1ESvEXaZxxIp23YSWD74vbtgw7LhXaw8v5Dza0uewyH
O5pD97H1m4hsnVvNzoqsuaAc0Ycm+D2p9aPRXmOcf3rMniwwFY9QQsDeEIiFIXUZ
3Wp6LlYEMxHGYSb53nIZfvFjwt2JcL4rNW7nNeX/Y54N5pS2s9XkiBzzg1KCriKT
/xx44qwbZAT1OCQkW74DQkydlNN71NiQflLCUGFiQdPW8Kp31EIlGcjHvs+ls7Q7
gi8v554WAqUnL9CRn7XrS/a3yQyf9HydnsOwY5sAwBA90sehJGU1pmETPmc3lCVI
fQLDq/xEHOIWaIf9ujDmx2fQAjBiI2ghrWrLxwPxBRQg3Y1y8v04gQtZojIy2h4W
w9VhqQHMhY4+7nZZDfFLa6pcvAzqAFJWwAiUq2aSRvf6aLm1a9weXwt0VuuxiMGX
zudtEIgd1VQUyCZpWg01H18C+CM1h1oD5KREE9and2apfzUsWyO6BFlJCZNX53kW
5mTlg9wAl7osnZl9oJFQmHl8FsciSOX8bGmdH5JvH75Cg+rWlTcD9D0HVLLep9ew
ORkgy+UOijDR/UfIn0OW24QabY07XZgGLnwvQRMtlyzPOyIS9vko4q45NknANXlM
D8k/5oqn4arkXlK5qjl8mcK6I4HyVfP5Q8kD/iTmROpucPNxBSrZFUZt9VjpKgvF
ATSOThwUxu+NMIzEWehWbV78+bXKG2L6Ba9QgiBmIbZqglXgz5GAs6YzyZ6GK+ad
l/25OaahDHrEEG0UV1U78Zt3XgzHus6s38VESl0xbwm35PsFNmzPV7P0yetZFvEh
/C6SMhz06IZV0F7YnmFGRfYFXKYwMQ5mNg8wYB5XXK4mb8Pb9pd7g1d/3YWBPUQo
++T5O+9CXxCw42Cr/fr5uqAqI1haF5z3IbmfhiWudhQ4Pw0HSMjnB0VdAbRmLrMs
VY5zS72pkIV4msT9lgOKtu0J4Q561K4piCoGqeVWriS3cWYPuSs9vBrtJpb7BmvT
pJF142hYEHt84f0LnK4D/UUn1pz7xB1VXG2+llBkiRzY8FEEdmT9vaf4ra+vaWjL
F7okYpqzBfPCQzYIC/DirVM1JLFlC46lZ1NcXtb8dLMyN/hObtJk/HxRWcck0Mo0
LO0PUqcX+Ygcm7mX/h+VHdzgVOSdLki60YAr9GoQh0RANmuRLUUNHHza8asYfo7W
JxrwfaqCPZQcDVSsrCZ3Ubd8//0RjbVeTN4+Zr8k6cfAG69A0pifzRIJlrEAnCwE
lEUyQneJurEvtGkLX5W9tGKdGx29Dt9EEyQZ8kte8telMtkb7bMCb8N3OLMLD6/Q
X1VBAVEv/tK7xRTlyuB1K4nZQl3VvS8lmrnVt/LlwJkjqbbN76fgR4T+Pd2zfW2I
0djukEJgo8c7eCiahPAx1D+yQCXHaXuObFOM6XB8laBlck7ms7lXW02LZWvEr9ZP
vagyJsfcqz/HPzLvdAt/P+4nlFKCbwwcDGNvfSSv2EJ10qazMkSUF7UcpsjUXhWc
QD18W+XVoZomjyoikhnioV67Bq+PjO0PAhQyNeSrgdi4Af2l0MV/KkL7Ivwe0TVm
KO9tIPt4C/QfrU9WnzcltLDAVrMx/qHodYDGaYItg9wobGqPedUyCnu5E2z+GtAg
6CuWHiSg33v54sRiMzncDfCTUm/2sTc16AEGZzHmkORk939d1Jsfj3aGogSlHglD
A0Zgu3ytDxnG9VIyF5SxqnGV9JviFBkTzcrC+IGwvVuCZrcCfVkXoiCnK2HgmFsk
DYZd/+whDix0jWsSBET2unce7oUc2IavirgCTczIMNo1pFrrSUXOB40Bz8JsnH+z
EeoYEtaqmfuhmcVFrD7leH/DNH6Y0clPNu/6rBbdcCA0fPLFuJEjF6YPW+rrI215
8uFD0lKCrGQIyyFFVGd0eBFAYTxGxYco+oi+Ms2h0fbHYm9VDuHo4Il5jkByeZSe
V2+wnMIozunx8Y5yz8RkfwAULOFP3hFmS55t/ev5pSOcDktvoLhkmDzEHnJIs6y9
NyNuqvuQx5t1onKwvW2V1+6hEghskIhEB3OpL5ktkcvcGooF6GceaBmgS9AvVuf8
RfEEKbVs+cmKHkQ6G3U77HwzGgTNssEIlW9wT21R/XoLwZkdBA/k3Mg+nEEBgNhG
97jl2U9PiC2aQvrdCCSpp+7OvQD929TKdR2DPLpV/ybIgx6hPzASjo4IHJb/vGN8
We6pPATYpDonVvU+Uzfuj+O29O/ZiEplabEzrRDrrmO41pt8WmR0NLlVlegnmJXW
1Tg+RWQEBPMeC1jZ7HMRikIGNIyPrmrcNpW7NuxHYS0lDDN8KR2fGyTOfhmCYcz5
80BBVRu8cOVZKTpevVpX0NKskW1OFUjHNCQLxkbc5TeuBc6dWB1MYmHa/73iqShV
7AtO1FD360gs+GP/68Pg2P3VbJmy1hJqbCxAeY0OD6pRF4rp4frLgWQq1MRUpRMs
5Ws3Twb+Y73UuEoPhEqWIDa17hyucdLQga+PjGNQ+FtwFF1fODaZF1cXeVq+kDie
lJJc4eE2kB8jNw2fn7ESSisl8e7lE6dydNCL79kdeXZdmgXHwmJUo54eGAUAFXPm
i0zrDPQXLYYrvV0U0EjvQJBptlGWOVeEo95yHoPDTS0gu77lF4854ge57LNlGuHT
wvajIuhuYCxBHrNofLAW3H2sBRAMzR4YxKmhfK6dBIcW04cbHYfzxgAuIJIdti3g
4N91SgX1oGxXmj0jnCt0DTlC3BKbMhnJptMwR+4FBA9q0RZYVH5TbVd4wmpVjjih
meihRkGftb89YfWCbZhSJcYvLBSXehRQf6+5YnNCJ5+PepQSjbe22y3RPtATlL2Z
+oWRS2cq6KbvBE/5ma5Ja66ImcCa5wbR9jWPzZYdOPTqIuFVstv7a6S8jtvGtStO
75QbJZ0idcRs4L0W/MrXc28+oKi0ddB0LExBMzxzA7SJENY6ey3TVK2q6kd0OIAS
w+dLMQsDrKS8O6y1ZTKEBtpYbdPpr6HvDtiejOcqePdGFD060zGh1t16zjyjJ6iL
ZLl72vQjrzVynBiUSYxmvHjoM5LD3guL2otd4B042voeFnr6nVBMKKKyJ1//Pul9
dOgvwn7gx3AKruXD5Gb2EjEEh7SjbiEKG4WOY8Vc99tdtq+H7gBnXsOeUi6Lij9n
mdeTttaPO8dLjqO6xPS9za6d2pcErvG0ZxgizHYs9J2yAQp9flrtQf0+J9+vNPUK
G8u3mLZNGkgj72KoJ0UcqPjDm1ptNs0j2MUXANljPn/dm1cWQkvlh2WeYG2KGrDX
Zy7bICKlI0ZzpSSK2E4+hVMJlHfzHK4s5h60blWlG9UZALMcBAXLh1XfOFY31bA6
bgmex0qI+QbQfUCelErs1M9NireuCyam0eBvAXWFF7wTbcS/39lOGNMloLRq1XsZ
LutuQ0c9Y4OSO6AUJXZQaeL7qb62+Rm4nlLPJrp8kfifAgi4lLLspjBod7Ewek8V
b2YYYxWjFaJRhhO+pKsyGertxMR/VT0CtIGvJv+Y4blCWLHWushBktfAmxuHo2c3
a4+U29w88aGiMgUvAOlOgeU+XFvoy+rPZiTjCxPCy2k04E9De9h6JBcnXLiHpdQX
Rv7m92voRknyZ1Q4Fb5mdoARd++h0CPpwXrkNQ5zszNNWU24L46Hv05LP9WrP/Nt
wJfsOAAPO5BlEH/fmiilRSjn++zgES3SlgBYyvYb6Gzlwxk4ZDsCzKt/rxZm7oKS
LpxdICKIcxSD1jxQq368JpsWEW1jXc/ExWsKI1xQnBDyBHPz1EA/Eqv4xaNSy0kZ
CZd4EBHoTFiRs16iwyiAoPFTIBi/JU1JgjT3n4GIkXBCltBULZevYrFs9nej1bLW
cGSpv+2FZ+TFPNeaYTI+XszDxQsjASky3YeLuSa4k8iKsK6r4I7NQQ/3Ny+U1ocX
WxCSbhVwgA/7F7SuL7tpSqESS8VPG+4JMVbB2BJkhYaldcDgKbET/yUc5K38HRRt
tDneS0S2CM68JnwNYIL3nuui7YVTUgI6thzM4IQW3M9D5g1PNNVYD1WhRjlEHATc
uYKy3PWhUYqsLDa5w7LXixxFgkck3dgCY/RJB4YCTByngkf381culob1jE3pA4dJ
8GuALnHdPsSJVs7RkuIF9oB/r/ovvwRE9Ezzc69lMr9r3s6Baunc5AqJGudJv3oE
ulGD610+OiMjXO4EvxiRcX0XKknm8OOoMlCH8rJ/N0Dwaox1pawtcltFR4ePOjSx
u69RrWg+5OhjH0GKvVSfwlwdVvQKCl/Jz6cUWWtP6tDgTLKLPUgpClDUFzKLE8y/
G6+2ANfdRZ6RQl5WtErJvw/YOMafzZ7btYaPj8v+IE0JDp26zMg2Nh3I7J6s/p5f
yYZSnr0hFBiLUHSP67rF7ZmMqttH4cKFb9x1Mn0g+QlK3GI0RMC8+NvCS6oeOnnW
qaNGXdq7tKMntbMfwi9Dlj2oMU/hOCi3JlMvBVIm7zHjJvfqypooxqEGCVsIgipT
lev11UKYrfUpDU6zw2ky9FXBDOGMBRYmNrU8eDGlip/FeOEGhidVRU8ZRnhoIHv6
2TyxVF6NBtUXIxDdL0e59rRu7peqNQuw8cEKPzFvm6h3hU+QHaB1LLdOReQQcITO
oeX3dMZAUdgDBCOqjpM3NfDXBXrqAcNtoOrKZOvye4h4cL9p7GI2ie6HsQ/219B1
65h/HfPRHPKNQnBLUjSLJPE/ixUxHPsVHAYUein0gta1gFMfi8TXJeUULSXZ/gW5
YM5G6SBZWDOoKpZMYiIRnyiHlaQEQmXniUe0dSzjZvpEfXHUFyimj6RANLw2W3zj
7yDNeJQCLg3OGFXs1xHKZY4w3HUvdiSNvrty7vBiHQJesuYdQIwfkdIMiqp7A0DE
FHKhYKGGCiKqsu3XmkahiJudnuJMTdHoZnnqUnSxLxYkOBs6PkL0OasZzPDjc3vZ
jnCPZp1D51iMC43yW4iiNbGlpuCmmpckLNYzoCMMuqVYhAgqTcj/k7R/gI2OzfrR
Wq/arAv5Mis6gsA4d0Y/0zDlelovbODLMPnLVq9ggAH+mx1+BaNb0OiYHQPtHYQz
NZThRaSk/ywP9SOuwtJdwDnS2sdL0Xg5QfOMdOTPtRPNrst8tY/vU+VpunX8x2oO
p5gKdfYhNnyUoSIQ9UWLbiu1TfQo7+X5XFCm1Cr9ROpjiKwY67/No3fkpe5Bo4Cu
NvNFuAPx0EHAjTCADkcMccxk5Yg7eafWC+eXAN3tbr96mjaDP3/+L1DNDPH8gpd1
mil7qS7LtlCABYoGIl4TrHbtxwIGoEDZgGHgBLuAB9o4iOXymt1ivZaXbKIl8X7r
vHJCLCgdhBLWu2U/8fa0N0UsqXmtI87AwCR9BKFu7E3WX5ipebzIkzrpoco2tBhX
D5ylOXl+Ys39MwUZjHBqQRINFCdYr7bOPHU5Xv312W6ixnZX+34z45jEuURXeo7p
XBPj0grdBM9rPWaVAfymUvCKgeYdYUp5B4CNCKWa8CzPaEeUj0UWu9UqZkFmSGVA
eFi/1+SxDbV9eyYB/Y18g0rA3b810avzA/pZcBYmF9hGvTJRwDZusyLZfhVVs3Bv
Z3W9LgCqJtaZYiZZBNelYhI8LH96WMpELmj+Y7tq7vLsXt/4mNH6X3ZKqQAW5Wy3
za9z33/9o6SCf7eLQCyQjpDaydr7U7ql9uGYdT4CoX6u0T1loRRtZwv5sYjt54ew
3kXTeIzb8M6jh6MCi5zhsuV4nzoKbUTkErPNxNErCb2r162leORDOl4dtCQV/mc2
nOeZoDiy3mmkyj9OEjfWr4klK7j+6l3UtB/hSZhWCj44DsRHAfzu/nnBSIIuqAnM
3Abz+aDBc//d0iWAYeEf+5DZiFCI9CNt+qfV0d3ih0TrIkz1oNZ/77m31UikxN6o
MQ1hrB66QV045Cx0apJ7KfZy4vZnmKB8JWh02RjuhbsA16URWApf6Kor5wOuJRqY
PFlCWVbzrbcX6ZwrlvxYcqAz4woLjqRjTelwXUb866ooKzZrIoT3HblA9XaVsoY0
p/SL7meSndqvVXIm9q9fURipsdIAuXqd1GSfNXgUDt5JF+pP6bjUymVIB8NIXISd
N2R0VPkjROpNXt3EJWmhbyuOKQn+TMt2heEQdkPNtfjE3K3sCrWomv+K+8dLUEVe
qLDbinBwF9gPUdVXgibQv54MsZ/kL69/aFzB0IOzuLm4rOwzALsv4XeFmnZ4n6L4
oEk+HkS+GeL1dBacA+nD5EQddhXwqGIXue6Ed2rF5fjSD16LsMkQ4bX8vdSDXS53
JZ9ajHyjD1I9ldXeGGrOsvNTOz/qc+15MTqNjWXMEagH8ybcgFouXfx+o+OV1FOf
SgZD/xuvUp/GgYxXSg1dwN803f8+NpS8BK68YtaBZMVyhiUIbqbsh07bFdDcaiRd
ndRhCi6unZsXEYlGUN1PCcc1lkw2u0bQKOjwWv04or+zXPk6/GDi1B+Lspd+mZSb
zA1CqTWv9jim4HLcEWT9wnnc4bU8STbltOEEzRfpsnBVblrlqpubb9fS+AI9/ubB
UFHE93mqKExNe5eXZ0Qlbw+XnstP8rXd0mdNemnMoKJEWA4DBHu75wmraDSxv7UL
8svklDuI/6QHgngE5BpbiNtcI23jgy8FWd6vKMpngl/JzVN8VICIh7dUa7JGT3uW
qZS+Vj8Csr5ZvHazxRnDLCu14FsPqhgknv8fDL/VW755Gvpdul13flEbLVv7fpUi
YX4WmX4y5iF2UYaEmfMRGwysVnffS7/1CYYBxgHMnMKY02dM6/dizly7SfvBMvjn
E4nKc7AdoMsBZMEVCMNTYFMjKhEXxLXgUd5ZPZbUJ9QHMn9nUhG5ddL0LmOgQSUa
yvePuFQpMeNZHpClz9AgHK/VaSCSPYejt5M1VkF5JU/hUkcCx/u2oVBmLIKCpdUp
BvYmCMrb6re2K2A2zNa76g5gbE0lDjC67RBWElHFdd+oWcGQXfzuUBvaYodGeiTV
Ss6+H5kD1zQ0qJr5iAXNWk/FlmvQL5nw9M1dE2fBbARYBB2S3GmR9YfHn8Oy9uUi
DFh13bZmzT1jn9flHohn+Ts558Rb2M0oyBfCI3VnHyOQ8iF76mrGU/JQ70Y+nuwE
Rg1IhRDD3Ps7vhYFdTdfOf5pVaP40368+fGw2eCpoAseuCsUuBRWvXqmU+/CSUy0
j2GfvemU2sI6T+7iBkDP7JAYsca46IjQ2KkKq/tAUb6u6rbuJISts6OS6KfPZMLb
ZXVpgFvs3DIQSgDlrembwj5BYsSY3/0U6ENCSxz9A2ZQK7BR8y6gyMkGGQb4ywyQ
QbFn0OxzPcPIUNC8bjge0Ob0CiqY2l8uG1oaw+t7RQ+3xk1XAGWtzxqDg75VNkRY
LgwTWOv7zuLA8kqOzfqpEjIiXKh/RVcvH+3lYGn5DW90zbGa5ODquTCf2wT4K5ki
389SSWL2DxdRgo9QjTQEagx7/jo6dXMPNycQrPJVKeIZ92ddune0fKWMuWOOtHNe
btrc3oQHONrew83hSB+c2aLESa4JWJW68+J01CAVL5grqUiP4v5qNgYIo2uzfG/6
HgsobWd5ccCmpXrtlE0LYDwk3NU39WkUQnMfRN4GngHFTQnU0mmXsndzmOPuHSF5
7xTeKt36Jo1I2PxC/IF9/XeyhmSMQPFX1Q0ZZhtMNUycxZlleeIA3K58nQLe3dDS
n1rkberUKoSEvT7nf+GF2dwVJ2gNdwfPdscQ5JUDNafND/dN7yjtxh4KA1RcfwoY
nRqEKzwGLSfWxXAFEIMqdHUACQsHS6dycHvzVEcsA0pjoRlMK35CHLHCMII+9v6G
6Y5qk/r9VPj2CabZUyQOeh7vpEKm8yDiIL5Kkx3Qr1ttzmvuUDnjhwQB1D4rUa1O
14v78UvEeQfgFYI98N0j2nHoVWuvR7yiA16P61m/Kw5ttV1+8h6/Ej6u2oSlVF34
UuLqZ/3FOqQKHeX0FdaXzilr0IvJvMJEuj2yaEbObSbuIyw147DJQR2yurrPLCqO
moXTz9oT+pYKt2mRFwmJqj5stkcjYurMnjWUH5cew/bM9TEIta37JaoDPyTyrxYW
rfIUuIDepZmq/9KLejvMVbn7SqP9xrnNwiATihwgFB8X0xY1BnXKjUyKddaQn4op
21/EBaDNFrH4YJMeP13mMO1dBzxCgZHlXu7yUnUy6yqordk9yV9d3IVSoIbv9Ujx
OOkYixIzIh8M5unkYt0vNfYtOnanA3/7J9E5kJ4XzgtR1A2EkalSYqzRFxwROoiy
lEUlobEUDxtCdIQTsxfHvBjPFudSHcH2kovqBbX3LkfwH2pNNxIB6Yhm3gAvjo9W
vU/X2rwilwYiR+coxrPSV2ORjpNKjvQWN9VcfM3RZAvZ8EaEI8CRfzqRKlnAOEYK
t+K7UM4cwUBoPVYijB3GPjdEmYCr2uu7YnPO2HF+LS/ZUdzPWehfPPTjg+ID3hyn
63bKAZzWWZX+3VcwJHzWhlvPUdJMJNBlBXUzxHsztVLGGjgGGd+SUVuexq66L8+4
ixEPeOgD/inzLbkFH8O1s4IHXO6vVpXfEglsSSQENdHCeoeCAZZLV7wDdgsiDrcO
Qy+oZ5gjFqYbefe/aEl1RSSEfviO25VJ5QIQoXmqdCLEF17rTxGRNgDuyEWMCKyo
ISsc4kwHUo9N3UEWAaooaRbr7YCWhy/AOAgHioT4CCXpIhZFnWO344weQhhCEKwh
aidckX0+aF5ZCijSggfY5ftjMhEvAaKgD1EiEAbgO+P3nZjr+TLWl02PxGkIUZ9P
wSGW6jJzVK6MnD4+MwafiWDo3IUSZHwWvXGtFVA4Bg+oOaGT8ZDzolbqT/UGr3Xr
qxNZJwWq2cRpn4m5knMJY8U8yII/ykqjl6OTfPk36AhsKdoTDsqp47+GJcSzsksI
fMsK9CSxZvRK24snjwqaYndXMwKghwGNCYpZv/a3q3mnsvdudvAu5HQ4eERRgHcM
LRHlZg7xChLE0I43bO2P/iVXrrnTouiW8LJMNcs+6Bj04qjx4alwTFJcOjcPHDEz
Is/HcOtKJ5LO/UFZFM9Ym9aBOldCz1ojgjC/aK6MUVJSm4AydIAYnRmgbuhQbEgA
NQKm5NSORA/hwVImzXq5eInS/06akzCi3rKxLEM2IzgHXP9crZz0k0CQLvQs8tjq
bXAWK6llxcbOHISwekDTKIyvJojyrDo63UmPanpfjKemn3U/IcjkvsBBM/l25qDR
ez/ciZ+e8PzxgyBLt8SlDgwK/q68RaVoTabnZNK34Ox9aHdfcKppebH0VkcTRemg
J0REgOY/vDDrYoGbirWvygo4dVGepB9ioJHJBTY3v8kuGa9QF5PFefgpBnYS1ZLx
Rhd8hpxKkYGJN6SMu7EEWFkFr5XoUEVqhA6SbDyS7jYUaGPn9n+/gnjZfF5ZNNxP
J4Nk8ZhRyvII3Qv2BS7DLZtW7rOtGLJ0ntiOCVvtrFLpMRHsj9Jb5M/BNBdNyEEe
SLwa7l4a0Wbt0WX+AJi9ZE5CgbzTp23v87ysXdPN1q2bnQmwLQS8PyI8gxq6+kgI
46uuLQRGFsB5JwHDPaRg8QqNgZoJuwzlQEgOQ9zOygrqv+gFs3bH4+uswOXRlU6L
RXzw+sAr65Wg0FWTBK63CfJqg9f9sO2Xi4zvxz9xyZaKymI/2D1mCAP4cLlN6vFF
256MZCH788A7r7BPvnAQ4dtgetlrG1W4ZTCHa0DDBRNrWupFYRkMqr/4GWhgc1zR
8/rj7EtahAfiDU/sYCT/ae/9gTHEk3ZaccxErv3gICa9cLNVUofLTu+gM9qTzGnQ
Y//dIV1P3mfiMN1TIxFHMMyVxtaquP0XmIKs/CB9O+Ec4M8r9CiZH018EDIoK9UW
U943y7JG0yOOg5b+hdR9C95sEmk2Zec42sJk6CYRfDTmRmd8SWtRk5A8mxIl+n0c
Cb4ubIlEFtPX5bCtdN+U70Qc2fmm+0LxC3avLMQ3zCsz4Zr2g6BwUu4/V1FOkZjA
fMzdEIevMr5o7WtXUVvedZB39e544RheWkx/2tz9+d0RFNPRB9bGMVf5Fb9ytkOu
cA6FiFNBQLQ6mnI6pu8q5hwCRHcdrjcColgmJJxv9s16o5me8TrEHbqCxi8CzyXC
/AXVPDIQs8LVlO789ux1hyvh0xYbTanMVuZvRIeNDBvlFfJKHTr+QEoBcWCrsbro
/L+DgZICAbbEhueFo54mmmdJBrv4nM55DJwL41NbBWSmDplnNMdIkHrlgEuCZqxU
svESL2o/ZKYMaOWYtqzSWqTP6aK2g+QoFU/g6I5pir8fyXe7C5tKgx3e6k+7uFC6
44nu6o6WChy3yQBP4FFfMsIfzBFFKoFa/MXE25oNcR8pRSNSZAsk9PUJi0bSk19K
pAU0JoJna3g6234os+E3beIt732EUwdEWZCCkf4I1KRoAtLHVWn58w9Jpq5SVt5m
lQs+P0iyl+D+YDVpDD6/6eMIswu8++8fwC2INE4HZzYqvQSFhddzD7tReQ/Xlfwz
JMw9FWMX5cT42mwS7R5Z0D45vtl7slxF/rmmGA2oqXcN8RZg77f/hwQXRNSrTzyt
ZBhJRAKJ7lpHrfVYwsEk4OUu3vzPJhKNmui3O2tdswSanqs0oz/vQmxtcItMdIQ8
4bLBJWpb20rGACby++d8QC5GS16Pc9w3rAdSfogMSBi5G24ANrMlguKW6+e6hWAc
u3orGv/IsUJyKG7aHDu62gK5VM2W/duxIWToD0x0ogd9noQZ+2au4GIUQUyvdx4O
P/EnvGdkKe6zy6WYAQYNV2fVGgSEMsDb4ViwZAzxuCJgcAo5rcMXnX++bAlaiDln
pw0WvwNUqCctES+8SqakupguEnSglove8r/2+4XudyGfM/WXJwovEKwgcFNETIDf
Qf701qxG7YtU0xqmlCpedLHzZtGjKIDPyP0RgWAaniLd0wXURcMLdaQOTH63a6AX
CY5LtPzjAWupsmOB7XNTfbQS/VYw7IJlUdaxkC9ZcS0aOsnx8+hY2eKh3TU2qqgt
DQ857mW9uoqH3VF7fB9R4HluB0kBGHz3rBc0mLTKGbTFhzuHs7JlseC81MkwbDpd
TXKie0CyF6Sgl6vNZLPqZLeu3nFDP4YGs4OIJqEzqrnc47u2h3HjAETEZR8QAd1X
I0C+BKLpZzu1SScFFM/4OcWoyKqQx/TgYPDMHiUtRYAyHqCtSgDPgZHZ1dn5F8qC
Q6Afu+0hylc66F5juuvl6OuAaYQce+vIQ7V5JG85YekgEcm3pcG1sg3AJEXRO6mS
eSruS72oqW8zwYBX8IqUV9tXXE1iUbjsCh6az6cE9ATLSLmkdLNIjMMxLOmIYW+q
HROB7hTVMr5iigqzA1gWKcmWO8u6XKbUccGeUf02EbGpFbQgIr/zWtpB2WZkyuuL
RfV5Pq0IfWBAqFev013wULIFU9z0aozfJAPbLxfNHoKCt1MtjwCpghiJGOHq1SAm
ABhoRL8knUiFg75b3srvi52ieFGDxIthALTwyfBEaVTnC6A6wSoL2xD0SlCehqBn
ohbvvfRAoPTpKg8mN5+hqs0UTULsto4XMlbw8j5apGozKx9WqqcLcvFm/DRj7DA+
RZAa/LXqtWG6NIcfxxiMjMtV6GNtER1VO+lWm+EaNxTvXNN3aY5wYVqbmJ2wsvbY
HHlj/TSSYS1RzLx93tGsOgbLxTQeRqdCg8JWVA6a44cZi8gmMmvg5vqx95ITGe1g
TYxnFILgkW0SGl7wIrUM6yIJWl71Y2iqFQtKUuB5w39CVH8lhdKc/JL44OacfZfu
NmZfMSyilgiU3PQa/Smvi4qqBbbhPV3IgWWnNs4iDRIUuy+6c/mC7jXdASODXpyv
EW1FFbCwRfvEVclIDKoD2Wg9iYEsdgg1VMUUs1ZS12+Jz6XEJxiikwcCCwXiokPM
jV/JNtCFovzQLLKOTOFUo2xkeUWVfyrt5irMKO+lQgFoC+dtlQg7USdS7A+/Ed6P
meIzeqIk4AkPlFkPHtHkB6cn9e83C2iQQaow9mWIeHZ4++LfhQWgeGkZEJdhYKah
Iz/aggLiaaDWXrdaUq2zGrY3YmcnE/myIwRQRYyglUl6l1aw6xdlUUtZ0aeATF3f
X59Kv3iq0k/4exUIR77+8MWc/NQENheC1hst/347MMhIdIU5JMej1lzpbFRARngF
455wuYNPU+Eb687eOb71cXwDID/CqCHO9UNriPCC+5q29GKVd3qmvcpdtFUN0UsO
QA+geJpr5OV7RDJFO7tTYmd2UF3Sz9TgaFSNGryfRn7R7IMfpF51KbB+xMfNdU/u
32b1o1tfVPUklKrZ25SVS8VT94Klz6z6W494BO68iEGaPZCP+sl8uHJ6h6b4x0Wa
HB5ACpVCW8mVmEODU3uaUUHhbKm19Y3tAUaJV+0kZ0HUeGULlcN77EJOf7WqUto9
EqG6tcyJr347Mg3RBeIhYXD/ah8+xewJA029nQ6v9JWQ2cocWUxOB+EFw/9IlDsL
Gat1nqlFeqneeowE3pyBag9gz43S86e+3+CfEXxERRBkUAuW2iaT369irsvZQlKl
8Nyf96p2HUehPB4mbFgMSH7t0KYl/j864Aw/yRKvmOsw4oAizjFJPxkUxBZ2bW5F
BtCRpXMf9dqeD/dN7lIa+4/4YlV13Ov8oQYDnLnCnGqzDlpSnv9Fo/aA65ZAtORD
slOwG6yZTRSTgE0dguJZ5lY9EaPnuEOHUqLGD1JepliVB2xjopasqmajJV+J/IBs
AU5UtjPv/9ypDEQ0TD6e06ZaKZqV9+dQdh3fbibBjgAEXM7y4k1I6QeJUhP5GowG
mmkGApUOmCmzRiV5+bViUHiTFiIwXkemDT5/y40GT0AQ1s4nX6ZpXkh1Azx2otfF
NfrLCrNne6A69f5pCSsaN6WgKRPOGDHAV0ChEZIHOJLyCYA774fBp5WgA8KB6yO9
fFNVb12Lp8tysb43W5mM9qimUtaS+RmMqIxlBjMxFNCbsePJYGHbwhr/90Lp1ggu
wl4cz7nEoojwwetoSrFEvEtR320n3WHnGmLTE4cQdB95ktD7O//xG0BqgOtZKF8E
w4hW50xLl0kGQQA6J+t++ZiFrCfxR3cAYA1w5lB7lvKJP/STR2cWaM2IhGyn+7Ra
ek2JtgvTkNvS5IUCNgzKTp/7UXGGJmLTlni+09WmR1c+HtgIK4OYugeAN074+oya
sJ+xPaIYicE6xfGWO7qWYn6W1zFroOJCB8UMWYmZcpo3ZCRHgZKiTEfIsMB1Q79d
7LyH4nxYSx8c+HuUthRmwfir1EWavb40vCWfU8+qHMFoDbQQc+Bs8pYdOUhpydNs
Iyj6zuga++Taq4TgHOHhhW3mRsHNHSRD+kOJxAgWRKUb90SZwAXv2y4kijWLBP+r
OzXdZR8X/79Vn4JHYL3SQtManFYLvkG5eHyqBq2TdapQrA8rhOY9lSMj15hFU7wB
1oOFYUcLbTsxtM9KaS++iOBeZvtV0zjzxBd483INGoAUx6OUL7rgtc1mzROo9rpP
f0rJNQ5MNDjG4jQ/zz/cHjY2+PEvRM5IlJjibhEUcLR2Et5WDSgtPfwsridI1iQ1
h6HrC5G3CesPIDV832D8W85Rpaiw1bk299jtv4DCUQLxkzyyZifN44eZX68fpIl5
ndpC3gtJ9v4VKJqLN6rE6LVKDn211Mhdp9XawmoJnpfZ5eai2wkDpl0Tx15Z5upS
Zeng3a180hsjWOAgENnQ08ax1Wmi60p0WSd2vUhiZSz5DK9wV57yYZcMfvxvl6E9
kyedP6fggFARIIS3WO2U/lf5FjG79aG2nh572qXPGh5yTAItPa2zHTYP7G9ZxnFC
N2VQ40vze9Y7sBEsLnBJMISd95jrLTIbgG+eRB2nwPy3zvCQ86v+y5PPQKEDr8iM
btc+44feZGMPKTu11BXhuYPIM1S60RDLI6P+KMLN6owsgg/71ddzSuSXkQHu0qVP
3wDEOmkvMTxqPAhVfaOX+HVy1stk3NgFQAd8pr6A9Hx/h8wTNl0WkZcrF+elHY8h
dykn5aKxV+BS7FDw94eVXnNnuKEMEouU3zhGgj8Ylb6Fag7wIhxf2zVkMm4RbIEw
rGIcn6w3C0EeUoQP17kysHaYZQ/wdC6KQ9FRbWyxNCGPl7ZkF/ZsQMCyYMaKof1C
6wfpTmPphn9+0mDouA4vszerBn4fbRsAyzsA47P/aEP8Fnzga1FWHf8jskefI8/o
gStleTbFP8UYQRs0+PAxV4POfiQHh4B/wFLi4nnjCGTMWacwxlVjHZrcQ3hLiHXs
Ovkk1Ft+FHqvfN/J5/u5mOCjV9CNk/yK3XEkMWwsEKlqYkL66DL1T5rnQPxtkt+C
0uyjhwclDNX42OAiVySghvqPZ1gXFudluPuKiYKEnqeD9sDvaM1QNm0sCnaps71e
hFxpkSTC0l1ZFq18UvEyvPYl4SpGprO2wPWYp4CPWDEcZUz93hQ2ad8VQKsA9Ifr
7BxkaAzLrCIGKP6c7LaHiP/iQFG0Z5BxMjffkQPlzJnpM5geHg4Vpu+diAqSe36R
y7QBQb8Wyz2+CYypEg3FhJvz6qRZvew1JjS+dYyrXXUT2tgnhGQy4mJvqkp/uA1O
p5fz4tdTnV7tKIJqfKBNDTDnzWRj7tX2ClkAIE1xnG6Ij6zaISeBYiz3X9U8re1i
yk8bRAnOFsLfCOP05zC06KIoejgWGyYFtf3NlM1O+FCfK2KfWY3hOW2Z8xEkWmFl
/rfwG9A778dVU26lIzdtiYjPNpYmUEY+5RqeGshE+i7VddStIYE1psrKHLxJoY2d
6p+9CyEXyoUs8hssBKGUpny/Uwenl+VJUSP817D5JLInRu1NLGWPDlZpZs/0g+N4
pK7HRgNcQqWq6cuVTauCQHPr5XLcsucm2DZigYT0+4oJdlsz/Fb3kJLQfvPej30u
jEq+y4Wr0cRUCxIKu/pLw0pJ/ikpi1dp35bHoaRjIayK1/E6Vb3/8Kc3V2WliKfi
Nubiv36MDmvjL8YFO0l/aof39DEj3oMHaka6uw7zQ9LuY+sh7cg28k8wxYn+JLy1
uXY3aCp+DKXw8a1/49LROcZ2YdntxYQ1q7PrAtZvpzpZ1b4Z8KJuXGXqqKPZgu6s
/PxbvwZiFvtp5apNcq4SXkiu90TcBICJfS3ob9p9HlL+9cWJ1o+siJmT8xh2xxod
ISK6sjz/k/DC/qmH7ANhFiuIW0/osumiDzOGGcD+0aAmJc0zyHPXG5HBFc1TjDor
D3RsPJnz4OmbXktVXw+kL9MhM42Ai0u+GwqOm/BwDSK3mkKydFljpiSGT5S+ZUa/
1swRPTo2d4fR/+iz991Co7u9vM2leuGIx/j3wtO/oiOLvwO7D0RFALe8ibZXqso/
Om9xPKNxMiq0KjEO8tjTWuO7EgS62pql33qjJCph7R/UusefA0wl0Uu9VU1gkdPM
ema6g4I7t3qvzeI1usBntXSPrpqE9Ir9rOldZ3m2A2W0tlL96igJpXxnsTl2xStJ
VicW3YmUdeVrurN3Mw0vvasyNvwrKys6e42ceJmPoEaqmz47y/DENKPsqDJCQZbc
pkfh3IbQa/tEEK/E+R1cgPwuY3FGulahiZSjv/itjjH8dx6s6Y8eMMDH/0sOLu5D
ySR6xJtnPV15S2ALFkkSDAlu90QIXEui1Ywf0z0laXMfwWEXsJKdYS47ugKgHWOP
OdhmJ3M7v7V5edk9XYiMtMex+8O8yYMkOVt06M7ymlhZ4ebE73+LwEqWEvVpXfYu
kSvQqauqODSxFsuNHcEtaGfKBMyEJV6Lm8kwRzJ5HU2/lIJRBGX+SYcDKkx1pM1n
Zc2fn0VcSHXDmw6mjCnfbbVU6pLToiACKjBNgybkJmgMRO/OCLDGMlbm2Ir6vdeE
8i/KtyV7Nln0A9FJpkvSUR/pf7rI6GO+kEd7U9jRHQWv1vWH16ADxBiyGikz4dll
+v0bPTlZ6QAG8M8FMmWWbSFTxIj7+yoQZ6o02HZe5kLTqjtR4xiD4KVRtmTXOk9F
pBAdom2TX2xXmzueLiy/pSd0ARDH3/CuZMDfKN+43vCAY+6TIbKU312XZo9YgyPq
vr1bEXMT6JopgtAIfP0GEqceX6l1Y94D6hlrXMNdvN2t2iAfET0IwTpb5GStXHOZ
aGxYLEbJZVAKzDZavpS3ML6VJSVV90NwbsjggOP6kA2k2cJtAogajPwCnYRB+6cY
wtzewAxyhE5ovleX68yZefFqU8A2bUW2TCYccct4N68rBDWUYbnlR9qc53HHijNL
WDVKrhqhdOUbimR3wQNbg0mX8Sv1pMH4TYS66Y+Tuvje2wM+YqF3Wrakz3Jcgk9l
Iq8jFr5t74H8KX9QC7oFRXE2iX/SHKORs5vsd+c62we+OEEq+6pyvftalqA4qWU7
jvaWdjeO0wqnRHT8hL+hEsdBnmk+cXQCqU7twkg2XvZ8nEVmsAoKZXgToswB9hA6
gUHHZPbimvidaFZyO4QnP0UqrY0XdFloaFrGkLI2SiQj38Dl3OoaE4rtGs2NlwHf
/kFRKOkIHqyZOZMn/w9ZVFszb2wwAJwT10T4p65phJrBDmspsSlE7+E1qBBL7t85
ZfsW6Gfb+iY7bH3e7lcn00HZPShVmpaczbwwGnTBH2U0OoVCRF/cdzpiaIgJCv8h
BfczbMiJPMJAxOovQ7iBxemA/q3eb9a5jL9VI4iO0G2+JU9SJufboHYkPZW4/QcO
jaxo0gjxbYANiYlRDXoaxubPunMtNebrGwp7ZCDX+SvK9UD2Juz9Ac/yjWvAJ9Oe
k6S9LbJBM+JEl+pmlYQtcDo1JoP2ACIBaw5Anzi4XvERtezMRlQSD6HJwjFdnWDB
6JEM9qh1+bvM2SeYbtoEpwsxI4i++4yre+Hfsr/od8GIEFkmPLZEqKIqoAnqTote
ILOZY6CHARsUDWlPQ3yme+ypWXtvIgP0EikD5UBK5vhC5gql9MtbW8GrkBJj8kvM
l3W9dR0bFD2Qs1WQIVxuPjZKefTy3k5K575ymg4w1G0UAOr9bK1NS1qkIKV1wDj9
NFHEUNkNxtZaOcKcyrIdq4S7fyrBdpjTufNPrO8HbK3RzY5ThIRAAxO9gRzMkjYa
UXEIEhqJV2sDzvGcNAwHODEMMv+LqmCElyVbkuSmy5DEAfF9ZxKYEX+l4J4btjq1
bLWB6VuULOkXhRXUPO5AbWsrWR2Fk34upwBoAVFB+asjDrLtDDV+JGFjIOTQENlu
NScxmGdXcsGdst1S7XddRrIw0pSFNdC4YcY0qcaPUCed9sjtJxcu9avX66eNzNZY
CFcbReBiLQcs0YuE4unqBNW6jEkKNVIVY2gNU9bmbl3Rv/sAH6Etn3WHBESQ7GRg
JmUPRPNrQ5jh9ebLyxA4oLktj+5ownTWWMxSDeLCekJf8E/GgJ4wvopPocUgEnH1
YOB3Pma3iFmggkbTsPYnDteYN6eKzWstfO3FTAUH4oGA2eD2hpQQE6CKwZlVt82O
zP5i4/bsNufoR685gSMM8vYR14cyTI+GuwP0eVj82yZNhsDxFmEKYE4eUUT75uI8
/mavaBP2kUAX3ZYdsGJ0nPInGBW7REAXURBnHHaYxkbVcZe15qI5/ZLzuu7bmCzL
wWypU17Mcnp7/+IMWXaNt8BFfIoq1MmO93TzvQ/JARxvpMCXiEnj7ObjwQwEgqrd
r1Zvdq7W/KrrUgfOGDbNihkzI81slfbfYt5K0Y6yo7QvCXf0653aOj4i62s03MGJ
eLolTpj57HyJ+KOfeCHSk53pwDvMV0Dtm1dN1FYHmKXfWT8tGEv6NgHjh5hquqP7
54lMTCd4S8cvG078KczO5S/byXO22ooescqiwMucy/6pV+AL26tlBQ2Sb3kKHfO5
8WSyfdfoYowsmEzyCzB74HU59iASsA2BxIyF8zJUP/Ft81sefaPq2khdvj8OncVD
rPdkby4uG90H7Y50lAEoavKZHlbu9iyPzZn7QEh/P69Sl6xw2kgQ40O4XjMBMKX/
UfrSeVvwaN6y49DDpdWSV9awChZn/jv+oUIz1bKYKvB2iN0wuB1omuOQQlYSiFZZ
MphVZ/VVeGYVGXBxmSQARlFbu0YCoPEmojDkmlxm/MetwJ1v70yheuaOHPLQ0TwZ
IEB1h+9/zN1bqEV51SIkqBRzP+C5D4A0gs7UMXP6HzYswC+f/w8Etd9Y0x8NJnf/
Gvl1k1KgKWVPFF8Hiq4eWqyI7NnUEvsbEDCVmOjED5HkSD7+GH4ZDb0bgWCeJBXI
GmHC16z+I2xpjO2G6AXFuLNdB8IrRB/k9KEzTFZUdM9P8NGWTu7XtWFl5PFpckF6
zwBsTUcRgL1c+DZjUPNM8XnDOldD5ibl0O7UDT9+YRAJW1rLRPfUhAG1Cym7OTQ0
hxToDJ9HanirrmVI61hwjYR/AYuG3ShAayHVfAiI8xeXFPj54wG8qp238H/2dDV3
RLFtjTv1jYE5683WCE9Nz1cbWxaC3tvH9MAJjOzJ4oTLPgL2MtApNrOwZo5qv5G/
xjkZXpiKF0+A5UI3JelW0i+nzHtsc5xUXVLb0m974CsjeZCTUEGsc24lQh8gO8q2
w9z1m2wFlcFrwAfbBytPA/xsirJFw/jxNy2TsLYpjeUjz9J9jPS+n2W384cltx4P
uxpAHFSC+TzRyxIYFz8zTq0LJA4EpQ/oTmZLYZpu93TF+dFwn2V5NLZv+x3F5+m+
SXom6spA5LEOdz4fDKS0FnodilemvuvutI8doKqWN0QhTRoRHHN8d5WSIkrCbvIW
hEnFRMghC0dvvMOITvt3fGt4qf+HOXyy1RhP5lt6Zu6jNPGptsd5B2pmnlzHmdrp
6WX8MJxawUx+9GtKVZ5quPVfnDlhVQbXN/McZSFvBX9074SNl6kZUma71TGTBnjU
dxOKGViru+zG1r5c78wqrROlJu7Q3REl9rY7+YIKNguwsBexZ75TjIbLQM4wwzVY
ZWFCWl/bkNHMG6TOB+EuQIp5b4bjEF6nA/fs5AfFOTwIq5YwsE5PedaGsi9cAXs/
Ukbb76NXvol8Ar4GNZMOvxOgeD+u8vQIMRqCRi/5KedLk2shwuMfMDnNs3ld8Qwc
cTvSWtr1Td+7pi7NkiGIssY38nt7t0eRpHtH6ZVLEYxLoQtO0KeuHQ6uescq6uAC
+1MRQdBL/7Gfkxp8YksDI53ZqVpgPXWq8kSOBkTo43PEFClQo3613Ua4GMGva71t
Cann4qdWYMcqCIbjJtbb+G+/ATayNeJTRWYlr9MWQwVQtBS8F0PFl6vWVtlCkJbx
/KlWc4ZAb6STmHdi2bogkzx9AVcLUAlTZAJEnGsqFt8kh6KR3nJIkNo9L7tvUTuO
Gc5YreeZjwj+iZOwXplYlFbcsw8YHKzKBSAbrdCmo6dfHpJ2HirWVmjSX+M6yTi+
rZDWBPsWAgB/lRsj6Sa7ItBvleLwg20PQ3M4JM1PDXTC3h70l8sz1FoTxXCRzu55
n59uK8H2ih6kTIO1A+3dg+JrC8+iU0fNicFTmVKaXO5fQlfpRKbvJSSbRWr9tUWd
eWZsCeeJFQXNkCEzWJuilCvSJ7yt56t/IN1htn0t46uR3kEg5e5y8qzaMnQb/A+0
WyxHXule5538nZCd9ggRi2D8A3CJUu1b8yFGYYAo7pUH4tOHnJonekBRDweeMVwG
OuCnJF6X2WR6MIPcmlPymB1qM6USpU5VMJGNvZ3Tu6X9Z17MNXxr77f1v5dYT7P2
5fTE1z2ZJ3q6ES8CWa4qpL9uP0mY8DhzR/iO496r3CopWu5YC6I4ea3EGiyGYmj4
ULrWyOajZT1iTl6KaGbsHfEr33B0OqH8HqGf/wSS6LfQxLHY7gsOE5LWz16DkMan
kxemIsWFhzWd37LPqstmIqaDwwRCZ8I9JsseQ4YhXDaLmYs2/R7YgsujoMEdp8K+
ccux7VzKGu8RtK0bNrLjkyUxmzZjAx2cx2G0CH8H3wffEEryHytjtgzYkC27LV3Q
zwSZgUJcXB3/f3ivujbelZJfpHJ7eAbpsAXdXLRMRkVmC8dNquIrHg+P100yaUjm
oeC3d+/1CwsvFbENPY5yTD4a4++kxK/exqaZlQfebL632cgsNsCQ01xb7Oiuc5CZ
bln0uD20AmYvaymAL6i/RAqbNnGe1Oj4+YuLylGRTJeQbjUAnlz5NoUBfjVEs+Z4
SwNT3F68CMSqadXEASa7wSgBmQ135FFQkWrmTLObE41ZcztxvtkFTHTHn+VcHl8/
CSY+6hj/hlbpYMOwkm7CB655js692CPI5iPBbRswzoNIecwdmpa1/jlUeMTL9HuK
kKOIhlcaOgpcLvOGFWAPn11yo9eh3P7AcuxPntkwtoStv8BmDLrCePboLAT/8kaC
wsgOdPKaFGswogNlO3LlQswSm6JNDtBhMQYGs65AO1hDEiTgNcaXklSxuulUdAOy
9Hw3xnfotu5kiwzEkqvUpsAn1TkEOTH1ndGCRU+RuHp7r0uVSN2yyDX1t0SecYxx
ZxsxYzLQrGANti7vdXhqsWMGiU1l+7F4+UmhwytJH6cNN9/MgU/Lunm72uvSsrt+
SUGyBtOiV7nqlKFYlY6L3IAuXM/D1lMeVrXS9mucZqk59F5IgTeoqilse22qDFLG
FVjL3ZMn6guhJQpbrOA+hj3TqzTN2VBkW7UbiQOis6rMkUbCmYE9FT7EgG2PB9GZ
npdMua3oqqZC6hMdMTCliKUe7dCwyhj9U/RiCIkcGeQE2QvIOy1GNyfpBxxtcGy2
2HcqsUwgMQeu+9h5EU311w6yoqL2tQySyasozsx58K2qLmBoJ/5v0l5GpYzvdWre
0QUqhccEqZWTv1TDnThuJddmnLonExvgK+iUEJfxT4PaVMyTUkJIH9oiLc57iAYb
GugzTprw53XKlom62F6+KXVXnGZ5rI4GpdT3JbYbGKIW8mEp9nYBQzLieQdMYRm7
zSjvm7TxanLPQCWt1lwj42VNRv6HAf/Twu/RzU6U3aMS7qOeyFqL9d03WUoO4gqp
uHDZYylZUYyt3h3qwrWiObCxhfyPEf/V45Oq97Xz4mXo6IJGWZkeFtJO0qdnBysa
9h67Uy9EBOn3aFPmeVWi51DspEUc4EEQqA/RPPc39YeQ09JnoAmSFc3KNHrnwli7
gCLO/cXuWKb/cHzF6nS6GbSk36+GrkzPQ+qgOgk2mO7DZW/PwJJ3SS1FPy2TEu3L
onPjiPJ+jyGAsXQSPzfNIXWXjbQ22iPdfoUu4t+3+WgTlWt4zkbb6CjwMBbCX2Pu
XbkbVQJMIf6Ra97YhOT8HUnZFjhy6W8hvDgjsoD8kdUTuy8PU16/FZ7Eru4i2RWG
vgQgTorop8sV8d1q9eoDcB/TtagHWo9B9kM4J8MT5X9vWvxWVNvBtDeoR7p84h+o
MrYMmUJ06BCBXZgc6ZjFacuWDprAPGa2NZvdP1HI2+cLbWI7QJBb126CgIEdPXHv
n8OIGsoBeY4Lzjij4XqP3KfM4Wint0PFVYbAO7pSON0Pti8UMzIVLxQp4LTVOVcd
lrys5d94CCyQB+jyR6nrj3L1IHq8mBA5WNcCCvHMl8tcaahNtl5osnwK3vwUbBre
NQxEUvWkabvFet+xmMpXN9y9ehR2++FUP+La8U9QflaOf8L0mpHVfe2eRcNaudxC
9LdHNYnpxYrUWzcBw5Lmj+Gib6mD9WuO/vHYFm9n+UptegyQlZ76BIfHjHimI2Js
4/U/Ad5BCNnexoLPnWMlC3Toyb6onFsYEIiiJH7BeFG9YcdZXvwRm38n6RWqce5C
wiLJOB35MwiFWc1z4DwXSIuWVKm6FwXgpdbF18q2nfMmKcL/ZYJX3tUtagUOLeOc
At6v59JHYS1YEczloW1y6JpHzNZFJydjhHLS/kLHaaulA+cn3a0OV5YrYMEQPgkA
2vAFPSBzDyLjoOt68fqR/Lkan8b30KzNZvesAMQ5y1+st1dWZyyoiU07m44u6/Bx
f6MyCIADn2PGOUh9i9vMN21FwuF+1NSYaR/O1EN9U8V0/Db/w2dmEhGaHsPFrO8N
AB3iHl/aCYyE03ObTtUjnTzuKCjpeXnfr+orVIFn2XPCp5fzsAQcZcdTQnHMv67D
UaldY+x85yEKTOi85E1F4luNWQ64P3XUf6mWQZNbN+ZcD8NY/1KretB9iXg0Rino
R29BoNRmCkFDutgp3mEFVqljzNi92o4wBwU82Skyf+tLBra2+wKt73TPaQ05iTCa
rg/GF6LnmPYX82e6db7u9HRX3ku0iKHP1r+Itphp761TmwuezHZEGT3h5SE1igtS
wohRhvmfhVyvJSt6tp04HAbzfCop+QW9HrVX1suRpNWW2FK5e3zAmYNq77CcK4bj
aYP3Cug5pGGRL9+6qEWJzxEPZndjQUDh7pq9e26WhEncgFaJs9eNjLQwwvaLJPh3
M44yfCIhCyEZp8x97hxGWutuBKlvYvNzw3fWwWCIoNmzb9/RENM9WjnxnLyT+X6n
IRPU9SpGifwfmRnStg283XkX1YKpkv7Lb29QgTjfCupOAOGDyMRS1imOIr2zqvdL
u4XU3den1i1+gf/U6P6AH9Zt+dF+9t8DMbi7MjhyVBlGEf7MNhtlrm92Od71dlEo
t4yT/cXhONUbqsFWDkZdZeInSdmvC+qjiuMIO8Q2tI1YSCUXaGmIBinRAFc6bBMF
dljCOutfteSVuPaXByiaho6YBTEKz2WHSHrzQ0Mt2TuK192HhkwURoyDtnSmpBwM
uS/FZ5axNxgOsKnvDRY8zDix1VXHbWijNtVzWvBLbuZjnuE0G/H7L6NBA9Sw0bbA
bM1U5RACwivZkuFfmd6cnu2R5ztwVijQ+aUM3pVLWpn1MhyI2urlSY2SrVybTm+l
YKwyaVFu2YVjWmuXMg1w3q2iRju8PZDP8HU+sJoD0r7iQb9gPPj5CqQSRqkw+gea
We0kfjaV1y9H7qzsuteDoyZvYWGW1mDm60fuCOs3b5wXd9MrWnKTlzj088qzGpPw
vw60cz+ZmiNJZ2yKSYHzK9QOD6OgZJ5q53F6xPAAibJzfbB0UMSoX40cmpTOG5p9
kLcF7h0dA60XPvsDx9lI+UmmQ7c6sPPw4jfG4c8prfU93ZU6cZzOHAsl70+0s07R
KTfqHYkTgbFuJn+4Vy2c9xH3HIV8HaAUkUdi1X82fJJ5X71OViiapQtJOz74cz1K
Uq/aC8M7po79FPP6Zi6cSvWLHhmUI7V93O3tb7W527eUfjS5QHHU4RNKLCxqUWRv
nuftl+NMw4E0qUoFcRDqG1fU+mBVipSVVrIzsY2LYHk3iLQDdiDacptCwjvhKqzS
54gB21ivaQUfAPX/EsWi6LVkegTN0L9q/KxOD51e7A3HqIRcJllnZHIbB1rUBef+
n5f907OrNVmfbTOd7ZkkzV3F4L8hF43PcdqhwlK1KzRuMStABQtz0lw/gUkEvuy+
pU7S5GIwuLWqP2biRJBkk5XUiuKalAgeeGeC82NPCpoVTyjmLRTc/ZkX0pxhUI+H
8XrhMTP5UbCaDeeYM3d8JFrLU3l/FfXTLSmQpVDlGhRmidewrDr4PMKUfRqw+IxU
4vl42pabLd7Kvx1csx3vQY0sUxgjY5CirWNtfhg0iWqyU6vv8OU7c8+R2EkBeFLC
aH5dBpV3/YitUiK8CCanvP8VcvmT0PiN1MyqDfrxEgRV4VZtj+6G3iqPHEOR1vck
OTi4fC/r9Asa9WCH4J/JsgwiYDrodunnWM/8zj9i38cBOf3+JMHh7uduaj+09XfZ
OAqwhVD+17aycYuhosUmfLpSj0kYdPgxDjjFuy79GjwBRaNvA30oqAXZh/hLPF9o
m6bIjkbTKZlxaAqrI6Grt3T/e0KkAYbrIWe+HG1Rva1rQsv/vT2uqSlmmrLqbhoT
Nce3PL0bRl6DOkpKqaKU2FHlMYUqjwu1o4MuF9zGKkysPaNZ1Bqg5pRIRM6PkvMy
VITXxmoAz0nvBzuERPj1tbILwQ7m9Qnp2Gzx17Zs94JXG1NGQWtxVs/94RnCN0Kf
iVb9QoQtsrLnDsaCrXjvCwHTIMgqrvFNUSc/QC6oY7VomxkWcYqao7XEv6bFDgB5
5ileU5yS6YcTBeRFSLye8xrIftogjwQLlh7Q/Wo7utGR68eMrK9Mgtzmpp/sXHHX
eypPsGygTy8MubXjmCxeik4nRT7Njt/grgGae/n/9UO5agoXq9ctgwJQd3cfQo1m
BILywN9npOQhK2Yqmit3C1SoZ8GHELyPirCg2P4xmIvmeAcI9HhlpgQPj959xlOM
xyeHXidsMTx2JwPcN74s5n8GbQKaSCQ9UNAIJOfwyGz6df8RzAHjXbrmy7gkeTBS
H3BlR5jYE+UX5e8A7xaDaa3wpuAj9hpMlFMfUMK71txETWQMh9RUmN7mWJlIBPPM
2z/VLWCf/IKToY3XoHdy0dx42ooaSwPB8UMwII/2flPs6dK7pEpyaCkoDC1wn04u
GkqhfNCfQUiDF12MzGh/ZU0gvjPDG+4/68iwhz7UGPpm3eQMt54Pvk3e/51EQuSv
C4+CWl27N/iOVUw2TOZr6V8lrm8lgnWwN0+LYeMd+rlpvytH6YJi+MKGIte3zuBw
XxdD+aEqkTlrqh9SsbHtrSsd3QIodCNFxP1g7Ac4bLlbSHmfzUCOoI4OIBAwyNYx
kXf0YB+zd8YY/rD3d6c3ngU9OiK+GcFMhL+5dif2CpAL1OuvC8473B/h0tBQFdxY
0UzrbFteHs4udKRURYxjfniwxrtBeDlFgiNbx3MXTrCQ6AfeajsM5LbHvWC1uwkH
pTQ5PiRQMBEgSUNuMmIoy7LojmrjPY9lrLNpwxuUj7NFN2rzYF+f7bHgRxxdeAEa
pPggzb//eKzg9u4CKnmfa7NRCNQKmmIoe+3N0WM7H+aBaynmG7Xtn4V93TR+mWy/
H+geZYUXOIzL44bCfisu+pQnkAorl/NgyFOsD4ZW9uwS0815HdbuIgnWvAmw51MF
9ylGjyUnlsiR8V1rlsOhPQB/cO6Cm7Uiwxzd/Gdpg8TVptDBq16sdLXsTwZ8TZCK
Pqt6bky0w0tK0PrG5hQhDtElEO8RBNsm/8OqH31bRx5n2Aj5uWu4st3g9gZHWf5C
B/0iIcts7gCGacLqCXYvrbC0I79/XRQPCJatK95yy8PW1ASG8wN5PYLC0Rc+TPOE
jX0pBPcQUr9rBLTZVntnJC96eKbtzoYCOtukHt39t7Nnki65ASuOjFEEoE3bh7MC
xokVgR9uakUuacaKi7T+fQRQ49ujOvX6W1rdvUD7U297NfwSAcj5m068pvSLTjyt
tI81vMPYE34MY/Ni5kZN5pb5WaR/dVpka5ouUC+mPkfSbkafT0AU5Uk+B5Wxsrc9
O5kHZUPQ0hZx1zdYE31exnhZOiS8rW8SRwLIthZVCRRVcxZp/Fhv7iEOYAQI++ym
rGlr0F7J3NzHP12mobNPNtogB1T7utPLgHbutlL22ViG1zObrFdI11iJxtncyRBM
wUm4hK6nwa0FfAJDLqBcYfttm3zmbzK4/TNwclpH5S7w57sJDYJrL6aKeeY3GpNA
aA3FD7gqXuoxduY4oH9DZ/gxEPsJ5sljWSbCWLOJQMBvLAMWTQJ3mrs4igXCT+dx
QA+4jY950j0tjUeL3y9MorsKGEP1FuGNoB+hcPwOtM9KIqmzqsR0Z6eeYl63UzT/
tfWkAFOwPkNd0ILZgqQPvJulpP4fl9vpkuix9H3cd+7dbAwUu/tgdkEm6Nr26Z7C
wvsqxxfcpaR94aVyU5sIawtEoj7TookBCOFNjTaLd3C1nRp2AoVYDgFooepoVbOy
tFj+oL4nlS6fU3/LiaMfntUgYIx1qrwjtNu5zZa2h2tzlsJLbYuPAIfzxg2X1BwS
sBxxh9nnyr8j1kfo2/EvEifUDuxu0kVD2AGrW1xOuhgI5fnx73M+1leVesvulmb4
892sDZXfomsun4s3ZCArvKtToTIw2elCsVHJ0Lv889wqkQq2J407KSKO6UyOkh1V
6pjbdY7I7foNmAQllqiax0pufDYGDPgks6yk1pSRifxnfbz4yFntRY0JTBMJ8MSf
IB/A9oV1yKr5dP5S/rphC/m7ASMfuWh/zD+tO04BMJWUHYFkQGuEWs61Yb8ZkN5l
SvYryjtkj7dvHH6Hx6lwbX9euBBtHOjET2GnTfs1z8/8DOjoXtuStp4yFBPSin2F
V7O5LnfMtwcIZVLyX0+OAiwclSBzYYMaAqvLdt3KkuYKm49ZEotStZ0dJEd5dSHI
nkJ9bX0rTmEEHqItyTDZUxZvvnbTybMdWXL5uaMo2wJM3I5+H8599lwXzRGIbHdA
EqFpBorMz7vpm1AOzwaisxbao8qujYITr6Bn9lndTPIalpgDYZjV5yfWsBRsIjWH
afJ/sMoHlM9nc4K7whyynyxcSJPvWJV9FYhBBfU4ENLCbHtUPJqa9JNMnSkq7AwM
cmlyKWC2EAkr/gCcFNswGzaO09afeKxktDRsnsLfVnZI3RU0zVPc2CRmw+FhBAGo
WYS3Z9SeW1VN0zpYq50Nbz0hjYiXtF3YLyAsvAJHEDYgx8N7OTSr3cdWDwXRp+NO
3AIGSheqnd2GY74Djh56bbeM7/8B6LdGD5yndasXYAZHQqalTh2t02jYBDVV2r96
rXc+uNG+B4RPmk/8BZScJ8fCgcMFsqKTHXt1E58m9RdwuQnIqopX7PnVT4YBcXJt
+M6Y3Z6Be/urmElg76MoeZfpmQCLr2yKw7l5NIKhIgpo6RZXy8nQrmW927G5rQj1
Xl8LPPDrob2VgdPIusFf0fzSkCzAT+C+dTLbPjNMOyWX51AGIN/H74o8302XPLIL
wqTOqXjeq5d4b5NlyYmNLQCZh9upwaHg93TugQ2wotslzCcpVDkZjpd3O8wr34e6
wTL7v60/vlUQHCqt70Ytj+X+pRy5Be4/9lrSmgxKWhDSPNbGGQB2gM6y8KX62eax
F3dU/uuV0FHXIluoiEYHtcuh7S06AdgzvBLaU0VYnlGDbRNZl9VtjjjaRhtkfDNh
Q8kcbISeFNZdq+hEgrgnSfCaElsFoM7vtUkN86ZD4rDshKEJivvlSpm1UvPVlTpH
nOwCisQAm4ypeoSp3Gao/8DqSShrDI8Gf7QwO6EfO/RBw2E+pqVJQzzm652ipQdv
VUlW7bnPlRnueRcolxkXAtWH5KWPbiOF8pAIEVLazHib6YpewUqfBEusTBG029Ol
RlKz0voqnXL80grOM0h/28NfwteqNwnkvTQJSEpn7WKVaPWmKweytjHGZQL3e1Ho
dpZaA55MI9TRDxdTiNzVn+3p+Mc9SwBHzl/k10QFOJKvr36hF2xOYM96iqFoRZk/
1VflxvfzcHWGzIj+yI5tijZuDcW2XIK5iKlQHV5sgGTiJPPk2UkLqRqXOS5ohFYe
Cz+e2HOboJ/jnaDtI6WdaM3OWvfyeOIPyUY1GnofDqtO1z8YyITq5DRMSyqjD08J
BabdGVcsp9ctmtv53Czv4p5/hoS+3NUKoogSEEGWfShC0nKuUaBNQ5yZ+0CiTdNd
PxclbtBMIC4HS+bg2lgQFovycEkT8eVXlDac2ujMbqAX1z3zBHHsjMaWVuy8rJ5L
ub/bOfqx0sDA8dmzaM+5Q/EWxQCN2h9vsxJay+yYmkmqq0tDbFBBFTKFdv2ZoDSe
exXflaWVlKDf/J5OtLONhCyrjTsiqlQ2W3ydcQ0SAKlYH/CTtmGAtneBz33/JOLS
jrSEiZijKp264EQ3+EpIJnRtFO/kqOG+kaEZepc1SbOuvEUUh69TIzwduOJBbfTV
X6tUUYRXLv7s0/4GvDEZPNsDviEGIRJgehGIblHc0GdikTSdBrRetN0FqPpiNpW2
8lgWT0Om/DjUwWqV20Mmb0IXahLxEgZbMiD8FTohh4py5nrprhCDdjZULvMIXply
TiropGyZAB85Mlf3YZzb63drnKgtOHDD6Zsg3xHEkE9MQqjGvOIH5+KbeMLF7yEs
W6Ei6+p5Cbc3tJgtiTcFHY8+cMP/yuM77m+l71xnrLQ1KtpYZNHzar4eS4k5VlEc
cPGNRoMENVAhUrhpd8mFSKNKUL81uatmiJ6SUSObO179XN/qoDbTjwCb8SnX81WJ
eCzjcQCWJLU7yASYv4Gcv47Cy5CG5a/FFJz/FXWKYtCM/Gx/V9fyRU9wzf6qA2ic
3Mche5zr/RJ4e3I2h3JR4uuFLiGr5nosU7AfziIsSnPTTFgW6JcCuiXa/lOlNFS0
XYaeeiP/pShTCyR/rKkbi67uivklhJo9FdnJkz0Bqj+gtU4/aTohip3xzsftEHXi
gzpWjOkhH3atOCURKEKofT5Y85kTroGsguEjoKpBWYO11liqa8YElHVbG3pXISE5
gvbPwWw/hZJPoZ1JSggLh4GzieETv/NJN41vD0tXwATpHHW8XP63HHBJpJLH2boG
HBuoVJCbLK9c14cKEQtauEtTkmzWbx/XozrMxxpXrtqDmf74TkvoIwZbvPrmFQhj
ZBe04FpOUXo6vZVaAC2KDZPK4WoICZ4VnsqmT92dJ6KEZlFn4OSWMNfaDe+iieFt
Z0gCMo8qzWDcXh7RgAzdwp9wxfYeQge7DLX8B/h5Qphrlynr44eegkJelr/ZmffB
VuHI2vuOuSpo/zmBcLu5xfpe05BBj55haBQbzJUfBKdbrIpI5BxQt/zFxNlNO4F4
hTDC5a+TOE/oOQaSO3xJGQycD5TV1DYXatbLWL5+sumGJrRJexKYcdm676Khw1rD
ZKAW9Aig8au3czmVBDHxjX9kH8u5FgvsYRfDY9inIYR4X6luevSAYojoaAEO9x2l
pHrrqW5yvY6jprC4sLzaNxE7d9JRgT1Sh2S/QJzusEpJifbdbYzbORi9ipNRAN3V
z67XeFWUE5bo2tpTYBAvAIBeEhOHGv9ybenuL5ydpaEO/JfqmWImik2vNxXVGKQ/
5OGyQGOpktan6qnLyziQ+hmn7wmDdKWXrW4ofd5etJojGK6TwWfqLQp15Keam7XD
jWRwwIosein06XFzlY1yn5Xy7On2MZ30n9MsWtclLlNuP7+gEwMpXoOxYGugllvK
0SahusRId6eg2xJiVXMeIRxFHRrZbfetEy1b3fkfEx+CW6hzrAYmhoAJBCrEtDdN
Msd0y824bpEdE5EJ+l5+VSTT8v0gTVLcdzysLBpHdoB+Dnkmx7XDHjuvVKj+QbYm
KSGi/NIos83/Rg+6lJs2mLjqLEFuA+VxXiZqc+PEFoLWE3TQrgwWmcRW9534hozw
puICP1Dms9KgnMkIoDxHk1OIwPVm0Md96Aczn4C4zHwUMQX72Nsm1MkGL5WDfWr6
KyqlIoWsPjZQoJ2cTETNoClgUEvhHHW+XQLY0Jriwkx8svJOJ21rlvrYFwLibKxE
NB7C/vZFc4wuXQVAqn1JRXjQ5DoQ86PJ4opdexQN+hxRnPNnbSvBCJCBAmEbJzHL
yxnCPKjp+2+t2N0gSlrncz0EWa5OXiNhNUeuDgQu973aF6DcajG6UDDrqML7ML8I
W705wUQlMnLFGrUj1+IietDLc9T2PLHQv6RwLf+j2BUNLdSEhl+51PRt0BwPZZuq
IeVCDVZRnqE/jMgK0iLrc48UNtqO1KsYsJdZb2XAWrLYZv91MrwLb+Ud1XVWX7Ep
v+Np3gPrG8GcQqg4TjAjiXhI9IeV4q+rt5W2pcX8Pss37OzJq9MHJ8OXF9+qfI0S
g3H71yahhyu2CEUGPm/YmYNuwkZ3VBmJyru6FKPupmBVQL/vQ3gan+UyxDFjJceQ
A5//xgv6XuvCBieRvIMP5mRftMIBDu0sJHpedpcndod3biS4wb24whymC5BIUPGk
lcyO7JhTnh0QL4qHpx7F+h8sWt6rx/3ZiI6xqQayeb2R5NqshLvf7lUOLpR8Bsg5
XMNtG5C8L007bBrOSNnq4Z6vcGDFGRezI//N8bVQfgAAA837knc6wuNVqGOKo+AN
ge397cb39IPoSHdcJi5DPsUHMfYDpb9J/bZDIqFchmYkXzIvgvVgIogtLEKVA2cL
uZ67STji991YQjlmUvN6OC/XL6+5NtXzyjAd7q5ayamJi0olqxcKMrDkGXe0JhTe
8LxJtGI0gn16/Ue+hN1dBVRDoxKQ0xscn+CpNJH29v4hWP26S21E3P0u8/NhJnUB
UO8YZ8ylTCIJq1Rgy99mTRearvb7mUs66b39qV4uFJ9+MTlcDcP51U8grlt2tXDp
UKOwEwYFkAwc+jYbylAFUN8N/wWn4NUP7Gooi8DUaNflkY2lRzpppSIMlgI7l8cy
cu0eL8X8VzkOzZnj8hLYQfW3VmEDM3P9HIMttp38XgKlcSIkfkHv4lgA06I+Ie5y
EU8MRo1kii+Ug+6Ps/Z55uESyTvAvrtEzA5IxcfvEaS/vCupIw/0c5tp0fZ6gej+
gC3qEtatg09qCmB9t10gxr5rsZq1EkPkQsE2TbYcduSiYOMjC4dz9RK5lbVe4wxV
gbvguvoDuXfB2oJ44y+afbl+vFfyvhET+gCh+9ge28GsDXmwyMwSVBEF+tGHOvQS
cXc+YRyS7r+mv8rUR0drs9KfpH9WSPNmqy7Ah82v3KjmE+p9bAoNBEepyVt7Ny73
ecCIntWaAfnKjJ9amFwzV+V3X9WfdBfKSp3h1M3xOcaWu10oa5EGWK4lyvwNd3zl
OxadruTQQI+aTNAxnhmvo4q7OmwK0N1/6qktPkuKvCQ0JiVWRbP97wI7alZg2qZ1
NUyaKKFtS/7/uLdZgL/6NdfSlTEDDoRG6A9cWS6IGbD4LkEikWPCqRIubiofA7qr
4QxbgNP9jThoKXSA+yP0rPgEqHIyFpDsRAuyBrDRNQwQgH2llNPCpWfVPI86/i0S
yzR73R/bp03k9l6H1ZBSPRaj6hkWYYeUZwvebr19KRfoLdvsmAgtGuxb2KwjJLyw
82ZoKf5GNiSs0W6LvZp51j8gm4WSx6iByyy7Loxnodm2M/dZg9oGOG+1oC0u3hBq
TIX758WDHZVlPnV5cAesXkZWAHbqGlVsEqkgwYqyC0cDiv+C3/c88jWENj5qHVuM
Bc4CCiGXF/7yXhf4VEYd/3r3d6AuZVvvM/KFbAymlR5bW6utTOTCw3l6+hTufYJO
LTPqnG8Pmot745RJ10pZm+OdAunqHvneqB0w1qD6n5FKoezvkSwuGxo8+zn0H7AH
n1XqWBu5WwHOQ693Fz3C4Hc7WKzurOqSPngE/ehrveUoNp2rQxlMl9xWfLFCmvsP
F7YTCExcjgDX0FVvMWS/UpuvsU1KsZlzc0TeKYRaCQuYitCEWMMZKAWSJZF/OR4o
NuilqKasCyyC7SMo3e5hXbB5G3k2KrEVI63ozxP7l6PKGEtef5b0AfJUQJHtnVnE
sfH5bqfSWMrQIfC85nPlDyxz+hK5uFpQvEYJaIxDPqdQd5R9BDfbawK4k3g3GuCG
dgzOQBLExsXTiUwOq3YqH6zhu/IQRUlw2mR7ZHqVummy13UOs+epCL1fQrr0bMUI
4wyTW/2Tp55dFWYItEruBYlaFqjCjLSj+wy5calJfkubhSOaOnP5i07qOpjQZ7br
8qKo2YYwoAEWrevKxx0Nw2yz7gu0rHQTla1ysm5IlzBKR6Q5rJH1D9w43lRJmlXr
eQ0C1sVWs+skgQbobPnRfpXms2oN1/om+ShlSgD94qWVQBEPPTLGw4l8rXOzd6Hf
Bg1zPMWoXNr/sJLyvUD7WlAzYXR8sSkVxhfrKrYLYzTo3Ts3Qg+S9DNwjysdRNHN
/IkZ1z3fymec2zDADfGzqvjJLYr0EqFZ/lc6ToEB/gdyF3MI28INh6r/P3z46yhX
h7ItRs4JQ4Yfk/VvqkY3n1W5G27Xh2JydokkkLlUQ9x2+Ph9XN2iriffL3xXJwa2
cvA2/nosm/OjM9nt0EVquQI9+ECTam2yu3uNq+K2DwIXs2LUnNtVELoc50MdgF6j
N8AlVeElUApIKHWmi61rUkxB8V+4Ib9Yz1C3R1VTtJrtVTThuzj3MAoXyAQqWABm
K9f53KIX11kMn08vKobAyXPCfsBoHcJIq5kODY5cf2gxiZk78P6OFsKv+jZUolDQ
JNZKHoC6T6gSrRx+1WxcCmRMm1dETqYQqIT85T1TvML/KHjnAfj4OnGKJnwEuPSW
JKGSF7UfOaNEwOQb0FcicFH+aD4QemVFg2MhP0/YWxsufAkCZmx6nK6ShBEqVc2P
HGXDw1zkWJiJ/Rq2kf8avYZHDOUwmAeZrQAgWtvG+RKIk/5ti/8/ZLrMaVDELjpN
on1/XtFAuYdzPQgqIsrDf/ectOmLH4uK5n2+fLSKwhUthC5W1KAZKQd34E+s/rV/
O7N5VMhYGlTHiUOLNPDXeFHFqP4sItIsvEi2V/rIt5bn9gAZmZRjCq0/UFGKVE6N
v+oOTgKxnflMyf86tWZWRAjOo3fcU7E9x4EffCRvyNk6rbg6OlhXfPlwvedveSto
3nDYifS1niPSsyresvdV2pzhgKR//ql6BpN/oNXNt+GRRCmsKq5nKZih/gVj+Y6W
PyQLQecekF5smcfhKp/CtfNNtxLO6FxmBd0BN/ASPgPpzaMUAxXhw9dmZKUaG8JO
wPvRbItwwF2i6ZUp0sv4NsZGJPLf/mhayRaEidlcVkUCZKREzG/TXVRjn6VgSPTh
i7HVgDZnPrZhNnhelHETsZkRXkd5OmnxmLND3lC8JNOZlQGA9B88Ub3qzkOASPoQ
DGK0CowD0e8tzvRD7b11DuhoHHCZQ08tbi/4hGVkLBwAfF53ZRVEg5t8A6FvjxlT
p3XUKz98vmDW2mgbYt5uHHba5PcbRM87dv+7pPWS0CsGlJSHWfNAkgoQMIHAvILY
8TMK2ukHV+Vo6uNHVAiofHAEuPAoBde4/k+nChZvqBrqGZkljyjizUZyWK5F2WAk
PnuXqQZtuX5Ye5zJyjoLj4VOzmwfyuZ5ef/S8XNwy0Ub2SYm5Xsw0zyOIpDa7L2x
L1JFQZUDpa1gfqpQQmWIzh0FplYXD8eyjKrr45uL7ky0Lfg/YsmYiCOR1M8qj5Sg
wdsxOK1euBtRn6JmQiHYxHiNG+5zsGmN+aF1EIPHviaAzyJgbQjdriFysUe11vcT
N00cjZgPNofnqhwk7Dh9qaqn4aqh3wxFXcl5QSjf62vi3IHJjoW8WFLT5ffyogg4
SQsVu78g5kttebGBLfXFNGgNCjeUZH0KNUbq8yk6kYFvRwgFTldZg6rFWk3fUuTN
XVBLGj/KfRfc3SuJ4UMAa5m9B3bwg/bHVAfVE11YclXKX37yspWLWeNCFnAHj/ec
BK1yQ5VsCPVeqK3ElwthTQq++3k02f6ETsCdGPXbj0rDO/r+6LC1rhfqNqy8h1Gs
MzPXBLnSj5r1YDYLPXH1n4LjS8hbJXoIGGiz43HtnZkLk1edgpImnmGak27BhL47
ON846A5lIaKY5U1/KUei5tQhhvcgF26FU7cVYHhSbbtULd9eupdjh/ulL6qmW8IA
0vz7tv+EeUzcDo0J1xSl2uNTn+v51hBVsosuU/ckfqyNWHULwNRoTdn7Oo4oSD3f
KEDMrMkF0BLeMMUm9ue8zulH5SLzhNzHUq6BcUMzUCuqrTEursxe5Mc4MU+xjtHt
8f9mPAyAos09IRZBE4XdRlXC4vPeW2z54DTSU3oQkQ9ndKvrohGFMa3T6Di8/X/x
x+Rt28XDwVsaNq4CqMsQNGpKaCW4OcJUHerLgt0blYctlWdHRqslHsAmxI5DPipO
coHK65HPTVi/fSIaof3dWPjQm7VXN1hPYbGAuRmcOlufX9ESC41Ly7CIWN27e8FD
ZG7cNeBHfWdZ3RTc8DHLCkdlERK0n2IP8zUJh8icthTLXqseAfdAFspJmMBY3g+9
8KosMTE8kEum2hgsVYz40QpjnlliRhKTK4KqYXmMOipdeDrHElj6c9MYFL7zGDsE
zKwZA6wBBfW2fe+xjPb+RSMcxuCQjyAuX8i6sa3nLEf0s2sU8uwvaUIHclYMYK6s
MyjxIO0hwoHtEKSc2AYnOs9pWR2gA+TKcHmjZGnGUFXWu57nSHuLXGrSWuDOUyWe
BRHY4WgPPnz7CsP2LmhuScaiXrCtnTxjlMOLdLjMwpdFDwYlNHLg06C6QJKjyvfv
Aw6MyFw8V5dw7o65qmwnxl/Zns3l9d/FORu8TZbE8w5qHiB3dnA7LvFb0g/Phftv
QjrKN+U8gFHwXL3/yCgo/jyTJVAlREDy4UyAV1VVZlQXYzdakfPghLCKRpG6rSMl
GOOO6dbku9ZxqivKio5m3XHO0pHp4ascAr4t9nqRQvEyH2IFzFDy1mkMvKw8vbgB
aAFC/vtDFT85SF5GFXYJtgKVl4ukHxAhlvWynD0R3O0SvSKADCa5HLJAD0weXL09
4MzbEQ4DGdCcODEyosnuQrG04i89pg6/AFQDD17MRjTU7CQkky6RcoN1Fm5RYPZy
k7II+4gZBEIT0vfZAYlxP41NkmkkDCa1CW91mxg0CIXQhCSR4aAoJOjKsjs8cwD3
/geiLiBr6UJHFsmS9CdkYPHFk6Jq89mKdnSQANZh6hfaMsDFOCEdexjNV/jfP2NY
o02mXbk50IhzVTk0COMrbqCkxBGYgLh6/u0yI1P5NKLBBoQ0SE4FxendjhdMDy3D
jEMci+FdGpIy6zu0Ml2IypeYSLWDlDfw5nPATl5rNOJmh33DcuyzF3wWsprpWIri
6nWmDQD75oSGKOpxQ0LQQlwnstSjCHWwYb3WbWkDwqa9Oz1RWYIdJsUuckZdsYpg
swjgPPVArALx85pxCibLi9X+ybgOkV81eMLchY+xWBJRfyNLnC8//1Lj2DEI5Lzu
uEFEUrxD8mYaRkkcmnWGwS3OBUrgpocacSsCT3ZXlTNCZeOv8EuzXCCzeR2t0+J5
4MbOYVURdPAe2Ce/Zpk2Xr0H0Ong8k4dPX6KSiNEb34m6Lly+EKt78O75+BZJjIr
lZ+kMIqb1yGJuClwDmyeDCay97LcbaUS4mTSjC7HFyxmR/se21bn9zds3vusmUFS
mR5zEozTCec9DbxwAk7V7MnbcrpBuvc4eQlsEeMrc3a798aRN3MYhPZFnpe2P94w
LafHtuoNB4QXwPxdKh/jkmbho5KeuAw+/1RH7P9pbjC5G8qV3Wl4wW64r8dBvKRg
PEpLuYT5b441c0Yz5GKFQm+p9Xlp3VjRcxyT/mz47b6B79JFcFMWuDK/u/WMAYTr
Duk0cwBra476I2t78Pr8JMmFk1TGrzHganyq5Fun+10fnBMQCZogJykXPKzDWZhJ
UxrTjEE9/Xi2T0gQzLQljPCeztmeHjUYVxg+5sWKNwchIh9LLAPkfuVtku3Z7E5F
KWeo8RdwqfBWdaHqEjTnXOefk6cSIQd/ZHEfDLccrNKTRk5rJ8/jrLXfPsEuYYMW
ko1ZN4RiAH3I0IUEQE/zCAYy9Rv5l10X1lrWHP5gD+wrMa1WLKwiYOG39/ijp68t
YFelnKo+fwoBFrkgTiHJBPAapow6fRMkjeGhXNrVpZYYKOxsXnyojV33Mib+uy+Q
y5A7dH5A8QlcOp3BdH6BCLr4NTSpgSoCBTOe+DeY8hr5xyMSN6Uh6L7Czt/B+CBh
Rc2GMgnUsUYldozApwpAGcD9OdbZn2GALCyYOPaPc7pX6fs0qb3FAVp7zBmz7DM4
wkEDmGXXMpLCq6mGI7u02/PsqQeq0tr6Q76qee5YVU7FW4btihQSmDCOJAg3Qd+G
6DjfQrguMIoegvsEZx4yh7PUwdM+mu/fDLg71Bez+YVn4zpYgMfAQ7kM+nFuKwMY
0irnD0sxAT/Xg5t2Xm1bvdTDcYeWcNuD94ivwIrtwd9tQzvMMV3BnGYTrzeaMl/V
+DvR+3Xq/LUB5uU26gTobgavPl2ldJv8xfD9CExwalqGDQTtFVdhdK1i8VxFhjqa
0CHDn9f8g8ii3p2iMHLBSK0ftqIPh1NGe/ucMstE9/9sYJVTK4U6UBPkxJj1JCw7
chNb//jxu4EKNJDeHIpmkiqLqXkOZAQV6ZD2lL2gqCqSAPT9BvCFieqq8R4zB1wa
gD+JaIPMDYBY4NKrjtoGsXlQoxwcfg7otzPoHtkthbVhW+xk4NvBsRuunKm84VV1
sTg9+uPs5x0+hrqjwi1YkSL+PcZ/81cSmu3lK19snYzFK1iXFoynQ6b/BPZPRuzS
4a56Sa1fXtQxPUPDqDSipDIUsIflpvC3fJxRSW4QGQcVT/upVOi8u0e7YOO5JAad
Ntv5uplq7O4ZNWPL8ZN8/QVO9sNPmMdN9R9U1sAlL/UV5T03+chgxg1sxxJAP8XN
Ma737D9jQadCemYJBlkFkrFBNA3ErCQB8Y/Wl2WyWvur4FydL1IcExkgfTHONGmY
NvFxODIhinJ4niPhGeGsW7gbCuy3iI0XYUp1wjJ9l6vEybJUe0+eahhB92YOnDA6
cQJuU50bXfQ5dSG3EN4gIDKw6zsDvtK3jzu0nSWzUsRDpHB+7i1cIpojCU9uYgEd
br9oEBKpYI7azuh5rbuKrMlDrrcEjh5Iv8HZ3YsSniPKJ+q6NSdcpjfv2W9CL2yo
/i8LoqSenS3iwuYCoSEfol5hPYKgM68BI/9nt5tew56OI/QWI+SpLQPFyphS4eGE
PhuwTclkud8fS+uM+YKLabUQZ5WU/THgwB109uLIJynsk7RbAwMfii5LMQDhidzZ
98lz6aipPFT7xFfQAFNPz4POwzvy7TyCtsnS07LuEjeVrxXQaml/uF3Nv6TKaxFB
A45CWx829cGz/ZTwj24BlXAcxTZIFwjZXeWGqNOnNtMxp29nD36bzbpPAO1Yg1hP
hjmqN859HsZFmowX4n1dy/xClb4deE2Zt+STFn6HgL+kt5NoShekd3D4bXixACns
wg3b9V+yBnQCy6ZMMKB5yCkJC54FZnmCA7jJTmf8GaeiZN33znDj6sMR9tddnr+c
3eET5Z2VvQoWX44LXomSDms8XMwE2YQuNDOCblMQNtTyRwjBixPCdPRCqtjBltXo
a+iq+KIzGFjPiuERvjzEMI6o+Ib0Cfgg6w4c6LRKFqr8/QnNIU8HyLy6u/0Lq4N/
kw6ux1/WTF0gGgvde1i+/zbraEDDxKiWEgMcaiMN+W1oLEITEwbVWR7P4bfalFDH
ycXoWot6zzz/pUMVjbm8NFGX3PaVfZ0gP9QRT5pmVhVyPhWl9+G9Hlc4wcnrXOom
SCz6USy0njXBV+seo+2QNsWL7TtWzL2IhE9Vvbq1UNyouSgXT6K7RR9rnR86GpoR
qPwcAsT2xmEfUAkcBHkTodShxYMhSDWmjjTIFQG5cQMXMRazXm5eXy5WPpqal9Wg
JrgEJ1Z5XeiMGYAAexqZcjyk//2onbTX7MXU9qwdSTIFBzpAa7gGCU/CKo6WqGb6
FkOq0KIGqFnJf9U04DD1xJKmHdHUEVpFDk+fjBac3Lcmhz9+TQ9ltHGtyUA7krbm
ROTmYPJfHAcoinal5yMsitz26TwTpiw3pEYY0F0yhJUlv3Go1CHtLLVtjPVniXQH
C+DtW37fAcVYIKbmT2vsFsrUSL1eRSkc4JKDoqpVB/Vm0B0yMyPxrXoHMKyHMOca
ocuzS/SmdSK9zTftt4BtgpspTOsPN4li6y6BUY+cYKnzkcgRPfzsf889UQOJoI1C
i7DvQHO5s/rwNMGiMip+vdQGLLqPcHeSrAPayzZv4dUHYO958cA38dzh6lxectJJ
trlDlIRyzPqs40itg0IzLJ7U8AvzcoyNVCDnmQgIOQ6mdem7wMa/fKfdqBx8BZmj
NKI/x0Um7+fjOKkOsXatQSkq2V4JyrSAMfT+NpUbcBrM9CdesVQJPBV4iREZ51G2
ZjECCf1ml5aP5hq8u3ZUfThvop+uuwCM4pfjq11j8DKMnrlVJetkFlqeanrZqdAp
glqjkPRLWtdFZA2LNOK5vqmVrcIjl4DZwDGqDAnHjmLyTSegaVXhxiIp2AGqNPVt
krXhGYiNsYoL9IdvpEPZ0JI/xLXE79pGZRCc4zakJkx/ZiRACTf7uh7yTj0u53iX
ewB9DzlGj2JQIpw/yrtJLFmzs//jJB0O1bg/U+QbAIXKXyNFNNCsnSW6bbUtnWrz
ITyFQvHM7kVCITYTRjMPUPJQoph21819LD0fo0xCkO2MNLvVbDdYH8DOYwpakaUe
UvfmpzvwaF9lrRC28laC9KzluhN/YF5dUYV/JzDyWUnBv2Mzk16I5sTZHGKNcGP5
psSa495h3jJ4JHRpAGbaw/VWE9hkhTbJaYqemszXPBjag+WmusBA6Tkq1r+FO0JK
i3rFFqRTb+tQJmm8e9IfoGJF55Zqo/oUezzSNVQDU71pchBRV2HvAwDeFrY53MW6
vxEpDR2yqHERZ11R1+NBoVp7m/yilxZxIIc4+V4+M4lyyaSWjLXCCRSSgNzpe65s
b12vo5wzj9AKkGM3Q9ltlaq4cNci1lky1cvHFYYTfHSgDz3hGvjh/1WkYUtQ/ugJ
TF13a9yHaKbSKgAz3BN6KAsTdLEjUYIJ7Stq93+5r2V5079GvqNqf7hgzhxfLYhC
lzdtiSMTeKD7y4FQCfF1lgbae5KO4ApFtUPoteTKkoAzN90qu2ARJilTKcAF/LZQ
BS0l1aGjnNouuvIz5AfKDiIgralZesIacXVEJl/ooYsCzGpW5ykc5BcFNycUaoE0
Xk+zJ6u+vIkoSIVxacEif1SPv6ycfEUaSyZhcfR9saeAMEVB3+uIaNStu0ffJpB9
H923WjfuaBK8zdXoJgh1/2UzaHOKVrqisb9LfdPgKNgJ1E59dv8ySZozRhA00Yin
LezwY/kAoBk+F0d0dzjhNMdBwYkcVMHgoQWhMa4yPw3t3OxbOU/fKvh4dscHMSH1
hhQItogkMRYMXGCrG0xOsBDlJgMP6n8m1lZr7XgqLn8U29y3ZMy8zVD89ToZxlRr
gMvuufs2hbz1rnKtZFHw/zafClqyf+Z1YoxzrN9j0MoF1TsuaEoKsIH+QndIuZT/
cvJnL1Cjl0X2lh8tYFpHmdaPWn19EF9dyqte7PkBjYbC/dXKx/IDuKorpXgflh2s
tWnJM/qPaHd9t+ioVuCxSu2N3/7bDORQNqVz5TakuuQkAZX0VF6l1e9MEHThxae8
WeaJ+DdOrF0UWDYjAj7tmWVmpSfp3kgJOwJEi7F7NjUI+BprAP/bEarPJ6HiM3Kd
cBib2WOYynLGNI2XgNY5g6JQpfzZLAb6oEF0z3/ltl9jzoW13QdNQsujs1y4ySwC
/pXoEb4KGsjaLkOduTD1aWKpKWlOP6fuKgHFVOLFmea3e63coz8C+nqFoRYzriiq
Fnhg2ntep+pQkZglPP/krBdOLD0/3Pd3BZ6b89Md1+Fp0HBgsiPD+kZ166eQ6fF/
UsM8NdL9u/8lsth0m0rchLIBIs7/9ToP3+PIFUp0ax9hCMp70c2X5rgreKVJctZM
SkeIrE9X5MOTLFNXH+/KPlhC24iXUSwvLwBZTKpfIzYl49YoZCBDOrgOnY0zAdbX
Tb1IjTgS4KluW9o02ajXugJIjHtd6SrbHvzC0rWqQ4RtqIfS50y94Wi+1CTEiord
C3SmC0OqEXm3GXfdxsBvt9oA8ItDt/U0SskdZJc7AYcXo6LvFt7b7u5pDDihoST1
IEId2vrtlEGAbUZF6srShkgmDg3g/LcndUY1/FLWvKLml2HAMGm1lYGUYyDUJgrD
KkalyjJ0xFJetYhmDzNbFia0mcLOSgOdkBiFF6yN7IeawJRTmS0h1M9+jLTAh4vM
OvF2hMHrPFe1P//QGscnDGGcvN4dzU6fD8MIFUW6NDk53qIpuvAezstkckyRY11g
tOOj9T5zGS315Kl6unuNFUj3f5a4qGwXYJVPNBmeXKP9p4fMTgumGBDrZtgh3NcE
P8DnxYFriQPgmm1EsQTuMUHJd+oYYWE0kivtwQqutfnRnrpd6v3yI+6+EpjMFgMO
VzNCb0ySpNXeOJh2RaI1IbWiMkMk5cbKz2vbnnzK+1Cy/DyFft82f5gcqIFxdpKI
rUTuOnYIeSPsI4OqJELR23I84/BRCEbhtIJp3xbnka4tvL3oW/EH/XTQWnm/4TxR
G/TPT/ArGADKtX8y3fop/hKRBE3VE9ya0tZDmClz3ax2Zzo1787KZ3+TTBCZOE/6
fOaRd+zSizA76tHpYGCO3+QfITIxCBTer0zFJzuBoZe5ce5HZbKLcNC52KwVEXjj
OTsz2YtePVXYuNGwJH3vK/KNR+1JeW1/n54FOQWQBgYU8MR7unZ/njIA2RnsfYiP
9fOGQeDQiSNdW/EHlN9Q8hX5XJOi6zLtlGZbLJOZHJItjZkjd3fthFrMKOjsvUXl
T7C9QAm5vdcmAA98S5+ie7o1Z166HXDhoR8EIYMxTq6nY8mJh1mzfjJQ7vl34PHN
qJhLywIQkH5K2TPijTlKxsnD/GxI6eknhhUaerbJypY4wnsJ2rG58mS5O9OWodb5
cKP1J1uRYTfQr9Fziqf3Cp/7dnyBUovLuT/6agd589ZQhF+bioZR8HwMZ5ICvLER
ulgHbyAl2CSxXcAEccBOYUHcF5HRg/oFiMLTTazfRJe0NokNnHk0NwkpmY7sACS5
n6JYv4buOTRe4wp8dndxGfn3XFm8CtK2JKJLW+1H3A5lqFazdAbF1GKAyL2pASVV
`pragma protect end_protected
