`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TkhXJLpBL4fLYn13vlnHssU4G7dO6TFf49nVVpnh5iQUmq+BPf4G7u9defVO/yJE
c8ROsnO/+xY6E9VfeEBm2GJNWzUwVpm2zfJw/CV80uBVxxiq9hE1Ai7q6YSUWHFX
xbS1KJLaD3qQKoHZK9toWZrxRFam2N1Z60dK4RvJlj8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21296)
+rcrcd3AStB1JyObq92rB4TDGJqQnigmnJFM/+QcrMfRZwDgT/fvZ/HiKcOGpTbk
rohZJO/VLgGRN6hotst2JZgsOux8VqpmRH6txnje1MzkcXRzP+2qKX06mVxgKw0A
d0J5KKLoPm0FXtH0JPzmJ+TDUJ8VY5XRzYdapLV0IrVsYZ9aRMTr6fBuxJpnWuzF
+ymSVSQ/3r6Yar5E68qf5te+3ZsYXdBq8lOR21KbuLfkotgFa77e3VUQA4SHbrK/
sSSRUcnPMVyTsQz8Q4MEO+6zRVcPSxPRLDouNkudQMe9RwofevfW4jAMH3swDvia
aq2dLlhrGXQCFhWzNE799kteTWxChcsLsjzUJstKhE4R40SKuGpa8r7LNFTqicHQ
H2YMOl0g22NV6Rd+yyGC6YfLrAsyQF88kMrpigHIOMDXBtzuE1qnHwjctbINUA4V
DnScUBI870Ws1tsw3WfejP5zj5v3i+kAAY0bwGhZgVkrJQA4UE/UiNxJ0lafEL++
8vFbmmKULkv1wQUdjMaWH5uUA8jO7FNWzI+4oPlzkdIKeK6qQl4ADBDa+ZpA90O8
R8qMs86DdH9J0Dl3CQ41BZcAA9aJ8bKNbiSe9LHjfYGHEg6r10rhE/jjHvGR7eBs
Cyi48kAnjNkm8NIUEQX0qhYxFJR3uHMPLkFLyoK7glTGi3RL6oppTUVwhwhXdVU2
xEFLFIehQxsPAatt9rD4RrufRGGmBWewj9UBFjkV4cJNJfcZj5F1JQQ8/HnOX36w
5WZh3mcR4gvaKxceRUnwjGZ/O0ZhUWos7q23ozS6hL3d1QGAxnWt9AHwRG21BEU4
TadGKy0Fpf0xPw+Y9HWBNhq1JLfcSmUGlQbSrJ41wmBWNxyz5hOEpNzf71FYWhYN
9Y9rLvKrTRcKlGcU9ORszMEqhQNEllqgkAn7i1nToVj1Ovjoc/VwtkY9P0/Osj5h
Vvqj0upLVBThZtmDJNbK/3bBxb5v+p/e+GpOUtZoWyxO8WJeAO3jmJFzSronn71J
8f4QJBPF7Yk1qHY+iTmsH1jQvpv66CEPWA/tRCmR/UFoiai0w5NPgpw5hvpb8x4S
q1cXYEJIaIq7C49GZ/EKIgYViMuCN7Gs15YdfzRrIkpnXcuNDGLQGB8ZD0UIM4wS
5e2RBSZUpjz20XZ2nBUZAXu+0OVZ6O3klCQKsS4LVJsQ3BbdRBG2YoPMqAJ4gJ94
yvPPmBa14nNVDnuzPNu4kVYPFIZRXzZz/zOxyoZgqWkZJeSWQNQUuAnRKq5bcBGm
VwGYaEZBWmheSupbJA3vqvxM0FfvOV+X8pKXBQ2nTOLHNr4vu9fnBiwij92D/XY9
BXj42wTyyWhK0Ak9VUBFansqLere0Y1qxRJfaLfdMex97O4nQjsCuD0Visum2s08
HFdE7JaP8+lf18aBym/BS5Tjjj/NJEPdwiz8EShRSKm5ZYSMi8ujRe6hPXOtLQYi
Uz/PQ+uwOhzrcnWlRktpOnDNgXsBPPrAh04pWGDuLHsG0Kwm0zLbH8KeCSLJtBl4
iErqQ/g/c0+rdpaEElJTY5jVzVuQN1RNjDgpa6BpDuUTxb2wRS1rdSkyWmRSp6iA
zMtsR7WDylGYwX7ptWWc3FWfYPxcs+qTFXec0x1oF3B6xHsS+v7J6IcYxZWGk4R/
AzUa4tVg0KmceXTMdg2TFtRx5XpsJ0iVL2aE8llTa0XNhlfCNkxLhhqJB3p4eNNk
mMezr8nWkbXh96pLsbRTkhLbJBA65M1AbNIiNinV493tZbIU0o6marPNzex0+iHR
vJZU6Y04ELiwTe3eXsfmxVmjriRiGHiwCSSIqWIFyweLtKGQZoOjxnnJKxLVqXLr
3jT1cGWDZmvjdmkyikPbZWl4E56twwRKQewtJmPY9VQx3gOIqRUjaEOQdIYgNAvW
/qesKQw+0dk1IaUvbJtVdBy3Ej8sefpspS5sTD9YRFJLMgdnqECjWMFG1KlXFxcu
X50zJUYYwzT7OofNtiNHR6Vq0MeMbcB73G/+anNlT8VRL+5NWsDGHV4pG35zuV5k
+6GcOvGOCcNxA4erREBVhhOf4RfUrSTRWLZNDQEKTc/PCqgV9sJELQs/BuBJxVYF
sRPlzOr2X4D0xmuZa9FbsqeBPUyg9aYzMgd1RnayJynNFZz6fKKRFzEZCse2/xV3
NZWNRKL/Non8Z6KNPCe9xYzEC4UzNHAlUdhMLYN1sKrqNBlXasDReBrhF4u2Y6Mc
LmaSG413VpjYipOCs44wlJBrO75pRz2X6Rk06FvzLPA+HiWseRhT1dPPrnBQCYtw
5ktJlcvE4PF40Gv/eeAygRu3paDBq6D3sVw1PK1vHeqdvv1+oxwziWDDcj4AqQx9
VxQBo8XYkK+ZuHWZwRqZtpaT0/qmwblvt0L5WlD6GlY31p9u43C1xRmbSMH5dnYc
cWV3j1KEq57M5D3vjM4y9cjUG19yL+8E03Dwrw/R8/s30s6/VQdd8nwYoGnMcq0z
l7OrO4c6fKrpLl+gUjQ4Qa2KtYbvNR2TKrprCL2Gf6vmdupifmWTfYmtz1QlQpdU
fXUCIpvdfRaWKnDFAFG8h1VSjh8dFEky4YzYnJJq06427B3YhI0jnJBjxXvoveNX
z+scHNTQ/4oISGEJkEz/Ma5N3dOfEiMaHor9XxrHfEv+hZPbWLPsh6H9cHIbsFYQ
H5LMU2uiD0Q8pklSsXQmFoEppmLpAxLi2sbZFjwjgU9BpHm6xW18iA2JF6pTH9P5
G0aWsV8OdTmLWRHKeFytiZ60zmXI9i0A+JJsciSb0hvuyUXd+hzx5KqRUfZb93wv
LjyH/9Ax/ydVU5BfaaAYGJp2IErWoSTYQ7jy8fDENFcOD+6NcP83VkEA5iqA40mU
Rhgyd+chc7CvcdcLBc3PS4oRfOJl3V7/GBix6UX7qbO27aSRrYUkD1vu+LjAwa1z
u5JCDM0z9ib6Lkq0mLjW33HdwNA2uML6tS4BXIwoeMwytWnMA1MManHsob2F0Hbp
a57Kr3ulXVU06HqTIKbA6dvTKF7ZWRIq/dNx3tbrtBQa6VNWxb0aJbq6XnGWU3wd
4dEllKEdELpCIJUhC80UJs8AvFdhE8GrKSifsd4ZhljJCubukSLGj7dzLnSw6BpO
AcCbHmKqnrm81Lwsk8U9TkMJCI4+jH7+p9mFRWShz0uXwlKGVQY6m/OkPdQpHwLg
BE6yYninU9O0aM4RuxSokmnvH0PhFHjIL1Ou7NRlwbbhfOSVYoakpqQkXiwGo4Nb
VmGoxIr+Go9aybSDzFS1OBK6zVKPySkDkCHV+e+1oe/jmEbxRO8OrhtzCj8oS8lP
i6yn/4Goq7qwjjMz4JDLv/vLN5Dxlv7Ir6KxEKHwIYg0C6a47u06GNJEbGZ/pAs/
vJWnO/e+nXI19jGZAoZven3OEgPGEoVZbvfjqRBe6RxGGL5kRVndNtx6Kiy76ni3
AGtd6xaqRHQRBIdRhZd5d1e1aXBf7/SCWtTulyRIOUEtSbvSbxqBOQjZTqaD2deY
VStYCXHTfhNjupoCwPKkiyy48eEWdciKV4wBm3ydhLfrfqZ9O7NkSG9v4xVTXQEL
13jkx8kvibiRfv4zZ3bY1Un2FDahDnqZJgl/fKeE0SDhp9VwVGjNG8kbp2Jyo5fE
piWkXfr72Hm4tfWbPbDviByokgaHwijMIrqhf76ZwDt6VCYAOG0A9tKurie/5QCY
I4TaWYS1TwqASz3JhL3aVkAZWDv4Tz1D2uGAI+xEI6VYQre4dtPCCm1DV7dl34/S
DtqxSdtfwlSdwOq6UWPPwWCtqhRLZhWRkC5p9Z//CeJ0SijVpHzK0iy9Db54DMjI
t3oSKZLU0BXmE0TXp2u76LIOaYxzVk2W3zqB5hA1yi3eJhPBZW1Z+qPjE5KBapfS
ShL8WQseRXN4zB/6EAuxFqu9ROlXruqEU29po0R/Sasl1J5j4HTh8LUbxq81svuH
9OLxXnubd2PMNP5+BRQsOIH2zX+wRfU6Fwkw2uzn4FykfYKKw3SJi/Q+ferfNj07
XSzH9YCz34wrEYsm+ry6tsX+mRoevjns9gH5tIgCcgEKTNBnnavxuggtD/ahwdX1
yznpOxRSM1Y77ibTduq9k5z6wH+dbVCIykVdP0w46ekQYX4fzoyCvH1cp+Z2tzCp
h2a2bmweMXajN08PMi5OqWq6aEW70nyoyRSZOLTFtvdBu9P0PIwxAJkZeghWH6rg
gJZuPi22GCue7jJOo89mqxp4gcPsLMd01Mz0J2NSRd5zQpWezlqlKzRQ2HHegUYM
zi/BIF/h5m22LyFrS2ElbnsVIn1X6MjkoxZHmmVbaHrPxXYv3RLN6n21bx5UGeHo
LwVp67sNhk8KwkM9jV/kMGc4/Fi+2TFER7lJ5wynNpv+Jy1qqX+OY+F3nbkYKuzm
ucZ0fGJPWnWcvELsgul9TMl5rcb6phBIABVcEnajNjMxVGRJ0Ue29cAgyH7Xjmrv
dJXRFIyf0d9cXxNOFWm3SWfZxfwYij1HeZf6GTBWk6ezuHn91WQrt80dwtBBPqCH
umFOxsZOX2cE2CiTzvZylEGgWv4XHnzCHH8FoAQ+N0Gzg5BBFkIlQB/VH92axchl
4wZdq4cEsod4N+7Z+z1wsHOhpqURyDANJRDs2A+wzbCCLMkFNbe7EHzjp6ZJil8M
QVckY5aO7wBnQaUjv8SwiHkmwjdWOh3yQHyuAErIqu88H3fUzyeEY36KKF4dqXwJ
6uAONV5qNb/zK6TIsumMzHH/nD3HJss8P+xQ1iJZd4uU61rOKIgrDvK/k10HGnTo
KL4X/KG4vWtfq568fN7zQZkTBoDdKZwNv9ln7iayju2ceqmhg3wHT+I7jusVHh8C
9sFCLAAVpGA+7Y5IQprp6qtB2ZA/9TEAu9R1IW+6SusWQfY3IIZrnytF4ZQ40ve9
ef/b+dgfMhiPkN2/CmRwDSh2hScSlrYseP59MFVgXag5L+plSwXoUCXKTRBgOEXP
pVLdEk86qGTHs5tEo9OG+LhDhC6Lc5cjfUbhb36Chokot4RjGsf7+mI1aTL1bYPC
NqBPL8Bn/DHj5mnbTe+4FEcU9g4DHQuG41o6LpCYdM+DpDCy51eJAKz9E0+W2clO
QJkDDTZEhRK4V2szuwO0MtesW/Uizoo2YUZqJLcyxu9zmQk1tMCIQePGGSvxItRL
HzrS0yKvVX1poE+NTEKmFkk4P+GQ6brrTaIQCb++Sghhbi/qiFlqZ2fBwtRHzL+c
pmoSNPzHghgUp0OseLsLv2qW4LqPeGq/3JQyJ5C2mzX21SWCrugiwhQ1sDrxGi7k
uQ5ri3kZ1BjgTh1e5Q5c8XPvgxdAy1rxiMLHlSLRUlc2kr/O1VqRSe+xQH+4aY6K
qY3a+QE6XD0rCJYxl9XNgpIqhCgq0kPe5twUi0KRStTUvcvYIEk+BzAcAMoJdVTp
TIlL/1jYI80Qtz5FowT63oopWppOYJkIJZ6JM6Oa7ncSqKqPmc0CEPC54aKvdYiP
Fax/JUwmtN2uaiZqCHCHKB9J7Eu0p4OxVMKgk7CJpJPkBmmvQoNSBe1+H0w/suWF
zC+JyiFieRAtu/vfQFsBUPp7HR1cWVvEOH0wNnR9w4/JDgegd/mQ1K2hP8Gp17m3
e63CTXKIOPJb4CJ05KivlLNeqJrQXNL5LDX3Y2Oe2uJyFOOl1ahpUXDwLDR39WB2
GuxlaQUmpilEJe09S8wxxxPhcJACEOKOWBpQ8Ad2qipb2gFY1wGAvWlZYkklUByn
6u4Y29B2VZLvHrAsDqLSS4oweyGX4SamqqzXqIQrIXquUTOUCD6Cm1x3jZlIlbQL
/CquVQsYLx7Wj37q5SoQx0x5iVqLbRQfHk1FNEXKXd0YQiOKKp8MRb/ZjhR2uyuK
Zhm2w5nZt78CoiOkWI/Cxo0ueavlg+fMnUZgls8yLuabysBoQ8R5otClaTqt1I3+
1kbSXHD/ZzTQOvjeCwnkgKwYbMwUguLlfk8tPKEV5JX3CmK9sEjr8gj/ypYdMkIV
BU4Q79qMcxuHtuwtXEImO05q5RwBsDqxMFKOT9DoFEEMjYU1LLD9bF2ycxRIWqbc
nbZh4EXbZPUYM+jU9O6SuLmu0NjmY4ubdV2VCJo16urQ+D/j8dFhMqBSIYnX6h+i
cZddM5g7ZfLTzGV2bpu3fsBHPbdzYL4G/rK0HKu04XIFTpXqwpjZLSjiSMknxcrP
mcm4zEoU9n+/E4UhoqBLzl6FjSUo7DC3HZtxZkxtzz3XZIUbfbfCE79vbW0e8Wbx
ruSrIXR8q512Hc4bMAcioySGw87MOl2Jm8SQKA7gNxcRh8epSW1ZZzQUAaSMJBlz
EuAnvQTC0YT5YWAueeIfaNgGdxi5Gfh/VIGALDnvYUff5Q/3OvbCE7PjCdkAIsir
A21nt4Ma+KuGaGZ/EFMGEsGAX3hfJDYTp0xWh7h9G9+GCwffYHbRbQ3Ga4rLpji2
8+Esk5y04v7ViIJqM8o9t6vg0owDFR4OAzEuLrnT43UB3mT9hqbYdzPedxtEqH+a
r3+Vkx9D+tZm7tv98UiR/hQXIini9WsoRc8gsvSQCKdfJTozAfaNs5oFOdq03OhS
2KyI73BxJ/sOvtcNDp3xrc5Mi0oFGdFxoxJS3yXLT1tXIpOCiU/gt91CGAdhPhVv
7m74qKxs2Nyu3U+6zDdcoNrHXrNkH8AjivBwclLs1uyMXSVOuCUBEi61C+jNwbGF
xtSLRaO2l9uRfi1uvTD/ZbJ3TSLdk96HqN1fm9crDbhwxGd8r2GBWW0yKanLAh+R
g+/xDPGt5yY3vEPP0mQ1gLTco01pX+MK0ztJAGFOY2LOG7/OuDRsAhu+XScpvNlr
a+XSC/BMuUrYdpfE30jR4kcur/YNQWXIrQWiiJ3YmJATJBUiCeUP197LUW9SCTbQ
lVeX1HSqfHK0M7QYdjFt+Hu8gIBduDlXt1KPpxrwjB+1iZW8K7msE1DS7XyMZifS
RiugZg0NF8cDigSaj0RkizpgZX4HXEWkoE1k7zeRwZCBTIitR7uvMffryz7d0MjU
7+q3FNDMu6lnC+z+t/RwodTwY13YHKCFLp3T0wJAdhwSeu3Qj6FDv/xupdwjIlNX
yfE3BiyOHkc/0dPHANz49QnvCPurHRs5GPLHTq3uSS0I+DwSKad3L8YwCfPFA32B
/J8xDyMw41I0WFQRnVwX4BEMlx+W+hCP0ZBuI5dKqGeII8c9spavDVMWoVlm4Tmw
FdibzCZchjD1a8XVfS7T/HwJ1/7iHMrmLRvjcE6SQteHze+C+ofaS8UOBEagOj99
t2cvUc/F681otqqpCQkx1F0tdV4Xrzp2NUveG0jpfPZgoZm83c/tRmmIQbiyxV3U
miU7j8eA0In7cFuOzZwI4cXzOp9Yt8ArTqXx92Jj5se5mDZZn6PRq4BMLhZOgxgr
bRGt315w2aWrXl/EdpGNy31rko6nmYS++8u9FXWTe3mrm5LjyU1NMY4G2rjwVkF/
ssX9YfmZ/1KBd5Kf6kvDPMYT0XPaN8rkJ3NDusegdabj1/N2I6C9PSC5Zy5Zu8XU
WCiVPMpcCNmqfNsMyw0wLPEEazX/NGIb4gOUcTwUlrERIGOHcqJ8ynUriFi9fuIR
DhrAD4/ylJJ+33gfvd7SjENvyVe8cNCYFGgC6ZmIj9s1YdVOs8zuMmvUWiJjpt47
8b3vPuFJRvpLlOkG7NUAhoxO7Ar0KdISYfCmIxzWjDMuo4WPBKg0XJ/OvA0Nc0gq
IZaKLxKjF8bUqURewFknYjlNUtcf4JBQteQRMMjvg5SuCos3pUSX9poAay1z19VO
RoYMMWnE7UYBMyC7hharKK2IOos49GCC+qMGFFDF+vZZQ9h3hp4+Z9UzrYiCW5vB
hg3puzvmW2F2eOTud3e0NInE83imQUZG0H0RM2o3B/+bu2dnnikpPZ0QdmOQ4P4b
RLhEjLlxVMcP43bOSJ1RMM52Y9x0PrJ4o8Bxg8ugJdP8AVi9Ls7kmHKfX+SbsGVI
6TbxvJMudGTtlkJd1kaLTlU2MKJB7xCAWYN4HSZ68bWzU4SALtLUCgqxtkZmRIVn
KCkzdqtoa2q3Jv6Vf0Qj2QvGc5fAkSog4oBuqCZjFpbOfLRwhqmtiLWrY+VciWxe
Y5MHOmcet+hjAfyXOPIhmc97XmL4vsbwP/G9FCYM73MhRw0bYoNnl47tr+M5aNAY
OaDkOFxKg3FG/qbyiIBcgHgHt4MaPPpasUNyBEi5XKA1vOcmCPTiWCyjIf6+ihLx
gpdNCx0xNEfXvK+Z4Xgrf5wJQP/CZ8bjbfVgGsduBgxEGxz1QxbrXeTn7ZREcUi8
NZIokv1QrG5oK2sFsnlReDkF+9AKH23bzrfMIzr54DHwi78ZG2uAnqhbJ8Z+QQCE
/IN+qXAFWKTzEI40QRV5XY76KbLev3OfOUiuq+f/040uqUgqLF9TXcG932A7B2mh
LNoNIYYKhEH8LZFlM/GaWKeNGNjRotAgdN7CBG0HRsAnaBLVLMvXbXacl/8eCfk7
O3zRZlnVYKM4WGUH8Mb6CNB6ihESE/0SMC0WUhQVFmqkiKtTH6BNP7ZC2a40DTAW
ccQqRI+eV20KPUbDykoYufngmh9Tf83KbPRMbA0NMiS3ohUiTxjX1sCPkDwukAsO
cG+7gf4CVkA3sYLRCQC901dZznAO9T9j5v943qtvU9Zaqie/8Yr5AMemJBs0kAu+
yRBlHZ7E+FiKKtHSzx+haqTkZmp8GQE5ihZrVMmkEnN4UsQtbcR8v/4bAToliukj
3AH/rtrHfQkyF2fGfNE7jBVf6PQW6Pz0tz53JGUCM45clNVQ/FiQk8cuVIbqPocL
qR1fDjpioym8D/VK9B+NEFoe2MEK1o1NfOlOPxXfbvI992sD7KnhQTgiQZP6XEVO
wCj5vmkVuSHhNnL5M9LYXSwc9W+cTG9HjfIxZ9CL1S9K2DpI0P/EXjQCh0wBp8cE
EdEAlAoiLRK/Zxr3fOYNlvG8Cpkc2Yp+P6tnPLrOl/zcVOE8GMj+xnLNw0FEl5tj
4ldh3TVokUYoDdtMa4kDJHY9CYc1BKZcwd161JkcY+8pBiTcga0tDkbukckpcAy6
dHn9dwQfMMZMVXmUHKRnBdWCgySexm9MY1+cZZ30tu3i7Y84K8aMJDAdzI96M3Qx
TUT5YGC86fX3madGmnW+Sv7hq4WmFDlqayjtWz1wdIlA43woVjLgGerI0GwhnpYU
XrPpoLBVHB1o0dCoqNXdZewJIVTvdEwuYzJ4vuIMZUiMr4/3vR98oE+iu4mxXv6E
sry0fd9uCk/Wq/3TjsZPM8iEwmG9K7LD7YUgNPiqVBU9FTcH8Y770+zDuW+hlI86
epJu6k9yjCahUWM3w2CN3dTjcntiE3T6IXN9tQy3PWpDQIj3j4BKXOpRT+mooDWN
6cvaittfFYQXF6S9cNriBlnHP/zBUQRlnV0TCZxoSc4wK6F4Hzq5LHdLskOKQbtR
1nQOhpPS6mZtU9OAavr43ByYHJaIaE2GeeWoEQBmKUoKxwXqElrPyrtwB5GA8vFi
2QxZqTCaSVkCLjRfnvXbIN7pZ7c7xX9JFxQTrBAmQfQEe8gltAaBpcZHHruJ7gaz
2/DGKNuxsLpXzxVZDBUznojFT+FKlOlYlT1BEtkmx4F9+AS2LDg70qJ9Ogtgl2lO
pJC4uQIIzBj4vpFz2tP/Ck9tTN2UIIDLy+2OZRQBqE+rmSKnbDCfdncysToKzHez
tKQKtHWhlD2cqF5k8Seme864GLiLlZ+fOxjxIELRnWhKHAv9tw2RIERy2sZNUBYl
xT25z2RDRKZiqDiigefsQSpemPsLLHZ/QfH0seeiBVMiWzKyyHecb1WrlZ50OGEs
JDmagMcV5M22f7FfD2TKNwaAszaZvncpCkxZGR2x05yfP2ITVEFkHKrsUQpqsobR
stat51RXv4adsZDWKLdu56JWxExk86MiuwVN1AFxamksqa0VJrhZtBQk9INOj+i6
ZqAmGS40aMMioDkLuj5//ld0wmJNjmquVDjCp4IpHIAyjnFi6MK6DB8y0k+9xd4z
T6WoK/0I7Xo3FQu20BJb1UgiuTLdVsWAtK3l4kpZXd9kRXhvYJ1K9YvtQkaWQ8D+
AMb6kgZ67ySS/rzClSS0Ri137wiss+K/AnVd9XIeq2S96t08d9DHb+lSJQeEa8gb
Gg8uVFD2x6+Y+F7qvEsFT+PSDlzVD9QlweCJ4jwXlyt/Nuys0Sl8E5ycLSBol8XH
g/SOYYo1ZDc2NAmHmUi03Q7Gd3Yh6Epx8nKJwzcIyJPeLCk5foxes+u2PCeOqGcd
daFMikXlG+X4mNehMkISFx7MRrM9FRR3E0MVOwLwN5h2Az+JBz27BHrhUacFsm14
gHtqJl3RTtwmn715LkN5aDEHzzc2OAVgn0J8oUce6/KEog4Dd1+3FnNwlrz+UzDn
qAXsMH9Hsln150sF1RZIkpvUkHPxaCvJ5HwCcBOfLU+goykqfXh2ubZi+PONKwLz
g96XsU26KKklLR8zWzkrP7MeGmAsG8+WGIYlB+u+27YFUQq6wVhtGJi/nuyXkj3m
q5UCjn9D2/Ukf/s99B7mB/MDBJKOFPC36ui8cmerzrnI/Lao1WA5pVxl1Op2/VvS
wEIizzyuva1zSCzueiqmUO8kVsUQOLly/eRWa8A3mfmUZHs+izze4Nt0wrHZw1TK
JG3jxdiYWbHU52Xo7hKRjUWZCX7Z4ay7IQvP+3QylMzPhvRy7dfv5MW+Rf9q7efK
eJVCLOlPIw2lbwd8ATFxtqK642C2ao8kX1IxLDEVbc2Sd/0mmuIXzrWAtUdJUCZx
tUfj5bLUVSTCIUxumEi9blf1RPIQVV8WAyFv1EIJQrgq/LtSe11/9AARJeMXTwfT
14PK0zfs/9uODaiM7Nny2jWdlxL3ktiD2kBs4/IqPdD90Hgbc7+9JSrRNDglvwEQ
U449rC6uOd0gaehFywDO2u0HzH5mDX8RoqEH5FlZpVZsG5bhiNpIWCauhbfkNF+5
hClpv+fU5TGHQclWwRzRKfKDm6Gwc1Lmdr4l400/JUGXCs9VRBPwr/BKTL42jupJ
thRHxnq7jJ2HVEXbu1+WNAAmnaigQNBkdkoOgA2MggG1JRJnlNalU1lAkopCjbiX
QqzOoYdsXYDG5VefeoT3HynX5iPqFJQXrSIhiO/jPigYTmDA0rDHqc1TUXUAWzok
c4TVW9xTIdO/4ssVNPWTIkEIUZywRvcJGGQan6tSf+NjQIurlX70H5OOpKfLDp0e
SVj7FUzHIqNUerlRrrngR010vDA5l/lVKGbPqxy9bpUHFl33LGetEaZumKs7BtpN
yQQ4xltsEcOUWHb1/1rCdGUPvySM8odqkD026ECW1/RN+qn+LKOwzJim5bUUc9yQ
Woo08tvFczw5iAmvKEO1RUOvCOY7P+Pih1+YrefMb8ixoiP7mdanEbiNvZ+CyN0X
oXsClaE60iMZffjrcJQVAeeneKi7Yql3bqMy90B/oMrNwGlHkhZyt7djcQFA65X/
T1PuNBsRSh38kSXdWo807lErWFh+V3o/HMxQgOm8KkogE6ke1ygcwrfdVJzuW7ir
UmX/+Wn+VNhJ4JYlyycJL+tsd7eL9v1vUxoGUhlGiaEG+Ijk9pyodtL4sIc/rBW1
6dNMeuqtyuE0S5EEylp+QkLIc65zrj0mGzWV7UsOBWwE/9a9A3xrS7VaZ+809mUn
mmdH9wkNOsLQ5JZgdxErrCpd82IK0s6+pluk3WylPvjl2PnEJTpfOQuZsBu40bIt
R3RHPC03mDVjFCMiVQdLykz3nf1IeFFJq8Z4dGc1+xqjgW3yZvv35Tw5J1ryiD2W
ji09o7Y0lyml7lXNA7AiRJAr/3eEWYfANrRM1KChEi3tqZiQBZM0hZYvL9dtTprm
xzoSST0rfxiR/XMkqFu3YOynkCgZaMTv5bG6bRRD/KrXiea9pi56kciKyh3HKRrw
JDLjuW5SESUoPCIROxXgsQ4CmSwuADArt3Iz13VmxODCwhEf/lyG/tqVOXU6ZEuj
ywkGdj62yy32xwNQ0zSY6DN+8qg6ffQ6+FE16vZ9XiV9V4b/zu5iON6EpoDYBxnu
fQTfdTJXm9AAkMjcm3A1H7SA4uWW9P+LIftZ8wJx3h3O8IEAi9drna/TA+8SL7Eb
Qq5cwJdyxpG84yfx2pZg3FNVM6e2QN/5AHHfFtBNk0vXeODQtDsFS6Wj1OwLbzw5
21YYOcdUOLJGTrBPqNbre/92GUa/Lk0JeiGKsGuTILVb91IalHEZt0rrfvo28Tai
caj8QmoVFYVoff8H04R/ow4EyvjGIYv+LBWD/0d5YTnRyyBnl4lH1Scy1n9xTfWR
vZ99ZO3igpijAEvUcgkh+JpMJ5M8xfz2h1pndgJ0bjaZCrpyMrR7tEYPoC2IWXa6
j0MpV5h5WwZFzznUhxrS4kz0afsaBYd3QVZMrQZ3uTnoFgq4b5Gu6KbREaPjiRW+
SpbGhuQGnShxKqHzwty9gx6M4ljwxZMnFP+Z8zBfhGNxmsrETOZKrZKSlEk0EGJT
wK2YWq15Gd1IZgvJW8DnQj8ida0Q5lCHZMkAFej9Yoo74Ypst95bF3tlwPaG+0oV
kVKzJactz7FfeatEolrjvv6gf8dKUGAp4Jfk9QhqRhTwC+ferANJ1af4obImPQI3
82Y5isyfnoy393FsR2KA7+6c7uI7zTmS4miPVZyDtWsbKr99f3vIE5PtTmWeMxZu
PpvTY21d6Wf5/wBGzMU9bkMgxORIqP32GJ2q2QCccmPWxWinjT6Dm2sWTpBHg760
fiao80TXkqMmrXd4Km1CLlwFQCX1bHuK3TccmZf+IDArm4RCwmpWrHvbQA073Afq
BkcPlDTXNeSGsgoV5frMYLfTyWvtDSd8KTrKyySYt61p1ZkhtywgyGcMBehCpAdB
47Oxh4S3vUGoInsuLx7EUCDLbP5BW2+L7wKDQEJF+3tNL26mgkWOQEwK6Kk0P/Hx
Ck5v1vIAxbKBPLbEMHds5+MTc3yipt41Z6Zad3eAARRTORbLzwtuu0j7k6zn3MKR
dMlKh8Sb/4gD+XugqxFivHG521CTqmAVOajTB593txYT/hmogRTGAvDNN6358iNz
lgiWBgRDZ6bcxq0C3F9639BGxKcgKiWy1pT753cPRry4Y4uy799RiDcTM4IEkeZC
tnspUSvtWRDP77ZhC+JVzqgDSIqb5f8SNB0H4Qko8NZLYwuHXERq7PsqBlIjI8Pf
scw0Ah1oXe0Qt0pH9xjPty4E14H/NIAZ6RRw1n7f6nx0Cxk3zndO7YTL+C1nt3wv
vQ7IfkQBDeJDBZLd2sWaNXfMyJT4IWglKTZ+Bh2EYsfMTr3Q9F7mSa2A30Y6MLZi
lGLLaPp70Gpv6VgQgfFMnDgrkTr5nqCn7R33HQvwzT3ulSjEjjmTN70LMv4ik3SQ
q6dhMMGWzXh+FF9G6ClkxrSIqo3aBjyriqKPK73zEM53H1uHoygFp7VazNT3igM5
WteQpqlxZG9cXZBSKj4R9cNeP8slot5wvjdaHfu/YU0HeG67RovvKiTc2EBcenNW
uwPz6F1iGGI4vOPkjnQBf50bNQ8rka5obhqiIDCh1E+VusqXuizX4FwRaCOuk2Rd
Mp//fN0ITGkynF8j/npqTNVz7mX2t5qbQB835Amtb0LaXPsiwWGt0u2sc7WIVh+H
ZMH/+lT1kS5Jq9YIkf+5El0DhUBC5S8Q5fJdy4eUT1hhvjiBysPzr2f7i/VYsRK+
2gFcXp3ficyVVxhpC4lo7iMix/rX9kix9aiS+HXlk4RLLywIkS0gVqSLFV0HoBIc
n9ynNWXz0STL25fw14Q8i+hbGhRwo9jVmqEV8iRpULqpoTFkg2rkXWPgf8IWAMUZ
0is9mVsdhWyaWSOceseycW5mbTUOiDJY912FUvPsAZPDwRt2q7Yb3sSiDbiF32UC
C8AHzJoHyEA3aX4YOxxxpxlxXliCep9vyLdqdS4BH4b3Q9tGjJYA7kl+FeZA1HHZ
z/rp7uXY+nj14JIhTOWNmx/8wY5mdA6fqz4vdmTk10+NTggYFbtRFBsXshPOkxNT
dBt/VKIoB8r+pccNDjWVGjMaM6cTa8Y4A3aRU8JVksuRoKvKEybZKMSV9FN/xY8k
4fJDp0YxsyX4JqHXyaF8gLtKw6wDOun/p5FQ0iFZtwf1ST/5WCE0hmxWBzCF4ko3
mw76yoW0EsFZgsHdMd9Cuw+ffBNLiVSoxQwp+viDJIB37uqq5MglMf6a5JfI4yGO
ax78U2csOioHkFbg7DLtHu6e4G5duJ8ypq8+lzRQvlXgMT3uOjWKU4AgcbMqejXq
sBwhJRdiuUIYpgG1KZ14maMl/TTA8e2w2du6p0UEpRV4gi6YCSQXtPOx/Mfz0h/X
bL2kPH5X9Rp4kHqqh+F6FlAk+pwFjHbAul8u9T0H4H90DGhXaNb88Zp7oUhK9Cpd
TV42+Jg8LfRTMwcYO4oBbWALc7PRljnSTH5x/QJ5FXTWtR+/JhsrHQtnZqFA9DSb
hD8em6Du3tTQUe3dHnjegSe8irGe6hixJ/Jc+LV8cF2AkivgqTRUFptFzYpxxYjb
eKW0BOVWwELIQcl5vrrTsCwDntIh+yPvIu4oV0EWo+JvDwuP30E6R/ZhTF/Y7Gud
4G6s9CZZmnivKBomINF7h5MLzv+wKpc/QraGtvY5Qjt5EFodzXVLEvE5Ev15XjIO
3aTVeX3lMVSZJ7PqSeRl6goN9BFTsmGX+0Kr4LPIo6AVR8PXVWYCxYOAstwXUVTs
QXI6YkWg4tRo36dUshNN0mG83uMiwD04EBj+gXKBQrvxf48m+ZpWdmrhbsMlGGWG
wG/3w6xBSb1476O8r5BmQqCTOVO+pLULtF7DUn4D434BFqHbPoclSiz9DOVzhh9F
j4TuhwMpGgRqujbd3gHEqCcR9eKNBjeJc/hk9mYrzsbx6WbDGn6fU2uuDFUyamqr
THiUNcBi5PdcKqgsoT+vg1D5gOLtVcxMSCBermjdxYtZ1BN4IlYxw7a1lVAXnoA+
zmsqwYBwWR9C/RUPCA5rHA43QCaJJCdY8lsuc3eD0y0eYxWSlpS5Qh/4eFxb/hQM
EU8RFmO0GN1xjgFW/RaWuUaK9nx93Y/x0UyhFAK9HpXdONKOg2wpla7k4A5TFUSE
w9KSJu5j/1BYMhjiayyGDSvEm3kt42s7+95rtDJjvvLx8GRK/6qqwXexakjsF/b6
ZwXNtl6wnuxvdEf011TOuoVsmdw1rdOpC+B0thazKSfZp9kyoldot0ZWuAYbGAOu
Li+1TV5i1TfGS4x95C93egMOwDJk9sqgEfhlH7hX2da+YIhFTFRI6UYVDyGJZWm+
TAG7wRvaw7ED+MfgJOhSrG/wAlU3FTwmrLeIQ69h3a5H97nAlVUmKFqUNQGRWjXt
IkKPQ/Xl4O3kgSHHbd8WKQ2R2OIacTA4RJHaSmOm8Rjl1e5Ybp+cMC0MhV+UVBEC
+KVimknQPsYBz/Wc1rCAiHZxNOPowsR7xqPGzPD91q35kyU9rCqR2QUxf0+/Ot5W
aJMbHiMVegSK8X7afFWzCVQkZAgJzEx9At2RRl3/WDrdJTpJ7YSQtjJWNF7b7vJD
Cm3bqdZIROhTwSohRb7ToemxSOrz+q/3YsAMb0SIFkMdHMdY/cgFGoeMa8NADWsy
DWxSZwh6YH0nVRdH92Y9eZ5Vys1vXrrz8/nlpfmVbemRxSwbDqeTt3nYX5v7XZku
72mFw/seH5C02mL0rTTCCIzcmXeoJd4tVWopTJqkbb/TKTPuXA2TMu5FuuY4wjPn
zKfQB46WYOTRMLtw/aNcBsvQ94P2iKcv2K3Dt6+5yobVsDYsZfQvB7k4/0qsJcRz
94VQHWk58GySCXxsyrpmv71wt5s+IJWZuTG+LeT4+ygvcfgqySYUrjvmrLVDmnyV
DTJaoOGaqU13fs8of1qANfzWRe9h0gbNOb8WmSo8z/lsj62/e+1YY4/iqEcK0hE3
OExW9QQBq0QojQ3E2qtRX8iXzxI4dhhUrLq3JZb7mN8W3mKZwWGDeOrTwvsSBdcT
BLoPyXx3SO4gTOcg8nlxkAgdQjReCHfBwgD++uApfzNpzgrSfVXqyX36+ICwNZZh
skb1Ov6iztsAvzdPQOaPIi0YWXl1S+YmNCXimlvXL/Ms+mTORbJ+Tx7Y6G2bNptd
mzY/15f1dZbMk+fMTGMU7CxTFWSDEL+l23ktRZClPcuTyPMlCdVMJWbooIb6kqay
WGCdRrsR5t1R/UNwBEkrHmHtQhWYIwwcEnO2g2xWrGm01dk+FwKb8FwcohQj1lWy
iUZr0eCP8J6Wiht7k10hxRFo80Prg5i5/alT+Iqbx6wh+LEX0opWWIwnpkel3/0L
U41WSqStp/ce6TrmSr5xH4QjXDJ9vXb78H0Lg/uNtnfcC/0YSJUh031lDWcl2NN2
U654nvwojgmS7DpF1lIUKK6n/4WxOUu18xKiXCvBqJAFhgneuJy57K+RufTQs5be
ZC3hL/TGsqnuaCWQreDedW4U5l/l92aBLItLTBeKwl53IYmcDsKiECuodct9RQGA
RbPepkV0Kmc9I6+BJFwPi8Z+8Yyhsq4dvBSTRXZRZGbgQh2TUw4pyw1BfuFlbyF1
d6JwLWnv/h8WTIUQ9WtgW1yp+lN3EThrcO/m21hWGu11IBri5qnvxb6d1C1QpV+m
zdHiBZ5xX7Y5FDbgDRozwsqXuDybVPZDzUTqaNpv47Ig/cEBbgEPpmQ/Ns+UGTJP
nc1hl4LzR2Br1LaZFXZoBtVc62wYoM1grz33CAhHhM7skTvIrxVEh6022zuYA7H2
OIz4VBeoYq6mNxy8voLUYQCCukGTabIicYFq9WHG5Ls8GtjTIJaCoyda5x8eSl5l
l4vma0tQoI9F+xmxSPZdE3gDy3Akn2Zmsh92Gt/BLG7kSMUcNOG3CUALOkOfC7oX
+uam3bu58nlRlSi6D/4r0XpbUt2Fx0bwOrfleDQlNRy5gtub9m010Ztf+TqgnhMs
bI+01PswRMrJCWKRa+RPngXW1ambAozXa6ZQl/Vg6bcmW/x8pENsiMIUcJNTI7GT
AKJi2b8SINz7N9+c2EtNqYEyvv0IJqr8Y3slwHT6A24yNTf7YpLMEI7MHXbORC7a
A5fjqiTxOd338b8MEi8xlYs/2hlfDJTKl37Ii7czhpezmVO40qurbjS239DeQ+bM
vzjJrQ18VJOsN54DoExQSe5n5ci+mVBLiTkZArrH9a/nGUYIgP07xpvzT3VVObOR
9gAIF+BMvkCMNUoSE83tPAfoBuunbic3iBPpkjl1zDD6zcjF8bRLapMpAz7X+P0/
dZaYyY5mPGFAju8R0D0u26uCctxCfTKQcWxL15EA2a2y5MvCgGbJ5iWzAlYDUWhS
jgBqTaJpFwOi5CVFfHi3DQ4StvK/Kr7xXwLBOlEiL+BJ34dr3Hj3/ODW7WqAlMgj
1CBSjiLLBq68xIXUusqvtTy5zZtLR/1pQQlR1N8oWrz9ggLLxyZ1KQveNqSQvaUt
cf7SAx/9rK4D1SU8COWCn+bFz0AGWWLnAcEU7OnrytVKL4e9nWLUssIUHENiuDeH
/3XfehNJXjy17wPGWm1sxYtBBJ3+z2e47jcvdCw1Cpg1NaKl1IukMiiCo3BuMNtB
0jC/XLQrp/hV8ZMQl0mWkPEd6y17gixGfQ/o4dZwP/+8AnbeY1e9dQFN0sQPB9sg
benqADu+nL/QrxTYtPVZ3slpeePNgJ1OcsyUjbEJZlILzdph2+cHp+GJAsscnH65
p0A3KHm/rV8ShXmhcZfwND0vzc6JOQ8sTcxD9eIR6QdUytxh2PSYohDhf4hgvfNl
WB09tR+gacCfwR0D0Tnv/rcvpruFRqOSJCiNK2sjoZjDCl2bVg2+g1ICFus1R3y6
IJLjNOuJOJ5ErVHRri4vvyFDU7pgOFZRNZiZEs//Do9RokTohtvshQOJjqHhZQwF
fjqLZHVnassP7w+IrvuMaBln29hW4UGXRvjnLJ/gHJhhIoy6mmsQBm7KQcdCz4Ri
16hO/glmthr5VTgU3C5ONj+YSKP4sd5y9FGqLwGmd96uEKe4ABZqYkEgGaQVNeXZ
glF+zpLS0q245NUPpe87Z9GB73WdzGYgWnEmJhQXCCzg3SN0EN9bHtH0NLsGYZbX
BlG+kDlh1FEqdG+pWS+JCdlz4z9EZqrC7aPDdAGcsSvvYrQX3b8PHj73oriEJ1Ot
vLharSUMPgcyr9R0FztfQAwtscmqYpEqkCdtcrhaGdtujON7l4IrGQPZIs2aNESa
7g17pl/sBPDaxpR7RD7J8grkfnhOMaA41ndA24TmOQ711j1JZX0NL3sIzpt517rd
KlVBsaS1/kkXu+K5umW0Kh4aDLli8Y7OR4G+vglcgWZW2CroTJjx7dJBs4aNpikX
QatsXIjaWAlY9vs9xHsN0ii/P8eTSaC0zWExfGLr/I88aO98G2WnHs7YhORIr5uc
K5cpqwFuDSPX54hVmle5gMU8d/73/xto1fpO5Gn8HarkgSlgu4oBFgIp5pRLU/xE
7PojumQ16Xtftw6uGfSxgA84HKDBAaSDJu8gI6FfFnuwS8DE59w3xFxCBWS03FEf
/PPt9unrHjz3PVmg997OcvEVhDZVTsIHuPoCgLR9JwtAYNXwtnNr42Jp93L+l5ic
1/7OLyBgXgofxOloCrLTWOh6+QVDZA292e7o9xeVpaYgb2ebhx3cXrpseCXYyuM6
e2AGbqKcxBS8x2kqWO1Ys88EVgoOOs3+jnvCI3Jehq/r41LCg/mwU4MnPVfNqVNH
M3kEIZUN69c8v0SyUG4WxM7uWf2D14gfZ/KCpywc/9z6fvQDSc6oSNRxYTxnlRJ0
S+CYKObm1Fn4JKrH0HmxSt4+016O1xScgVOUf0y1ynEUwek2v7hfbza/7m8U0ora
9IZwhzbrTbZBGe54T++APWLD4xvHpfEBFay6VyQyINfm+jJcgza+i0H7ig8E2OMs
VHqo6BRSng75+0V1vUp5HF+bDQe8myTUpnh+8FxGS5bWd7pKmtG7qzhwajm6uos4
uIZRwr+o7uP7wAMHi2gxfYOAwkTcMWAh0Ph68DS7mooU+mlwWeWY4IJXsm8nkjmU
EQJkZ5AgL/kbcDINDrPp7rLcPYbnlMxR3zg2tMDP3wVRrGOkZ9Y/J6mpM2DLbHP6
NrkZ8tzuGYVUGFO+LFBZmh1nqxHVL/cRTJmU0QrGMwY1Gk6pICy2ZsliJkQ3glAi
AakqnPEq60AQht5fEKhRz+q/SWB6BVd+MM6eGHPqvzD2tpc/HmLmaL66PLvajGCl
IwfDP7ZCbx0ilcaHJgmzpt4V+9xvBPhkr0FufYxV9g0PM19ZWOfceKkJ7YD1oZSA
sMHNK5R11hJ9Riwnpu/tCihzoGlIgYNnEEEt1jV0Qd8IFpfYErc/1N8wV6lUs4qa
KE2kwWnQxsR3W3TohlzBVLlX2lnyysiE/7sfflhoJOh4NvpHzwUCTDjhiQiYYyPb
pqD00kPjJkJsW8e5pEbB3+mkDp7cS7G0FWV2t5UfCs2JZ6WjB5Xe2Iz66aqn0ZH3
7B9hv/vFVnn+r74vSjrKvz8gFArzm+VOLUU4XT9N6VvA6PMscF+yY8CvDN0xCtbr
AFaBvHF3+IfBI0Pupz3tgeSjW4rDcmxFp/7NSxmud2IWa9KpkDojfzIxwYMWdMEV
nT4aofitd7azrZ4Wfmc+0ZlMCKKA1h2hbgsWNecHBqZE1HXZGzNE0iRjlCtI0+Zw
Oe4S4dFmzZ3xIaMwtUey2Ei9MLhg3l+AJO3ciOFvXo2PKAh/DQjBaQZQ3xT608V7
FUzpCbpT8wnNunnAhMaU6gXvezR6xmp/pUC6aE4AbVVs5T9sxnZVbrQsPteGmIwz
oMlrYKJoyO4SN6GQkNTM0lzAwmplddBhaMYDipu+HphZ20B5WSO0yrehl2Nik4nV
m4Z5qxnqefadQUdTxjOqAgbwR39tp6GMbIO913B/REb7+18XD8ForCE2/XDvu1Yh
wAW6usHs9fNB3Qz2T8pA83MYv0/samobYykLxCpQrlv8XpRtiF6Gve/7d6ZaYBuC
PobcFpPsJGdLCCz+1ufISp6osOdCg17vXeXh9Obo5iukVyZ/zjNxa75dCYaQOxHt
PTY9BTXsK1erVJd2E/RfrwBu+XuWVIhyOFKNRSP4jA04McOwmw4gDtuiGkeCjrND
Y+201foc3KcC03hdC5BboZyjrfmTUJs0ByDom559oThGPfc+rycmfge0QjoTt2LH
tp3nxOY23enIny9CQXU4zEKX8g6XZQzOHyk6TsEWHzlrKyBVA16uAy4D2H67pHNR
QGqD6EIhdvchfcgs2G7Pat9S75TKX5RkWEqkTJkV+jQhseCAV50eAWDdsd+ZgCwW
tGNVGc/wFJGPx1CNVyozpT1Z0NLHpauCl1YBJgMp8VXUmh860l5omm0FiA09E2lf
07We8c9PFBcki3LaurshDj7lIoU0NsOm4lnMpFwx8gF6Q0tAoGxgzmnrO4ruXYfv
3K5zUU9zd8kFDmHpMpOuuVvhszrR8qO4ehiZJyOCnjuenbxqMpeG6aCLmtF2fr04
NlsjC+5J9QdCQvfpfFxx8WJ+w9fOlcy+PxzzRgn08ZC52/3rb7s80bqPAd/Vp9n4
SMCMlRpFEAMjhhpkS6syoFvGgdtSlul4g4tjgpBPb7IDSbkV+UWgYe1QHxBFvoXo
XKZEFrdWLzl/TdnaqsnWJXSnmNYyARYFVh4arzO06QO+fBOEooUE/GTKtM+2HAof
licn5hfp2yVnZsXHTlHe/oZP0RAi4obaTg5w31lTY1zSBFMDufFliFsh9rp54up8
YPC4bjMkqi2En4S6NMb6Kz/IuGBx0W0PgmnbIqiemd+vKXz2Q+KPGSJJozZ/SXR8
DSFHHo7U/05l8n9/LLYK4B1Ue18GPmbKYQUDnNak68y5btOODB8kWGrKdnqE5+DX
KynmivqOMgajCZa7mdB3oJMHsvf7QWtQHyrslMOeAdo7JmnBD8X9bx9PYja80Pas
hqGq5wDZpGpgS/8EwIb29+V94PHlGEzWVRPkoFtiBY8aahjdYE5CidPW1YZgDozT
TvTMcgRaPY/GksfsbYBnHQKLZqW0ibpSrgXYbQITmdu1wloF/BZO0FsndPu3Q7ii
THijL8pjaNwAdwu9THcOgcbfyNXdWYiChT9fkN+BrKHHv2Wdi2tbAOgTmrMlm5hA
7ZQA0SaASkE2C4Q8cOpMOqJL+EZ+7HwlhlQECS0XStXIBi+sn7zcpbWQn8CI5PKr
hD+ZRVbuBuh4zvQ80FcRkBquIZV1xBqgA69lyTm0CKgxoGuG0OW8vPZYMBvGDwVy
6ds5ukDWeElMvLsiiQTvsGd7DdWUp/pur0kurORarUSsUfKF7spxdqmS7+5duqKU
0POoPGGg2ZYv0zvDfW1YTpMwsGp6Ep5QCX9i9k7qMI9KJsj2UD8F/QRyOdr2yWFN
X5w8GOHqoq96YHl/Kp6I5ATkrtWSC7NGbDHPtBi9KKuP6fwlAzQxvAihvoLCGxRf
uBNR+HLu6gxfgs/qmfGTHnld9xzhE+heLHZjYDyCRoycRG5BdDIilQjDP7gZ3olZ
80QRy1kncFox6DksxRKX56JjmTsl0mQi5P/xb8dlfMeLplvXPVxmKaPTasuP+JZc
FYrVtjUN05DzcDkDWNE+cZq/yKtcC7k76RaAkij1KaUQV5aL3wF5tqlR/hTygtPe
UDdrvqGW5lMeFATx11yCGxzs1UgydO192hNetws++NEHeoy5GlOqmMuLnwg28HE+
v/4wVnu4JzjupUet5NShVUbwqxJhnpGilC7Rny4/4pCSivBTBeAg/DSJhIrYhXq2
xn4aBCcqrlsnEGDuZks8ztqWRLVEH3lAvdPOor4iDCt6iPTTYHN4mr1dVEHs7Dgn
kTNolFmndJPNaq0U20JxDiEq99JgjnrBQr+Hv/4cM+GZN2LzwZARC32Q61Ie9nwJ
RPNni7YkNNANaoD7rsRUGR+MnOHY+AzpYIltnwBWGfH9aMQZ+53Q6VIJK/CDdbHx
Gr8wa00YBdLVeGI4SSNMuqt6xFTsiegW9qBrtd541qryLHBAXvYBBinQjxHOImDF
lMx0a762b04svm3flRsO4vMmm0i4bSIUxNF+6K+yhqETq3/U0DvGaLAmBuJmb6xc
pGJyxXlXmiyYCJf4lYiYJKVrOMxBOTo/MoV1pGbST7DJWt/QN2GiTLiAsvkKNGOS
VWXg7lFSS2cykZdSZLMIsLj7sEM9UbnqjecN1qRvFD7agepo5crSOryBTKBVNJ16
Tgub5I4gSTibaiUvH0IBjz5YS6h+Qgm1zk//7xslMylrgtu2lC35UdxEdRNSRHcL
3lu185LkZojNAJdMt0FjHsLjLEzJMzKOeBrgo1xTWNHCQIEkrk6spfv8DpWymZ8d
OkP/V0fX0aq6I0jhp8iRHCtErt+1bhcZ81w9x0flthwCjrdk4ksgJduGHyIaEmJZ
6/0e7F4psfNc0iuZcKrbp/P1SAKxkuINvfEZmjkvG6S6p3n3mE+SML3JAoH++8FL
bQOrmgs+ZhYfN0V5Aepc699h/HyAhj/Vm0pLA/Af42qx1H1fa3RV+BLKiJVuXecU
KhMZAdfnPl3NPvwgiz4diKfQ5QRkrC+BgodZ8RwHpkGgHGIAXTI9fDfLk14Rwtux
nVDwZlMo3O66gcsGptDMvsAJYv88zGPuBf12sbjB7q+UyQXSqUbU7Oj9d4lcjP37
SnX6WfslCiYzBBS0jUeIRmZLzHrlSxhnPPZ0okOo8tKidHtOoeut3DoSkmuo3ewz
nLOfOlyKT3xGl5aGIw3CyLcZhKqwgbpmKINxx+ASJA0K/qgGDlJXqMHDwKVyi2Sv
1wQXEttkOd0fQvWSDgbJKkEXo92pnzJwRm35RNvEnXUiVVD4d3W2nXyXTE/cqMUS
MCnmtvcCDYME9DwouZe4ms0mJ+zvPc5isr4wXg2lpDPul28ligqaq8c8QOvpXSdS
VB6WwrQEz2kvdIu1yUSdLFPnQimqCLEreV5Q+K+slx8OIdQCD6krhu/qGqb9NnH3
7TurSzMOTcDBYVIRojqu/L64RMCkdSJM3xqqz7S8JUd9PjzVGQlvZPCJfm+9CrBs
tCtaYSTgKoUPtts7ZEzetby45B3eADymMheCh3fNIHq/MVNruw03xQaUVj54SK/j
0XzeFyA2JI7B2emT3ZYzVj2NkkwT+rZ9eMiAJ7CyCITGGzR39DjgV0qPACvma1+j
hFDGgO6vO/EmL5AKlO+sAYtmsc6vHtPHyXoOZ92V39sVK1wXTQbYnNBCuFjJu7T5
EXDbz6nvVH8XqHbc85ZL9WePm9Lf+Rlru0d2AnCh1ic9iGRDiSXX0dZW/UrbmUFF
U+s/mUFeYjANm9NJR62tJFScBAVWoSOUXbk8Yb9M4qzUT1U/GdH1vByj05CWLyFd
SHfjmPJw8YRSI76MdFniC1Cc6ygRZ6mUro0itY9Q5kkYH6O+3sxp/+z2Vg8Q5xMD
nz3DH+oagTHO3l2AKsORwWsrRVwr/QNc/u0t11uDMN+vf0LzQTPlYMG7ngnkhG0p
mYB555CDy1b1CXQ+xL6ybQf/yEpDgNpb/bdnsWO+Mk4c+jJs+VVD0l7i4CBXSpTi
DN+3v+Imoyc52b6TPO+pTGxyYpWWUXlVujQp/KKNjG1TYT6sNqoRhhRu9xEHO+YE
eg5KIlSh8CLfmk3Ad1K5vJ/htlddI73+7IeWv3PrN+1P7EA5GQg/pUEP6DSMqih4
gXTqyZbjwIxdAK9fWuEqqbalHCJWgXHDotzufW5JK6jliMjlXhD98Wea+xKXyROw
Abx26rpM8WxFLZnbS8Og4GLmPdq8HYqBgzNrHD/h/9jEcSDr2aV949XdGrRLnszN
L41GZaMuNy+KJV53bmcENo5k/f+k+ofCOBgHkxEyYzmF0azjLTs49QlBrqGy1oyP
QQRSgtYp+k7f2Qau6Xabu9c3BxhaRyayrI+rAfzSnohE0VRYX/Q8luu7yI9GmI3R
0k+gNP8LOuY/YW7E9PC77z994nADeSqIY+VqTOwH5J+HMfQau4gVFv5fJVWZyvbm
Xap5agb2yzhakxB5aQ3qQ+XDwKvI42Sh2EQ8REjuK84Xh2XL90cvOGJ03+Ssib0H
YShZFtFPCO7F6PuOBagVl0BHjPAtptkg9IKPhtZERl4WXNB7JPQLDz1vFDtYkhNQ
PO6N19PoCTCxmfOXvLtb5pnW7mX/PKGng/GVo0+ajYNowbDUzZ7zPM+W/v047RDh
36M12Yj+5RA3GkVhivx5I2szzLxz1//Y6tgBbYzNek0/GkUjngigSs+I/36p5XTN
44rxKHwJaXlJYxEggnpYqLFXUNrlcduwT+V17v1E3zmfisfNVgeTV5grsb6+3bOv
z9VegR/yyeonr0XJ538OMKGz6VyBLV5js+B8/IuoprxY3virgTDkv6UPxz1amAGi
sFTTd/COhDZJ8O15AoTtv1j7YdOv8AZDmitX7fVgT7TzczHn76ezQfRPtY99BMFy
gqdDjEO6igZUeybfYwx21zHoQgc1kHB+abHgkUlNhgL2sG2iFCWSPeLCBY5rvyfq
2noO9cCt0a/rxYPBOqqonqyUIIWBQ5gnJQHQ9Alo+cYX7QqAOejqMkTB4tnyg4Fv
KZPJy6MZq4LHSWCbEoT4D5bkdQKomjLHg7cCItUHd0yUjsbmvtShFBG6U4+HWoa2
WwuKjJsw+/u03aCnkTnuzhuiz0hjSDFsx2sU07L4nkIAS12Shl33WpqR77wcZi+B
YkY2/7ThCCo0WUC21RNN5AAPf/ryfWgw1sPt5t/3ktH1iOj/0gN+4J9A0sl3cVPj
IuMPUCf1W9xvM6Lr8DgGMDYjv1yuqgw94z+fNmcRlhxCdCXFLcyW5xrz3mpMS5XD
03mtHiH6i8ctkhHMqP2XQctEOQoYHetV8ZplqTi9zX8yXoPmqqre5cN5edsOCEHM
G6cnc44P6lmMhve5SRT8YN0ZicRhuf/d29hgXI7WBr33ZmsJF0eqLcdeublz41Og
2kwWkF0RuQN7uhXiGXkH83V1A6AXhV2396F9BeDN/ZYFwE5xFS1NBbmv8HMbT2wr
3I8KhiTdvtI+T/Ng6f3qzpOoUZ3wiYKCHakGCwWsySihXk0SauL6WFwmeEFrJ2NO
yWbadn4d5mcOKmfTfSPMoj04NVlk9SqH0dj8pqVlcCeyVjpfAO6rD93juRBuC2bC
wlGv7TL307oHeh1FuDsIdSYGIXchXrBuDqeKKUBoXXCPCz++1FiyHcUQWZYmfijX
qhUY6+QR8o/Jr1FU6qUPDht31qRHlRrqmdbVTmAJappkdRtKFm0pa3rTVAmTbAt1
7K5q0S2qX93eIjNADvB1MOQX2c/kowq2jDlrCyIAYimfGN8it1iFtpnJyuO46cH7
NwFNGdPip9fQvulxNcf+4HfMRRojQpa1MSi9m0oXuRCVUPdrl4N3iZU/UTf0JbKj
oSMzgtOKXuTf5r2wlwPlclW3BJVwrZYhuhgEKakZNatarbx/0rFVZMEXp/gh+U7p
Yn3kcykwaPZUJxEBw99xAwq44ptwtrQG6XSBqJz449QWNl+MHkrpKkXKWQnWUAhL
ntXEP5ZbfLjGivIks9ycIxqNRf0/rfRoJwu7dWfostl4QzhBYCnIplpEIUOsDMJv
VS2GlQOZvbmuA/aINooTDLT6OJV5nMTUxUvoE+h8Er7CCFmNErG6EO2dJjQ/VAU1
xqIWSP0fRK4p7gWOJex5j6DXzXsrApqBJAjFfuRlVAPl9KyA0oej6GICfrl1cWjE
9hu85KCiBxXSTu51EdH0S5/WHjDGk9kVsi5xJ62WPcHLgs4X0d3qT1Dmq9TBvks0
Mhb+48ehVCPI0uV/Dv99zMww9FprMI331DemuPeuTc1+HJJmeir16kLz64CWAFxt
aCPil0zBZFmfaZgFo05YkXvK9bQimpu19adn+C0fclEivKdG5Tp2hpvRz3ruHnVP
vxJuGeNTDzHqZnYT64s3O+1B9WSd6A/8mLmYPizFrj1Jcqyf3GcJKYlBVlpESjlg
QOtfjTWuZK4PSvLuulspZzoOIrkF0DNE8gR19wgDGDkqghLSrwR8lzCshg7pSx7t
ONFVQVbA204e6aS3EwvmSj6u4dubpBgIxuNNfyG0gbKGHFL60UuM96nDYlNMbwn+
at0OZbRilhUVG8nuZyybhszDDyxJ4gDK1L9ERYDsrjcEiSXpD5PIFrh4JBCu+o0f
G/jeRZ3OL3dSluoDU+VyTnPe2zCVNumeRS63R652ZadhttczzDJBV111LVmdDy8U
t+GY7XCG60D4V793l+xvw7yx2nQUKgltdWGXrKuYbcG4ZZpLtcA3mJuwq8do/kq2
6UBoouzsRYLMiY0UJVQo32SYcCvcXpCXyrEfIg9nhL0q7LL79x4oQakp3s3+Fz1g
k1VUVoR/m3Mwgyzd0PKg+Et6amFPTzHfGIkdfzT9HY5X25a/noeqR/2rzaPHAoo/
Qjkb2VTQKcknKWkL1kjpS/o708SVj4fK5r26czbaoYdTdS9iLIfXX+GNA25KuDEr
sobZydfRIU0eVJphJH0Ngu9wb/3MlQUqn8AZZhqZP1jiyGXpyiXYfu2cl2MbnNYp
wwI0fZb+5kuBb61pziFq5gEZc3t6cuWPrw2z8GspRrtRTe4irQZs0VtTMhP7y5vk
V/DmynIkTVA31gjfeCoynhvAhGBRlltV+f0O0n4UBqvTMfzh3gXXDlSTy8PPqW+T
eRGsViKl0VPk1HoUHrMmCE1JHtoei3IT1bZrMgnqDLiGQTfWIsF4O570L/Jgs8mg
NOXaUx2r32jp93u56zZkH+4aY5eWZgFGBzMVl1CDXXy02dHvqxby5CuJzn9/OYcn
Y4/1emKRKtAJoRMnOacMv4P4VA32U+8l+wbIdYobIv4PSuKbQuxhdPPQDNE+YJpB
OsE4DJNATtJa0m6fPANHKs/zN3CNBzIxDs3aTH7H1evMLcRPZ6WUa7YnPioIwprT
bbns0zgf9tu0AKDB9fd7rQ8aOkjGc5snXlpCQ+0uP0AuqnFNYduErkF8qNx40KlU
bLgDE2ou/9RwuQSXjj1sdyMCIqJSDxcVfrq6h1anjQz83WlxwfROX4ncTky6EfeM
LRNS20l6xPy9N8GPMm8X2peS20ERUib8eKK8hhf9oF4hVf+NGSSEUTkTkD4P17PU
sRukZE5pQDHkad3N9QPKZVNbnlFQlvVi9/oRVvaBX/A4XHd7WdT4UzZeKYOh5MLM
hWgWol534SUcpBk0gBeYE/7yy9EfeyZTXakOt688k6tog2PplBjN8ox4a+WUXE4b
YLrsOx2R7fXVtFAFuYuYGRl1R5FRlQ4hfDUKkU5i42YSgTx5bXZq1DrBggm6olpE
LIMlH3Uof/tMknBIUdiEm8Yp3Tj0wUSCuSGVUOl92s6op1IMY8sbRlLDLejDUMxA
aG4mz5DQwbPbJktocazjxF9E6bbi7IT1e4zyx8svST4LoVNQkQsEYPZGo+2f1qil
DjcR/UgLk9Qz4N57Dt7UHfbRGNOXcJizrbzpsxHnEr6rNv0qLcb1B5ADEL978a/O
3CogLtL9FlgkVrDav1oSoauGh5fSs29OLN19ae0OgO5ixp/1M4ROFxGG3UDc3p0M
c549m8quR01OLbImWGObWbo6hZIyzjEQyMTCIUs/jstgXTOSPeSo2di0JQnXWJ67
PeATBehBsrS0YOKiOJOjKRhvH+dFbv8fRpOIzlB1EH158HIl6HU29zG5ZDozNrXL
kS18upiGiIMrNZqObamj92JSlQSZSNdfyuDA4QrAfhkkQIZYkquORYkO5q4V295d
d3dSypg9l2KmIBz6Zbt6UZF+947AXRQ4JEm20bJBrQHTp8WaEyMVfgYLqDCENO9p
PiDcwbclvrC9udVYrX1gl2xH6ppmBavZv0bRlx+4T4s/tJQrrqBDxn+xvLAR3cHj
k40JMgqsynMeTqvHss+b+VOQvJ7ioTtf+/BaeWxk2qr9OSYHq3vsMQGqVjBJJBR3
f37F/aDtZXjOf0SwIBVh7ArCWN6LAPS05eaQaWWHOmDzuKmzcmKq8oEUCyABMw1p
R41PA2EeGZGA7mqWxCB9h6j7X4akJVbv6UqW8dcSEUff1mfu8Vg8MUQ2C8cpl77X
mLyChrsv3AL3sd9q/tCoEFOtymMJk6pUYulqBtcymG3Dghw8gwGFBOLLR9xdpqb6
4/s9vPpxrram+EvTbXjK0Jdcepn+fxLs1qTNC24CkkDFq4CeCPmB6TL04MRm+NTZ
0y18baJNjNN2Cw86D8nb9E+x5oqOg1p+0opiQheUE0A=
`pragma protect end_protected
