`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rFrABrxN8WBODres9Ow7HUD84TPNxSj/lpFohf4OcByBOUAUiJBc3djTlrDAfZc8
qi4+5uEDF5g+ZQRn6ckJ+H2+J8jp3JuAYAeAzlMtobNe18XxdfEUi0dpomMLx98O
pr3JYNh9OEUCKT7Otx/YBDktKPPE6Z3/FaGdUX72O5Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3264)
gULuud89iWRLzHjoVZ02soEBf667L2/450+ZaWlE1mTLiDTItjDL8f6tltg3Qs4Z
4yINT7D8EJLBOTOM4zQ6kgw620pZU0J8jTeOdC0oLPqEqel09qRaPK8VR7xqy789
r130yWonm5wDIFpOOcxdPhjwrtCrm9d4CgtsiE/+5Z5vyvXh3z48KUKx2gpYhIfM
bkW1b3A2UbzT+NeIX4lJ7p5fKJ+tHcAHScuY2obLlvU99uNkWTcM1l12nT60YCVv
+ZW2VI/GfA8Lup+BlvnaO3c4oKQ3F5mgMngyXn/0dLeMTPZzbZg6L3k+OCewPeIJ
/hup5K7KOWpS1LbxE/lpMLLdOGi4QyjxcT1DaST5QHFHukD3+7ygQKTpxL3os6E8
1FddB/NliYDyFmjqXWc/Rkue69Q6ppRWFTnzilu6NE3Lq3f7PptWZkmglriTIYXC
VEhSd4AUzfPwJKf+IYIaukBaqFehTtQKKDWgZoTMPu3xSaje/YjJnp4maCJg1Z8i
v2Yh45nJTECwNLqDmBwnQzQ+gYPn4GlU8ovGYHPTqhkWhjyTzwXiH//OQ1upF+LK
nMyj/R5up3rt8fJSS+xV9I7foykOO9R2G2OIXAUxEyny3hi7pgYtmeweBRREN3FM
5H5oLnP1GmxVmKNP4spUQeTTBdgB04WErhyYVSiB8gy30j7j7HFWzGFtVhIh/MHT
zZd3KeCPtbVNxJAD9k594tvd9FNilx1qO8WV93inmvSzmaNLvxW4X1AuD/Z2kYlO
Wv3wP8raEOywVDRW22b7fbzqCVDe9N2q9OgI06yPpNAaryIlzVtkS/caqmpQhHhX
9f1bPi+Gz6WRbkQxmMaNgLgR1s/n8/Hv9vPMS7EvBZuw1xJEbxFHq2JvTI6cIrJU
juaSAMqqAg589KRooasSeHqhjE7PvOQYz6j+WsQSWnC+0azPIg0xrHIvz6kh+g9y
xGnynZmH1mNt05sl6/kRlKxM4DfHTdijDfqX7HD7AVG5B2xSiFZ6sI5amN0zNOoz
g8G5fZ8aE2BLJymmNZyzr7I0KeHHkN0qYHxQCECAa8G+vyCTW5pQ2NieI0MTt6D8
Cm3JBpNLvF89VFuIK/mscwlSw7sy6F08E0FaHhbSoqaIXbuvg/l8zV5zSlxBSWDk
rEk1dkYoNBajcqkUpXMJPz2gpw0r+5jGTZAdh/qDqlmz1TIOOl/lqYMjLZhuOnAD
GoHGe2zJDjilazVvkF9rvTHCcYWCKBF3s5u7mhS2Hmp1vuUvCpJd0vKmmUrvLUhz
GLC8klErJj4TY9dDdgLmSeQ2WhZJ6uvm2+5Dw/G8Im0VqTvBTi9dGtPHXYItjVCT
w7DXqlJXirwcSpNnRbhIa2WNcvpolbXwuhRmfG+xAH9qambXlO9ctmcUSN3lwImb
AAoNPBBIxeAzWC7BvYYzNQ4qdpu3LGhfvZV8wtKW27rRjMiJ8TO6z8FBtHsZGgi4
FjZ8oRYohj3laG+RMVMcREQmUqzAbwLKXAcOCqooLW3vmKLhnk/y2wTxao4Xuida
nQQYkarMleKGjvmsKE/3sQBOzZutY+NE1aAaG+bRPHvnAUiuYcLgns7jzBm4XuT/
hZKVDAWqE27QlEfsU0ZUCx/oCIekVa+TFNxJEVIsXpNzlheOF22mcHqzy3831lKF
tf+P7UCbXAl3Jch4tCATzAOQaUehKyuOp0xAAVUnq0zt6pDxnvlpDElhcMB5MtCj
vYivk+4lHVVqInzuZjNNQZ55giAYkZYWvckVfMZJICublHCPcrXUSilft2j7ozKE
dNSz99MKiuQmF3qnTUOZXtC92oGWasnI8oQU33ayaUnawwa1vgkBqeyI4Obef8Ap
Df36R7DWeJN5/N4p57H95NOpMtB8r0hZHexuCCa0s/tpFzgIcxiPPKu6qQLDNW/x
rRHVGrYEfvqPvhAyoZ4uCkPKwPU5BAGArWvH+I9e7jQCA47b10+jIOUE7nkTFK13
GOl4W8XiMeq4jK1TggYkOYoIZPaAsAUcAtIOP7FBpApPRaxz8cYtYera4nbOyaDZ
S+DIc7FXHG4SPjythZaXV41FLyFAdaXXu2YPEWx8Jvqx8wZm1s7Kip8wgqvwUXSn
HEpwN/wNuG/qMLDUOaOJ5apKU6TEA8/N+T2b4SNG9QBGKglgWLmqYgzGtN6FR8Ek
KjmC8seq/nUXJ93XKms31/FURdBorX0Z81biAFu7vfnhMuCCZffY9WqEsYwXVMdn
gJLwXEiY8AYYr01hfZP5fP/tS9hkatAYB/6vWdp6JK8L1C3aw9PEf0s7M29PY5aZ
YMRvNzXKbX6oQUBGcxOUDG9EjQtsprZE/k7v3UnNe6AmKSGetQJ2s+9R+Qizn4+r
avV6iKS6CrmXKylJfnE34XtzUHyI4Yqyv7jf+FERBZ+RTaX5I1//KDiZcHMDrR2N
OOUat0nvq0rWXZSCrn+mW3zY4EmOIHwwe2KRv2j63U5JY9W/ES+6PdTJ8AsbHRjx
OhHDGMBm35LmSLhE0w5ArF4hpsd6b7iTVbloWyY7JZ8/DKqzieyk1d6LxIOTZagA
TkmDrbIBzGL89bd9rWvnJcng/ePGxLD323PQ9qlhnVJedxVswHg8HEaNwogrlIWn
pO9M2DNO2ylNxGO/E8C7OgnjOP/4TuxOQA052UhOUa8q9eH7plF3cTXtrVcJihQW
9DrugtGOhiiSCUapPJbkcSGsx/fi9bkAS9l7KZ50+QFg47Nz2xGu7wtoNkwZMb9I
c7HzhWaOI+Ofb8Hap0XfnuwELeP/bewMM8gvqfYz3X31hir2KpV27HGjYsIG+ZZ9
lLItmODCx6IeKfLGg3QP5A0ZBiJH6nIjVnnvZ2NYnzo/24wKyM2RFYl9xFRQf7pB
X23wkDUoILuBMWf6WppiJZKe6fjTr533asyS7J9N/Lbi105SW78MT9ZYX4+m/PpY
TJ/H3uHSs8PvH3cEvtyKQodeMKXmYjmoptXrEDgqIXv2t42gy1rP72x7pwn+1P/T
R4T9k8V3vJMH+NVut4EZ1wG1Wu+rLAwwB0+FHKnR43hjmH4xjtF7ONJHkMI4Hs/A
pMpb3FaO+XNc/qu6+ftWbkLEKeGcWHMxcfyr7hO//Av2MZe/xY1MrVYNGiZL4ssc
4Jd/n2Jrxj1wZTuuTNbEwCVgUnjnxmzWd1LHNKBDVFOITeOKB3QI+M9tjjhG2OHN
Rt7qPeeVrVifWbOWSl+/AW0NfkG61Iskdz0Z5xYlVAIeqqoQdUHGAMElLu3/v7yz
Y7FF01+fqmMzG2Kdj7AOFiUtETs/F4soUN8iLLjGdRumhVluu6tO0DShmLKA2MhY
TMyWj6d1kG6sp+SWZj3s5fJhB29jEV0Uro7j8CExMGwch2xoHWWeiz23L19eITd1
qndpryPZogEef754zWitOu1IEoDusNarpSjJmP3r+V4X+pLDdt2id3bg20XY5Y0K
Oj+A+V/KeRrbeor11ijCX05u8hmXl+pxO5OOfBlyoYpp/q+7qp9DF4ZjRw8OpZh2
TOqch32R1JqvSznfjVaNvfqGpq9xVmlx5fMS7nNz1YDCNKnDfze4q4gxS1HVgX6J
8QcAM1/34w5b15qcdgmCnHkg3UAgOVX+izmz6pgh92ltu4g7Kfq79TMRbFK3XYkJ
2FzQDeogAqNTG3a/brbLcUyJECo71osRrNPC0oj7OHWdCpazW6T2YJDFs+6xeUOY
NVjgXZz61DTAvWooKCjvFFIC53yM2phV6ijKV/DyAg0zinZbHlSeGqNGsM0/Iexj
VFSeAQG0+3Y4AESgK2l4op733EjdjM5+KiVZYMg4Cx7gCdERik218KU+AQuQtpOM
XSbhJ5KtXhnBhf4PXxrAmA1G3R72Q4+fBHvimyJMn0/2/QpEi9XuHktaQ0efHzto
3qis85kPDedctv4BvxgP3w1yOq/OeK6t6fyj48TI2ZmBpawY9C8jg210LDzr17ZK
XrMs2nxAPb9HdqKkGUEG18a0Lf+nj+3kdd1VQgrU3vKr/zvJ4x4G/S0OlDM74nG5
W3YdQtKgK8erlepioW8a5p/ltpOYmnFSeR3SvKDrUS4/R953WfQhaf3xQr9cA4RG
sb9Hztiw7p9TdFw8CmZfouoPYdgm+prAaIRgXU0npVjOUoFe0CJyx576sfrO7V+u
nP/0RAPtTdXnAX8YP7KwTUi6jb2+6b2pkkdz52zPDmQvVhXVDn9CihQDt6CDvNTO
3Q2Xet8nuMxXFZClIK02whfFHUSEAQ5SQRxIP/c0kpb89o7WFIBiSIFWGZIM0ika
SsAwfiWaEsztBTK4SZmxpzOFqgXw7JKd6UqGzzXnWFN9jK34PQmxnQ6wTkDND1ll
`pragma protect end_protected
