`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H8cWVpGf32GDTCVhshrfIlxUhvJuRLEs35JTl8aNDKKyiAswJqeWdvQsetzpSq+A
10f4Ia0rB74nuVaF1HO5Q1ILCQCdhvhZoIN4OQhQAfOX+ASoJIZJnuJ4DtL8JO/K
0QeBPQydMVImJVFxcJjS3YWYsNecDVgkQxdOyQA58MU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15680)
tf+If/aHIBM5TwV9ilf5g724hy+18Hd7kMUq4pRkvC5/RfFYdqo7QZU6W03hYgnV
hay5SGPxRNfBnPAQev5Ng8GqL4bqunY+PEOKYbGvTaFfLO2mzFlA/4A4KSs1pCx8
5hMJBolZ+SV9bABE5tQhZGgbI38AfTxFTtadBt0Uf/4n2eRRXLjAXp9W0/8Wjofb
9drP358KV9n/5REG3MPpEz2FYlm7immLt1r/Tx0YM3gyJA1H7WHJswSq9pwdg3mJ
3DhCs+I7K7oSW1zl73pdRszCiKTylOJ7EdE8IL/yiv0X6qrv8dcYZ8Eib6RfMz6C
FrcAVByMQnUJ/zf5zKw7oL5gT6UgguDgq92eJSHRER2gzZEEaktJH+TfTRR8J/tC
NKDD/v1db8Q5JaMTu1PMc6tnJzoUY8D6O4Q/qGvQixGDhDUS3YCB4sD+Qlltj4Dk
31uklIGMWSr+ALGOCUFBdf4pUObCRwhVF/TBk04ATe6OydCdIWH5MnDehhjDg33M
hGAitINHpfDJtjWCfI5HEOzANxzhHUUC5nHOMIDg9sx2MpV/ci+kaJ6rOz4zLDUf
hHhlqvwZtZIKGb8/9K7CZ0S7iiSVoyG35/7Xpa6yfGAKBAtqhl2jbW4WJbIG2H6H
01+wJwsTO9ltlPF5nHa4WVHFbUs2XY0RBvoHqMg/lqQ21qOJjWsp31aAhcsGG+B1
MqNlIdHS3b8Hp7qbR5CYaxwQlqT5VckHF9DD22m0mDJaW7ylOr7O2YVhO9XyPGM4
PGt89wHQtRc4AePV7l5N+tBGNy6WokW9x/Wc6k9wHgOdiJT9gl+wDhnx2eTq2/sO
YnVZsuJFI1Gz+YLxDIm9f6p9D2QWrcTE7C4vTBQcD7w/OnnqEba322Sk5jJise44
79H8n5JJFLIvxsIaPdWRGw/Bnc+/MkX9uxCYEQZw1MGOf78wPQFY994etHqD2DhI
QUMLrG7tXX1eYRYojOXDeGhLdqlO9SDzZ/LDy5ElzRspFZ7xnJ/qKDQctlYjudLM
v383F9JjepUZN9G6uJVF2+2Xe9iHPff4xcv+Uw+p0nt5cS7KLfIWiJwksixqCwpC
SMvInpR9No6IMtoBqLLGB1PjgNAybn1in3r8H2fzmHx1xapvHeoubRYvyxeWE0B5
JHrxF70MqUrQH+1KDN0G7ScsWErXK7NDaYUzj1IbQR7lpshugd2mrIh/ua4O85zq
khgfB6kKJoGpMOZ+3r8K/7ItxXmltt6rog1VxZ6ITSgYkRB13zim6TPbmzYExTKU
GvObChOfa0K+vMu8M5S28bkpuxHDBUNQvmpXAWL14smIpPlIWNYmkYaHxHLHMG5e
+iHG0hXIaaf8Epipo0sVenUoKf8dJO/bodVjt6ECNcwQ/N/b/8IISmeRFuvOVrok
cvHTBclzfBb5BiAJR/Bt3guSJ0AMciOqa1FyAyxSPYS0hkkBvPFCxpX237uxAu+9
mGVmk7PZMMvwgTcWFyYFW8PuaxFAoTCmYhgciysrcyYEX+tMBrmmLI4j3IuLOzI6
gcZ5kNPpIix2cldy5jmKG+lDm0AutJcNQQVYRo5LQeblxFYjuPqQQc/7pz6h4ov+
Tzm9LTAWdDRHdecAOtdE5CmdWtDdnn3kIoJe6WOVtFeFCHNpXWF8pv0ppBQpyRDZ
ndriiPxbylH+BafKKVCdgdD/qW83J+MI0uIYy05T9RXwVruRPJPDwT8bQUfSfnSS
c+tf07TH9Iso3aqE8U/WURLCNwmajlzyKvU+Pbmuzkhh80bFzvIAHjvRwQRCnTOM
mQMxmkWoNkePbrQBtkHDC7I4Rl5TFWymhZMnzw+4XVDoRVMnAAn291DHlXdApHIA
jF9U7l80iNO3wkNmoEf+1T01MvTUR94cGjV1Cd460naUKf25HbOTrC/ayVfLDjDn
jufno7toaiJBloqD7C9D3KmmF9h5oiW3tAnO95npjXlOSXjhczAnuEsYsizgXQZd
ApUQZ3Rpevcfdy1TKNyjjNqw3WZAziLhQ4K9TH6soJDYuzB2AnpgmVCVaePbs4YL
IIASHMx8G44vvAQWQNIXUXLC+P3unX3jF0KOKmWrvVr+fsEyzK7VwWKfNGe9x5zl
VLAS7txrO8r7OKMKQwrrV6HISxGiZKUIepHzq5tvgUPAyLxiCnTz/FZHS2NMnpre
loXXRjDATqS9VxqfEjq3WHYzUrTmRcm+9FlYt0tAIxFyiZldm0cMxG5oQfuhvAff
exJ587HZJOipV+2xHS3rwQsixfAZLkJZEF3+J3yrA8Vsus+j6wzIcv13qs92Of7C
ikQ/RmBDRmKVaFhMCfFEqQqqkzXGIqp/0VFmJCcBC4NGnNLMvLt4zYbrJBIwT8gS
nbLB5OqIfO80cy9TQLYOfgaAwN/b4Cd9hdve/6eTPF8cHsYrFN476tWup9HxlZNf
8XyN1hm7UYv8m+qk93yJl360DUsLJtunlEK5mg+EiG0XKbepyp9nngvLZ6feU9bc
W46ESeKtWzEl3NrevDlxbnZqh9yGs2aizivp0u512nnTDR53d5yhd2OlmmvoWg8T
JQ62i4kxQ8N5uHYYZ8HToV6+VZ6GdDXbIfUgeIgOkyS3AGnOXLEk3DdqzluP8Cv0
Qqv52e4xjlF48Gh9OkpC1xTS6c3XosERPf1SLSNDxDekUwoJt37RdRYfq5sNZrtj
o/nEBgY3GZvj0HNPLVobZgvbVTDfJZpEIuO8OEOSrGGM4R1OSsbzYRPM1/mdoJnG
47Ahx8PPo2Gy1/GihlW8FX3MfGl8jISGzmrfESj+t9QUz7COEu1IaeQFlUmgkeJ7
UIRbEmdDD41RElLX9OCkhAm0sK49iciNHyKeh95O9vZKvH4u/yEsSY3omfCF9F7P
+Edgjy+ln1jvJUEO58cZ9TnaSSFHqqmdjoHSaSxEaoHEeUZ3bc9JHS/jKcHREay7
5JmBbffKHQgQHm3ecf38XBlrvcMOngfKu0IIvDuGYgbM01EgfV5UgDCaT8WCMGYt
l8DrY7JgHwGLsUAjagZzlm5oBhR26K0OygiuNDGMBMT0jLicwidx7KVnCQYX6O7H
1Zl782e1r6wlIp8jZj9O22Ia9bWq+OUVVbfaXOOi4pXmTGUndX3goh2N2tAUFP3c
KGaj077jeflTiRB+HHJKfnx1IUyyQoVR8mbngok7QO8LTGa0PfEaVZUv/UP65jnq
GDsNv9+Wo7zcQyPon7qpk0GooopS3aj5AvIawkUyTQPflNLG81d0Fl6jQ3zYOukS
4kpJuz3SEtUrLFVEt9qqD0KaeMYb01vwZZz10MAzbYkDdpdRYDfevXq0srX78pqW
Q5pT2Uhj1F2yLlGpR3X8pvPcK5MyXO/L9fIRZGcaUGy0C71dV/kwmd50lGj1qm2o
pDJgnoecDXj5gk0b7ib0Dn/Okc/k75XdlwnpR7pUV9hH8zkcfaAG1X5uZcvqcHRN
KUwd9ziolg3o8Dai0/tqRzagtPmJ40kxqrLu5J5WgXnPR7gj/671hdPJu59xVaQa
tgTVK63OUBd+Tzv4VTF5Y9Rb3oTW6GwY8nhfhwfqTjtln8BHvkyVX8A5nhtqcgFe
3Jq9zhLTPB+c/UmZd1WLlxVwlKJDOJgZ+5hRLLdtbYWMw1mZWyPGqwOOLyn/lVza
q4M763KBgBt9/oQQo5IwFoWmtA6TfvaaW6UHrTY0UZ3U3aUBE3oiby9HTDMjnXt7
TwF9UMv4Rn4L8y1od5MhRgaMGtMg2rP60OslRmDbFRg76Dbn5gqAv9KpXRDuLDhy
/rJYZoirQgMujpG8z7Z1hXI0h9VX6v1I0MZOkyOhKXfCto12s6m0S94E670VGN1m
4i+8I6R3hZ5U0s4ehuvbqSHbi0uMAzeThCfnnLYpqbRbAqKNnUXXWvpFQWczKBku
Xo02tyAyP9pL51vx6/NwLYqEJM32EBDKSMuXfEeoddoihyGIQVzZweTd4cLrDuQZ
57TZ8bB+2UMjLnPSoF3CU+8VHHN7qKGxpGaQZjYw291V9kqV36MHa55NNTvx9xbz
1ECT8kheEMWxb/dgxlCQB/VsXPVAvb11pkUoMUTZSrFg18WZ3VjWIq7CPauc9O2c
fbRIclK0uHaTpBaoqJfu2JjVxBSiC7tKFrvUx+BORu//RSuk8mj1q/jm4yYeOoWh
9Y/vn10GJM8HaAPAtrpqoCw+2PTeADue0cCrcniLxj4APkRYd+TYyolL2+wTJzhd
2dNo8/101QCqxa57jEBXb81r4aMW5EvfKaJyRUehRug4bBlutUQ8nhX4s/4m1IsO
ZeZl2fhcLTYGlFVQGNBz8W0t7pOU0f4u6xUV4LCHTaIi+3o+sni0NYfnQV7l57Pa
xBfx+TI6sJmeKljU37Xs7Cb24AaSlxkKQMRiWLqMHEPQ5puQWHTb2ikkPFRMKCiQ
+7y5Oq98eCQ7vSXpxlgmrdnd/JlF52O2EoMSOJL4noAIschm+hWYS2pTB6QgsoG2
HoDF61I0qbXwpqmYP2BNwFXl9jC412VeC6JPbja1ZdX+2k6ACtPPmijZcgKXIcPk
Zeb2J6XksnckiPY93oNVWljoer11CgU+Y+4vgJ4lwmZAK7IADrXTZFHE0bgVzfSn
fFQjOy09ggF3Z1lcbM0BxagqVcpKGx9nA7zazGOo7x+pxFHVNO1L+W50iijjAXMx
4QQASqoyiEj7Mr2V7fBMDXuMVbbbvyV9PFAiuyZhRx55hq7OLRebLTxiZHtm1Ve4
yiCPMqamumcUGoZo8urUeJuVbQTay9tapr1r7v0I9roOkCCqkS1mg6r9Jne9xLfW
PoWa8TwaGlhVEY9ethWzG4nAde//wwBu4ULqf3jkIwXzWZ4E2XbXBrxZyBUlgxrA
1Lt+KZCPTy6IOJ8n/YMCy9YR3aafjKWuUlW2QhYl1dslyMHOSdpx/61cYaNBGUvd
TxJiT+WoSi9TyR9m+OGrYtHJvOQNvqqtiUdSxPZVxH/VstUpIn2U7RyLlmP0kgbQ
Je19bjekQZrI4ggiuZX86TKGJUCL84byclq0wFQB2w15kWdtnZ5vj8NJJ7RxQRtn
5thZUJ3gCsBtbSFO5BBj0bERt7n9Djs0aZ5nkfGOQWQC0joAlbVRwFkpYjWhHrfY
8OIIl/CKWWiCoH6qpqNRBoBO4wzu/R7LG8IyzbXitADjiHGVaKjtzuwGweqcBdsA
mJHXZILGwOrkPJfZ4FR/hVyl6fnuYkmHKnqBvGV4MF7e98SudRfN0qWwpKk6498X
Sp8JwNQppNZy2TnXTF87J5306r4KCqfGlQ+Uu33mnL2QWjL6ulsNdZW8avr/nxPW
I9nItw6J2RjcD/tqpObWdkqNaW0K4p+n/Fo1/pQ7c5WaVQHZtJxL2LYjn1VYvhgD
LpEP6qjxp4ZXp0kNJSHK+3O2ggD/cWWbgBNfjexIx544uvj22/hUOQatSVC0T5Qq
naNk4sollwdoh7WRZhmrNHQxdg+n7TKO2RmKXQMdABctBswOARSdMM4xJ8ZfUxw6
toBp8Daxp/7AKlhEv8yNOuxmuHT5MCO3E8KmFQVkGucErP7qu/8phUxOdfiJbG8f
BhtsYEzCTyXgxNhBb+FIlcAdWeIOH15FRIXD025nVAVo4GJNRyQAOgVgon8lUhA1
S+Q7OqpJ2KGJLaYHl62bbuyX+GVLC5Mycq1feXrmq3EDaYrwOe7aCg7hgnjrXAiP
QCem3j941/R37L3uFy3AaVKuOQ2c8oQQlpA9SEE2vn1ZouqvdV14KRkLfs0npm8y
RVM4yEZRRgbzPLWCWUIEgTjX54kyOpvFZwg8IC0M8B7bTqqV7BIJWhBnIR+SqFJX
ruy+dWvusvCOoTmdGBo7AZ2rQJfIUGlxNSURqXERjkDb9L1aj9lYXsxavXWKodum
t3xkug/aEo56Fv8yMUqPVtvRkryXcQFGkXCgACD/PZJXXP52KnG8ynd+v1a9yQl+
rzh+3b2McaH7z27h+z4aCl3n/5mx9CfK5zcxr/t/5EOPYX1sv7s6bUfFuHG4+Zas
kw0cszFTguzOrEg6lG38jI6WgQWJ9erWyV+xv805rTUaaZVvy/rDKTWxrMD03MJ/
rYJnPYSmnZAsXNNUavTMVG4PLePmyWPYVqHORuD/rxW+G4oniKPPUfFKwiwI97B5
nBxJ7Tdwil5t/ul8qRIeNM6yAXH8eYPbVYvRnJ1GnC1/4y4xctSJMTjpavgK4V98
Dd5oJgJ5KxTR1qDl0gXrByCHehQ5uFza7Pim+IOVAwXZOT8wtNjIRlRnv5Wh1Rn/
J8D0k/R7tQTPUtvlwGUxlLb6KzxZAXXyFi5gb59FH9ZfzMWOUbWK9h7dAs9b0OJc
C6VkpVluPYUlVFO9UOwl6WFtYDlRhaagEnnI0hjsxOlO3pvsp5rpa+b+EmwJDUl2
EQKWtspObwQSsNW7cwNJGE7zE0VNxO6mYzsg7am24txIj6ytae+gYCkGjSokjzMK
0JdHdlZSXpx2F5JDzd44NmQrd8Xp7l+urn6BddIbYIB82kbV10T14mFcECTvhURl
/8SckPZ4qUWqIMQMVOXoXKHpOhjjP0PEzLqEoqeOAVzGbRxJun0LWZArqfTZdXSF
mWSPq8Ps3mJH3ePbdERci2ygjN4VfOYUtuZgSCjfgRjm7LhckXVp3OCRodf8XRqY
7uEIBzSII6oN4OYMglszCoWXQnOSa0tdzvtutr9SsmB1IS3tz/Nxb1trNH6U8fOn
QYfdiCgVzB+aqw3RCPvpDbKHUmNVhQIplQnMT+nEYv6csnJtudkR69KOKUH9/TSv
Ss3hpj6mf9wS78lL+zwa28iefmfV5ey2DDzmmw2/3LAXx71Ov6vZ5bz+JT5S3/P5
mdredaRVjEYtIy8ol1vQJVceSQdQO6ZvPqUrRoWq7VFtaKlTWCYcnNj34gV5KLKX
yUzC40lW6d+9itmJy4zBiGS9BVDg7lZPuornvcoMZrMgoHRTO5F5TazmNZtsJq30
xoeEAjTfBXdFMefSmROlxju0bFk8ER9/Nc5/hF9gwyk4/epCWFm1EHS3dJJC4o4R
LGgeYHwueN3PSbd5sMLHCP26MFy14+gF8SK9FFym0xXq1DJ1yMVkUjiIvSdtgc58
KRzRIrowZQY6jmgIk6n2H5Y1XdtEQzCZDRraOOgRpRAX79e1CdT74ovAi79EMADo
OBly1r1mVXITJxSz77y8Hxg+TvdZVYdUEZhHVmXII82P8yAGsI5g7GSCYlfAMnM7
KD3v2StzB/UHItTeyoctVyavRsved7Khyc0dcZKtFb+gGXJ1xkNVp6bSJYy6VwqN
CT64W1fVymQ8yNBB0TyWe9btweTTz0WqyI2v7PaVp2xVcIzD+BHRB8vUiinUo5Dt
UMZ1lEB9Cw0r5n8XdOZY008Mn3CQZD2682O2Fk/HEhbpVb0xUnhanfKnkDKRovKq
V4MFXsLNWtgeRKMhLgNxwmenaE7B9TV0xBHyxgzd5+jHYQHShmPkE99DBIyTwd7L
9phQ5rbqWkb/bF1JihfjIO+1ly62Dj5SLcb329nfKsy+4ggQbBgwEY3HrMM0dpFJ
N4vyzuwVzQjCIDQdoWAxwUpLDWd/NgK8E2VwRgXFdSoqIVG0WQc8dUteKxVcsebj
5CcltWJNZUiI0g0cR/sA1a2bduvata7JMyEJ+urQx9/qg48E0AcAOnmbaTKN4i14
xThZUkztMfr/Tl8ji0afMpxWVpYqpJsDMqjY6Wj0ANcNH9FHdQ2O6GIUkbo/tCj6
3e20/Kc5SScqaaY067xMIwQ+xaro8Km4zr0UeXWuDL+vbCEZ1bTEd8k64e17GY+B
wMYSVpGs37SPk7PxB4l9DEm6F/j2FRmXIfALFvSOYHWy0R8RY4KvynWFwiV4JtcI
CMiofH6p8qSxXVXbc+XPpql5JCJOWzMemH8vgCoT01n9p1H6EJaLM7UFyofrb7n1
QugPwhspDVajgEYU+yK6InJ/by17AROLwpq9//JUTe+slFqmrlU8CGikFzhXvxT7
uD7xPbpaCzrLShq66haWOfxZF8kbajhdZKpbLt88olGg5jmEmspxwZov2UpoZL8w
1WbRpakf7TCvyxp4+b70117XbHjgByJW/O3dubmVPzpKQCOGwv2CZmxRNvm/zxOE
sUwDFsQVs4KsHymSsmNs/tiq49jI5PiiLlldzN1nwGcPDy8KfnS95FS1iA0KTN7b
8nLhIclDuMqWSOfbVxydNRqRRI0Lwyp/WEj96aC7nS2IHc5YBIaA3aiWnTK2ms2R
MunICTPrII8wKE9AJ3avIVso2U9FwZK5koK8Ma478jzkIT0q1vJW/iruOjb3v3tq
PNnVSpap/D7+AtcWwuBGbHoePwfxzQUB8OIDaFdLwEtsRgOU56QXbPLec2WcvknC
lULjtg2vawzrhZrgZ4SobWpz+el7w7XCaoC1rTQlSs/JaaLGsM6dC7Syr9KQ9doN
flHYEfm3PXQuECjKsx0VfNBqwPBTBovwuyyJe76vsMtUiMb0DIA+VjvC1dr9WCtK
O/M/TOXfsiX/9DdT7w8inHs27PhCpo1mSOeX2hFzEs3BrEeZaWULeJTGRPYmSrFy
IZU9bwnGrmRHw44JRFN+Sca1Ejy8qRbU/KxZWTH7nOKu8DK2ItlbcQ6tSBompDOk
qiPlu6ttIro5aKYFq+eXLUXAlYirSMhjYl8qF3LsN0W6WIsVp0LnUrfVfE0IK2OT
h8FHAr5WDNpl/nPKni8ozciypEsN/jU8Q26TBvg5AfgQam4oDqsyXOrOdHDYBvYo
Y7wd+xO/nWmq2vjRx4zKp2h9suGbvTL9aOCsscQw9i+VD8Y1saXo7k/9yt5Bd6pc
FZty8dEoS3SVWDfZO/ItCcwWlQfouo+nTX5tiliuRWLKQ5cvhtJ49IFzxDxErfJN
pO8jaHhUFD8pCU9gUScoMUAy2toSMZv1Yz9tH8LDOPioa99PvJYiUqvQ+BFUtR90
5tcSHekKoWrgAE5jwSFSXfe5pwyhSQ0vkg6cGh8s8qwi5AR4lPgemv0Qlt+2SUyl
GDAFwjzX2KmW0lHpg340RAnii1s2ClcC9ELZ5iUHExP+l0qzqa88KCj9qhifCVZw
d9Ibu3pZQBY5TUlZkwXtxhk7DMotq7LzxrJDPuowDH6Ju7CcgUKUa/tRFUfStyZI
T8STvbhB0VLN55NwJC+9sUELv4HZqSGqVjhkwld9Xer4VsUNbSAAyVwKhK5Myzrz
OOn7amSCih7qYkGZqbLq0RQk6qq9Mlf2CFo6xTXRQsywqmh8mgKwZulk342u1gtX
2Ptszrg7i7Ga8NjtICbrTIa4uuPyusK+LhRzHoaj+7juPpmQEnIvXhjFDFUdNcY1
oeQfTNJKOiy+u3tSKNG28khrJUlvwkAkHl2PulNfZdx1TAIJh75Em8RtsSWVb+2k
EHfr2DOnTHcNIskXIcIyL112esXSW8Rb52diwBEdwr29WKqwz1EWbIkmduR4Q86j
bU7BL+bK8LGGG7hO9MSez4ir6o7GFF/6swUrPIEhsZL782sxbHymj9xZipf5B4zg
w7WHgd2aMuawnIA7Dm3jEyA+HNU8nIapgWGWVFh+sqLHfao+FtRy3+rvWBFQ6mke
W/yRXULBufmV+mYaoBtepuWdh0WtwcwPE6GihruM9DaoV+FNIrGSNp9dj3UbYM1H
DL8RjBUwF/IBpnlb4DpC5bckb/1lMScSW+rcTASO7dIWoHUVzn6dgZu+lUFnuHzb
Ek14ktlpAt7U1kyt0BlBWUv+yIDNVfIjbLKUthkESEdDMTX22T44N88YoaeuxTfR
zBWAVoHCemyjy1ThzMpLJgLPQZ1sc6fh0wzZskStqq/CzFvWALSRfi2GpRTwsGWb
YodERUyAqyIwqnBTb9FYrVQIY6FLBTNQ7zEE9BdOPv8OoLj+6izTVSr/oGnH27AS
IMA1aQQq15q40i6Hpc4J58LIYfHDrcaChk7dklucpwsGUKaW0hHvm7mFGdhwfOpw
JWUNGm2X+8BURQHR8W9BMMeORAwSa02TmxYHIKsA3f3wKvg5j7ihMHFfUQUsM7Uw
PIumc35jKOLD+yAlN6rnqcjMQ/aH15brE5UBrYrHIYL5nmtag8QqlV5zhDv3y/Bq
ADalPE6u/r6yu5QkgrgPmM1qfgvg1j7rpWI2x0QirSjnFHsNvmDtaLfBGKaphkac
zOC4nYuRwoJkb1qa+50fofE0asxjed+U86vSlMEJvneTSMaznuWCf4bMoHim9TaD
ZUGVOLciLbeHBAbZz/8cvp99OvIZLlMDkVWt+dhdcQgEUxxtH4VQlKHB5XT1l+un
ERaepHyca+NIifVAnogyo8qX3gUbm3QL/Gz4qtozwrrkgUCs2BTlXz416eKWX6iz
zt893x1kF2TN3FbB6YKCAvQ7KrbpbWgNmvSk3fApvT4tKBkyPd3xEC5L4JrHA2Ux
arB2yr/pgzD/142YtX9uY5fFi1ssbUDGKQl7Z9Ntwk4TTxya4nM77t74GrdWlW+G
vZIJr35JPScmmkr6ycZGBg3u7wCQSbEy34noJmAIGpbVrJas4ZK9u747+aolCkyh
Rw7yBbjJYG+qMgGq5WI8zCdC08+hZS9XTjX3KoWg5x3VI9ZMwaC7dkvIWuqbg1jV
ETNYRi2J4wFEQoOBTAjKAK8CMjqE+u45ehia3OW0HhPWdcsN0aTZRxF0na3B1VRr
vmorrfASFNs3rZF/v/AMBHlo/dPBwO81P2Qx8RFUehImNrHNmPD8KzicCN/L0YDb
CdgDEg5cbOdLSj2VESv8zloRw10bPZrikTOFwKKFQ7++2nkCYrf93otgPzpUBQhL
Y1OGHi0+eMOBhCt42Mg0pLkLtjOR3indLdfB6ncwSh2XlvFUp7rNWHlrw1KGdt5q
y3tgCP67C6j0og/WaccdqXRIPu6/YJmOiINdl7wJMlQr+sclCD5G7zJYJo9a3vgn
12+24TnzdBScKNMv9ueb7skXsda4MFq35AVR/R6TGcE2+822zHT7/ol6b8oBIAJF
dJRaVA/aTb4GrR/69e9En0QxUw2yV9vd66ZzGpljQagJTRlrgcbKL7qui7usjjtJ
qNARHqJCb2h0XTUuFP5nlkDxSm20Se0PyzYECBFAJZnhqO8ckD3XyIeNNF3/kQdU
nAL0b5A5VgV+wDdg18HI/EgauZeW3gssIHRQYRUN+LrRZPFQ+x5ydMtyGR4h2WbN
o72d3UXs5PNRVzN0JBehohWaFdVwXWBt1R0fsiV6G3BDLToJQLT+fpd/GTTX/4SN
NGl3cU5YycZYUQTw8pdEVyWVVrLP25g5e5GzVdYL4GrE74YdqAO9iflN2RRVwN7H
PsDaGkD9im3GSeq18kpMKpKWWi5nwPlrqY5i7QqAJvNqTTJAiJsZaD9oXs/9eiS4
6Qj3bLkWkuWEQAmlkHRr+1gZrOxoUX3SyIAIv3/jhioXn8FXGQ38ICMUH2yMxGzt
saIF0xQp4SE/0//JDaDceU5YUPwwDqx7i0TyT+R/d2jK8qOJ/OvpxlhMTFBOhYl1
d9HyA1PipCNVmGUg3h+mPylZI/v+aTavLh4AxX6iw1ty6za8zFMqL0DU531rG23V
H5ZfcyopjJCCcjUTOc/U9VtbXEucIleJ6LCcoSVJ4OtC+GLyA6lC/cyAm00773VN
a0c886yqsqoORe9wDg3AfjVAKFCBJu2YBdX4koYB1W2f28y72lTLbtWCYvz8yqTq
dD4q0xC0SgvTJ5rRFFLcS1WPDjAvgU/bH1vhghEGXwL9x+NOCB5nOuWPV0pROtMQ
CuSCYpcYyBBDlX6K1pG8LqG77ye7xyfy+bkXeh0ymjF86RLpQr07VtVjVkwuSPOw
ISG8XWGohQR5HQdR4tr/da9neSKprOiegyW00zB9nYzHL3g5w/ox2ks8JDFCaqHQ
PU7OlUQ3MBx6vgUS7agdP2NBffbJNqVPCfdFTo21giYU1xegbS4iyr+zjTEq6Gwh
nOWfJ9P7086kn9TMqYfnbyGt+ggl7XNDdQC233efa4xd1ebRzsMnr3yrEtbTOl3V
PfDb3l+AouQcZ007NvA3kkGsggZ8SSzmJC5NQXZQK28NdEmaG9JMxUNFKd0vcNjK
y1HfwG7xz/1tNR9qM6r44ll2X4RkuG4lIyzEzOi29m1t4otkQrncKiT8Qor1Ajdn
zUfYqAdZ7/cyDuyzikYA+BF1UAwcDrS//ZpPLFBkOhcOC5fA2BnpGM6jG+nlB/UU
ivGSIW/Sabh4XpDhQUNGlqBJwFW0b+ndM6/4CHZIdwIeErrunhMIa6y/kOCh9jRU
uDYa7eq1vMCzz+rjtfiVNQsXz2DYMgq3sIkHLLHmXXfFHv0DGX/vrZq7FnySxAps
i7+evqu9448S5fX6vEmQ/OoJkO6BtT5579rfu/+DIeLpYVf+FM/th3TibjFDF2r4
T7LYU/NwKnAHT+6OaVNBBUt8H5Dns1mKe19F/e0kg/KqY84mYU31gdTASYrGfvgC
Tj0hSOI0vx/RvdYrGTwMWiclFUa665ENC3qIBYxAE4g0LCgSD15J0p3R/6YtdTLX
ae7pdd7gajnBqWiQPZZdNwluHt3fOMZb6g8HxH3CPCtBYryuewK+JZRulTeFpjTw
e8bzhsWIcqMDQRofQ+lCOxZs4H91i3bCuJFfEVB3jOmIlTPQLXzpShElUz0ffjNr
zAmaf2t3RbX3yXTBcpxnSOBdOJTPfVCVZFfWHOFpQ8bZRp94l6QToJmRGiSGc+gk
Hwb1v5MRTnUF7WQM76LjSQ3GtCATQMYsLETyPrKmxlXhJNPrJbdCpdCK+7v71C5v
f/TW5KBSYw3dOfG4utZxERCOWO/UWZR93oCzPRFmsBFWTvpj8tj2O+TOHXlVxfEt
NKRsbSGbvw57Hl2fwr9YjQGt0+HiXsu7Px0xeMv/EhCqCOFpjJK3icjQFsjpK/KA
QXhkwDu2D0xx2yOz5NNlcWpgfk2c+oTP0kNhek5Ju6KgvWskswhVjlTLAGLiMB4M
E+qf3f1i8tU6XsvfFGR8pMQVHYR0JSdc+dzEVFxX+bh1EJCa5WYGDEG5LeedGaw7
ujuyblP8gV3ZsOc0lu8ZytI017HjWjrMg9QbkHhRihsOYZlA265IYTe63FlmlI5H
OItanjHM1SSprv00OX7n+/cBNcU6DY4oGy1BVHaXC+huazzIlL9KbKNXmh1y0tav
mRvE2ghPpQFct/ZUj8ssGPT4tUnh2UpThyE1HzHtriLb/+Iceg50obbmoLUzVhFL
0sU9p/xVrkj8uBB3EJUNZEh6eO/fLqNxZ5flbkzPPYInOcWGJZnsUp7lKJ+8kHzd
NIKm03hQ1Va14O+/OyPpatN+76aEVxVPmjFkkQPmpPetx74uFx0NZlnEZMbK26k3
oaJyAv+egpRuYdblI7xn+ZreQdYBy25A5e7GkV5WmdU67XZDZoGMN5ar3yolFbw7
S/W/FLm5xdmAe1W5kykcfu1jhIT7m6FxMoGP4VGan+fHaWeCfBS9IF4YeZJk/EMt
6Pkdu7x0NZTf2nzovekn3efY7uTpA5qQB2YWHk4E3MKesLlKTjNpQkMw2jHcrj2P
othWOnchhFJVsSFAtHqulN6o1Sp0EgA+tnEzeNMnIsddTrQe3IEfbjVZXjDM73uq
z8WLVL1YDUNw0JeYvt5sUW7inaZTl542TgrGGuKZAs8USMZudfPuy0nG4VXYdYje
pNin3Qn2pdx8yFbDteDHBWhsTrBSbGjovOuZXu6ZzblU5+6yBoert2dOmaUR18hn
ccgsz7xD2/CGdnyFQxXulGw3Pv1kbsF9FraficQxRq2PznpORJiIF2vImB/dSGy4
Pme6ds2KJNpkr/EnnpbvsM3PS/RMbgrzEQJJAhIT306H2R/0okynIJe8B4wvsagU
cc09cOpAL7ZMxB8LnQohzcYUF7MAwBSfO6r52N3ycvirQoMrdDtJu+IR4Iujt40f
Fvc5aMOOs6181f52dgZvzZcH5Ci7cj1KHtl2qMGHDqbCjS7wU7F+hgrD8e+pqh8g
iUtsiY9oFrjRuGZ3NCukVmwVgU4LQFwWhOTC5NNy9tZI2TqbpvZVFfouMvfCirnB
Sz1jue5C/qeuJfUFxBgpaf/E/EN1X93I7rp8M2QlTFxqdGBcPm7b1+50uQJ78cYE
ZGYcSeak2TEt+RJffibN8MffrVEAfkwZU1gIRTTOBdUoBj+YJgaDlWJnuX78Kz45
EWDyYthgP+PhklznEINOB7AzBYt8kZiaFKvPosx1t161EQutNSaZ1GVEAFiQADTT
NK+cJSyk8DiMv3piUJZ2b4yAY7lvkPLfVBM+JD3nNTOBmaWuJXWPk3YQe8cTWbQ2
5Ia94eity6wzWsBWyvYMcqc5WgYxxQYtDhgyzkxH/2UUmy0+7cJ+nDL4VoM1Qj0Y
CHW/EsVsEL9M99++TgSMOW1UMrQjYSykmOUejc3V/b0eGq3kz9LoHGT6i0Z527bC
jbBUmpPTrgUV/lmtpbmIcrrgHGFVShrx2Jj9CcHGHB7uQ1meBPISjy9BywccIHvX
AzcQBNXNTEET0+UvdPEDa01gmYUPZ4y5/SWPFgQ29PtvwuFC4OQc7D+7LYOK802G
ZUICxPZAVLAthCdNhVT8OnP0kYkbJcx+WNP9WNrjUE+EJUxhHdejvbURD9hNPXbq
nKVqO4CQyGqXF2MOF8dmd/a4ASfcSkZu+45NVwtD8Lfn049bfsx9+QZd3DOyubpX
UwmzYpL/y5AyFS88AK99C1YQd6oGaCLpeOAHC+1QErVJ6IsA1L+dnPf35JlFClZV
h+Ec2KAScsLMQ0aBsanGVO+VzW7UyfeelAzEZPYAvqUIh9PqIkKnIYAVhvF0MsEo
ZACxj75/6WPQ4ohYSY4CPBbwSQXoChMKn8heAie/HXP66dx7mrjQ8P8ASqMBuNz/
1ApntUAQfRVGZwLoULUGpXYFCmoBxuoZWseTNxvoviu4RUw0igiX2ngjrEBeALLu
fV7CuLyZKgeBsXBZP0oDflfOSJou0CKBWQsvF9RNu46zKSPhVlPYp2Vfdit0kGQ5
yg5IIbG6uMOLAf2MONztGQ9wLqIFHs8+38QamPhDPcgqrtuEW172svaH4XdEdyre
uGXYNhhfqc5yySkEGV6PKGFi42gJqZ8vC41GsrAO+SZWVa9+bLoooRTXdarfFfQz
XINQz+KPRfVeZHh5cuU3o0XZaFkazUX1UbJ5uPonOPDPYwMDawTfOSSXNWNODnxu
EVn7l2wnCOtZKB5rEvaAfx+FD5jhhXTfI3+n97f34SHG55r8T+B+byzyNP1RYxTQ
sBjdob11GTgrnQmaPdjS38w2M8GjzTGPsDO2Z0+C28iGX8/nXVGuFu/0IssPIHdG
KKcC3JEgIO69CyrR0PzLQ6h70ORM2ZJGivWTlNBvCtmzNYrZtgI0pp+kqlc37GdH
M6OLxBCW5iegFele7VMGepFk6rPdP/PDTMeg/AZn8bgfdD1XBJ/WrpWXUGAMoAxo
HMUTzIhWuHXeU9WFed6dVkfDK+LH5tzf43vFkM4mjsJhLd+5R0ZSnl9OvlltpcxA
cNKS7dtRDzvSqvafm3DULnEMuMP9Z9hu5oubXk1bdOk5Sr3HiEnyn5Yt+4DoEogJ
tKxNM3yXzoSM3SsjmCZb2koea4zG3SlkLRly34Dw7ME63WKFOOsgWNa7XhKGSfcv
BRC0L7RCUNZr+0doR4MtWFqD8uCBPLrO51XQGdDkI1VFz7k5Xpc1VlvC+tEfLJeK
G2N9W691HY2LANDXKcgov3YCY5XMGkkDQSMrOKP14hBZnfSmY9+sVqOq04KRNILW
5SYZK1dFttAE5JwmmIfAApGncwTFqXtxv/Nni0jYXLN+2gnipf58AanBmBlDast0
82QcPwB2WhdP4RFdIT7SmP//48hf8ZY9zDSlQNm4a8+b/G8Y1bGzyZofUT1SWU2I
q1Y9N1cylfiyxEwrqVOjJXqElLKTK+6euaM7PFMIhf/LRL2yACXdB+X1wahWH1oZ
OWNtLidpRugAG5MXsNDMGScQ8Gfiq+R+IKUmFJnDWpbSUXRjxkFh+bbGgDFE9Pgp
cp2vZz0ArnqXxKiO+hU6fWioP+zJXVbjJZyWyvqQ/oezWY89hiMoFh86Ar1kmJ0k
UAJwIswNP2XCY4IkHx94Nvej1NaOrx/I3sCs564Cor/XcKti32zE64r+ssGwMCsA
Pft0i3KWy9lCbqfdN7Y/4Q6HaXdj8eWlE2BQUXC/noXI9JirenNGuV+hKBEOlFnF
Ix+w9I/eAv2cMSNZ9a4cZdmiK1csfBvd+2+jFOplWKCcfTg7C1NKY5GX/HeFDNwd
h5NbmOpAqvsTJzf0N6yI5Lt06AhKcqaTt9ndKVSP1avaqA7gFK7fMbysXotbgRWq
rKQyxmWfNz9kcaXZvKlKwDU/i17ZyxbKWt3hWkE2+OA9d3xGrmi+ar9Gudrd1xhy
0SflgTewosXwIvUftXDO3WoxWb3Cw08KwfofUVh5VThPgLDkdJ4E6JUeu/3Cmq4I
T7SVNsBbyQJXHnbzymltLOiP1eIudd57Wt2J0f90ZXk54tSJc83qoGbkKDGT4vf7
6YpVRx+k9cFSOPx+2hxNNoKpif4CUWIXWZ1XEzMtFlBVVrYgDJDbvW4XpgNS2/YT
yfHdQJ0i+FotcFTnucZ0HfMbFChHaW9kb9xa58J4znSfbg4D62lBoEEOvq3MZTk+
oGiOhJK70isJkWWInU9ME8RJ2QhQihO30+khzTjgpix5VRGjDS6hpCYv7AIGgmdX
bFSy3yCWXE/n+lNLjahxrvtC0KRga5nFSIdugwDlJIEBtN1ZMTmR/2aQKQM9RmfX
gDQLVWJ/TuSWvFbe+nLJiW6ISmCwXhKZhyJc6+7e1sY7hWyitPFJsUwZcpQDXEGp
dxoO8BRVFLvHUf8DU5CJW4ogzy1NxkGXcyKFPIeGEqIfJxLLT5AiaXHd/3s8FSqy
T0RWvqujv+4vfhmlqPZQNzO4nCVOkWK9htN+bVlj3KhjGxXNpqozfbviNZDD0S+a
nAnl9Q03ALiRHrrpckbNLjelvxDx96kz5vbimpjppawUHbrqMTdOZ8qHilKtm+lK
qoHJCq8ENzLDQY0iF/BIiAAzmzn0iJjxx4GxqHGeq7VLQamsWAiUlUgArK7dIdbm
MP53imQM33xuuopEBYioHQJdNgDwXaJvdBH9EckQs2P42RUKPGtqmF5bBA0cLPLe
xX0PxUm67N8zStT2zx9ZKd7obymIEQfPp2Fc2R8aICcbebnzanlxquDNUsamcG+9
yPfdTh/TWHkTrMgo4jXXnYZnBVyIysldyPIMKt7ewJjxtPxuvIvzMhVhjB80Kbrb
am8Ss4KjvaXY3c279UFYyY7/p2kf38fqnY90LrwRxIZ3XcyDlPl3ahfGU3Ja+Pk4
oei2iuAug5my7Oy/2qIqOQnWipa1VEa8kJz2Nn8q6b76CohJ4FjQBpsxeESC2O4C
4lEzBcLSNPCPt1iNIiPEC12Yhm3kPQ8FbSB3x2jVw6JNSvI3xjMkBhP/NknTbN6P
OncT7ZqA9UQiK+TUCM6mC2JihV/xm2Y5/KMCZaDpebAnT6VIfIP5imQz9w+UemWz
NJS29MLrDV4OY2q7/1LK770Y7t+1fyScxq46BcIQ7aalpHFuSd+FPWMZu2c7KUpa
pc5OH0Od7FawaNfeEjeK8+26dkYnwc58X97d3m7KA11b7IF/sQlx9DLG/ahIBpz1
k9L/vh3/dNBMsBWTHWAMqXW2ll3seWIzXXs9dUoicIFrZM5jxDrrQauhUME3LIAE
dlEvft3Km2/0SwjQxXh5Znt95bNDjOlmm70Jf+OCdbGJNg11/V1JnqT9sQmHvQ5Y
BYI4lOj+j0n3bR3QXv5ktZzJODTOy0mXqYa/2oWcOuDfZvFc5cBXpiOHGynSYC4p
Um7yB4cjhBtWLpHFEuHFY/TQ+zAxmWpkqvdyTBbfTGzLJ7GMUFpFKfC0P6VfFnar
HC5w3e6zYFqSNkkxardJSB9Cs/YSfWirVsyP/z7qJBirR4JaIDTVwRaJuKb3KYyK
RJN+zfg/RjzAMKJBAw3Zp9oX0w+JyPMIfQ+TkhCXG0yRMKKWb1wivv3pyQhOLzpC
frYbhV7T42DYmiIDv4o+oSruhmjsqhjgOFnoY5jM8K+r7GFF+MeE49zuMDN19v1P
trUjphwVzJvh+in3x2O+Kx817EgbjVTgWJLAn8I+pXnALJ5IgkRqniDojWAiSqe5
GFo6eGwApHsBPESBFDvfq7KDJZq9RMGmMnQWpqTybe4qB1pQluu+UudGbYopjGob
QdzwqmzR32SdGENNQ9oKhI4gByxJXHbiwX4QxWiToXjIXND9vXCauUUeCwbKGyC4
KUQ+ujVkJ9UlMybjDArgdqqvI7hp0ud/lAksq5JnsK3uvHRYMQ3j7YoUN5Wp4gOB
JteVjsp/vsmkOjrJKmHkukxNBO7FLJIqCMh7yEmxuB/8920c/OQJoCOubNcPys9A
NP4Bol21vjGtdwoI+6TeGNleLhQhfcx54oZ7446+nDc/PDvwLUm4KKk1PS1skXv2
GwLJvTy74zJ/pbQa73yimf+49KBalY4NEwh4Aspegaz2TRYz66SbhkdybaWv7Hhl
+HaXHWfgYT3ImB7hskDI77mtda51EQPtv9IFgFQEqsxsD+yqEB5uVtO3yFFblQg9
znCYM0vuH5WeA94GEyQGTdHhtb1eWLtIaw3m26/Q+G2ARYksPLgXYiheRpupEaKo
tCRTp4IP64+TMQKVtnU5Gy/X9Omvx0Ggy3Y70R175N+O/1zpXzd0WKigoUQ65Wkl
v8d4XAsa8MYMbRKCn09PM4Rh3OE7ik/EEzwaobbvRC00yDVPdXBC60wZpWVaRpYd
6zA/l/s+KBnSAWj09Wss6aBG7I31rZu/jATjnehNjEUf90EpwQt/lmjtn49tG+X6
ZLdRYmTCzlmsItF9KjM6WDRNhUCC1Xvxz2DKYp+X5zqb/eXwMZZjz6XVaLTWodxM
BVbWaeX5KmdMQvdij3ujN13NHinE+GxWfLCZp6IvxfOnqDBsrIkqRnR4fIhCyiBM
girTxqGFP0hWO+SeFn7BAQ2bTsOWkf3p+zl11I1XIgxcCbg1y4QxJFoZ9XSyklKC
A2/ZEX6vXE+rvQy12ZnFvGSSrGQdtzy9MAF5/F4Uiu4agaejrLAVpHUiRu1C+0YE
9Rgfye2Oo7qqhwVuw1avMdHRM8ljHdao7TEtgQ0w558Etiq6LBz6861/UDLmPu81
m6NU0taYYXtdSMAJyCZ8pjMlAze5P6lWUHtP5xOtA9VXzXHjDo7rnohg1tcqnggn
O2t8Nv43xJECaXN3IyF+xAKPHwnYoBCJxDyfOlGNy7bm4JvyY6pqGUZvy3T5S4AB
qJtORV5K2o4YBhU9CYSJEu6eNa70aCuH3TavuHWsrvceaFFXzFeythABhIffOFWp
OJlV7+23DZBgkC6xPzpahFe+DD+YQU6qmWMeGtkUXTxb2GaiT5DWl/pSRpHTtKdf
DPV+yUKJZtjcdOBil6d0tgoY3CXasxNH9NwDNwWs9g8mJpjCvUichgWjcbH6LOz8
ibUQ3jVrO0qfrwXDAiVgG4qv9vHDaZVWgXRVhcdeQ4tsgOlXtBdAeTqy6GqI9f/0
OjeFGlptuqalk2/XTVz7mWuVo1aZz7MDp/xoNBZNaSnQskv9zFxuM4cyfUEBolkl
2exOYBhrSsaNixr7gC98DjDOfJwkSn1sKMoP/nQaFIWumn5PoiZAW0kCCrTdOewd
I6hGnwgUadrX4kruUBavbzu+nC7cU74v5cKU8Vzar4ACVymFxyd6+C3Tx1V38uOT
/dF2DVoLQ9csfjj1BIXRQQMpwh0QSKhVebpAgS9JlqDJQnrHhl6P2feS1EfyTmhX
KCup167PvRbgtlvGb6VHY+l46c5zL2JpQ5aKETDCUtA8qEJWmKicbxVTUwujXr2y
89/kbZlCsl3m9OCFO+i2K+mkSEOpVnYVsPuCrXM8hxStIRcbCelM1jg1MRc0YT95
o+Jwcvp7KrfcmrpMUyWHx417/xa/Gmp1tPZtHKzmk7FidgpICD8SagklEgVdeads
2naZ3XbsfzddKaLePxvC+wV+RhQvu7cfotCgLHcCsH9KcO0tdVy/vB4Jl32O1EST
EpeRmTu5SLJxJ/l2qTkQsD0rU7IJbeL8wogPTm4aaQ4ag0Hu7Agzb6GaXWEyeSNx
hlmfvJgvJBzIumD+TWGE4Rz1wCraPi2JxcVftUDFgcjWNV50onXXYoQ4uY1xAVzw
VKI7AOrNLvNpv+054BcYJjyO0ic1/uo0KfDwF4+EQAoXyAu0r9JDSNCoNzdVQ4Zw
fjxjdjZ5PSHQ9NIx4SZHOtEqDQAx3/TNUhuaDz6dDF9WwFdzRRNWhZ2MZ2ioaHGS
/iUbmpOvn5TBpeSNeGQkrpaQ8IPjSYoydhOHrrEo/4UJC8BVcUpiO22SsKcU8xHr
3E8AvM1nZvoMJRO6z1tS/jiAQLsLFpdvRxeGvoNUpQrT9mfvFMrjf8KhigQqn3DW
pSUISf6Kw+Tl7s6IV9DPyMa/6o108nryId62V2EEo/V+ijbPRde/RUcTGi8uAL7Z
v8GCOIW9eynumAxbZ1CEW7uyW7tafniQYoS2MzgPJc+peIkedQShFxAtdFeS6Y4U
yW9gB58rCd98CyKPm82wmSDHYBSoRFwugYVOoWxWgPu++vcErkWZKN/1GCdziR8q
l/iZyaNyEQgCz1Ept374ciHHBTPvesn9Ct9oAHd1wVj9a6cEBMSwV+pEVWQb1a8V
HUZVOdLh92+SGz5Xd5fGwu9PMWPJqx1uFKeEkcRgPEyT/1rdH+m0Gg1BvEiE5bhZ
Laf12O+Tu4/7x41kTBcBPSUdack/Zyz7bdkieub4y0A=
`pragma protect end_protected
