// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ScH4WY1unRue7jQ0AjBupqNz3rUnVVcDjahwc8+ptnyzYfoFnT0Ey5JrZuwvn1MTYPFj8b5mUP3i
rX5NdC/hjrp9iEiFx+av9nTkF1aZag7iqmGrgztgITSpcdG/mHntZRdvwiTripUDON0XNjtAPqLr
mB7uELIhGr4o/6OTCHAFx3eg2Q/2t6yroM1iXeE6ZtJVzJFd8V1HdbVoXoHG9fX2uNV5xYqdjhP5
kz+sS/hgxbHqcZ2yOVQqEW+7C7nPvjap58s2f3Ob7bpwoqp0mKa/2dC4Ad6ZAEI9MBS3FxvKi6jR
Kwkvf2bVZuyEwrru7SlPyDNUV+wX71EKUh6Btw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9008)
BAwWCOaEm9obnfIrouCjLL4CfVJqZ92tBK7EJVxx3MJmmHS4Ifd8Jrp/RnK1NHQQiip4WTma5p/n
iEwZqDPoX5SSYD9ncnlkTFkMbw0tbYqt4u/drwkhIcWVonZspuG5OfVhlN3dlR1Y0O+MACbepObq
3vQJaRevQQR6gsSKXHTx1VKSdoW0JmjqDPZ7zUwzrHm/7ENJoxtUeEv9sQ+UPio6WxhDDeQT6qWX
pNBVCz+9iiVZ792HBvKeOo+8m6mD2UVuMI4TqZWFSX7s7jSTxFBcz6qg1Iod1jP4tcYK9WR73adk
3ukQj4GP+L2ubxF4toEHgRW2BKzPqZnldR615TmymHcNxu/dIPYs+bnGnThVcsLbPx+ovpjfh++S
PCYfqstTMRD/KNIq9Hd10un/9PFK/QEJG04Obq3Vt4c2yKMz7TZIsYr/y3b14GwacoJ6nkHcekkb
58IaSb0ie7qzrPAaPIBr8VIpmsDf/0vGx87soCb/qdmFs/75BJKXX2qe1SqLzH2KUGt4h2GXYTaZ
sP8Rn0mp/F1ECYIg48VnPPiLy4l2rrINvajU1ueKNCh69kyXaQF82URxlZkX1s+5F8E5HgS/OOVp
JrTz1+qJtAnuUiF1mwrgrj9M/J4o909STANftqwts7crGlfuiAK0GvobqjvX0rYZZMhxSgig1njO
zTvYwZCbxSIy1W6j7aVQlEk3RKo8illuHCpbc8WXEG0n8yERJWjN/uZa9vYoA8YwxvKOdTiTGbCG
3bd08qdJ9U2L/IUXXynLD11GGhPYMTCQKfBOOsuVRtsAD+HF7GYtoCWBr7KFbLF2Z2zEnoMZkQog
cxKW3+nPz8kiOp0E/jgkPvnq8SAn4CBU0uFlVZt4GJe3j/wX36aixEuOzhMqGbO8FFx6FcdCz8yD
eaTXa5+9SnrCoJ/hdVvdCeyAPaHq9mKH+Xhaaa6QtfnZGf53ZHWkl7dMT2uZyFV+/Ze3kIxzg/c1
v8rzx91+NKa5rGJls7+S+BkqWoRZWrR1NNIon83eYoYlmg8vzALeTTdd5EjL8Mw6sdeHEq+42ua+
XH1pMq8B1VKGZxOcDaeeIkaf1/IDgMb4OKbtMpH3ZNX59Dzk3GhYJlD9H3jH3WaoVs670A0L+X5G
hFOp8N/WXbF8lzl6/AOGB8BaYBpLnpLcY1Hfx4/i5fNOgSXbaTe1C/Jm9JVXb7rbJx1c9Enn9zsj
ogME9pcCIz05gnHACJ+Cfb6i2460lpx2K3IXsMHdT04qe/CJSKr8KcjH9ebzRUSTIPEI7Wg0bKQC
vaqJqYd4Hv/XhMe72JdZBfymacgvO10rOCh84LkfHaugnLRBOHb6KzRznHMTzJv3ssxQ0dDTbaf+
eNlQkoNW8eV8h7T9gaYoABcdajloRmyfgdV60kcmG2w1ToqQqfo9opaNwAKQwxYdtY84wZTWQsOv
nECtNmXeY5rdauZps7QEZ8gumCs/LAB7ARPyzr6uDvevElGRSXZKwvezvmNp/dXG9CPIgsuOxur8
CmurNOk2SZFqZJucyu37f9858PN70IrDUVG9e114NSMZbLW/1SiWstdUY1nb4XdHZTt0pq9mSY+/
wbzOtRdC4j7OqFrEQCcMVWczP2XOJX5BfqP41hhrVUrMbaMkhDTjN6OjL9P2tqmzYPnwdflQgeUS
K2obq7Ibt24pPAxwArpCH5iR+QxmZMQckW2UkTv7y8kaCcVMKCXBwQCSHRcXiR7djxyENAtu/Xkt
DERg1sy18Dy3TRG1TptuYFVWCfSIEjLAKIJuyS7K+zKZVVXcdzw1igkgLLk+nWYDsOfn7hNbmW3P
eWPnmgELUzNq7+YWnaN66/we6504OFNYpHupcPD9w8A5Pcvl3YkdF+pjX19kY2C5piemvGkncZ0w
5jlrEtB2Fx/LagGuJhXj5B0RKkd11uBylprkdFuKXfnq74r3n+68jP0p3TFAxt8D1d+V+2cjyt/l
wbE6s4dECTc8NwlSEeIx04OXrXNdqBGX0g3CB8e8fl4k75kTVuO5h6j8ai8azEz0lMtE3KqzLM1g
h9h2j6GEGJqIrhpzrT3DviBEbX607P4eofkkdlrvL02G+tm+cnvQ4PKK5r2+489Rmxtdli8/FRx0
rMAlD8lmI7V64bnlwZ2HNbDSslSsEkFelSRFz46FX3k4qGa6CBGT0bZR2aP8H0WJTUwWDfxLcDNa
DS3GCNAVH6y/g21/S4DgHi18plYtbITlUJ3bquoAPE+2xirVhbdglArOO/8NETHDw/DMYvs1YyBP
L0KlZxviIr2Fvjd5BFbWjvgZNDqKfCnZh3Ti8wcE2UOOTbLjNYi/3nNz0zNiEgnGYGCSpLQy28hJ
oWDQ5JRp2RpTXrbTuKDv05dpY5K2K3gmN0/ysyb1Jdg1TbXwk6+EMICg7pnnJ0x9LpBkABvPjWIs
XQ3G6P4Kn8g+PrCHfbPFqVP7V9t4PkAgELbOYwG92x3DfsAsjQtF9siigq0kNGOUQrQHONIdok6r
RoZ/qandtMG2ZQ/bnAdooTSvbfYI5R2Wei23wq2cTjbUbXkfNoGwHkm08PSUldBDcIs4hsqwewGw
irp+fq+ZzA6+eWjLUZvEyYgzAyxT/Q3R0Tv9D72OJhOj5NUfAoCghYyFvIJU7v82K0N7bkqRXJ+F
L6mhEy9PJMCo1Lumui9a10piM7+CeXcIYRNFEt0aa06W+QIsLhokBOSdUUvScwdZ2DcZXxig0BGL
ZDI5/7eiZyniqZuNsyJ6VL1H3QKiNsEYRKOzViuxZ684Idh9av3Bk/tpmq78Eo2incnS4aNdwP9w
0Egy3+9/HW0+C6pRa0B/EgsY8PZZaOeeRk06NlAVZpQIxKzqjHrN1dGwgzzoQKhx99Hey2GD8GiF
l3Fdfn+Vd4kOrtJ3iXmequQXBWM7odIT5mV+84oyU3V+Pz6jkLG9WgqDgVAhMrY39t5pKeye/WXO
bCyblulwE3szjlLGCsK1rKoDfWYv5aZHVU3hIXFE9NerhDjT+698HBLQp71oL8KTgkxZdbWX0haF
umVSIEc1XTDnMSrJYaGhqBjhB6/HF7DD5PlBoNKJtKtttLaipqtvVccblXrWJ0qYTEq6YU6iVWEh
YWSlOXdUzfTOhqNtMnvvw6w+xieU1Hp6OhoriZ1BceVWZQPhhg4QRS/z/3211+5Ux0d2/akWt7ZR
sxJRZ0TGYy7jpd+D8VmblIv8vlkkDpsokaLxPZaXpj+eA0EYLKHHmwhvvjFenfIXQ8WP83fTnIgS
SV1zuz5aLYAfVYMw7hjK3+Z+bZjGcHvSlUQCYM9SE47XCCdGBnM9rtF/vRhLY3lJJUVxNlE2eaIy
ATVjjJxSbrpz75q43eoBv+VMrr265EoO1qL3koxdBOHQiiRwxE4/wb1E1xgDayCbgsZtySgwr+7o
nzpKeY1uY+Co/kcQKAAmtfDxlqcLlA6Ow1Et2jjBtw4CMJM/cvKOnTrOOJ6P1EYsfVhAFL2pdgo3
yPGF0IEYvzlEY3p6oqESIcNzMlSvq+CnJiJHrx6yRVe9lL9847VYKON4+P+N1kJ07z0Wgzo0KXk8
IeMtJ+RYwK+fOB3AxqRtpxN/3tjF1x1zrLe67VcuZS92VgG0F6groUDIiwpBmBYxIIzw+3ImhKCP
fDyB8acYKVZZXFm9SUt0zt/20bcJRm3HXjPEQLejfSX9w6xI+HlRZ+/9ysJ9pmijvheW7Q5jB2A0
ZkFwt/pBqGpVHBnqyjH9la7fYHD/5rjlK16iBcndTi9l4y2kslgtTy59X1i5XbIc0MqtMcgtMyQe
COPAS1eEUQvLdkN+z+UDi6MAJ9BvhKHpjQPhd9aNOfRxeTpGmnSibBaO/dD5tgezAQjHQZKC6XwK
WTqivRZQpjG6T6fVYsds+WtjDO5RC+V1e4J48vE3KAGCjN6q8/6ATi6EVnn2ScrLDjnHYVnh52NU
MCMCGDC5OItvBS8Tfqfo/6Amoe3MHwrbY6VvwLvsF/hk+uFNOgC3pFA6Lc2KzLdLvM6+/VJrGpen
880faMwGh3n1Ezc/RFTQZTual5fIK1L0AcLcDgHI5D2TlL0p5rJhDDxww4Bej8J9zGymCW7wwHZn
OVhYX6PszbxGWm2jRB0yYmwFxYPrUiR0cnN0D9+fjhe4qpTHTLzTQhF3QxYx5IQCHvmJlijktOV4
znXWl5WMXWtYPcvNsVxnMjr6brXOiRW3AAbG9d9WkJxacElPV/0ALR7gAANrNIp8jEkq83K5GxVs
6c1aSqknz7MGqbHgGvaFAz0AMdIL87exPJNENn197WItKNQtOCZO9rtU35NH77W2WPKbzgNSxSH0
5t/zbO0mxJvW2SN1BHg2f6asbQHytKzDYfq6rfBdjo4Qo6sdqfNRRkE7N6cVcHOgxQ49yt5P7CHZ
2tTJFZedJUkh/THpasQbYmVZXIQ37ppfN0/DkmtIkljY7A6LhWQUNVBa2GpABOCM8W/qO/OnYYLO
ChNf+nVCTeK3cItRlJxpyT7O7dpHdZAZZNSXGHcSOfkV24UzWMjA3jJxcpsKoEtudqMlVEI6/+xe
ISD81dOGp8MNU+CCMtXsn+6rnFf9abFEoZhGxYQNs8wlDzJn43qoWvKmvbhhPc0CU5HEpO6IxQti
Me2ISdPMbd9RWMkqHC263aGdhpLt24oZascie8xRFPLC2Xm50uczC3GOJBY+EDv+GcdvmlMnj+YI
1Qeq3vwQByJkPQ1b+bTr7SwxOTWtwfuVboZ19bZSkEdFPl2NMQ4h0NqqyxK7FAEeXURMyQdvCP8t
PjkPu6dd/7AfwJEuttLdoAocVSpNLpyr9dgAQpO6HUntfV+LpxJyDz0EJpTC99FwAXcS6Iw3OFyX
qyd1YotvR0rS1jPBQkr4WVARLNtTn5yCdPAuiJWhJdEd+strDHMXnSabF/gOQpxIDBErhhN8iek2
Fy9ANlBJfxc9tt+xnC5dIAzxqKLrergkpqsTsHQDpBgKvKD9XtmBmTG8ZAP4fK+eOZASxdFbIEEa
XfWpN9RpPBq/IXQxMXRzu9Ge+YXqHV4EWerigKRemIAjOCxG8ZyWXGCIusG1H1yYh9uNEw6vuFvh
rvMWPkYSONXysgSGXtdsqCA5yYWxfVSDw6+a0AJ+OV4WDkjKoNm3rGSkCfpy/x3Wjfsiasy94MWp
jUVMy38/Peip5OJjD7DpEZ7dJwGYsWWKvcbu0BJhLRez+XVkJRw2Q9aiqq8WriT7lNFeV41wVgfP
E0OLi+6uprxCoCOueJMyRmbeDsMCSjPAikZDeJ9B9f/epfg8NMNRSB9gV7DEO7f3xWvqfLQtUG5q
SCWxzNw3WFYkKtq3aXzWeOC918totVvaONCdeShOJztqUMm6p7tOzsdN+rR/uNFLw5AwIc7aUpQK
yNDIBTHaWJ2RPvzdEHYi4YE8KnqDXyjM+7t22NU8TuJ5flja2fd2m6Uyr5vytMUNkAtMZ8MpMIhw
39rY1cU0hJWXgy+tHGPQvMDRKeLD24YAXfaEXyodz9xkPmaTCmz9PFVmMcghAiIME0hpJA2zOlRn
X4U5gtFRGzWqRo8C4dnuXQRAqKQEpcjdXmFpX8BpfPKoGexZqw62XkjdBYco/qQ90ZT+NepF43JD
hzCKh1j/bpPaTROhh/frNr39RNICd1FOG+CFCl+XwMX6SKy1qIZbWtcsJHw7L2cIh+CjRHaZ7iDS
W3Bz0yiJO6w+FLYEGa7z2BmocMfuCmmhGGfax4As9x4houRuG1TzrFkXRqOgFROYSOSSalB8hWiC
iXZKOsBysDFVgV4gj0bTY5Blo/hleyAe2bdGINIuYQvf9EyThzilUGjOpXbkT9N5qLnju4M2E3gw
8ZI1cg1RKlUcevqLRQ81+T4/1UbrldUTiu/jZFlXiCZcS8P9bRWM1hbd6R25t7ekIvxmTMVKEIlo
1sWHMcBFho4T9HaUZkNUWJ2XLzBa3qV4BEgIklj1MFHyVmKoxR/GvJm/bp4v+lrPj1uw5/C84JUX
nnGk5g/qCnRlGAmmu0exYN/zvAb1VB2BD6zxDUR6hgq0/JkAPcrJR5P0rAMyPmOFJ+N+W7VLtR3T
Bgl9xZmhFWA3JcX5/gyKO5UNiY3sL1uzu5cqC8WfANoeD6BCAt5aT9/OmpjlSykoHLZveCqD6sUb
EMKfUeCpLBWQUg+215iZC4pxKX2tflAHIj92REsdAAq9J22fY/MsiDWyP3Y+tkRWrDksPvz4qPHc
HKxBUP4VItSrazxmRo3BTcvV/8ofBP1vQQLzNM6C19mtRw/vAhopt3wwYHgx9EPFmDCZL6LtgzQ7
hk+ZkkYNSPbPH+NsjDG/k3IeCPwKp3bJLAlqEhIDssO6c6P05qJkNdtQcQx4Pkm4NiyUv/ADK5Nn
DBMF15twriyzeYtmfFS7UZWSFdK4VbNzHQg0bkz7ZN1xWaFjSVD/LJ3+42Jrn4ZplY06MR/Jg3xV
Bm4UGHb/YeNQwszG5u0c9zPJ7N1RRfeVhDU3NGJyyRm2+z7soEVv2siX7q/nUhTF48Qbh8Zzc5RQ
Suyhh8aUYWTDHNGasjghMYVOWdOQ5KIrceZAUkWO/mWUQVOTBgjABfQhvs8ziySuZDtVTNyvwegi
X4LcAfgng1LvZAdZIlc2u1A7V/2hBWvEnShWoeuRTr/PD2jbCU8ylzVvwBupG2Uz0FJdITxEC6Xb
Ok+j9JlV9jssmBt4fyCHCovDzCHpdYFs3KPHtIHRuUGwhXQcvmmT5lDBFbkthFNOwjnf3Ehb816/
ikTf9X8NXdvYnJRUpqNO8uyGeb2XIzX2dDiSnxA950Tqf7K+1Bxzm6eGJRzSnPjWyYkXYCRzdlH5
oxjKGN3uzisyfJQRCvWGVGq7R1qAcZXOcb9roCKijAqVR3VPZfBbR3wZfnwkdOmxymeEUthaigkv
1dCo17gi+DuNlU5l4ZN2yfxfQ7XbgN3y0vQskz2zoaIyJU28zBFSwoWzmXfxjRVbOzkSMzRVIQ86
f2IwII1Lt3tFgq/fIe+Xlmx0A+cx9L7DqJHnL1g0G1TRu6AvQy4x1Ii6S05cDfB4IkfzGWN3xjK3
PDxIMbcRrtTvSjcykC/BKSCSZbnBGivuU15CfV8NXahfd7UPV3fWx30G6AohxVE1wcMoQPg/QCN3
k2WnY4A8wcCuQ7c+Klbv0VWZQdkieywCNvOHG4iEaDIIwRDrzaHz6fOkaG7XsJ82tBzoA4Oa3s2f
bwe+fsKBVc0/fLbhb2BzgMWW3zHYW+ZtCx/+9LXT1NZ34hYUV2MEnGofu7aQ7fBnAqyW5vGiz77f
PFnROqn3GbgDWYT4Cu/uSNBGIEIC3Rs/lsL6njOdJzMtOJc7yrzqO4tYAMgK1mgKhMpn3uph79xa
dD9J6k8qzKG9sqthv8pYlvpKsXmQqMoXLev5Agb1jjHMEnBN7IGcR+hrig6eJA3s51qihlZ+Ezk/
t8Kbhf48hQtB3T7BHdwXVqL4+p9rUy1fljaFumXHU1vDa1988wAhL/V638WgZkNhYpsICNKsouxw
D8SQbr19dCA5cGA8ksURyZvRRC+oP0475qiZoBg9txe7aFNrcJ/aRtSMkmOXcmxPyK1pGxb3SctB
HDfd+onHGuGzlPBKpxiyRMCF5BTAn7ynyR9ppPZdyntva8D+ruOwxw0DBkgl+izUDxyX6q6zpT1q
PaUO1a/X7Ibn6wIb1FL3bsq5kOrd4ZqWpWa406m8leM5TKpVtL4q8veHcKvZJRUhSDj7l2j1aIDh
THD9jfTdamjIXdvIEYm/oLUGHumPn4PpNWA8O8UsO3CAsbCvsb6hCpl0kNV/8KIbZ7L1zZGKGgAK
SnMoDbZI+VBWckZlSJ9ViH3iyrq9c4c5iCtKxZvUfe5k3e/KQ6b2+/K9syz45rtTqn0TbZqIh6YZ
xg2fTrDPxF9GIPEVFL6DaXkjpxXlGoZhSknHLL8gY6b8ZiWGIhpqIsFfLYPSxZy+Jj85iyaek/xU
IC2AsaEUBCpv1KekFKKFsQiS9c2gW3pivFYMCTyLWJqQJs4KVl6tv2eiyphRcJTh/ccBn9hS4Psn
2qE+Aq/xPCOgXebfVKSOVFH9KAv7/ZCDregXh8so5VVsgvvz82GTTcHz9dCxf607AOKqMxrtzImq
vfAUJLxzFNQarXZa0zGiWd5Cq6atYE4R9Qor2SOlCGB8Ct6JAPrhGdngDY5PRQm6LZc8Nb08UNd/
EgMrJt53rASde9OnnZ5vsQF3vB3Q6Nif1HFY9gnzIT41OxlVlCeQ5nleRY42vfSB83gRw7+18Ywb
pjzeSLe/CDw3MHsO7dSZDCWdp5Ag64kc/VdNB+BEp5tIGhWaJCQcRsZDBqthgf2Dhsbu1A5WLwrf
RiyVoN03o2f3Ngeo77eTIgP9ewzJOxCfVY/VKPBTQZwrGohhwCZeWfisOGkAItNFrPuNXS2MEIc3
UGN/uhRblnjP2PRnIpiWQDt6YZA3xHLjgGsb6tc0HwjughAOq75ItSvq1ZBwB4j3+gc40DkvfJhG
E7MAChK4FjidZhsjni0gXg4gipt9hfobWGrx6vepTc4bl288+Fii6HN6gxe7WdsWmLcwH7MXWIwF
yFRhTqqgM0oIa9sZOtm5ZbqiczHF46RepzLK4RGKH/Ro+R6NEbUHqZ8kxHA2g5fzZ/A0qLqpwSjx
cIXz4L3OzikhvxCN91OZ3eASxAvJdYuMjqjd2kqqyuEhaiZ472h1Fg3/zsCuzVZfBsDwNJTF8oCN
xydTzBJ26OVesHY4qstEi+iiu/68DTzlpsxpm4Tuyw2CLPL2m334D3Ofg1BPRDG9OSy3RDd4dQ3R
qX4n/4+4WwJkgRMaZe5bosFatBdyCJhteu+6HGkz0+fxvm5Hyxr0hCl3ojZifHsq8GlWsNA3PQXh
tk8pB0APmM0RJUmnv1XFYDvzi/coEJL9OyGWbozOXxGRgh04N0YAtkIDQc3G8x93ApthtD1dSNIo
PTOGurkNN62wLwjtPlB3LsteyZR3xImrrvQQnUpl5bdkItZ5lqYJhNfAa5fG4LfJcs/beyABu726
wHO89CbUZSrGzL52JWGkzb7m2ChO1hnCI2DDb5J1SjuSYuvdGIIwpdgVWM3Jveyvz+l26PbbJxdh
GrJWo9xYQSn/Gu+j+EUGvUxYAVDdYACWFdIkeG4HeZmspOF3Nb1ZCdHR6SsB5lUQF1/mTCygcv0H
/XpBMGCm4AkwRno9gVxKDfnSCc/fwumwiQySp4jDbt43t7Sj3tK4Vp8heZw1N/moiHJPLwRujGcV
SXxEftBJTXI3FyLvXMin6Sjzmce+2bJBVYprHOUhVYcPiHxNQLVYW4aUlIzsR50zcG/zF5p0rYjP
jYYqkmadaw+9fUq14lNljw9VXBz+6BAm3UYQF4SPQ2GV4sTl++D0XKPk8s1xZvpiOzabZC+P9UR1
GSFfe5+Lqvj/+Cji6tktvgFDQ4rvnXhlPmSxnWolsSYeu6yvigWzURX1MIvGP1KPJsn4Rc49HmMo
nSBkMRJT+H0KGQ3H47eTwG0WAvmEP/yQUwcuZ/1en14xa/OCudC5ebUO+iHWRt2b9oNT3jE92uEe
VRpx7xPDuueNZR//vuEbajae0c3WWL0Sc3lAtguE9QN2JkQO1a6UhbzoxFMFtc6FQQOVIoyUrEUx
tGzMr+TWvKK8jOc7PXL9zRLXt1U2JwzkXGnYi7TxyTboGMvbKWzY+AQQpmKBzoVGV/WTa/skALw2
KPVVQESecJt0zfh5tXamtIpGZgmTIFF6nR1vPYqG7pE3kl71FqgbaNqmS5nYFheXTAjTVDEZSQNS
o/J/MG04BEBwembSmTLDm30SWvgvu2oWXEilKoMrPqdXKgMJnpg+rza6MwiCB6azt0tFgkjVFZ2s
jKn5SzUFs0DqRE4zlsK5Je+hT8XnoPBWoIY7QxTIdsbIuBSVO+kC/lx6C9Q6duEzT7D1MxB5oRRl
7eN0z1UwxhzzbErHSkzfAfOhAMmCJ+KjEv65FDhqTGaY9s3dvVp5Prf6DDoFYWeyCWImjkuZ0tKQ
L3G2wbbKPXPm5gc9X0m9O+7POFGmqf5wVVzIDcYYxkXPK+qaTe9pRM1G3H6csJxv1EbDpDqyrCTc
vw5NHz7txFjp++UV+GK0lpVwjlrwTbeOcplxnmr3+8kuaFzQhdDzHvn9Ymdxk0O2t+Etkp7t5fig
E2NyzJWEWY/0BbZUpyKhqVuZehJBN2bxOwoNLH5Pi/UkDeGQ8CZNWR6nS0FtbwrfFZVkJSsd65Dg
TXmTwYJK47LdGvZGDrMnD7G7oZwBFQzxiA58ue2vMhN1J1YC3G+c2itSo0x8xhjTT3XVdP8cFeWG
vr8OGQ5YvLgQqS2cDkZnJfTDSMoZ0CJd10Ljo2pKNhiYEL4ppSuL0o8c/E7hfPRmgNoLp++6NaTa
hveC3cFGj0CNtH57Kmmqgqxi03GLTSQW04B88o1BX7EZZzGgaTrW6aFtq+cmh98KOeNGEGtygsj4
t+/6+yjCLMcBgteL/tf3H9b/4a0GJfaJVUwXPWI81swI85xHFD6pdwwTFuFL8YtUITJBEWhCLuyH
i0wCVRmu+2/iOsYgcQVlk6stdVbmesSebeLQ7PkT3SiXIxCEYYqUujAsh+b9QZae5gpjmu2rwAnQ
1hxDObnaWvcWghHkx4ILaXcs3DG57Ts4mV/CetGppL0yPwtrJoSv+zU8lL++bMefrkO4EWAsuKAZ
4e+APdnzhnuIsv0OdCHKNop6zlLHzV3NvDUSUITA1Tly+C+B8qaRFIHJrp/OY1m9cY6KuFMHQ2/C
RnEtZbBxOTRKtFBprlWeUlJEyOiFuHWUTHI56JUmBeHFMSZpqltP/kJzmtl0oItbbl7/MTRQUQcv
ZHDbkYYa5FUuqd7e4UV2XWeHTw0XeXgocjhmAPqFKHFaU5PxVYlf9XfC+X0F7Qa8k0uVifgwIGeH
L+BajIeiNvwHa35HUb1ZSCxPagtYQmdJIwgvu3zJi5zPLsNvocj8wTIFidi3W616KoddpTrpekpx
qDt6mZ8IeegiA+Y1zi7bsaPM+qRdPRn9V/YZWe53Z9quQ3ibtSwu/dhB9t9vOPumSJw2oMqUup3t
cRGA9R/Y60twZrV0KWmkmE6pGGJd6O+2S1Tpm9brALhN8fSfb5bb0lheDXqNpqMvKESiI1KoXugQ
hVbbjbcaFHyYktdE1qQROqw4SXHao+BxpLiHHj/eu+82KmMbdogyk4ZSglLR8IGMpvEN7SDzE5aN
Z6WjpL0KkhvwRVAWGoFHg2rQr7ZeWSq+WscV/GeDAypNsIFCJntkiuBTLr1mxpzm3zYEfXXeQOG0
l35rc4ui9phZ+6FqJxa6ZVxhFARQwNqUxbRcs6rWR8wydFfXZf3FOEJo3GFmIH1H8SWLztmDkndP
sPNWD6teZGHPRSwnLb+/hDTk9A5HDIEpDfK3XOeVUzAcz7F5KrBO0+LDDrC9qBDYShh6kBRUJIZa
b/HqMo7p5lR+LWco8nOquGkQfWDwoph9R9TfflDzFMhZ9WJgLKphV/R2xcD3VOMAmWsEdilYK1SK
TCUfr3ynTY/+865OfcHnYlT5L6kxa4l/fUg6CckIMyPotDY4DS0g0k3uo0BzYDpoSXiVPk2G5PEW
L4OrmS16JFCrmcGNU/a8Gul24aW6H0sO4Szb3ndIynbXcdlYahRrVtFayhVF8g1ylpk8+7EyN19P
8ZQnpnpK2jej9vJdAI8AjdNtwDH3ykChAL9JTcM7LvlEdQGn8H+onfzQ2ob+2RSMFaHgIVNJDWuN
uJntnx/KCdG58MRy3EayWKPoB0BO7kjyZZx/3j5eExd/doVWzajUiwW+KsEebaQ8vwn5IvO36ger
wgHoIZJVPlE7ABqHm4di4O1cJth1eCEUW4ANX+j3iQAJv503Q1MO+9ufnXZQVDZdYEZvl7CLZoJy
1fqJvWYGaS9hRWT148SJiZeBvXaPHNOO4VSC8rdnFZkWRRuLBazXL2sBCNP2GjaaLSf2gaZmuGYN
F3o=
`pragma protect end_protected
