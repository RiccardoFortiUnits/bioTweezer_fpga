`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Q+hcIhzIk4q10aFgLJzL+/DPoEkiP39INSyBSaEAq5kh/Ltyj2sX2X5paVppJy5O
zicbsxuSu4jKPUEZ3PPqrnPehW0fOQIbqc92H0z29LxZl38S4LXKeo4AIdfZgAEP
BfWO0FOSl77SPGC1Y6xnNY6093bGOrS0tf3kGBWKpR4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
SM7EBAO4Oo+bsOzzYDLp4vV8F4eSzXLJTfSRYvJ9rE40FPKbFXDOEG3hikwWAeMO
ATjhNJTLiwdYzahIsXtODf8tcViE6bOsIMWFNxCEX4w7/Ankf9RrGk3KN3HrvCoD
qJn0IoyaayjpiSdihrs5Goqty6/x0jw5lfER1C7lcs4LJkrpLFLLe+t59xP5r8bd
jLNyB3AvY339NFD/zmoDBkE8AkRE7lgDANZ2SDC3YSn7eiVEHP8k0gpEpMXErtIe
+ajS1AK52ojOw1aqB96mhB+o+PDD7i94vatrr8bxDibAjdtYMQkKQYllKvWJDA8i
onKQLJ6HyfcoxSEKPKPhTxBSsEKISQ4wpecijDBuu+HxLUaUIGcigElrUilbVU7Y
tLevbgt4nHZxWEXU1Md3tMrWuaGItd34JVE6Vn6jTECkhvnvQ/rc0abSYz851KYP
dCQD3XTQXarhQKvOYJuEcVzV6UmC5RJ2rA3qUXng+kHnD83Ny3Rx7YFCTvVENt1i
L022LNhRFqhdbsPdrEFDFxIusTAL8gXDuWekoVX5lu7QZDuG10CGwa0IQFcrZ2MZ
hRMV3KgC/5xDbhgQuiPVwca3527+xUwZIKpPlK1vmONid2ODc2u1H0whuySaOUO0
nmdkB8Xdx78XEWOnXHo87EI10/gQibuLPUyqnRncsw89I2RV8hu5wo3uZcsrPQ9m
2+/S7Kr7MGtP+GzONF38k3a3JXW2WjLNrtBfw6DGHRKTvIwpJdePoJtgfkDra/kf
X48r9OFiaJmqN1QlFDMOGfHWV0t2t1YeTEJib2GMAjGSaF2pv9/GhGGK5xpkHosd
qcZySnbLG1WOcOvdRZryRyHgXMKUBMM8GLZRp4yu0fSjt6OoZ6NojoksiHgu4T4X
aHm6RENb0PoK2TvoHXd6j1bGvLmGsPLzXQBEKJGJKUCcEqp6g8fCeF1J7gDit7zr
5/sFceTsAXr/ulDxOs7rL2deaJ4gvDEjb7larneIjiZo7Bh2ZpbraAfmbJW/Gh7p
FnwhJgBsiUrha1TG5YiYUeGW3jFcS3AqKrTJd+rnHzqK7J2VcE4l2eqkXbdGtcYC
NTazuqr5JVC8aychdEsuN0PkJG/YTMxvVXBBVqnUYqPB1bdg/T51Zxmsh4TALBng
uuPe0M2TZp2bp8/JltzzukBWEWroGssbbXm+N9BVx1pLlgTvh9vexvm+PnEKiqu5
8kpeyQEYwcuq1aD4fncm9TV/1rYyOgxcS8/2RSFsrmVRnWMqtsC2cKRH8bONg74+
SlF/oACLkU5xvQqNIa/eAnf+Y9TC+OEqSh5a5jxylSdhrV/xJFFhPnNrBE9M1aUN
kt+jrsBIELpvhG14UBs2wMtJ/7m8Wnt7OImryUk2O8iFTlq5KV49aqOk5JExBfp7
NqscCK5TdmvMjZZEm4rhoHrxA5XKkj3GIke1gnDwOTMXVkksTF0z7ZjlxixGuK3B
GVGvnjxDT2CbqJIsrj42+uQXwXF2VYJKTXD+8iGS8I+3aLOudXSIfODoAYpOn24L
NRbtt+ncRcFqeF/6/pPk3xrGe7dsJfjWeIuuoLOzjoL84wJR6QtvYQeRWm98da6J
AycXNGv4qDnK9mB5PpJPTXNvKh761P1L3ss5Rob9+yFlwmz+ypahayMrwyMIO9jw
au5lwUovQ3yDFlQDvBb1ujN4xmQ+wCa42FPbpSJE/7dCjKjtPUmMw2muzicPTRxw
rw12qz6CDNuogKSeYUFFj7W2lCRVIYvLOJORZJTbbwvmB2pGRbS6d+z/UZPXDKb2
O2K9ZtIfc+ReBnKmjlax9QahpWgFA/IVBvRQDXYBXPaPvySt+gnIa4U2d63t72oU
ZGKez2zfF59IcnpC9mvRPAqpK22aO/FoNFvgURRBlFZTzZ0ClWpMTnVEFJZzM0GH
YBR5afGOKvTsHEY8kyr9alYfIt4M4CFxS7bFISo9XMOFYZnmE8PpopbhltZ4u9j6
J5FIJKyoO/HqfTOEN0d1WTgjdU/hCshfICQ6zKxg7fmae1Sx4Rm73FDLTlxzDqwM
zwXpZ02ZTlgP6jsZxDenUt1uda4J7pOCdt9r84RH3TRoTHrq2jxd1n4UI5aX8tdp
t4Har6K5SUHRvDKuSV9TUQ8fHiD/GBSA5D5KuvKN/Jhq85mLQB4TbJeFjMqxxom2
LxlB1EVGHurYbQEGzC2zN8GqagLL9Lm4T+ikN57ttSfMfEV/+V71S0lBpVlHKK4L
1eUu7Ht1eyShWLZ0mNs29B8+pvkNcu7T4Pgj1DbqYM58iSHa65FFlYHqw+Wh/McE
ow/7UYtqE+vOBLMMa3tq+girViViSHNRgBHWnd1p4KwZjdCmKzYvE0hAWvd0XBTg
2bw9TBdU023DzDcH68gHQevZZrB1QASnu8/N0wiYJpzzYGFI33pcItMOqAPUQNpa
L/5k+JCofYXOXQkSTy1HNLNhIa78YCho0xU6xTfqfrYvNQHdB+B3A1zRGReoTMQP
dNEFE9BJUhKr17SEDwlvZt3s72Wfc5z8CcEY583pRvaqlw5OrpLAaxo+CXCcNbE9
S3cEdARlfTgYvs8ZqstBg52bduB9OcKAudbhvlmS9Aak5wLp5AJPy6DZ0xX9B2nK
q9YClzcmYmSQnpFoENWkjodvR5wOd/CVLIXJcRLjEaRwrgMTH4Jjk+rCrCxCtgQV
vMSlfOoSEr/Hev+NuPaMsSq8Zt28IIbNJVuyDTyeHDcJMtO04cxwSYhob7nLgM/K
fOi1agItTsGXHlTUGnSNcB3MisT75XVauoD+fiyNN8R5Jnbtj2B0TiWTIv9YxhQB
6aS1d8Q3lVm+GEEPXFlqgE+fMxf3LaZrIMziM37FFtZVPg9ryDG/MyibOxaNUcWX
hjbvyp/T5ZmUyRx6kaPoNrHWFu0hRLfLaXnJPe0WQSkOY/wgKEACEFA4iztcvnkP
AvuQUeBXwsSbhzgMMeU4sjnF4GiGfUo1IrcoChemcs3mx5zf+eHawLI2nvmTATV3
NbrMLMSM1jgXEdij7DbOoLg6Debnhy94kGXL7niRpcPnasyurjUmWD5btBJ2wbl6
3oFJafV48jFXFXWJEBVyRgUFnghmi6LcMFJYZ2VioIwnH5ggMDfpcSzRgappdA/n
+bkA5jQLj/N0jNsYws9oICy8SEmsHwHpHaVBh+f561fnWzUT7Ev8uXYdKxTOaKV6
oUgyt/UFTzspJ7mkA1HP8Du/1ST94jQM+fwohtQPfk3ykGau899pljr46JuMi2fl
N+OXj6Lz0noZqNiwzjnebUATeHHIaANcsNFAnYuTKzsbaa44b7bpzl1F/Co20WJ9
wkD2qRde55GFngBugIx4KrIvp2IYel4t0x5pxam1dPvXxXMeTQI/BMJnc3t/T7P2
Jhp262s9GPfnmJoRZ454fUoCLPqsYmpC3MMmi7gr8iBw/oj1A5xI9WzJIrQP9bUj
Mhg7XD+masKy7P1kmsitUTDAYPtJ977h8tEJK+Ca4c12YSOz6YBBTZPYdZeRTGaO
dV+XHKk5MZuqhe8WmDdCey1OXK9XIrJGchBVhmmmbIbcfXQ7Hq0lel1wpAOUS5CG
4ZFJL1YBDAU4kHvdQTfX3aLdmVXw58JB8ra5FHo6EeAj4std9zuLWMKC3FJ4plLA
5RawrVKqDTMAQXuKRZrumP2uMq6e4110/9SxsVc2b7OsavVbUUASBw9SAbW97ZUe
pUGqDpF2j66jF4SH5ErzJZBPny3ILGsG1BC01QH23uXkaJqx80ns89nUX75X0oWf
THR2FI4OyqDhjYeyiel06FW/E15HPX98z7RBJJNlzz5MwaHhRB8I/d9b56ojq+3X
K9O4CrbniGID03oMf0+Zv/h/PBsAGT52tDSqOZBW11q8sQ2BIqhtkoYgXUq6EZKM
ytsekE6a1qRI5vSxzHApczW4+uSlddRvja4JJOQ2Dhifyzhude3UsMUmyD4TQJ89
oGejRtxrR6Eh1Uk1918kz0Xl/IF1bEWswNsSVahFOQgjc63OJGRrJeetQV1CFMHV
xXUeBMZyMJ1PKa5hZ3yLUXbjZpy8q9BHqEH9x8MX0lGu3sT9wKbHeMK1CD0SjNRM
OFtRY2tdOadbE9nf6VQp6R1s/GWw1at5w6gLdm4v38HMrvgnN4kDidtTbm8dA8Ze
fSTTsJ2cxoOo1AMMKUHzEHLvMmr9LpM5GfGckoXHJ2jtDuWGX5mEx1yJbTQ+zSJL
PqpWp6W83iof4gcNcKmMA+9yVYAx46IAmyNFS8M4kBJJtkVvdJadqx28eGh+RMyW
wlwNLvDmgeD1+uReCA3UUZGdWofpRpwdDERFQwYAwQ/oRb0jJjO39vz8B3rE7Oar
l0QmtgwKYsUQX8zvsSKLbkFxDnZb7R2AmsFTB0TLkoSm1g3JfmvSPpfvY+E91dN7
njfmtxLSn+9zdBQTn41QfibAfSu/BR1poPPwWYf4h272GpuQ/rr+OXk6qB7MTHKI
QFLBM67+oaNtP9M9yd6FNczUmBrBdyTOr5LgTH6V7rCT9+eu/BAsXRUp+XCizW4m
uC3+ZzjI8BflwnCg/9GqHQkqoqJDeNTlDrS9x0UC2b22jq6LiDorDYCz6j22SzDY
l0HranEZWO9oTlSfkSQgo1EIzAQ9MDBstv/050NzqEn7nasrD0spB8wX7dFLpYOK
tjaH0GUT63KAAMDmM4uKL6fmmXmfMn8MyGTJbhETy/gsH3Vvm5aRIrQoNYEDPmaX
uRaSBbksjGBWrpoXySUKXF4YhJphQ3Mc8unHdVmYYSlwo1Qc8m8cuVI8HvQ8tHrg
UQhheRZD4apU57I7nWbcOG4WpW+3FtwsBLfNG9bPu3FL9fZ0K+Mpz8Pm+POB7JsD
QaPWYHaGDyGA3gaeP0amKxfmETiRGyYd/qbCiFLeMP578ukSz9WDX6a6MTMO6NHy
aYuCfG7k1CZet3uXwfG9Xc26JW7TbJUosEPhRbimHossvrVkvVQ1QXqsNmZC/FvK
ePDfIL0RgNjyn3kfV3WbnKd/SeXf5EnFg8DrY7zqR++gkOr8bekwlHh800khFIZV
IlUiARtZ8kUSC6LDGd9Ayomu5KHYk0Gv9KopeZrkfTZLw+3a9xPxHtEOjpk4NV71
vl0gilw7wm/AB85ZmQDWFfivTrgFbD8EH7LdJa66Q9h7/6tD8NbampzhDNnahS6V
W9gJZUDD3z3UdjlAIxnLavjFGgvgFirPyoJC2JKy8ZfEuommcb5c6i6NzFFLSElb
7A/gQKfE54ZEFp1ZpU/2IADpziH24vC1Seqt43gyhgUUz90Ko42r9rW8tV6iJxnB
ihfaFdFnbtOikOYe4q9vTi1Dt17fj1mSNW8j2SLTgLSbXfWHlZPrqkrrO+mbqHpJ
brXZ8TZE27Dei7Pd74212A/qLnTd7GZAAZ7waQ5aV9RmIJtIA8+2SEQ14644s5R7
wLTnJh419Twr3HYVHeFYoHspHe9lwbd8ub677FINe48fbyIYD/UHPstOvwhxZTxQ
A826PTsjIYsHyGyrJbJ1TeJYWkj80en9yHBer88zph5Mvqrey39sLNnpmSeYK8u7
xDxDmcLQ91TQou5Dh3KN9TB4cnQ99/oF/N4uiEK4UNcUzwFQ92+7f/mfbG6KGnqm
m0VBsFnY0/Gix0x+6uIQvw5HUA4GdxRK6PxGYy/Hs00uG1bHJNZbxRpQ9jRpa7en
j869naMrZEhAv8rYGQMnuEQTJUfBGx5hr+CX8ShngaxBlx79w+arWsCOGWG2Eypl
lE6p4I/2YRHRjBKXn4FtaRKcLCLdHK6MX6aRVSim0BC+0DBBb8FlmFfX4YN7jmX1
ksmzwuJNZ7lt4KeBTlNQHk+uRr+2OGZGfz5+ivDkYd24Y9CQQDpRfcEV8Z1JAnLx
XwVx/rUMWjhNHgu27Nn5mIyBXRI2bBkAhPaGl+ZYPjGBk7LdLGAvTm19NrZjGYeb
iK7mXzjgIoocR68ZTvdCEFAQ6XGyS7BABrWz/4ddG7dEZcsPCKAih6n9WC3cvMET
yV+ID3Dov2DpjesK6aTCvlat7IOh5hA2vUxs4OkcqPWoe3DDj81O/KRLQcRqZTPu
c8Q7S6HHPKbUSi88AMGU8H2549OqFXu/LnxGF/rKTLVyBuEp+NZ5DrYDPxuNdITU
i9ioLafveI8d7nGDQpLs5UW2BBvoZuUZfYUl8NU0qm+fP3+yrPmE92qRjW830PnG
R7irnDQIauPQDg7Chu7HlasWeZ5XJCzDqWqtByjWXIVQMkmjNaESjVUHdbC6UXUQ
6rlsxJ4DqbUVVa8n4vUk+5095A5UK2bZ3mECYW4IYjDxFGzdh3R6ZBuOIfKLFLnr
LAeznOpxpR5PiYOTtYbYDjWyfrQc7KlCiC8UvGHFi+ulIOhjXyArRif3dxib7T2m
XbVhGQpojAG9MR93koOUU5NLD57omfbzcDqLZf7s9C0A0oQ4q1BBTqkRPy/o4jEF
wWCxyVkggMeUV3vdq4CvWXMbYE5oRYwQ5LKG3yHu1jahIkhuOJpbazBPbMlhJnes
8v6qvkoniCQz/+r34YCKsJqtfvfbeXDggmtn3Q3G8xaI+RePTUmvjXwpFzCVJp33
atLUuGrguS8rxZQl2UGnazbpMI1ZQManM3/S06UnfOj9mF4kwB3ipoVrAi74CJ9U
8+zWmFmBBQOh9okg9rXnAcyYtYPvfUmMQyT1CQxMUX/pllGPJdNlz+02oIvO71Fh
7QwTIug+n7KbtaMLanit55OsE0SF1E1u3L8V8a7CKNeFrojoX4IysAR1xRVxrony
M+5L5X4kj7ViBGQQar2RI81M3BCeC/nGjyjI544qDMpzTxoWdxWnEEgy4IQUOgfL
NoCw0CYGUcFihiyBbXr+URdGMge3VDOOFpDnxdQKGeOTUXtWeFnFEBr5xMFYyZ7J
KBxYlA89/ZYBv5CfkSa3lRPAK10OVsZziKu6DNjpW7HtD4mAAHcuf13DexrnAOKc
chLlk8IHo+gVwWwPq+zvZahgCnfwFwFfgR12wjG/5wkX9rDQo8QcuRYjZDNuFo6I
DMjlHWg1DcqYIKDofs4xj2vbBQPSRzoyYoA+PT9uOx48i04n4wS9YjrdJDxJyA5i
4g6E3d9uR448Z3fe2vjJJKu+H0FNs9jasS20uUBtc0O/Fwuv9O6iHyHnHWQH29rW
T3zbFL64ZuQVJWq0cb0Z5jWfc4Kg7fHNaQOHZQl9sdLG0K7scBFT4s5i8Gii1cJk
5V5bi1/v6ab8GRi4XWhIDxvEAakJ5RsL7aRjdvwRBQVa+Aq6jRaH7eScshj6FtiH
ezpq/hbzrqPHm8ywXPqFVOX7lh0pH78HmJbL0mAjH2a1jXZLIVRVHZOmwQ1B7hxR
tGun5O7KnhiQSqegAgAl0r56FSbUt8b3hJH2ctrWFSD6NypCe9+wwXBfWEpemLKR
BVZnjwRj4YQNffZsjhPbI1cwhblVBLkbAMLx6Pn3nHj2feMrKmWm6I3NCoU40tuX
sUac9hFpdmO0oX8J8lR83ilK1XEQosJneJDcppDzlrAvUtnv3WwqyniPyaIBmy+P
5iJVRs6PkhrD7BQPejatZ6Rxzob7YiI8iCAsA3L+FhqOAWcCInEp8XV6zzl4TtlA
aeMBLPHNxifAa6HSJoTZHXV8+535bGf+1UX0n4J/fqd7FT6knOudCoyZzk1cJ0R1
TuzOrdqzsv4mMK5f+v6ud4fuzxP5f6hXQRqAYMAw8vrN6a3j28WYcsjKwCx9cHpS
Jt7A0+UuZUTH4qKzgz6BbHecCv+yX83S9g7acAfVwshf5//du/W+bmeoBWiZBsPy
pBjd8vMG3vd4dztkKO5IEDQsKm7Y+tG17nmjOkvE/NUah+nY6yvlnLkHkNNTWWTk
XqBaF5bw5A1LK1+ozNtJfXtKtnlZ9pRMejDWox7p4qwF0gtAcs+cP9Rk/LvmqBeg
s8A0luBzdXzzkK0rr6HeaLHHlbiuEbirGy1CeJB+g2w0H5xFUMMhzobQAs9cz+OU
VDspWH1h4njvyZ7CKSY05fh5MmoZmnuhKNLUMJhCAuHZM9O3q8A3t7e5Gy7hklfG
49RQzeqwR7kJGOKXn6eykMZicHMEmI24sNbbhUsI9d4uYlqRxaXP5FxOSnHj8I4A
EIwmei+psXS/QbF3F/9J/40e5NcxkaMVWzqK0mpxCE2iIdlPKm4vBczHGZKsxC/m
HuGJLC3r6nadqDolznNUndcDwPxltlw/EVvqCISAoKSYwvZtmfvDAjDjkS0dFtpB
k9OaiGcWCpkb+aFGfJyocSVPWJagp940nwl68JuBfSSWt6eNuIoPJVF7XkebhOMk
lJ3B4Xezjel48IVxCsYlktJQVxh0ShuJwo7eFbkep1MubP+6dJZY36LSyzH5Wd8X
PFR0QH5bT7YADmrFqPyEMFzFX7SyzY5+O1lfR857kHKBlmXQM04DQQsfEyQuj1z8
RT6HuvAWSARKIU069IoOfHsM6pHG08yzont7qxO+kkPdbQNXiAHu8adj2FgXG//l
A8vnIl8Z0uVVJ5MuJTnkGhP0ZD2KniXlUmMP2LByBs5s7CfERkxKNUhWXKoRBEwH
pZbisnNAyW/7qcgc68TPBjykAFnmNbi4XoFzJbrUCmsl0uCtBIpOC5WWicVsaA1z
UUoP/95avZAzaTSlgU8cA0J1DK3BDgN3EcopYap1AAK0sFYdnIJ6EuDmPE0lbgRI
kf4i0Tr7r9Ypk73Ns27LicI40oQH0MOSORXTJiAMQm8uz6PkpixUT84FbHjroslV
5iESB7wLdt49G95NldwL1Y91qtL1NN4j7dp1UZwf4jzxw4/6Aep0rkY3hLh/R1le
DsGekQ1gmqjC5Qfeskk2UsQYawDJtQgwYEX5U7KLUSgOtK3lh3gRI3mPe3xUHz0f
K+sIuF80rwPeaIa0pTzxcjHFO05heqVm56LOC4cePMKb53RWNY1vTR7wWRf7axk7
wYgiYuqFlE6Yg7S6sC3ueWHrK6SjRQx4nzkavpCxSfJHwluSJmY2tEKvVyUhta8b
x8IDmBi8ykltzgTSlrUnjJe3yMvYpk3hL4AAUwwvLkxYINrFZKCU9ZtEh402jM+c
U8G2tMF0wpmOrJZjn/WEAteh3Gk6t2bm8470hCLpKLerlKeVMSSLWM3WRCKMSLUT
pR9CmfBZ/afD49k52Fui98kXbvqdxPEdJvk+mIwi58c2NK/9lVcFZG0kIkFvSdGE
G+FtcXs1Hf9JEF6KjXBjPLi8ml0UMAmWqKKt5dJl7uHI1kL+Eq5qYaGhhQCXVa3v
FrCyhPY8m8BdfpC13YGWMC3EG6reEqYbNGVug1aiHXOQhZ7qsUnJtj++FCZx6Yio
SLfVQUYsJa6jQeSUqTdNKQdNKZMUBfHqraldtZTMvgO4wvu4t434Xp+ENDnvu53+
32fr3orO5zrXfD5hkcTSnD1Ql8YNGT4t+5TjoeIXiNjJXo7Vuy1Okmjsu6X82bHJ
bkQSU2rBHWieD5uhLSm26uotDYjmHuJ9jdvo98zOKwn0ls6slI2eSbCQWRzirCpU
njpKEsKs106EiNmYZZfY7Tb4tlPWEUlHO1xnSnukC/203mbg2oIWaGPHLBF40BIe
n9PqZHLg31XSQ+N2e7c65k19TegG/iId4rmMIxCHSRBRvMmr5DwxS5AeTrr3O5wP
OfYXBGcgVdYOuIb8mPL8k7fvkAl7vNEhFN3qxg8PxrW1VUFHSruFpk/T7FZo4uLc
7WUKSmOtywtgkU/g22gWiT2Cr/LSSyStNh/rm+lLH2fxCInd1xhtQcXlKMP1Q96w
s82eCNmwR8va4jpqs7B4EWDWs1C0havXOeAyQ4cVesf72FaaI2Uit0c7eAvca3nI
N8+d24V1fwt4U4EzN5WLdaaUBP2pjMTnOoJvWbKOIsVe2G0pfrWu6Vx3wWp+tCx7
XyUwQxR8JilXlQ28qjkUKd2REHJyUQwPgXrkrif6eqsGR9ktFu9x2rJ7/Zvyi4c3
rhbGWFUNIa5ZV7WRi35x3nKVSCeqyvT+mYY7WgnHWeu9fkXKUYePkt16RYBoEMsa
IhuWvIRUT7fBtf7BEkqujGESzf3j+LulXh09CbA5aiw94Qc1WSgOpcfQo/dagHr9
CXFs6qgvjt9SBAQZ2zzlO13MetGHP/21CWjX/I7k39ip+ciCnvR3Tppdmav2pQGJ
TXygPtwP9btnunZ9yXRk2CJMrtlAwZh0s2mxee0c/CTp2F4M1sGwqVapbeTRpdgx
2+vKV2s39B0fZAwgg53ez3KNjZhX9LoZzGYNiPi3ELPifsatPB2wX8yJe+Ht65sc
aAC5SR4ACmuMmmrdOXJTIrg6yJ7xtNzYv9RrmBfEnxrxYRlZXp5aiBAm4pUjT0uN
dudw8ztsdNVcVqh/UXLaQrnHXE2ELfGuK260BvOKqJ0hOvefOaO369r1SJ2/oYs9
Y7M6zHZWQQsZXag24/0HI+FlvvHmHOOdjLOHFy/mAncQxKaia/aKurDKtS3Fhf+z
GTJnAHpmbW22QLxMZqQkKfKYLXXXK4+Wq4TRoSSAP6HUiM4WTC3x6G4NS07FFNZ8
qiTPSZX3Tba8Y3xt8Hfv7ew+LbtnB0iUYivXng4wAa71YBaH85zIFsS5lqyOduIE
GLBe2/quRiENaTLhPTqZLYqTNqnms6zuGSdPpOssd6tgmK3zZfb6lus4hN0CdgBo
6JvYSEmoGwHaq+pmYmoArYD18QGW9WfhL+kppiJ/pfQgpOuvrNuDOhsQZ1FChlKZ
XHwm3cEk3v6ajNwEyanfgdFU/OWj3hPdg4KMQDC9BGrd9O2YFJCxVh1liS0AgBEM
aeufeTH3yLUfabl141DXDlfKrdsTX5nRuylNhZ+tCs++ylyPpWz8ElhZz+7QrNRb
6fZCJ85bIomffiyJPef2FgR9OSjZRscVeq9yN4wjvrqUXnL26cNgidzJmsLZdoQ/
ZaQoEMwGCJbroFJ9zOKxIPqZ5prCJTZib64U8cUshnxp7aiK7ba8Zbrgnna2RFKq
ABKpG07B3TWwOXjgswkDBvVT48gQcL4I2NYcndoZZ5v54Hy3vVhfgUtWoPjWWHT3
WJj+F/0GAvliQaCuwKmYIPMdgMuZ6d5xiZp7jAMXRMx6Sy47vaCQjq+axeyrruHI
QkEkSrBk+e2ceEDIuPSoJV9xQfniRUDDX4djLlzqB17dJgRZx617yJU+bk4B54hG
2mgF8Zm9Jxd15BwW4+MsO0DMhgBA6xmZgb9rqDAUVS+j4uR+ztZu7mbIxPLMsEYR
P5/XTPgO952frOx5uUz60Vj2W/fNPn1m8QXrPnAmszHdpNwlI2r2xyqkavud3s77
IsbbQOxX8fjmPcFHv2Uow2QkM8ZG1+Z6PkJL8B5g6Jq/Xv8mW2CnGe46E6i/qSmR
2/ccjCkkE3pEZ6KF2Qjw7eW3x2pLV9obXk7XxYTkBJ0YXQ53CDrYIybGrxWhm5n/
yPvA4yl+cKQBDsPZH+s7wXyvoGX3IVZN8epbXl0VYh67EuzoEK80TjilOdk9SQba
pNkeFz12azkXL3hQbokw/NnUvIOp7ro4SuiY9qOAp7FpEJtrq2PFaRAvXHGbedls
4mqXhercMnpe1iqDiQ7UDduhmN5zgxZwqMnDkfLzGIPXefPrijZbD9vjaPUVW/7P
NUryaAOlzH+TNKl6qDlyUOjO5Ni3UsNYbEDRkr0BRaQU4EQ0SrnTsLEIQjDWXEqK
Aj/kujv/QkjyGD4hejN3d0Lgg5J1k2vVR9U8ioGsVuTwktyvedPgNXJMFaf6nIF6
8Uq1dN27KkprkxmqzSD2jiazgYRbDs8R9PQ3AXX0KArK24qSXfIbz9EbpelMB/3E
6zZJcbjbpy4FS11XG4M01My4KofgFEMKZtpRTEu/DUV9F3IGfE9pYghY49ajnwlY
SrkD9dQU5tS7MMKPm89uE9tfQbG4bkjQnwpYokLh5kozhA8jkDqAxrhg4gJkIi55
USClVVRZ4aT0AaTqx3Fr62UJ3g0kfagVAWGujCY9+rQNYMZdXjLHEar0manNptbM
/nkbtWVLZKLgCpJXjWYQFL7VRYNS5bhNAD86EaoAi2IqM8OHxV2a6omcjsNeT8+U
LqUXfGdS6iBYJH0W9/6S34TDBfAjJosrqfm/btKJ8M5G+6ulvPJzVtWNORW/Wutr
SxncctaQh8YMh1c37kVXDlIrLw45XgFlCM22YZ1n6RiTV/oW3dN9+815HAgB/3G8
AdG1S6qI00eMWdxXnK8HJ+CbAn6CDsrRTkCid/YoigRhrhcmm9VvLCvYkFMy7Q75
ateVVJXayp6U8o69oHDjQeu9MEBvnLK69fDAklEKjGG9NMFrQO2wbxeIJJc5FsmI
5AFpoejf+EuroZq449L/2E8ni13MPDidcXWZkMBpZvH9JxHIctlfqakYKVFycvDO
Ls91xsjG5KTAVFdIpPNWC2iEa7WMlujw0yrkci+5FqQ304Z/BpPMJdtScoxgVvJI
Gh22bjJ2w5KstJE1yHRVBrnvxBwIOWB1JJMp0E29G5HFERmADTk/UWqDXLLtfcYU
eODDs12fNDV+wb5aaCeKiQsEg5VR5FF1l1y9R1/tCH1xi3+5id7FbRJdISQHZ2/Q
9RtT62TQ7CAXVntucQQ9NznArCDOF5TTVnUucH50SDRLAobqdR9PP3LHg7K7eXzv
jPicP78rgUozO1sfoU+x3TN/GVZ+oGLmqaBMY3alHGg2qVp4iRH6I3YMB9s3HslS
9D/q3e+DPLBbxCoLH8Ka8EXwoyw9Czmnf9LZ5QNryIxbZn4eXmncy4zxEThiMQ6j
6BnfhQiiWTXlB1c0FHPVZnHocx+TdTRsqjarLFNMwjj//NJBLblYcZxMVfVJpymH
vMHooH2BmnHW5I69fZ8odEisy+zsiqiridzUj6mF/H7nPeDkmiz1Il7Pz16ufDe0
6wMQzKbOkPDlor4x2L8xm/CwZrqPtnnvQ7qpfaPl6v50fx+7JzjVAgQLQnVxTMR7
GJ0XCu/vgkGsZ/i/EFZ7ThwRCOsJP9yPn596DRIojlQVV54M/F1w8TzqekBPGftN
oWYQGaPN0SXXmc0G5tnEii/XD+q/GukHDJI1JsXnvs3SpBnywK20WwgheaxA66Hp
1qMrjBEq8JDQOPPg8qqUHP7YO9TBdm3gcO+TPDN+HE9Y8+ETESz9JvqkhJu587C/
3O9qhBw2bjPTbWk+uJfkP0QNchkOjEpfQ+euZebGFOt4Rov927iRAFSdtU9Sdi2E
p7bcUSC95+CwbKcR3P9aXs+JkGgiEF1LXs44Ch8W/hdQkII4vn/Vl684iUVVryx/
n4KTsplc+6Yj71V4nAfdyH9rh3IYFWuKnqdLTRCs1fJcGCN/Nybx4e+E6zpMip6k
9ssGkPH3aFs3xeB+ezdrDB0VTlOM+tky2FDxqIqFqit2lxBOuF/kJAkAmVeXvkfO
hP/pQpx6BDbMw5V3R+U4qygBrQnb9wav1hc952W1G1Uc3Pdl8/AMRVN7Q5HBuKL9
M7rvZ+9E6Yjdi9wUfAazlUeCRafhiBFR/BXV4e0v1+8ULjX4QejauQd6NVVmPQwm
EFy6r3KPRSHRXY7JtA00u2nZ3uerbpOtfAi2JUfc6Pz3s0lDQ0ZAfivwes9ngNM6
60ZEpOgrAAN5LAoaUIXiRuvUJf66PPkpeQ2JJvkoIhvJcUkjwpttuZILYYRbM+wE
Tz72syRFjFIS7hNR9jso0jGAClZkXK58293eUK0YDunjuoNIqJWKJwqiWg6zXMhM
Bkgy86ptgWO0vCE9S4+CFOZaOjxWyV8tthsgYvnL3hHnJmYnVkjQ7A04ioZlgkj3
hdncolUgzTkO4huo3vK0CnJD+9F1t6yUYOU4nQfT2y4bMmWgVOYjZKXnWMb2ZQ6L
SJEC9ZkTJwRUy50eyvxHlyRsnEQ6haFdN31sBaeRHSl2ACSfyHJ/nOaP0gd9QR+2
w/CF89IAMBHBaND5i0UM9/cRE0yHZk1uWyhbCoI1T6R6iJBxFJUJZR907BEomJzb
jkaWvcKW5Z0VvsA2e824iL50oHrDSt3KlIrJTBSbYEGZZAXtJvgGyrMRRHL/QZrh
Jtidfe2UWFc0FJc6EkI7BYMWdeC/3V8Zz9YF25ud6oZRHvXUF6XytA3/J8KYwW8y
QMLEIpm1gEKHAQklhIUrO1P/NH+PFlh4jfmsRInCR5dp9pyI8vFEtAuEIMex6Dfe
n9dBFZjAOjzFxFX/CfCMeOdiK8OyAlxzOvSD0+dNA5XE9CIMrTSHVUDNp9crdGUe
HtfSOZbCBkVNbTB8fbIJ/GmkKgLCAK8A4A4OJwOw2fg3HzXqPxG/sNDzR/TlWxsR
9/fbKByu1qhIWzPPPP2QYA8+DwpiVerR/u8zsitF0tdk3EvsQbfCMBtpVEXkdzKV
TDkfNF0Y6X0/KNDdvmSFnqcbj8/RmmKnVbQCQly9uTrqQL6xzODO+/+Z0RYyXyLB
iY45A+HbP9gbosTg3vbG2X+JhsSAGzZ+xuRy0grwwqvcCAuZeBXB6GmjGmAKxPg7
fnEvD0bBiv1HAn36jatGJgZ15kDWQNVa/KdMavprmroVE4pZqrSCPNR4VqRpC5IX
7EEDMF+VW/HXirdVfLuv+1dykthplXKINh1brkALo50PccRoMFuMjELnRTmDD6iD
CvCX37qr+0rsVIJHicxwTUpzgfjtzR/mprtmgyTyqqayDi7LFt+cqcfiwLJw4NM8
tBlUahPm0Y8H9HA+wqmyLnXA8Col/wnecA+WzurO1YJ49ne6UZGHXFNNDvzjm//a
83CgO5iFIjug+2xhKaCP5ihpXZEiXb0q45CGu2YT8zCCVAm3RUEobL6X/wjpQmm2
pIAUBlOBp20xqIRKq+sobDhyFP7QyMUCZ8X5nXxIuSV7iTeM8cjSF5d2J14nmRw2
UHMK2rUkshxjGquLD61OpFg+2v5d8VUZR/+OR2C1c39ieMIYQpcdypseB8hg0Y8b
cwlkk1AxgTyrotKfLja6QhgzCEFLWhYH0JLW26Kl0A71rv1tnf0ZQ0e6YdDs8d7Y
PovZix2EoLSJRT7OA/JZiVA0f1AM74svEW2IsLWoSVW/5lSF9OJ4ZcpXVAnOS2HK
wy9qtRy2p4w5rXjd3iMX/CZAmjv12mMaHhB1kKHoIAHI3GlRselUa77S/qVMx8zN
GBDyX14P5hNT1/nAP02ZYfZ+PNPkfeD7XD+MkiyjrFRl8Gu75hj7wcXd81v3a9vv
oa6g4xjJb5hxV3pn/GgfiBmEojIMzyDH2IfQgXoH/vIwdocwotOgBjU3qSDhqmpz
vVbVRcQHWnDw3cH9wDLmZz7PhsfOo6TnvUdIJw6h2ZIkIdGXxhnOW/rGe82c5AfV
8AJ2HzdgOFXVMVhkCjW+P5dIiYw7Kcq7XpQfo1BiwgM8GLjmePLWyUtizddxDStV
qF7WtYdfpFgf4RDsDazuwYULI0jaCbiT3ldNnnkjQD4K2H7ep/GYQMICDh7DyU95
gxnguJ7+9hHNZlOLJxl6ZG8pKBrKxj3kSHFnaOyPN6bymK2LAKSVetlK0/+Pc9Iv
2n7DaFx+ryauOsMwtOosFFuH69Qx0ADGpcXL5vxM5NDTy2y9nZZvOaPH2Wv5LxmO
cmNSMpyVdNksVz/KBJBhtzNDXbkXcJrsePun8B6u/CL4lccnlutGwwjO+P2Zlelu
BoUJCy0Vf53WEg/ljhyIrOsFsKXVLiUe3oOfjJctrMxCfNQgAMzlsfG3lPfG9nlL
vxPqwMLDopOsGXVsoiExh2/o5FJYW45VzsuOjGLDtGmOmwdTgm7uPeItH1PYsGft
IWqZ0NSPOzcnSGywiP3VMfp/EA8ODuYNR3RU/rdv7wHKEh8nX2eq8PwV+FMrGhpd
zXM2rQfzuV+Zmkwmkik/NNIuM0W96YbYzKx3iu/Kf6wU8v1KGgV/kdBXwFZ0Jq39
uHyWR5mBlqHNfAKUmUdMFYsTQtUm3PliGFA1oc+0a8Tls80zsTCYbiNUJiNqBk29
cuCU2iAj1/8zJdA2c0PX761b+Goio8PiiUkagg8ru3DzC7AVTt1vQiWwOadJT04b
ntfdyE+S09JAcc9JjhcM4EakvgigAhiyNFkYdpPJjt5ZuWo9OReiezRK4NtjrLfT
9H0jIQksjVW78DilDqY22WHxiSmJvZkeOYkTiKTQHdq+s3PNimbcVTCwBHNzalh3
7pjBqpc7qzqMzGXrrOcDQ4Jfz40NgVCDIgFwKjHdLWHMEQ2T4SKN0nMjBYaSOFOP
rYhMVjoB3k2guwkfIgxJ8ZlLgxrGSGofDci8Hl/0KoU2qI5DVrf8EFagspO5h9gD
gwaeaLG17pXypHVK8WrckVlcjusJoBmT8tbF7NYTSc/TqhT9VogEtGv0IGFBnW06
Z0mSFlSUVJtTr+baM84tLaWSYMtXEpv6+N0CzDQBBkPqQK2WhnTUaiHcFOWkE2qq
1GPLZtZa1a0t28kXhyA1PEtRakGAcraS93WslnxhuOhqEZPEZsm0NK/6Y9YGxhrU
HruYN6Yejg1Q56trUMFtBONu8bYXTHA14R5xlU5Kissv+EajrD1eIITXGF3wQZ1N
bTH0hL3tE5lLWgAsl6N9qy+JN8TwueHVK2gkwKjLPpz/fyoIIjdCLJLg0oqvgHFL
M95aEzNqhvimUSdvBUx4fmGL5gcQq2G1+uv3Bmfwb28c2w4RMACHfa4t8YkmTtNQ
YLzRhOXjZ8ei93yQQIuPrqHkmS/eOL2Krndmu4LSjIJHd2UmMSlFPk/cF40e2BFK
R8Vp4yhcuVJmCReERyRcThXhNoGIp0RHuCd80miC7nHDvwlOSYdBmkEJrx1QrJBq
o3XDRYWqzy/4ZDBMIhe+d1kE7b1tgm3whmdkZClkhwRpoDHd7U0goDtAqmkkRgMv
znGqF67H55PWmTn529oiPMjDHmgoaxpTUPYAgrij6aNepBScRZ7yQ8py7x4MF/lg
M2zt6xBOkfzzx/aS9iK7Uiz912/GDi6rAzZyO+4iVf/TA0kFJmeeo/5488gHQN3v
8+XgoepiIPtOwgrcE+adpoaN2OblpUuXYQK1AcrfD4PXeX2hoNIhFk4N4wApKkbr
d4dw4a1XDmnwp8th75Yn5nP3GRMeFtKLmBEoueu4GYocx5riGM15LQEe+WCaLhPF
NJJFveXBFQPMuGJ4Nb6FseD8WPwwKioS0vm4t03Vqjv099k1BtPqo2x+rXS4556m
Ci5emGqx50aYz2/z7gxxgXGse4VnHEicMEKcncq+nufV6TpwnTvIjkCxU3Kqe0EH
eI3sdXLDmpak6dHgsc2516yatrGdkapuJc98nPuY9xV8gsMehSNe4W2tjgo1Gy8D
lsaklPtpBKX+kmdqoKhlt0dz9h49u+RWZzWaPS+vBaRIriuwbeNgHXO2XUmOx0Hw
wxT9TxkokSRmbNTToyczjXZomL7NKa8nIbfZpdanBrZcfK4/gRNrcjekqT4Gebuy
Mr5KPLskc+oKx8X9qJxwh2ooEFroWT12GJV3Bv81ht581PM7Fr7giilH/zNSVeDi
b4iPTXfiXqc0zXdY6QdqHBCWLYMiqVT2krE2RJSfVbrHydz9dbrI/yv8FqxgKo8P
CeYz07LmxlY6PXQnbjqjrsDLJVMxKlbHx2D48ODsOlh1QuUs1UO42KjlMxAVHPMm
Vl8zVxqxvcWK4k9cClN+byR8kEJARk6TSLXJ8Ec/aM0fyuWcTP8pWNCambIGA0zI
JcxcST6JinjpLshbMJucOa1P+K4Cm+X4ZzTfUKLcXizsSMVbSUyuLOP9np/poUh2
OWVSg4VQI0Zc1tNyVW+DAnxsLBLoa1ec8H71YTlveC0Isxallk286MFCvaRNhUW+
gx6Xi58ymDcCQd9hkErwOSrDcZr8f/p0Q3LqsdvZkI9uL2IiI5BE1ZxvMcvVnQEf
n8pwWf+wqdsbr6biBhCKrpUJQV21Ge5uKCwCQ5Nu1t9bJ90Be8oFgOSMbkhATTdg
0hTfW19QU9A+ohjAFzms+TlIh5oBN9V+fEbIELDxRaCkY1HwaIP6E3+EfFmHg7dk
tqJe7cG2gI5mxZ3Fpg5qVprZN7C7GjmgSwjELP7dLSIFVC7117qHIT3yjvJ/Q8kj
JVbd6PgZoAirFAL09le7k+QD8gwdDpwxNM15P1ynIPeZtG6yZaqG+uGr2KTHl8rh
choHUv32DbV7B8DeGoIyyFovFHCvSuhk0dbN9TBIljCx/O9lBpUlyUUwqErnaJse
EM3IvX8NGw+NS57eC9FPuVVGLHEyoRLt1xMPwAZzr+F725DMfEQyE9AXS+jszDeT
zx/44UFa/tS3379j+N9VAHqFuOi74aQh5K2KVJ7HF6axmkuqOr1Mzxmm27s0k2Hl
S1rqFs8Ehp78tBmS8m3lBDNUA+kYnupnK2NTqTA3Pu082FQpqfMNo1c8sJw9dWrp
GbkeSReLGUpNjZngXgrBvAPebP8ZHnq35vqq/TRNhdtgziKWliWQoMUtNKye+b7q
BWEyTx/ybu8X491yGifBiZcEYKAjaoj0+Y8EqbKOSciTJC7S9MpRpRnEyqfnDY0m
OBt072lbMAkNd3bFGrXvAB0KVvDS2tebaoK4D81rffPa6cabhDHd9bQ8i9lcJqfh
N7bddxDPU07Dc7ykXwqDp+0kssfTm2c+J3Jh65BEmc9nAT22FNPdRhpns1P2r7ic
Hl4O0W+wgLcNgaPYGqilGVyZi3wPbiFHJV4URonwP9ucDp0uaRGkYj8sM/QR/N+5
Yr+qSGm1g141tq3C+ixYVfAHpzDkPNMy+qIkUt+33tjc2fFXFH1CjhWlGZpVakdG
691ObeVFSK1SQfaEadJVFc9I4fl04dgsBfdkpB6EZ2IZCg3GlxUmfBn763N8tQuU
GfPWSRlXyT3ODkhNnOyltypjz7k/dBHVok+nPFGNC8i1kTJIXACEcPGesd2t/L+u
IZeyYIUO4Ns5B0i2sFCA1hDHG9l9SvF6tt8UPU8CC58KIFPAXyV7EtTmOeOgAxch
I09fSIUhYonf2RDnelTCrXzt055J4iQ9pYYRoy9uBaTyQIbqcyICQ5IMijW97lH9
LkcwaCrJzoHAMsVNOMWQa2Va6GSX2gxHbFG686TIU+rAIHNwvIKKp0R87sUUxWPe
2ZoMbUySjwBmxxBFUBnwgl971UZCOLibK0LnSzGfVyLf93ek5rQgHBJML5ycDAaT
8vYjg1oGVhEku1MB55quURzJPWjBGtD0WyemB4NIy0asOMYKfxN0GH45nwyyfbjK
86PpBJvjrCch1SK7wpb+WeJk6I4e4idpLWMeaQVH9G5QYZZeCOEtk0VKtlaUhu/G
aTdOkQsYE3G2kYRMXx33tyNiOuOurJdVbqLp6jFSGsfBUjCEXuvXY9YxVVkV0pvE
XfYWTg12gE0OJODz+c8pe8vrZAdmfnKuEvihuKtwlXe+WYNTY8sNLb2iQc1n/7C5
EXbDgVzY4Phzcuaays5FVmvp+//dZIMzHWms1s3X3hdUkSchcF+u3vhFUH11bb2q
wgzShSvi5I7JcdU4p+oNlNkO8fRBaozcifIFoI0hdxmHceGDRFdHHci+jIdHFfPg
3rAXokv7KUet37c+LpqzqDCjYJxSE9Xucqz4AcgfKtNHEu0waJbJ95p1+jpepvaD
TKFAuzJXoG/W8N1RC5DOPo0HBd8vr7h2VyOXXidRt6xAjfxggHjkAh7QAKLfZ/54
Y9rjUDKLg9RuWXS77D1K9dgmbtU1H+F9LZovG1VW9ab4lWeuqR/4OIcT8fjD5gs3
i1dT1lhRp3/Dowgv6a8QQMo1JIEhrxSHLwnNzJyFjR8AyLG3dEW8cwgVnNPidnaa
zDtMABZFkeqkU1K46h++RuwWl0IAe75HrK+IH4x+1kNsdyOyA016TUlk7aPxl5eP
a4/cxvB4GFqqkB4XiEZA3jNH58s9Z/U0g8jeB0X4cUTkn4oV9ZFqN57aGJnWHXy3
hSOPnCG0VE7sSFB2Zd8qKHgGkZWn6iWGBulzhqNRlRtNeswXTxcw7JAZZJqtk4W1
8/e08GfUi2O1vq9jlXR6d3XnZ2TSMtKjuRuIzBWGwHr+Lp2B8VhoFtkZO8TjBjp7
49YEev5tCuosTWySQW7Z00PRyAD0obhQn1Lpo08Ht7b90DbCk9dYm2qTtcMngKDd
oeLZjX4E7xuT2EZLbHtPslWcGHHAZl6OaLEwsOaKnScyTaTZ8BznrY66fKbMKtY6
0Nkg23v4hnLMc0l3eWA/2Ygy/KOQUtDq+rtSqkOvgwPcovtVznfE8QVKq3Ajux/S
JHta9eTEhEEu/bpL7C2oC8/J0DUT449njQzljEE7D0ACGx5QeyG2ioT2wa4Tbu8a
agnkArQtovzB94fwU6N4gSoFoAkXqS/451YA7kmbSt0lR4hXk+XOQ+mM10QurwXy
CzSgah98uyKSANRV0g181mTypQe42yMSUGIZdswEyXzgadNkCgxbqU/ooJUN8h9R
oEQAInvzw4axR9ZE4TzOaACSo5RA4oh+yhdrCKZYO744u6pHY0Ta2uyvd6ICqOTp
5lB8JjP3soE4OUOPgnjlAtP1/tSH3kQ1fjE0MRyfotTkXdjOZ9WdNAHn7iVhrPe7
ToGNcHLN2OaxAF/nTlJfymIJf6aGOjRbdy1/2R8EH+cqyU0pX0mRD0sAnR/p1rlH
LSAp/1ruGXiGKY5w/aEuln5xhz/f4W+1XqGgyfdtZc+W4fYPIBl4swkyterzI/wC
YsfVO26sTCaP6RACse8mEB9Tzdndk9DgtAO8ANPYHU/cbzgNjFo5VCsnZK/bMwgq
Mnx0czD3Aio/UfqWfWE6uhMqz/Aka3J0b9CEtj9ivAlN794lcBiUeH7OnUmxxQI0
Wzx7R0JsNe4weUTstzUOHbBrFvGzfHqasvJG2iVCk5IybtQW0xurLAevzatYDlPt
HOHbfrtOUOuOC8PHEvCCPR9FPqA/63Gc3ZahTzyyBkTcJ6zbvnTDSMspnGoz0lfL
/Nwev2mibJ9IgdjfwmVbVSfwzmsjJI5zSl3OFQJ81A+lTWL9JAZv3K6pLk9vgCRW
oyhV6a89kqJDpFP+Cj1htgp1XbxbAvLCXB8chjDDUZFLceyEKqqgLF63V9jlba6X
lLR5ZnDncg3pzudH25aEfgGUzA71Abd839zxP4ADltoT8s3YeC8P5YkrHqC2LxAf
uRt8F1XTAsWkzJUYcuG+2vqGLqKjczRMTJer2HkiWH0gc95SR1K0oISVf8diwfYW
F2G8RP3M0cgVXxX2hoAxs7dIMfwyV6N2Tc4BRsyveK5pjYmc437teOwMAflwzNkk
AkTbeNxbw6yeuVZtQBRA0v63PoXjHs6lrtcJ0bPYyWozoXnGcBckK7On2AiZH2Nq
WqlD708iPAatnVvDqGOn6j8DHaRsI1cEBVe3ri950d+LzljtrZ0FQKU+TeovRNjM
b1rTz4qzWMxq9WD8uubruxLySnr6/BKEAGaHt8jps17j3F35AplHcGzBCdk9/F/f
+wrQQBU9qL//cmguFqHVmq1UbjeTB2+9cqwC8MgvmQfTHPzdLSzyOXhPAx9NZR+2
G1Y75OrdBAm/axNpaY/oM76t346vClzCecvX8lQcZ6f3RNXYmb9elP9c8n0bhAhz
r0KGmnZvpaG/oxiuUkYkJ8YZrpSLDvc5WeE4JNpCdOnIVmYuvw/cTP46ERMl1GgL
l/Nx1yBQhqZMxBDD8MDsrU3tQVJzbT0pivxbEe0DX8i8k7eT3SZghfrjsXwpD1OW
trfnjqWiOfJuuST+k+OQSVx3GnrnNhPxfG+WLB4V4ofLsGHSvWb4zKnBpSUvzaF0
Hy1DnaZ7AFyH36qx4lElZyOHPIadRBD5JYm1fRKJmRGcKA2mTcSk0Tx3xEewqjGR
zF42GW6GlCFcPuMKPqkP2ScAXyRD4teVnhu2DR5p/J3HBtR8eYpDQrzk56q6403K
BJrMnHlnY4oyeS7VmDoheqTDiDiRLx/Rx0CFIB9R/x+zHDrjBWx5xJJfnEN1mDEm
IYBnkpUwo3l+5jfyaKgJvRXUcmM1r8Ah4XJ3ZwWZmBz2VYe+gJiy7JpwhX9OGQ2o
HRjiMn7d4i6GVeq8zUKk/dpdHXv/JFCRkTm+0sJ1sm2ozQ1YZKh3bs323/MoXia4
lYqkqIUyIk+rc5wkpsEgctNhe+YoT/BLwxUdayS7Fz7do57aEqwFAfgndAEUy5St
2oFCrzO02bUsJmzEmTvWlqazEGOajz8d+/MIfGmeB+bz1tpFPINW612K0LUwe6Yb
cAS/ZNfpi/t+P99955Kq5+VCLVtndpEFgReJgmlU1a2N6XUMwSR7U46c0WyTI7XJ
hu4xEyR9M5VKCLa0a1SQLtgKKx1qwkjJkFIgjQWbN2MRJZY2j/6Evw/0832eqQgt
LCfhELMmDi5wOQTv8QxlZY0h9JofzwG11ARvchM4Bnh5+uHywyYGTTyNvfqWRhby
LjqPTXRYFpYNA0PgmSknuA6tffcXMduQr6ZSTBoQXP0sf5144tQDcFeLNAPTaRqD
Ycvuj9jGgJviCyHT7Co7GoF+dCyKpaf7yhgGi1zvGDuCKrqkWQQqfvpF7+wj4ktn
QsL/C9taa1K5TRD1jxa8gbiaxoloLr5DGOD14dzn61NQ3twRATzG+6JKtsVgrsg8
iuFqNh52eiz9anqsRyM79fEK1tzpfPbJwYXd8ErfOpTbyWwyRgnJ8nG/Spt8mL9L
I9Vvpk3MouSE0NvzWB77AKNUAqV/QzFAM+sHyyDcq2F+4LwXXuf3PZjhGbPVV8WK
pevjjLRz4dOS6D3hvvyrl+/2wZRgaRotNTqrIvHVerfi9W/EpO+COCMf7DiELtWw
Rij+fnS3kEHodya8aSK3GRvg9IH5lxFqryXZYKJtKJ8/4AXfSj7IwxJMiu9sLi1a
6VfY7qJxIdakpy47AUbzhz0x6znWJC1aEB3Af/vgrRlNLcATB4Q83cs7hwPLr9EN
0K/XGb7kuWfPZh4HdfCU58KAugOc6onn23Zmima0eiQU6SVEvGZcxZzBDi5H3piW
PKgwMykYx3+0S7OZ4wCO2zUS7SKm3l+/4RyMyfbSYl0AIxAwKbxOcDKtyz8lDKEw
Ygd+gOZItc0y1Xe6CosqOWMuXQiOrD1JKNlGvovGB3PVbuguaK3y5DImYMDWRRxG
3s/07TEF/HUf91D7COxSZVknE4qKxwfpJ26cAzZExGtYfQjdTLiRqMrYlMEy0NWz
giwTmLDL5OgOiLN9iPetYvr/Uzx4zhXKs/WSNcaIOUyzdskuoibCAXf6XaPmlWdU
CBLSeId+obSSwRtiv8UkBAIHvthWJiKfzwxTgZWzikRNszj4M99NNR1PyTIqd15P
r5Q/fKwAvmxYAj6UIMeghuVZm7WwcwC+NYGVFi0THbcILJQpKTfQJ1+yScMEgqQL
8J/dJx4C42Sy5biDtoutm7Wg9rD++SRfrmCr85ArjWBu3DCatzOLs5XdVs5NOYsi
PuG5idaz+/HUP0U5PpSouPNryc2gQJnIMka9eMG8Q47TgR4SzMK+Lez0tceiQ4jy
nv3Yl9pa29g0MOPNDlEkWP3Po/lA5ijIdqdegxEZsd9TmILoxtiyJQ1vMiC0dJ9D
oyh9GzI8Mi1o87uUMW7f5gOjw2quQ7qyO+H9BOVmGdjPi88eR7Ygem+tVeIwUiwz
lPuqhYutzOPr1T+bHWocyovwd+7OzPmn/kdnv66nTm2VWMA8zGpFHRxE4B0lskqC
LK6WYqsPik4CdG7fNZTOyQlt7483c9dKiesxRaMmojee9A1VqEBbjX+XF/N3wxAH
vXz9WqYoe3VNatuAbFMORbvCCjlK+LP770KBPqOHz2UTVpMtrgzxStaXxEVKL6sm
lCE1+Vg+fl1CCkEilCyp735BIPKytr0UVWubnEh1e85WphDSflfrC8KFWfE5KcL9
kREAKUQMmg4qO7UF0wUEi3Jw/KMYaPZdVvPbcH1tG5+gN2vGM6Jn6m5WGA0KltXX
WZqUFESHPT7Ce0ht2rwkEOF8olCaIFnkkeAv6sVpANUk1V2mI1OjSpdu/C4yhZ7y
Zl/wZQzV1vmoYw2fPIyCSLA4Zx8zspqu80e6pZRDAmX9TpfVZSdw2PC3ftjtd0gd
hQcJGtKLaFtgtAIdSU7r/0XBJY13Mwo87QcOXBQgBtvBQhX0oDGhVmUOhX7PeaFP
YYW2451W6f0Up/jhTFyrHW06/DH6GwrDcajCNITUKRqS754Xa2hNPIF1p5g9L0ms
rD+BCe6jv3DvjS77PP9K0+BIqogsmKGqQvzS3zYdrryosAEL2SmIMdxGW4eU4QvI
RILwFROyFWjvaFYMKH8aH+5KNr+5Rr5DnQBLyNJEScjYDjhIVK8NGiLbURBuioaP
Mz/XMnynMj6Lx8s7oC782+FuzJXlHpyZiBUjgAk8GFsS2Y+cvHDfc+GsXLmBRDSk
ZEMVmmTe0UZcfIWcH0TL0GMq53Kiziqz1dI41KWK8vwM98ihJPJFlj2T3Tm8gjwZ
5uUD3V1z52StTmLmXFSeRfr8BxB1czIAxR/Rw6UEfe47qoTK6Wr5MDKbdLiaz4xk
Wvnp0WrrsNmdpCuHQgJAfSto4XDsOI2ESy+x2SNZPyW4ZoiUoBPDkA4LNYHq/CTw
rYjFweNzT1ZiOkYcgwIguEggn/10RHC/XsJaAFfrBU0E+FMSKYHQdX7KYXqiSFjO
P4tgHmolrvdVFM3nJC1IpheBuL/7ubWlyhwxYAgCw8meP1/QwqaZSmeRzQ+4P4Lt
VDJrphQV1LSZCMxmjKT7XYkkFE1yyu8htAvUIT4AIkZBBNjq2DwTri1brN2rSqMY
OrK2MnwiHHYX+r/HWBjtlibYlxlg1k34tIcrECLrIGcPCe4UaPrKU2JsxgBf9TIP
gSFYRpBYzWLitNBORA9SEkeEZf+NnxHQHVGJYtcY7AJ22rvsnZ7UKWejBm0fhycN
7dxCjG5dgAwXdgZLluggjh9KhPLBbhn86CdUvkcZlhSktqBDstUNHYYfvy58SNXD
v9ByeLSxs7TPnr4DVNA2efNxtrZY7usqQ5meCcbIz9rycrKzrg5zzz8pLmNoBNW3
cdK5LT6F8iniDScn2hy+b5aBbKiT2K3lThr3XOYn9Qd704lWWscjst+CBsJrfoZW
MCLhnXR8C/zgwq2pHyAEDKJWwpRZViPCXDg74jqXem42GhPy17wL4cAKTqbm3vIE
Amtx1JJR7qtWQKz5juVxOxZ4wI5UTe03UR5R0o+6usZU82z7LXal5hw76t0rokaB
R4a0t5xEV6w9NcrXrxlkHbJyHEk/P5/00NTGsRwJrFIZM2qRdGC2Vyhoaj4s44Nn
RjS2rNg0jpWB3Q1RXBGE0iLeVurfQRYqBGr+8FAYlE0qNo+EWaUjgirxRNQ0r2Jp
euTnpbzHnWfgPAryxTd4hzj1U+BolT16WuPrhuey2xBdJKeGB6qa5ojqDbFurOPn
HRZIlO3fCVJBRt2JM66Ft3mtnHYvB8BVOr9r1xZhrqV16cLjG1KmHYVvHosrB0d3
on9MWu+OsGlrrAfHdeQW8Ao3b+NAfWOZndZvBUBbD1iEgW2AX6Qn+PEDkiCJxXxB
/g9+0AO0/GICfESNGl/A5DFfFRWXAPAqJPNKM8cmN0Q/uZD8iXiz7aFxro0nAn1Q
Dp9OMrlsWDG8o4WYj12ulQEAWxdEfC1QDIMpztGMWFTJqg+9AAGl+Jq2Q8S8kuOB
o6WQxHDWPzuV7c+PflitQVQIQxdTrbmWLRrxhJJRlIUsOdlUFhFjdImQbUA4y/vP
JFf943lS+dRq7DiGOPbom5Km2EhracwWxBJX6RBSEf0jlzrcL1V6B/ytJDXIi1qX
fi0JH4yxnPOTapPQhu3dHqsBeHar7Cr5pLRA7HZl/2rX0/qgfsBqE9YJ0JzFICfJ
Py7J7LDEUy/s65tv6xSJhb2OWV//gDU285NvoKQq0tJp4Zh+0mFP9dsfyr1GepOS
pGNs49nrjbnf/aXwklyRdOhg1KnPbm8i358MQ5CjHhbv7HHWqr55T8/OOZvVYbVm
mGQiGdyCgs9fTRdYhVi6od7A6zfU3Likmus559rlt7GI20h1yH00v0F0GLX/eRYm
diRLCxKrFXMgSHlSdoxZ+hc34qxhPrMvgWK3Mtqdy5w=
`pragma protect end_protected
