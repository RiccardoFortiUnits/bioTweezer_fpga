`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AghXxPxougjrtQETFlsc7TSZY7m6OOoV4MLjtxLsbv8oD4yufvuYnXKhSVPSw4IA
/1eCeuTJjo11t8PZKI6MqUS+zylbYyZYC6D6GI1W9dyMv902fy4OEHy3AAlG+jA7
zF1DAdJ4c+Njc/E9jOHhCdN9kTwuSKsEqPtEkxIEB5w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20976)
6AGz0ZFJzJxEAnmMbr5yVctiI6ZUS5WwCRFmPHKhvPjgmmeqPq6d+lIQ+omNDdBs
10Q794oaltpMaEN10Wi5/j7m92cVGtq1tzpzsIHHsrIYPsbPhcTuV0KF7i6l89L3
TPea/b++kVNaoon5mGBM06qKl/I7ZXDOCdLt0K9opY/EptB81JdRvEUUzg9A3VjP
Y/1ikc2bnpWLdy4f3VJ3tLL7jSOQHhKXHZoOqlpqi6vPMJALFgUYSXJ8z1kBlCxT
rgdXc9ke5MYZ+Nrq4H6PbssIRpsBBKkHFD+vLCIlfNAG9zWdbVHgR6GyKVe/61dP
NPiyrde2DA4T0SFhPlotrkPkrglnrvzA7N7RhNlNmjojyiacQ2YzMTIXTfqWPJx+
8XGWQxQrsNXZTFjLn6ZkKz+c+PKfi1qlh5qJtmFE1c6xU9iZKVh8Y7pwn7Ls+WoT
igdAle0G7wPLUFUpFfal4dQ2/kqXqwo82qqn7cFR4NDynCzYzjufOjIGidTOo7G3
5f0OvdUlH0ak38+ciWl06kLT7zIeTIjln227LgDempgzEsY7ZbTXdHV8xAv0wB2c
mCWfAPOd0a4eD7xBCtJI+0+DOSC7UXgHORAURoaYubM2i8Ul0n4chIyxfbvTytMg
uh4Ib5x0rVAp8KiOLhtn81eHAhJpD024EwoAw2m7nmTwtdXgW1UVBZlZxSakJevj
Ee+/OejUgzQneZh+Jr7qQlMy60kSbkT0VV+ZQhg0fPdYv7bdyfxqE1rPM3XsWn+J
K9um+Iv4XjBgc3w9gVbYqdffo3oogfyFKB85MxJ6g8Z3htFFsF22pl7Bx8eWJ4Ri
NSmfEgw0Hsznt6dAjf7/Ju5NTsgF4Y0VY4EGOBgJRif/jhgDd3lgS3XlNcTR6OQr
cGTrUHthuTOVjI0evgRvP+QtuFP07VMOhKL/6Y7uQuJq5TSFJMwEd9a9VluPIsqw
OykKUnH3DyJNewHpsqusLN69BWSZ3pCVnuJ1RgFE4RqDzQtICkE3aDRZLMFeyrZX
McYAroFqKXj2tymKTxfs6KLApxWqSWwoY4BCD/oaRQEh02k59SwraCFZZE0vjYtG
ldIypLMSmKQirhUufhwPDQwUcXy8/5gxTCjU4nh25bEhUCJmJKAKshx7XrGuMg1h
wYY2WiqRMZKP3/zy1x2ViVV/7HKOyU5c6B9Mx3M3ENPyatg7UVlUbTUOjKOHHSsw
nz6qgjjCeQtyJJNyaHBQaWYLrsE3D3Bbkt1z7OmJPrglDaE4FRTE4LMHraFUDNFF
PqmbtT8dFnUp0qZemh/sj1MT9bOhYLHQWb8F2Rp+saUbyj3QpN/wPxWZ+kKdfD0j
Q7rZhrf2/FpVXfsIUIaK/RQfLEsTiKOp/KU4jMVhy/O+8RnS6e57+14uMp3x+mk3
GgKKC98m3vggRNlF7roANZY6T1E8mumzpLU8B5qKFLHDRafwk4hab4PnBMZiO5gb
oROj9snv7aPuYNE/e2kVfzT664Cmlj6AzaDTKEqyLzvUD6hNtXZeMPJB/9eGUXEB
TG0UPWKS9R6Yqg1BfXTrJEUN+7IhReZEkJtycDRMoyFfQDyTqiBvOWwP/aiXW+7/
j9fYDF2z9zF4jFmK441f70ogww/PAXqQzIHGfQ14LSCZfOT3nJ0XpytRC0pCD3WZ
ttGw6EECcHT9frxdgFZ/x7v4nlQc60VdIhqIvJuUCekN8ZaHEuiPvuma2KgEIDBC
kb24f7J9/KlRJVtwci62MPqB6+B294VTiBqFyxx40sUzzp6HuCyXKOeq078THA5Q
SbEIRrajipKCm8NGjnOEu0cQOiGQnRwMVtunIe0RxmHiJwG9iWMWoYAZw5U+/cM0
31XzmUmpm/M+iG+EWObVvGrQTtEyJO5hk7S7gLDrc6KLyAEBZFJ2PG5SfFTHmw3U
/8LXPp5rjfGpLrYRXmiNtXyDAKjTDmfo+fDvy8WnMTKT33uxZMlzc4SAJmwJa2+C
USzEZtzhVBvtikbBsLCZTUlHeeOhfNEUhLtsg7WwTbVvjryL6ODj/1ASfcGmfzTP
ETtw/lpFLe2/BTEa0iXpvl9QmUDyhNmn1AHRxAqU1aB0WlskWlb5zeZOaNRqYFAI
P/suW39153WhbLOwSLQ8CQj2COSHozjZObWZuya6bpxWR7wxfsXhuDnrXG7YA9Y5
dO1KRhhSwrkrLASr4K1TCZrdzrZ3qKVdHSN2fxyIni09sdetFkQVs4yNormDpKOH
rlOs+2OIWVtfrTe5B1xhl5FJQdP0sN9a+avsYmGfqBLXREWyu8kvd7+fq/MLV6oz
9aO7GKL6YT9ysqvoMK9pNFJxb8LQEErrLdIB+Xqfh53sYA/rRP85ztGHnCCRa4+P
HtlrmWZX8W30eFt30TsUNfHGftef/o3x7Mzskqb60dQ1H8NLeUoayJDI5PbdZ3c2
Fr5rWnhTkrKR8WE1L5ji2TN9PedDJAiULF8Nm7p6+Iv23hjH07TxxrAF97xphtGJ
I1XWn6JGwWcLCc1S/uX1wOqLoNtm/c0fiKsevCgyIl8oLS8X0FK8W4+v/R2wkAw5
e868d1QLt3o+1qQ5UTle7hCgawIVbwJgNPPs5pWIgJyZ5UkzBJGW47KjuJcVJkFf
CpTBmte8xzt2nh52TzuiC7oTp+nZK3mmYepWo0zjQlT06faVtDVK6kbQx0A9tPqi
mrJxuhDqKG6gOSUIJIzXu3M3ehjvmg5xDA50tsQA4PNSdmH0h2a3qDFgivzdZ7aU
oxu+KKrD3u31trkgWmiFTZCKcEzVkWbCFhLBYiVlhMdK8F9jIDvgGOctwccQBHa+
i0qy13Ml1va8uE4g4sbHjaSJAYq6loJ0U1++hWGmXdP/46jfOeAUIrpSbNBoKEK0
Pn/s61WYDpIADmwDxWIQArdNlN7R9UHF4wA9ErmoLP6svi3q+Weo4UBJJkkD4PkK
dYmh9AY1fo5QXoUemlAyDxOpaV9NfhaZCECm9ArXhCqLsGwvGXocmBfj7AUBca1m
leimUWizDKvPOzxpE+7XKZMZu+UYDNFpKUU8tv+jy3H1va8chK9O2hcoAP5l22FZ
YNS0C1MzkvaYZCZmrQRPQ39AqSfQGcgUXumZZ2x4Waj+GjrolQsSDr0nkwpTJYFU
WE41PIRtbalK2QX4KCGzL8uumYSOBZY41uLW5M4wjwIaArLaN4tPpIJ9R35TcKJK
kTLrT5X2xWe1hiw/a8dkVCgq/yiNy89iMNrw8Eh3XqrCPpSqAaB2VHxUINhi98aB
kUXHIwg1nzRD6dtb3tZEClvnBJRwNhH2V754jNGXX+yvGmuMBrHAqrOaA5tM/xeM
N5vjn0Ab7svOnh/kb8kcJDpxzBzSWHG+6Krpa54yDEkquirZmUJ1zJsSj0db/CEg
a4GN6du5apcPOCQvKDtft/RLwtp9d/vxyrRXLa958YlopDPMXffF90GsyOG3wcCj
h4kiRCJYFagEbzqLyJ5F2Pr/NMF5iI2ggm6rmvWcxY9chBnZ2M7ezkQ30jHvRtOt
gDFV503AsgUM3mFuCU/NgaF4mc/Ve9D7xUFNWiqvjLck6oowCuPqWDTTO0Hy/ooa
7owUdQaFe1PyHcuTa27GJp0X5UBz/CMAanOCF3IGcfiv4oT2BCtWFqgrcpMV4tcm
7gj5vf5eJM1DF4knhY5RkOugZvd5zcjjuueihi4Vr9Y8Euw7s4WGucrnSvsxCp5o
1MiSTR/x8C7nkBVOz504WARcz4JNdP8y71ZnKEHxuLgHna2zwJ3/YgyOG+TO6oVw
gSQRfcNqO6iWNaxTMKGuikysIgKSzTdtYqQX4Kjr0A5X5o+QBywZ+K2ZloPpFiZc
FublRyHKglcCSqWNSs57y01d8+HXXbhnWuCDVpv4WQxMr6BHxglrA1UONF3LQNBk
NibWedYX8+e1QsWCuzwf50/460WSQtkTUXjZx5OXoEKbp85gajzVISdLVsmPgSGM
L6ki2Qc5fvdbzKwiIs7x7oRRlbWyivDjYeVBvXuRizc296eIwpYXPudOR1zBUVHs
mZhrGRdn/r25iS9aFEYa+tdByhLcBf15U/Er1LzwfFjWIx7ERTEe903ZzFnHab41
gYsciRsZyY4T6ldnijyIgkbQd4yCmq8QbU2yxdIfhc79LuhXi3cicPNqUs01y2U6
j8PBg/NRF0TvK8ptIyVR6JPJqgPRKlfoUMlXpXe5bGjWvCxj4nBuotYNJ2435r1K
x5r24Ly4JCUQAebqM+uUGJ9JgX61vTvKALZS3+rfMzb5Fmydu3WkxNasYLWikabN
A93EJGW1NrxpsL4Vw+eo1/S4h5Fi2Ts2eoWJ9cyIhguDLnQHL+zrw2I7jFaiz4WX
XTb2b1oXCHMbe3kvXNdb4pKK0MulZiSA/eAS/dRerb8xnIiGYsgAfxqm8k/rC46/
jnEyUNIYvoAEU+MYtrdOVqanoCCdzIXAAuT/TmDrrwytAs7fV9EuhdmQDRPkRwW2
VoP2rOn7k7uWlqYRM/XutWQwbJhqkUPePU74u4woORCV4li6Eoqzmj3xFXJfKEWR
WRUvsD/PyRsUVED1DLGqT50R+RrIoWo039bwZWrGZ9Xc3cG+jzXEqZAbpvWUfo/v
+0F8/1R4EyQr95yFEHXmBTkPOBAOWauxnNNrOfBIg0Xb+Y1DdJa7d09xVxsvqEws
x32tl6UWNST4zvcG76A00Y7WeAPJ6ieVS6slbIeG1u/Hmz7urlw4flXHuuAIzYo/
0qKa8T7qL46ZB4494rRQwLpSfasmHjPYhzfPCJGGzbnKGor1iFDL+uCD1xxhOcLU
EywIfzZbf025+3L12VTh5GaDGROEMOlxKtyh92KEgwNujQ/1NPlw+Z186B/0nEAn
4HxykoiidVRgL9LZPaLwVL+82Nm2SuF17sgwbzh6wjVoBnhww+eATe1ZkXFsOmzN
ldlYGOVlcwHICum51szZcrY85+oD+/XBtduWq57vcP5h9zBGMXIEwDTKQ1ZkrsK5
yK8+EUxbvDwFu4Lj9dUiQSabuO2k9dfiNuoPDcjfKrLGN6ux3q/B6PDrjWvmZR7A
BuWmtQWqU1ohKn5q8RpALP+6DPAxiEk1flznuJZdZlt4qdE0QsTWAzZSr5iyvpAz
Uqtowsy09mtSu9L6x96Epp9RKMi9GmP7na+heqn7tSbqkNvS8+7w4pGZqtoHGNmv
LzJjaF7dxXq6miLb1juSmA7DqriafNHMaPDxSEBz3W2DdhsGsSXyn8UhijSeCiZi
SyUoTDWs9XmBPbzTnVu5McTp9suhgkHm+N43YYX2RQbSZHrqjZ3ImB7cJxA/4ZVK
2X/KeGk8F1aY/YJ79tl1DyW3TAI1vVTPvi7Oo55XhX2nU2MiYdqYmSBxVI88M46b
NjPzEbge9HEc4jNHtcnBWZ+VwC4ART50P3fQO6Qxg6XeOT+/+/9fMOkMRg/BhCsu
cFkW3XJ87iPTYqWUwTKPMy4prXDdHlDLUNNoS5Jornwa7r/jUVR05bFsZq+eRMTI
9Q112xZhDd/eJyMw3oYlXv6NQvt/Tw8UoNrt8M8KZElTYMO8mrPCtiIQBzj1RT9C
Z9dZf5tD6Dn40x1IG6w1n3gjaa/2gLyjKkzd/XZSm97VbeMntv80i2yfxAdU3N5I
0/TTuskSg0RUi2H1Jc4a36ESBKMisnLucJDi7PPxN9hA2NwqYp+7kv38ISNGFt7d
iRT0p+ED2HgF1TLVqBRfewRsGIdhhPvWBxQ1AyUtWYOebFeuCipULwajb9zU8Lfe
OmwayDtMTwYNyvkMlmu5mUSJq/yH45grXpkqfGLjtKZjiOya68T107beZXNVAMth
JKYQZ9np3nDORxV1Gn3fSuQseUu7u0qerpuK1MG+GY/qM5OVDMQBGWoGbaAiwvSg
NrBsZs63FI2UZE0VbWuJ37MyrrSkqH0Fk8NzC91rMRJtEmcSNntw852f41sN3Da6
fbcnje0FII9+cSVVtZGi/VE/8Z/XaETePwjPB9akM8xj0nAOjPcp6Kb08DkxWrzy
Py9DfEkOSTDxR/kLSB08/jB2KXVSssanIJo4BY2+YzLkzVacSpLv/f8Hw8nWypGJ
wHNU5qUZ4BGJbl5KMXcNm8+POJ3RE1tagVVxxAfW5urn1Y6jgP0xXOtZj8K2lN+W
cD4j7J+Be82EHMO0QzHsWC2iiKeZbw86SfFP8zvWV/3Kg5YMzVZAKkjuPf1pGb+n
HjkrFnQ3Y0Jl/FY4qP1DeFTTnOYIhg0PT/mN881QqmB9f6ZhsMEj3YGM/JFqjnCJ
QHMQZbqOvIhOSUzpDhbE62v8vAmhizB3z/JrnFSErXA5XHdQqK/4y4GfY8IshIhH
m9K6xHXbYlBpQWTc9csi+WHjIYUVXA+0rdLofMfFGz75BZqlpupy6qr6Qo0xIh16
6fw9FiSsIDV7kh/rns4B+Ylu6ZwioDS9m7Xh3Tvk4ollB9si3zJJLDtH9AFXd6Xv
YokMQQzugYT4OS7DWfXuS33QMNLkdKymhj+HCmGssCK51WNOTHIhoTD1iHw/cTy/
TW3iSqlgKDP2BrLuzaIS+NuUdi9P0tueD/jR9hK1hjc9tb8llIdAC88Pqcirfbil
hLvs11kwsdgLU/hNEylaDfmED596O+KlcOcHIte6dtps5aDkRxUyZ9yemBWmDbch
b72ATaLrE3CtWfrc9563NfZxD9KrizjNxPEHla5UcjmN7aPWW0EeLse+3ckvSliy
xwIEMFNJNi2D/ezG50EbCmQ+zBDPVzKWdxif/lYBHfWcE3u9Vcow+nPLfoNo2Se/
usSnLOcu/wufmgM38GwQQFu0DpYllDghi1Usro/ZKYAKImzBcZcO8b6xxOhz61Qs
z+h2AsguFuVsbH9bhx0H+vpNLFjR4ePrdoFssORHoTOcX4vIvewr09p2rWFNGM10
Vcmc7Iv6On3wByyHZbQcTs6+DySHZbTCV8DGJQOTGUXEOC8l02Sg9CwUOOCOjMw7
vEdDyWOdaD25NQfQgdce6QWGwzRzgatyErsXixm4A3iWUtVA1pHA487DrFhVz9PL
d4QW5VDtuchF/7/PUDdPW9ofWwQSq1hJQeb3mM6AJTlC4rIa3fRG3rxGRQOtLtog
KVYuaioZPx6U20doR4ZWGAkjClhvzcOXhtgE+z7Q5WDkpe8zAue4wIeLpGtyqSIb
Su/OxI8bZLU8XKm+Q5gnI92m6w7c/tRXjnPfNDF/2PfI1CB5LEN9Y/1r6UIC+D0F
wN4SsJJ7ylzUMVh/do02F+t3rsGR1Ul74HtXNbeb+d8yQXTuZ73AiCyCCBbI/Y02
RiBriPJbGYH7ZNI8CPf0V3EnDgKfL8/7/+WmLs8yojGHrLj4AWqjtiRXhIpBF0g4
i2RqFLeAca+XHYYvAFJwWthdVnH4dYmW5AnCJc8NPr8dudt24hwFPjtCpWtDVu6f
4sQNYvZbffHObm12ZqOdeKhFbkwpOfI4TRQY4U0r78DHxPnKMYRwqWSCv1Fu6NQM
f/uv5oVFG3rpF5nc+9TztiyBX58YcpuEWynyX5xRDN9OH8L5cxmQCB7avTp1xxU4
SKJtA4DbqQv+/9zIq7FjV6IJXHaUupnGYwTXv+Q/OJLdHssnJK48frEC5DqdW4pe
2YpIIkni9ad6bcz212qdvcsDWG+q4i57uUQnMPSJ2WDeoP02WYBOBpLA3vMBHs2D
IzDF30W4uhA+mVl8eb62no5cRuQZ5HrSPf4GpmsnEqUGgXyhmFVoQGfAMaKkKQs5
/Z8TFo7z+hoChrzOJyAxerVPWe12bJSOR9SvvpUGH16180DeB92IEnyejm2rM2h2
mjTSFalcg9H1l1tTxiqP6GA/9olCgNc5zRK6yopT4p6dUzz/SWNi3nxQc/wvC5um
OKUcACBJwXD7YsuV2+eBg4fyKIzrrkofrtLgh/XmxhjS/Q4FNy1aDFDoNLFptwsY
zj2blcAUuVal/IRUu8ZxYoGcfC9RRH0XwKPW0yRE9wX7+yljctganIyAuqMfzKhf
kNXZ8cSM9z9YfsnPUGKdQjVGB6tZM7fA1t6OvEtB+Qg8Bs8yVozr/d8f3QQJRBHh
uwC9LrZzoqJzq6wNK+mU1xniDPZjjzwopQ3KkASJxUJZ7SzwJPPKx7c7IYmOPgyr
Q++1AzkejduNg0Y4cHYgB14vunx5WZEWDXAJ/uqMFRlegv4kJHbrc3mYfCfoLEMp
YZYxzDSasLkWRBRUlX0u3E8Ai6WP7dLkzktdMuJft3kWAzpq+lm/j4DLR4gzZj24
addOIr/0+OYfnl/XzeHSCCGETlwA3uBk8WYn2uHfsaOuJngZbHYpUoM0cDUBYJjs
PZmE8nxxyWBWVsAJZJTQkDdWf+2wX2C9FR0nvPnanf0dNnvqZ1LL5KOOga8vlwzL
uF0IjY/dlUgkNazjZ+/K9nY5m/kYfnbdr70Kv26NBCdMcH3aHdGTsxJC6s3bYMBK
n5C/ae8u26d4PWNz61w7V9PfvbIoI+JxXBAEhXaAG4DYroJfz2KrAk6x0Dy/FcyW
ioo9eGjexz2ligbc2telsfTiNXOmGm1R6tQUxF/NlWtDZsm+mSRDCmT5R+edeLjR
EtRUvTOhnKhkXzcURoQgRKQbWz2NPIt7P8xwQpphZAPrl2zJuI7McMlZMhlFV+4C
A0V7i6hd7iqeHisOTh/h/zxSlmMoEZKCH4/2O/ZEfGBZiMc8oGXHxGRl7ruJ59NP
G48Qn39vqv9z6mw55i0jdqsfiv3Iaz4xRUJJslo+VY/G4qqAdjPvXy+nXUl9DPUz
x2RluYwfzU/csRX5xR7IVRam69ssRVjxS/d88JTKeYCkOpmb1MfJcZYmj+G5Et61
LmsywfRK7YEouP7C38nn5kCyrRdHphi40pNwxXdMCmiNiirTStCl32IFYHw8ZwPW
huCVB+SM/OMXFNpFu+oB1fzU4X//wZYe/NgfpQF3czZGOvYcwg3tzYKRWTSCzH39
8nboJmfJ+vcEgekGB4uah6+Vdhce13Sk4tuDIQfi8qsLmwfpoCl38mi2ny/6TODw
WT/Ps6dNfWwe76uavBvwBlEeExqY8YOdBLlFVlHn7eWPVzSAvu2RxQgaeJE74Syu
1219m1n0kOLmppipWxGZSNkSuTZ//rtBxXFP41brWu27cNW7PVipEIhd3O/dPRN0
VOJvCJKC0RvoQm9QDqVAFzE97AG/AteUfzLglALFgfsZnl4vOsLfM7V707tN/Wf/
YdMfdW8bq0097l/gOx0Xiun6hBqlhW5SmCqlfKH0S8hR1Qgd6SXMcgoNgd4tefY8
hv1obl/piP1bnfR/299xT1YPxW+1y9AfSeuZWoMfvAPe1z1dnQLIii3xeIUaHQ/t
N/jZxyTB7gSxfIA7FOaJAcGYpJ0WeHjNPVYmp7Bxma5D6ogoLGynMhMy9ZM5RiNr
QhMMxy0cEHuPZq0RdBujcqFC/L72/xWlTUduJEa3xl8rpfa6hpbFn79M7W35iXkH
e/SeDiPV1Hhr1iN1Bhwm9OMMbvqyRlYuN6WmaxxDJUxE4VAz3GBDM49Om3RSnrJG
ZzWE0pxS+gYFI4IReYOFNIKh7LCQsl1d9lR6hE+zLwwkpFKcVLLXlS+M1u2NFZlo
gIokXf4NduLSW4mEMyhlq0cpxMixh/4XtHmIrMPwpyxFydSXQZp84u7Os9XtHD1a
AxnVNWHXy8aGFkl9nCOHLzvwumdvWCp2Ux8e4Wb5pdbQd5vR/bQwRYkZXfEhUImf
l4N8Er7HhuiTGsum0UBmrQmsDbNUzI4WXBSjmeM59eb6DXiUzMXXlOG+rqptoXsn
guDWBQG4PYK9i3Iu2QH3EjKwKSw23shjSZOlL3jMRgQNzgtNE4q7kFWofgDy59w4
a+a7QsrddXZaJprvKPIgX8M5Zady6vCPC479a8AvaSJs10rbrj7MxjHHhXpp+AMH
boGFNgoVmO6iaki6vI4zNwoYUGF4I846BehqWEm7pFtHzKic0cyuITSybPLEiduf
Gv71wGgdh3Yv/MCdooWYV0vmwALLU53c2980YYYk628Z3pFe1PtKD4CcnMAGvs71
IHlQQwm1u6mkbArTcpjw7tJGizylRlMx086V4cRzeiU9VKvS+qy2l5PzgbKMkx5u
rShc4G3cuDm5HN2g/heB/5mmIr7E91L4/wb8xoB2KstojHPJbXlnlfBT9GmC4Jod
238/iCpnClNHf20cbMHSU+Vz23SytlyJzQUh9TFEA7RJ2SU9sI2vZgiYhu8c0ci6
/T1i0NctVe+5WmM53ZxB2BhjqkDrohGSh10T+sd8Ze7qlXUyOfvuoZjMuLI6EPX/
a6A57yu+abgaeNUErQ7QTSNftOT5g+Xt390Yg6jNYNr8ORg/psgER2xf8Ss5kHyh
dQcTJWwp0xgCHFwCu4Lp1moBGqA/h+e8FvXH0ClIrc7mTuYZYG/dfdmMUlMQKE2K
VopUracRGtkaWAkIhz/V/Wa1GppgSCtNWe7lvkdzoCr5Ws4RTa1rLdRADDhICbVg
+VCuPt1suvPYA7Glf4ngwxmGKhjdNqBHHxqjnIDMASuKP7amtjlH7U/HsGDCNSDh
zocIRjV6cSXmpeDhe5hKsZn6J3aHMNQl6k8PUhmGvu+Ns1eWRDRYGfJgnsEQK0iW
kDq1ZBlC7yt2R3dnF6WCcxn68FpG7scohxnZhNTnUSsByKf1OhYY2u/1z95O3kXs
lBXRfuB5ibV/seOmmb9h6LXUD0d5UvMF1xz2s6HXV1KyJzacfUarUfATtGQkod3e
dsaZiz1R/4/10VspgEjJQkeNG3LmgabooVi9ml0FRJXlZ2GqvmKuEkwKWdwCHzNw
zug2v3003laDlsy8I9+krCOdnxRb3QSpVTMu5AZens2jRW1z57mMUPDzKbuTSjRf
ZUshp00tq47fxbCbrhg1N4Hrme8GxG7+yewqON0RLyfk3DluJuqpHB5uorIeJyvN
zj9pHvJ//Cc8AkzktJhg79XfEV+mk5wc35hGeOwXe3keAOzpc8/lrDdsKubftB9+
mujeJrE88cxLLOhNNMz5DQmhQaY0H2fmHNz4gT6veBUr0r9cSB04kkF2Fi1bCNpe
8Ypp6I5Pdo6sqGSpJX1n/or4zcUeJiAXrCydHjBS0jaPnPdgHNGlttOKxURoj3tt
C23etwFGNDct4KXF2+bbY9IU4wa9wJjdI9V5DDje+ZdGRvgfzvuIl2c7EXoAr0uA
qH9O1FPZ45kW2D1lwC9FIkssPsc0xFp0TdLkKRyCheCUBVB0EmQ3C6cXKrCbUzoR
eb6i14JHgUgDBwsxJlNWAXcvKcI/aMGGKR0lXzKrnWsIhkwyy9FBrtGbGSsswt1M
IIK4l9w0Vb5HYIj0BJAuI4WOL0i/aeFLMyKkkEz87aH123MTMDWSN6uTzjw8ZZFo
mirXwVfSVScRshBkpYLz/M3F2Dm8++zHgVp1Gk77hX3NeCOzw02JUPx8ohWdkxDx
w/m8WsA4Iwm0X5cbqNCpaSDjn6zHl1FsnNftO+9/wPUflUu4hNeo8rsZYAtJHB4E
vIeWNxhPzacBp8SoG214iUqxkcZvJQRnJn9xCb08ZO35T9pS6ejSfuGyR7OMlj+O
uofjKJ7E8QPEyPagjhotkZP66DjVG7WyUGgoVKFKp+Tgx9pndZXHm0opJsrxccNp
RZhZ4P0Br51QYkfolS0NJ6bRL8bDp0CZ1vqjTiOuHubXE/Bxd5RYc3HO5PShuLst
gh5kMS6GBmALy+wp1QNOtYM7DkNqppFanfr870vNHlgA0WYsJ/Dq8w43dCQAAg8p
XVlF9P0U/dvb5t5G6nLr+A+c8GHgNuKHzFfvCd2hJlA/+vp/f79xL8gSRJpwUdpr
srXIWLHd3og++hhY/IePPyA/bTBPu9qOC/JSYODxYSzZkgi4cSHj4+k6+yY92aBd
NAXCsxMmxVUH0FQ9VNzo4Y5wBsHNeu4jGXnXhJbm/A/uZ/7jUstD6ld6Ep8zww36
hupugSrD88TYwrFBgAtqcRZaMa1zMyTWRrnv8AxAy79NMPyi6MkMU60fPgzaafvc
HdiEKXpSt2blY6oqZQFzltCNQVBuZVfo1nhzsbHl0r41+2OHv1c6VYWISUcTVH7q
cxLplH1CbAQGUSwn7jeuhhr54Tz33TxslwmWJAIz+bPNg1D5kBSQy/tsizkNadb7
7M/FM2XMjW6hLeMewUCMRYJat6U6/nqej8Re7nXeIqhWeq1p4R463COwYMCsktMr
c8aUzD4MNIJ4aNikxDuvDijex4pm17DDzdf4BO3LKY0gBdgfPY6KgNKpwpcEI+JZ
7FxHp0Ky+MEEiwIdq9t/VYWq1hpCYbkTOSeMZG0Bb4BucnammHTBcfHg8K6WJi+4
HFA4lDUsfB+B6Q5LlmA/JxgJXAFozveiONN772X13nuSiVOFTtymzFXXtfoVt6HA
uhMhdF0cLwEkgqhtKdI3DhPQdp87ahSeSx301VuPUSqYEVtbRugWLhQSNlXe5EHr
S3T6sSPtzVRIPVKBEgcGIX6DUk7AUfB//DlzNgFVuHYWdCRDgaIlM2OJYeV5QivN
XtrgqmmiLfRQ6PbUUai6aRUqesCFXgOxWxRUEgQE/54Nw1tU7rphAwBVLPMOg5qQ
rPsYFZy60mx0OuScKDqm7vFpTr2+WHBT/NzCfb9I9+FXL6XGOMxKzJNTew+MHbz5
xDKag4ENwX2/S1gRllo5sOGRILF9YlnY/PZ+SWSpLnbZXlfaOMjLEbZIsaaLRNXT
eC8HDBPvqTeTotb4oFH/fyHc1ExtITyV3VCyYVOyq5wVdoF2Oz2X2O7ninIkBn+1
biJfqgzV4wtsCS2f47IS9ixt5RY3DPV7TbnZz5HtVuEwRfp67B7kRgjX4uFPqjlQ
Hj7CSFsFJ4jgZ6RMrL02dgRz9DLAIozG8FbnamgLJZIELkG4Wjccm0FLg3oSt0WZ
lYKLBcDFVnq/OKTG5WBelKC6c6vzKWOy/YNTQKGL4tPy5YB4KqyPnl8+TQueHgl2
uqzyMJA4fDeb6pRAm8Iz84kwT/IOjS1nUbH0v3WMO09lUpjj4KP4gEY5Ns4aRN+2
654NEwHzsI5xoSM3EiLZ5fs2kvzHCwGoMloEAs1ce//glPNCZ4YHPZ75EEhl7xv2
sjEW6JZswCi2OAIjVaM4feg3i+i6jqE6zPcqgA/dLWzLeUk2FRs9HZ6eiWFkZDdg
w+SvCayod1G1Gcn5Dq0yLrEpVff0EgaPSppnjLZQtR26Gp6GJ1WSLYdabYAuhVnn
9pjjIIB4UJHSLC6exN2ohUQmrSOBOE1ViDDYMq4gcFpMYAnDYIq+EEjXkjAbSvqN
BbufmBg9qD52WA6fh0A6eBmk1EU25CQP9nAOfeQClW4igCPP7VZRNxPVAxGSaWBd
FfdsYwfV36pxcuTpmMNLe+w89rhWScdqK82bQ6zxTF0EY+u8KHumN31nI+7RQmrF
rIBfncUV7UB4ec+fz+KaeCXxN7qHf8Eaxq50lHOxlBq6OV++efkJlrL6yypyuua/
IxF6YTr7UULsT90js118nD6mTEDaMnLHf9sAnBLKtpx2RGjpgZnhWlQRlq0gv1Tr
zQatOWDvWbAPfSIynm4q624qShrCJqCzraPHjMYbcm+JRIq8Z1ePeZWJimcZA9Is
8ieC8toEEus3ygOLnQJ96cJ3aK3/xpfj4pkhvYkYunUpFsGsysCx25C0Skqa3EkV
HPnsYiXdwugVWoDcN6kxxDbzqzQNGX9bBvbhaG665X+KnBVIW5v2W1sijOITSp9w
XY4SJ2BW6r4pnRXsDzgMnZR+REumKx2WcYCEuxQt2y5tB5G8c2AUT8hnHOyJ49WI
i2JUhBQcR4bxsFbeZJB36xRzTgyb3yS8IR9Z9yTT93yVDoE4cq99cCAvwn6JPeoQ
d29NPg3OiJA4LFT7Wn2gz4N6RUbuNoL7EpZvSGnVMm/9CurD6Hp8hFCUL/Kvm38N
aRQCSR+uuAVNzXQWuNZZe9jkglTnPneEq2TR2WYHK4IFVGLAHEn1tI7lPYkR1lvZ
8kFkuBuLCuz0UyxKvWKAzZRslb5PydrHqAH06nPVzTWeQdzTDgW2THloimzUjloZ
OTXlDHR+VXY3/KS0hSMT4bummHHceWJ45dw0YEOd1ly9E3mBS51VtKvuQQjlzp7Z
Yea1Xy9WXZz+M3he/jvUAf7PdNQA9KLrjfQUKdkUL2TLgqQjGqIxRFzKG6C5Mpqs
JVi7qvVU9XJTn4KkuFPnHVoUl3jt/HvC+kK6HZ3Wu40CRQWh8DEOggzBVWtlvlHg
WhBRRdXEXxhmiitCp+KTQWqdN2GylOEj39BNd2xbz0WTg1O47V8S7TC82UicSung
PQ1fsF/yLVx6eyOkoIOsJjYfmSQle5xftLdS2lcjBqiXasEEoYNeXlbMxYM5+eUD
0UT0clu3bYxxo6pnjGuF/I14h18UeUNGal6GlRxT36ZoQI0kD2tIn4C6ID803wUw
DiJEjiqDrZ0eK65Oo1Vjs4+dG3g2O44p3393dSQgigOLdrQKI//6/Q2AkjM9WsNy
a99xIPkwE0AVPaoRbKec9iNFqV/AbWYaSSFdGm1hJ1h8HrH1+RB4OBQn5Y9weegS
cPD4uavZhR7y5LIVSKSL5LOiHzb49vi36rmFvsXL7ixvtIGqCK0JhspwTdY2r0oB
saHCsjloz53uJ6/TfyL1G1OXcCEGmuq4hleNsepHBlXmFBUDltNLbeKHFmqCBgi0
oNZc8KcFEAWhs8+lg2zt/qZLkzqcNJjopDhGO4calTMrh8xMU84pbNjwlovSh1sJ
uWPCQ02yM7+X5KjRQCq205jboPfIhj+9PoDWUBkkw7W3tGgH0/1OLogztZIyfyX5
9GB9VCqC34zcXdURvBgvglUbdG4oT9sD9xkcQX02+dGJM2tiUkjSdzBl6FBxRK0i
QHF2TMFF3JT/nCgtXZ8fWyhah6whM9c7gVJ0HT5SssfInKeNzDXKlsP2fVPgM1b1
gW5b9QEhhcekZ+DXzzjXkHbwec8FcqldHbbg0hxsKEzTJe+OCrjJjODUST8gPN4w
H8q399CYe1K9rZWxEXUIJ5ZLTsQaIutVZVLb8nT6qGYe7BQaG1yNj0ULYa50cgXP
1r74xb/mnkLKN6chwRbJuc3u7uy1Z6JH3yQPfd7rvCNL1gazPmmSkO6LJGN/7rPk
CDsmPRAnNI0MStlMk4VVpPFotVCkpxNzFQH8dQuqp+xGH9s+APmwUal8F5BilJPT
sqmsntIVhX4ZF3tYAFhUt8CYqwjQRe0Ifi6aF+/xt/rLyNpTIvFeDGkoseFCqb0S
w8SRKDGJaHwuZ3Cm0HmBx3149i0Z+WiRkQkZpsslhbilL72s9UvOtxE4vS8GvxNd
d7APujYekDNZ9vsLLrKXFn6rmeywoQ0rqQq0Yuyx/MaY7+GRRRWhjvf3AUpnIjrl
JQQ1FhKCxtl6scKpwIt9d6O0VrA7yqHMJLG/qt+zelQj9b5PMvZkokOjhodjjmhO
oZWIrp4V21oE5W3HEjDbn3U9nxFP+vXDQF5TPxWJkSB89z9rHeJz4Jyp/ckj4B4h
I6S9C8ZMnvy8aBiXh45xd8d9xMXuk1OmcUn+UgJR1gGwbGpC4KH02EgAVcRjy0UY
t2OPSwq2y3isKE5Sss5TUYRcL1dY7lMX9gK7H20nPP/mF3k3oAfjNjrkr14/ZnHH
wKiIekK5IL3uWsVDHNR9+a9/9sp8zoEBxTOnUBsN0zF6HK5+jYVfiW+q9rtIlJCm
Mkzeu7wTMc/t+FxYYagz+3WEWqDKfzOMgZ+lr4AoSKH0wgG+YmJjyR92x5PH61+7
WoD6oJzo3CQf4OhpgmSeHyBBu8W6hwhTL7El6Ndr2xVmG0A5aykVGkGAftSf93PZ
qDIo3gU6FxY59LJ9jeRuKrBzNyFyEYoPdaJuMjMPPcJVJzpauTu8x3i0mSk9whjx
nPJo/TPbp43VQfCzFheJRJxAKk7ERH7bSboM5yAas0YZ5WefrHHJFZ35TQ4PlcaD
Cq3vYBfOn/nk8Auc/yKky28LLuesPwa5iCpV5ggJHeLOUy0wh7JGG93CGCWjnQJr
9bGYLbZ0kF9nA78CUeGQE4U/hw/bdk5Z4rW7aYslbRf+0LsCAfi+3w6fgEhkkUkV
TT9oMKk45BLxz0nrOJgMNd7zukQP4brhCz2/ILHc3/JdPa1u/koFIcXZoHOx5g1H
/NERRb712O6cSExhJrEMZxkVqreQOX/IpCfY5rRYq7wYwc8avw2+QjMNE4pd2JRG
p4I0/kMa0+qydw+s47bnDugLDLEdX8Fp4hb7TkSGnSBwARdbKUTkckHrtlxW+sJM
L4x+OQ4+20orhRNg8k9v7ANM2hwxd9WnVJX2aVeCBtdT7yUh9oDDKENoSgsJ1TLC
nXio2ctdiRrljaAKtOknPTmlhyfSWmhVgUbgF5Ab9LsxBwu4hWU++il5G4MBOvGM
9WralTLG22gcECKLgGanIiQ88m47YJdMSnwA0Kl5QnT9TWuB3aIYeJHKucjjFgRm
8TuNE13uMVUYvnk7NCGDRbRvuthSyxirDAuvYM9lDPssluLrdhmIBE0PnzaWk4sU
fVirDHnBBDkfEdMcMBNU6HTpBgCXyPmHX/5/nEhBwou6cBYj0Sbv0B9bSye83tAx
jgB0ZwqJXekaKIn1wRGXb/vAY07lpEUcCkP0Fi9r0D0rM1b1jIiSq3u5o0pMcPFw
p1L0syO8OqH55Qz2CzXy+rwfG6Adq21CskPxIIojj1a+69T59V24kv/U92EpnxBU
+8PBQMYPZtwW9Usne+C/lFDuLHwH+TM2ZqCCAqD1RcYhTluSYJOkew6/IOsFVwl7
V6eW9pg8rXKfCDxeOrCET7gJLJyE4FIiYCNq1M+95VV0dLYYASima5L1GJhm7Ui+
RR683ILqadR3uNvFrC3jhb4mvKWLdivzbPTu2KjhkpXeSg3tPsFSodUkyeOun48W
dvMwGwi22LEegYoUACzZqmawGA5WMZYYYpiwywzLyAe1Tt7zTc4YeeM0kHKaFu/x
3HTIOFI7CrYQSs3EFY9Ga/yEz+GdbMEkuUaqZaoLQVBMXFzxLnitQmNJl16YInox
L9fcgHKoHFXjbPQU2uWoXF5+h2DUtlc+GJJrPkKR0zwJmcFxWPtednLsUXbuR7LC
b5XNgZZJmeFlgCRnHm+rVdHj1K9mID3PmfeE8U7t8sWCgwQZzYwEVPku0lACWK7f
hSil/9vZYUWpQ5rjCi5CoHzwWC8UWqsoq2o1OkNxCJZ7lkgJSL+RXW8g6cw1utX3
kNU0IDtOOnGRPQrysDn4riK8PGLBKZsGsOiDyhBXqlV1rmCvid7tBPddnQtu3f+C
JwbqmOBBq4c22Pahy2syfbsROv1ftTv016meri+Rw54GjfiRivQ13t6eU+Jib4BU
e/rzskqZpsXh95QyOW9uABzm9G+eSL/qV2aXc8f52s9R8eKSmXzNxdH52ee5wv+i
Mm4Fc03xusV/j/whkssaWSAX2j5Jz4BArcQb3v7U1xqUjfmjuVnCX20I4v6/jk5M
f2OsPFBlWTBlZ+cpUO/IM2rUUAieGctH7Hj0l/lbJCptTBWWJ2VKSDg0Ay0G1Nfm
8E27JikVBrFrAao3BH7rfrRdVDLRwWQ/wTBh2swYSBuiH2hM2CYRopXsW2K7XO9D
3q2cjCJ36dRKQBoP6+CZUXFVEKbRg0g/KCrtExCn/W/nS4bDRa5ccK1ruZptk+eP
qpWmO7vcNpWYl15rYGKTkSHo3DmAESIYhMi+/Epl+yZdfI0l5jHaM5P93zM+1D7z
DcXtsL1RRNV6wZznBEj5y7qbeJIQmdQpBdDqFoFM0ulE6A5MoEj0Zx+b2qigcNBV
y+KPrfkIHK+2ikRAmTWYr5I7NON4STPwqOSNMGb+0OCOOPENZnSg9694hX4jOIII
1wIYDB6TM/lul6vNkbwGBAOCFn/sqsNfghPtgx0Ggq79LRXBQk8puTiaudPixNqK
nwvjeSOHtNzqaZvwhMd4/E9D1ODVqTFXl/Ait4h6gOI2Vgjr0EY8nzyuOrZv9N4R
LhrsXNy14YmxBndvkl2pmnJljMKf4+Z2rwYfVIH4i5RjiUWY8id9WHUui4PyuTkX
vhRnTV09681vEooEdVf4aHNI7dDSKbvqZVxfaHyeBdPb1BRFLgI7tsFBK90d5Bpz
g1+F4TJay+RezGD5VaaiaknQdmoXlde5OOaGV7IR0hW4wrSSDYEQldUasDkWVzF3
HjHCIizoUon1B950JDbLGQNLxd7Uaek/oaXpXmGwoWh5wd283cUtpVg0kMiD6wu0
ygbJ8gB/THMv4WQza+VSGe0bmu7Wzuxs+YoYfi3UFz0K25nXoQE9/Gtm5lPTbL72
17IN0uhmXbpeSOlJWRcx+I4AsLbg4/pWISaY4hFfwEEfxBlbbzfMHdqowjqlYDBB
doNaVTZhfaU6+5nZBK9C7e99+fPfMI4FW2LQaFS/Wowjz/PwhFREii/ZJJLigAjD
2c40A3c1EFIjGGa4NphP6UV3aOtog8NiyR1kt/bktIYuz/Yphblka4OIq8KWUB27
Yg/LEBBGkPCvCpX8obXyWCYKwPcFR3zb24hAvOQBrgrbtvvf6pWUImz5RUwcbSUj
c4CN4M9pCnunNOX6Vb1pTc+0OkbivtP3y6Td0/myawAIHlpTAELwNnaAVO+mJdng
AKtEuOYd8zP4S2Bl1ju3BdFLsNx0S8db8339gEGRvZY6JQquyQQgZeXFgTXmavvN
Xd4IHXIPmRcKYHTMp4Y1vrN4ThHYc2haQNmdl5tQgGp8QzyLA7AgC6YHZmFRzg5+
jhl/bxS4lTqGvysqfW14oe7t7N0m3vs7WV2XDC4GvnZ8ouJmc3dunTK0j6Je6oWw
nw9NGI2Sm9hP4MpkVTWlAEW1nhzkfhGLXSSSS4Rj0QA9ZFoTWo8SpNzqQHoUWb00
Tg9NXaS10rAZlRlP7DTuN38WPmw+FfPCPN/W7VOoVXqReIejDqZHx6MKjGPUNsr0
R9BjH28ED649zcLaUg0DNS93n0Y57MdKeRYwgQ19J4tdPnFtJBLnby+ztm+Xe+CF
jKESJsx4PhAbzclstfezGRyYXH9ZbckxggsxaH+pAuo8wLc8eAA+74PCnbfVwYk4
vmDNEF4qUG3XR9/lWZ2cCgaKpgbPxF+MKPlDL8FthXw7BO5J6wwygz0AEIuFAjSv
RrLsLj/W4LCuMmbmF+GirVMeDXDPujvs0GFreREDJEsVCB4miApBF2tJT7kDlP9k
+XjHiYga495yKUI3friXQthBB18yhL5UbsVFI2mzrjYRWttKegchxYkz1r4GePpz
EW4q64hPOmmOxOIX13oIXXMrE1KDn3h+NVI6gBxXr2LOt5JdDi+N4mWPAOrhkefl
LawIyWeLAgIhKLIqoeBpMzgPAeDPDkzVm0L11KNmucrFGzOyDaQ5kWWXxeuBBdMU
hqiLzRSaaXqfLjow7oj8biMe0dg9XL2jsj5byowA6OYde210rhNdHeDoDb+1HRX3
s2UriKNF0keb5w5wa7o2pg5pOXCAL4RQs5vWO+hFpZW16FDxwa+3alFMB5laJaNd
33JucSyGoxXutM2ZwBoX1OKbZGtX72Wz5PhOvaCCRCgLNDtixnOy6fJS0YL2tTGT
jiTU78JlmBW6NZ8qhK08f1IR6ptO1+UOSeWxTTdNd9hby9JX1v0ACiJg0STSWXTx
w9vJyNZI9NxxRnbD0nT38j6HM+bxqRu1VRU9QcGgHIenqqMVOW7yiPzLKZRFoI0o
EW2ocIIrNQEa+W5lvwwVxrEIUCd/Y69tD51+yTBhCFj+q4gAnNQjcdYTkv3RHi/K
5V/BP5xc3+qa2LcHgnyEvIULTphjolZlmzXrewpxghwrRo4+Ke3tE7yvE+7dWyqX
d17RNgbI34bZShlT3JOlbeO0k9kxjCBTT8uBCMj77BZISGWmx4GCn4A0yar2r0Q7
4TyiyrNibQGz6eqlewq4xjCwMfHl7r4+T3l3XbRo7WzyQlF/IchjpTt0gzOwkQuz
tb8z/OPuIc79OLqCm5olG26AdNs1skpypXNHfQ5OWUMDVrWfY7i647xcvTIbruUf
sBLajxU5GRM+BU9iUR3O1cxeD9B89scl3uiKVQZUdPyslygMkmvscL/+s9e7AGQE
xuubuRDAUaPRpmMqEnWwplrUR7vFGE9QFoJbPi96fvn3z3VHfLMlA23EB/r0j45P
8rdehOA+7GLm6Q1grYVmfrLSA3t8pMJDx7lZhq1v1hw6T+liNfnAGwELql6X54hk
LxS88Sh8SOopF59qmxh1WB7GBCOKj0gpQ6mZtYs0GiC+Kot52GLHGwwDg9aeCp85
Y1fCVyMSOK2wIThrRd0BNSsT0SZkV9KAYAdZst8KSRYRvJa3mYTDJLQTqbDuNV+S
4i0Cy87NH6Px5euKIr9s0ta9XSdStTmI7/J3Vc8X/X6MbuFiWJ3/QKIZV8+PGiVa
5vUyZZ30zZmUz9HxQTmejYaQiZQlFExbVQn2wHSvUa1DgxwcYttu06QdqTq/8CFf
buPh/TfBDUsHZhgZDvM0/1GqdWSsXengmTIfq5JGokhrIp1OeU3QLuofZjCyhZhl
+VjAjok9qwZiaEKpCpdrARPa3Q84GEfnoDMX+H21GzUfNKWm78osqjlqdTw/xfEX
fdENRXtVpgCmo5j+yqnQ3SlHBcXISNxjAnki71XrFBxahDgOjR9v9FoxwN6g2LhL
KFdJJltrY/fEzLAn0UXO5ZKwC5pRo/gsOpLTAUp36mQXRzQqUMZmZ34BMzTvMEdB
P6kMn/DHrteafSpa/F4mClq/GqnI3MjspIAGpnKPej66xEYI2GPrH/RhFuEgOc5j
VTfi9pblgEWAga9XJxWbDUi+fcwWwhoP2VmXYF8r3IxNDrX5VIT0VNlclRvCxuD3
Lbq3u3d4E/9oM3kbh86wTDeM3RzmSkVbVCCR6zWqs4m3r7bzRUbiNHsveSwZS0DP
JRj4pH9iDf+oJebEBZKxASBCAsG0hrsG5647qV/5bSzKJurvXA2fr95fP2HgEL1M
lUv7Cy04sD+b4zR9Zh5nqsugbtB+o+NixYsQ3oLiOaxBfYgbgE4r0QuQQU8thJQe
R3S50CWg0vsyUCtgjdBe/1yB+FhPqQzysgz15Qwp68wHoZ6qkJEYyM5Fw4iBDlEZ
c2jbOKQSfGcLbWtRixiayTj/yLovarlCNimLDaJZ+mqQ90kap2UEOICJnw+fihOu
2q9D++4vGjfJ5qQTCz4QCZS9r/ETkghGRHGUsQH5+eDRks5udwU5pxbH4TwmeLLA
TG7cF4UYMiMpg0rXTUvwacGjzUsAlspFCeQd+ma//xX0fSUJMbgCjYBNOTOx7AWb
azcW587vfDtkImNPL2Ru1XgvBj8K2hkX9qByXl/LQ/SOpiWlPIMIFrTsTOyyMj2Z
mfpt4oqTR1VVjEwOONZ3tbcM2J+/ffMBCWBmwi30joTREDgz0gISgnId9/1672nu
j1RQ85tldQvDSkGwl2/0cHFfuijaNvY2ZB8G0tP3/GTgeWLhxLrBGVfEqb1ncZQZ
i14Nt6ns6D1RkmK6tRtNI5Of9Xvrg8dBFLazaSXHlQ+VCmIXF+5F68OaR8kVNpGY
cPL+5IJF7FNLYT5tULsmuBlTqPJx8h+3Hetwb/e1MsdXD2Bpbq3dN4IcmI/b0nla
k3oRebh8HSp+nlOWJvUwjYerTtDHu1+j2XMS+iRr1ygQjnsE5aWxtMAqJGMTnDsw
1CS3ROkb6mLjQv+69kxFASTdxOIir1KiTxF4Pf+1P+hEF0gu4LB5LSgXfjQLFo8w
dQK/GFqORpJNgAEpQenjSni39BDHaxmfDnRG41VXcwdtX/JqiWF2F7QIMqlhK5tn
YN45vLmWg4uPn6NFsk9lPe5l1n7TsfVqCAQzcOuO8VDxd1Q4kqnOvEHZFWPzHmph
yjyE/Y74Wa5GRkHDEOWo4CW0l5xi2tvpwAB27fdMc5BMph959aIn9zdrzgPSBY01
gVZxvik8TYdaDHDHqZ9kEzr4QNokbwqE9EYFM5D2E5gJRHUMp9zeFMDS0Ca0dXh+
AIc1skjSPYvTaMQJjwBIYqJ5BZ6OCNCU7c4RS5qTsHgpTKrPVKQLlqL5mNkLfQWV
x7f6hVQ3KEKrIF0HkNjT0d1Vrxv1mY59PhRodYbsydFrNFcO8qSJWfBZ4MYC0y7e
rTbUs8Y6W47P1XAciLSQser05lfvtM0l8hOvc2+4RGVS9VuDs66kXlggsa7Lvnwb
w4xHYovEqkfxVBLZ1l/OlPfgEC9m5DB8Dst1nI1jk1NO76l178wMnDn4eLDSL03J
4ogOm708ia0jUYWUfsLqYKH6mjWkRLE10ld50JxDfVfHc7M9DdQeesDjPwuF0Ehb
xYwCDlvQtZwkVp7lLzHuk4qZ9pJrQizibsoXI6Ye08zcCU7RTZEptT0LqLsEPcu/
NiWMLmkvdzHVR+HdMCNJf63Y4RbtE+8SSaoEAdWQT4j57b/k8/jggcdVmSqJXPHv
pnrvbRw1hbJU28mCSB3MMVPxBEPzBMCW5x6sJVGoa3KAh4HbvBntuzW0BQ7vFToV
fCVK2yZ725eLzvfN0lkWRIbh0d+Wk06eXcnx51rhkHsBkii7AQPWOHGn92+6mfTt
FUwdC0VoUC7kL9zySTee4U/O1GZqoEb1eqEX7bHcv9rYVilZC32WM942PNpkV9Ef
FCZR0iE055Gi52+MtmZCo78GdtA3VlePMyrH3j9aW1RoyKPczC3YF049oGPfmF42
10LQhoUTZUS1R19sMThWp+GNIDJIWqeNRAGhPM6R6L/bvmWxoNfM4Vxze/4lyN8T
VCFUCZxi9pEreg/iyx1FkxLCvoGwi6nlogNAV4fAjf7wV+OEIBROYeu6Q2B5gSWt
JRM0mqCVl6JZ5qGbNjqDVdZMxJEJo36jTuqKHW+fJe+TVddfq5grb3D22vSif5o8
siVvkmMesBe9e03tx/f4VJYm62kZfiaRtZcMsKWv2LpHk3aUyrRw6EY9hOek26v7
JttaOvbrMF95EAhZl3lUQeCRBvFo4+TucBuQpLrw8lmLU8Z4/RcAJRqAJgfOsRhO
rIVgR2oWp55g7OvePmsqEnhDdLBmXdJuj+nqqRYJm4fJLn4n+qL0Ru+YqC8WkswQ
mJnaYp9dJr/gYpoDaYs7fQvxawrqsRxJzpQXcKodTv+WpHlSUl1dbyIzuC2s9uMR
ER3/HAvK6GLK36XGbvnL+u4f8UWisZLDOABapblHX+FH6vjxTbjUvQd3TBgSoEPu
9H9GedWjgdq16S2KNVfH7BbJ9Em2R5DEQUSWHHIdGBAUc5tHWMA2N//oHLs9xI3m
0O8XUupTCefvCgjBGMUuxlb7oyAgtGU6j4fzZAuZ672SyEJLVXyc6FRCznfg87n5
zl8PNJ1ggqioOWiw44CdLvmIIIsHoHfkk0X+pDwrwI2bAVMYj1OaSZVxivpDXjwf
KHskSkQFB4ahkRK3wWXSg78OZWsZkr5IKoFAMYYIEKpZIv7kzAnkfPCFS5fADq64
KLCqIX8rMl531nM+kFui/vARvHJzxE9tcxtJ4NIERIYzhSUQVwO/zOxIWSKLKd/P
045RMOwSRJGQl3pWUHdQS00wqt0FC0fi/7CmGPVsoXzfTqu07dDaxUyWZwqi9qTn
/NuuAyitWexLJG7prauL6KwRCDQSm0Cui3S0CtJoGnzSZq9OAvDbuTQFkmDJ3qxv
SSxi1I0Zi4ezSp+J95QkSuKvtion/g7I7bW3P3KnARfhPqV9hobBV8CUXGOyjF/7
7VAOPUDJXag6xl6Xl1LajJxuaqAb4CUtjZurU9yjgmmHL0lrMf0ZhxyzvQF6i8vU
z8vGVN0/iVvD9qp/39cTKzumgD42u6T/RlZBAnSSnXHnQMM3kPdf2ilD0uyPDGpy
BcF5JC6oV6G9aMMUi44Zx3yDLRtIKU7Zx6bPsoUyYUY1llF1H04ZMoMWFxW8JfnJ
Vhsm0YF12AGmpU+KVhVVFtYgyIFsrQh0Ft1nhNv5LtknBkUjUOywzPJsnsOqe5v1
XXA450sg2jh3iJMwaDjJQPfaS5+/TvBn8c/Y6BLhf53ijD1xp7LETb1abE9h7/vX
5wg79wiAkGe86TbG1yazfk2yKgCYA6Pk1Nuv8rfbrbVdVzQJFq7NjfAGWParJNbS
aK1pzI3SNfJMfOnkSXF+P28M5YJ/+qyvUL7hsPnlsOFoYe3cgy+/s0iwyH/hZBEm
AvscIzG7m4lNW2b4ZrHm51rt2bf4fULQXeB1mtfPSmm1cMhFheQ35DThmQ/7h5Xp
Y7p+rR5MVA5ExJbhK1wFp6C6Q72/RU5UFqhOhdilyx/Wej9Q7ZTmfQTTy3Yk8888
fdOWyobo0wA/YDxAUErYGyZwUYNo5oNluzR+JSir1UHAIvE0FAbJSLKssm7DuraQ
OE00y0NCD2ZwRAvMj+s6YUbkkPQYe7/u38DBs2SdeT429xOfrzNsQjlmn/13aV6D
AHT82IhDpkxJxnGMTWPmqMv2MiGV0lDECsQtHrmLIL3xiyuWSVj2xbqyNX3bDlj2
nC6elziE9PW1G+QXpmPf3NxysDOZUm1fDoFh9DdmvqU9norGj6qx5w4KEHErCu5z
2uNs2zy1l+TomeIXBGHx9U92IFDqKFHyw9Lrs3cuL/8/dmOTWzgyXqVA7s2UI515
QXxIpv68tKk0DzMnIdSDYl+aRzgcz2XCf+wKU5+w2nhIPtptFQ7Wz6t3lNSiLY6s
pNZ6ZSO/SbaMG0e5wBcEfFUSKsnsAcf2R96tiZ+h6rTKIQu2/a9D5C7RNnKc8uCO
I+1D8ErP2pG2mJkHAVmvxZOujvDXTGSmvJs/Y30Lt2B6saVFZOuHPRqiRmqryH24
7dKTZ7/VcerrLbBbJumh26/8waVwdxVHMDjquH+CNcCjgI2Q4cnro25uMD+Y8Lrj
knMYwRVWTdbsoXXF0MnVzlYE4MKy8voE5S5wKhUdfQ9FY1rJ20gcTth63bwc5Otq
fAZ7NRbVtvWqqVYlapE9D9yIrOXnb1MVrGqANncyelQ1kS6V86JracH/TbSw3Wre
Nq7Zbu+B6yZdA+gtrfnHV32JyQF7iwV98BbTYtBxXrY7A3ahAHuzF+PloGn4XCdl
a3d39GBqhtwwcuKLQUwRp0/IgvTmza9T4wkS+jFs9iK1ILWTnDMap1F854a+zGWU
xmMKWVX/S8aZ9XFPyP0oL8+VeSL/yUwbg1BzVKLu5pf479mD1NDPq9ppyYkSJ/eq
v6wvWcklLztcfivWzaAbg7SWsWS2+hfWd5Lb6Fm7NC/vEl55uLJIy5zWen4ym8gC
qOPQ5ROt+RtJkY3BeJWRIXCQOsNEfo1Xm6q4SWmtC9JSH6FiLWfA1i5X/4+nSmYR
nL/+qh3Wf9Xg1YxH/TSmCqSrHXfXacfZ1HHMcLAqfQ9wnKLB8JIrBxKaEIGZRfAr
RCVKxFjvdyI7eF3wEWJz8qW9fQH4P3mc3EAIZvrDgCogX2S/+DUacbhKLqIIa46P
sxsF2IXLcXqb2Cn11yj2gv93AoDstspS/j3z/GDTaM0O+QBYRV4QfS8Iux1go2j9
xKXJIPUEOxzOPjOj3F/bd0eCYYBgdvoXiurTC2njbsFwYQsK+TfwPSID+5t5Fsb1
2pHgGLPY/qb+yn9CJrE8JKim1I3XOAOCYc2ok47/yXqo6Ruo95bU2g6tgBFmJkRe
1XK5Nba3pmRdjgq+1Z5N16C63EIB/FDNSGBb3RZvUURZ5YdiCW2Z6f/tl5iMl85+
e6iTkAU+bfptUwt8GMQhtpzI1DbrZ2IBQvPXTFsTqvXEhUasDKVHnkZoLhdTloU8
lMOYtukw4YHQq/p2aSXNmYyovZEqlGkSuRIIwxvjGrdq6u3oc2XfBnTVzOWIqHfo
pBTfRC88uDJ2DWDneb2lMhy38j4mBU92qdcjxQa89IWodk/lLc/ij0NvkZtEAMgy
m0MgM9og4RGtrPnIzZEz0ss1M6Vua0VGCuyq51RkC2GML1pKgzVUAQNoS+IqtG4w
Q5h0+2QjFsOHmFYhVyZuVsS/LCRXTmnFPTvxPgR9N6IoEx+6MdkDVCLTUfxLfcMm
+rmZiSzBkV+nQjNoXeBPq9HhzTnz/B8cNxozhHH2snHIJ33TlKILvRs4pMoOsOTd
vUvSnm7vaw4wedQ1ddN8ANTLuPaFXY5N+/Bf3wEP/eUEjKyJYJXc4PdIBIMlxXWv
Pqp6pm49Dz4Om++FYgmhroagLCoupLtAsUL2SVIqShr2MZzYQZTBsd4ck+28Gq4T
quTolu33K3Bmw3gHEiJ3Rdxa9ypvBp1Ubvz0YYawi94qk0I+vYkh924ZaQykrmMt
EhQSJgTafoQyB0AFZh47tn0TV0SraPKChhSSuBWWIvD7JEhyBC5cm1vm6qP54voP
7DMWVf+FMG3UdhbWK/QWc7PB+s7nY/nVAHTEQYfbofIWk6oKaj6bidQhykiR7UYU
VxjcZZmiVHNMMr40gzHVMz6vy6oDn8RwmlB8PbtHOqajmbirrzhPNvjpmhxyDjmo
2nJkZ+SI+zNcUdHuTi/nAGk9MyUu3yG6pek0cNu5MSp91cTW7p+IpehUChtiRMqX
jmBb8IOTwJfHFpiV9tTGetaE9SSKmwgGvFylPehNQdAmTNAA9gVeeKCJdI29Ku2R
dXT1XrsePzd+kcxeB9MnfY5/96N+dW4u9vb3CVxVM8fPC+bOpcOOrTADDnMSmhQ1
3qrI0I8mEd/JkDMOrp2dmvPM8emyFGC558VChzdjgph68GS87EUfaQxxSDfjXYMJ
ptAdNrlquMzIYH161KRMulx8Y/NsUvGo1JpyOUBmLV2ICdMeTYGWUKZBKX4fqVp+
7WwmaODH4pYcyjwIs75XA3Es9oVqWN0HesTwpQBol35D1AgIpf5PugtgUkQda+Aw
jbfycKeq5tJ3Id5jQWQ8lQ+DXk8BE0xEzwf6Q5rU9HGT8eskmYMX0GCTen3wolG1
YKSulfDJuLhpkn+knoatdO4+3nrK4tTzDyNjHiXNytqwHBEpoPTotwqzTW9r4NDI
trIefANm25aUbR+CTjnJ7SID6xcbLT59FCmxbSAHG41BXM0O6ASF0tFowbfah+ox
mPJvuZFujhfmjcsQ7bdKJIMGF2gb4Hu6aUSZZDfCo4QOgKtxyqZyW2boq+dthDPZ
NdsgOLA/q/RcV4mPkKTXmf1mXSmDJN6biACvIQdvPCNNrV0e52AU7NwRf7JwEDMk
Sowvgc5cP6h1+obINJ88kgP+PY03CLA4I3lXIYdf8JSYsi3gCG8H07XEwmigYVNb
jqEJjAbIku7TRyr+Q9gvqfD3ce4kVChYh/mxitjtaNQSU3hIkByNY7yUEblG6Jfq
6JIvV/YW4qFakevItaVCzbq6Uhgu8DWnYmk43Pw8NaVJJDNkKXcwz4yu3TLtlt6n
tsbA8FanpRNh+UPJphCs40V6RgwBvljQ0OK0OXA4LFA6uSyBJz6VRTL9IhlaiDHD
T+Ey5F5eZ2kD0k0ny+TB9nyq+G0VSf5358BkCVGtd86Aaadc/GjDnAl5MfUZqrmQ
R9qoIwrrLo0ZMwzSEsV9uDmiEkuShX75yb1ZiELBA+smYSXuFwYtyMGid7yYZVQd
DPILWNBWxaLDaLz2DbV1dSa64WtJQmuIUUyjptNtze3RkpJXvzO1c3MYnMaaDjpN
HSUUmK0u5nJM/kOZKb3vI7WPWHl9TImFo2/bUj7VxFvzOcNWid5RWcWeS3cTpl0K
7ewjfLNLbYBb9BW5gMP6AolD6amVYcIk5UhR61utDnXulaBNYBH1V+citPWgeWzm
kHTdMSKFE7ZhdVYId3IR7dleuMlpAGshoT4thX649Ckh9vyzv8TD0F6cDSshfgU0
jEnIAXyMTRAag+oLj1KT3hL2BIUvOGGb5CSUvknj8XmDBOHfVDnz2QWwGDwtxuBN
`pragma protect end_protected
