-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wAGqNmU5PPMT7zwzHmqknUNoZiz0EFAy+IBa1etuCtIQcD4+nfWdFbEFZFt0QGzkXkUrbe+TpQ3W
i899CBMIudQK2QAkAYNylBGqGiKvEngkf+hd1X7GZYsvQ2JXWWWDBEcHmFQw+ED8ZfW+eBoEZJzM
ohjhgKfUz8DU5LNcPC3uhq8wdBq90R0SISgpGU5OsAPtmMlS7gCIAd6UbbCR+z3a0JS8zUu+i7SI
0+a8KkG99vdp6mYmr90hCL5sNn2UBLUGeRbXDmWjljMA8EOhzqHVRURoH3CFbWlwuLGh6ybl0DfN
kaPw51WmPeP8jekvGBMQOiH5/wesmPz4Hz989A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7696)
`protect data_block
lOONiodncZ+Bpo0/aucN2pk49cr1MgMvILMTOOUyzZV57JjPYGK4zxmXi1uaroAzLc/B5mjQJttU
8YpukQXucxvGbf80rhjv0NFHCCSSFItHtH/wtVDjW7apifbkQIFh1fnPM11qTWAFJy2THaRVxw0y
YssR3iRDFJPTeuGtYy9BjGSwjrw62MTJA8K4d0l3AWGdLfWsK5s0szS0wq8UxaRpdd2AzxrtuLsl
KmZa7IPQzSJJbNsnKNoTR1zI2gb/NEYHA8IpKKxWSzFMqtzMbmVPXTtYWfqH6mxz6udck4dVpAXm
y0Kyqc1+wzxMgT577B0jTaLiFpwtE2003vAMoOhOHCzyFAsocD9rdwODAdmFkzx+QBGzN2XpMdLr
6MN8Q1yvmxe+KrzgKopIimoLCbgqFD01U5Pz8KbhKxr1WzqB6gon3Ufv4QYxAyz5lnarLfmqJV8J
BvrrKGvHCoU4RdF1k0IWyAstXiLLLLWz+F72MuYCtaaEY0762hIpOIslTpE3YTEpX04UESrS03Cj
anJC2+jbgVEi9QLeshfQTGRDQO4G7OnvmWTCrCUzdmJOmzFsoV+2UB9lNrkadXo+YNTafqIBp+QJ
cTszMBNB1MvZ9tlBLOUuDzwKLG10081EqxLnVHhVjplYqBpEX8NfPdBatw9yQjI446Znusooy9po
tVooVgn++lpoyH1KUUGuokRmxyWoJQqnoI07/87W4ZT2y/mYSqtVhRi+gx5FzRhwm+nWx963lNfm
XLH/DhAThNoKu3eBF9rQjr44NRZu0kNoI+KEVcLqfMo/A+/GgGyfbd+F+eBgqU9W2cFllSyCUuDP
8pQagOUKY1rD3Orrn7w1T4gmDfOSO0W8jp00hD1LsuI2VVqw2jmviOMGCzgOKkRnLg/+zwpzMpe0
Ny/bGFimdZ0+zgjowCmzfgo68ty9d+BgnCpiQUgIgoITZwE5otUcG44Lq6qUmYgEnt11abMbRoe/
BmMCxcgyqSAHNBZbW8fgi8f/JwM+XNJPjypUZnFwgATQi1G3dnPjsK/M2TzKt2mW3e2WJ9rmxCve
XGhHfoM7F0hS1zRBNLxxvaOuIzUSy2DP1W7tiFFsLNI4++/lR6u1X03aAgK84QeQEI0tFsLeR/tE
zPZtENwsmo4tVPcbHIH+UsgweRX6jUKVUk9zux6L0U5N7autX+b5oqk98TBLiQo9h3QyOieGEvKe
XnqMEbObm+gxV9TNyJ/wFe2SdCu5EJR2kgTUlBQaigo39Z3tmgz4KpXaW8tkUQ1kcAbfCuDzOqxH
FyX9ceq8Xjm/H6ohqhSzhDls4qHW+5VHvdrVoETiM+Gsrp1txZYyylEgmBzcCZYQQ4zDAVX4+q3h
QnR4xnCvICYcI1GerXHxA45kRRWhrkbGJ7zonJd+Hv08oB7rP1OYm3vAmIF2d1yT3RY94juoBCUX
xKP+L7fHnB7GYK/KkIlYxgNGxcpew1GQ85WvLBao5te7dO7QtjqPfiyysMM6R4i9D8yT5eh9sejX
xGPN2DYodMUMGBvdoxuPM6wf2QZNnlJq4v0/7klrN5FK5DCntiukt3/+b86bpbsUM0Ia1kLEq0Kq
H45Kbi8uIJcx2VK5SL8ovzfftttnuBAjBAXhrP/p6qQylhqhiVzjhP3IUfDhZ5xUjx+DOHPjCM3h
C4VV2mSU/2G+4PzoLLJlKP3vTMSr6AzwDDBwrHMKzdFPMzuFnRUOG+WW5Dkhn/TW1MNiULkariO8
5KYM/dNYbD7CNpAv9yO1MzWg9EKv2nkVI0XuZzdHv+IbAInNalfdeUx6XwI/xrNAxvaWduvgZDBY
HYZnm52g5cQ0FTQx/FnI+skTbSuWdk/3u13yYLz8VSSpIgpnz3T25JBzf1M89iqqsp6a/A7gGD+L
NqOlMO6uvLvIS1maTkfpHKTs0AvxR79Lm65bZrzYN/baDXkqv0sVpzW5kYT6X5MxjNKfm6BB+VxK
saLWJmadIeyeyHU05GZS+2KpJ56PIwCrgJJqtnPWyf4OUTVNmPk7JWDdK12ZV9wqSnzLg/TfXscP
83CTGxirB35EuPjJ5vcj+65m3SXVclR5OGN/TnRXq/+UETb+UZpHEJ+uYCK5nbzGL8FD4lBkjA6n
T8rljiPotb/RKX+ZcQk44BMPFhawV7T+chalTG+OtEA67RYcbKTfxyhgCmhsn/uxaBnyWfCvqBD+
Zoi0E1z6JSZzI8678rH7iExQrAR4x05K0h5HJ/r3Q4Rj2ROhLQdpq1E6Mj3JhFVe2st/dIR9sfPd
2x1S15wMBYcwzdOcttgO7FgjQLyAcr8M4f7ddsWv4sg/M7+T382qd7oQ0T34Wskkeh0p5VnyMSlL
A4KvVVDpkU8OJrCyeEnJYRbrJR16XB9OdM6jZjzGfRMrt8BXFpfHj8k7qTsKnrSXprKMdndPaxod
Wd5z231SPMniItJjwJZJ2DHFsq3dRw6EopHSiOTAzqseCsAo3krKn3gA4LT6Czqk3oQRtcifHc65
F98ISjNi6rELg4V1kzcr+CUgbuwV+i9+dAlkQIptMb/evkmM6vzZNGqQldipfvfgozBfGUVSNw2o
6QEa55xPUk1++pf8APdhtDQQQHZ+FJly0qSmctk0Tqu2/mq5TTVOHq5/INx1xNTLq42omvYOtFdc
VbMqWdsqr95T6zfxiyHOIy01Q30dOim3PL3aWCtGMOaeksQjdS1CuTmrgQoCPbt5z2Ai4ljujy3A
ff74kSrO2xJR6sC9ajxxOELJ6IEh4qbz/wqC0BPI14hK10XnalAysMYi7SGCDgepeeYW/Cw3O5a5
IWiM/943GosL588TELbpOgTwChieojxRXytkiD8ZlxIErL1moTRHc3f+FDXa8YJojYO4gKKmjXmq
8ofPIXkWFaQ+aQHw6rlhu5yLY5aXwvV7VwmexjdTjnqSt5vVtd/Ik51kChPiYrlQamivxYVPGYXn
Wmw69gsu1V70JtI/fcgnvNPgdOkspO88TEtQ9/haYulNSDactu1l0WIrBwEwd2LMZ7Lx3Cn4FlLB
NYiZow5gtGXGQDF7zIzG7g4Wtn1SPqEJSEzHje8k+5XaFwsKQaxLB3/YKqVwwPsPA6nEaPRLtM5N
udBXudQi/XMToLSzcoM6CgV6qe9w0PTM+g67YSRFwOLlilrBU+RQrZGAPxa4gcKTXCZzsEl+rXX8
dSDJGewc3f4gx+ZMpM23C4nWQfSq5VgVG4xWaqoYoBozdNERIDJOWyx5gTOnabGUjaGfQBw53ckO
UOJTeEqqdKlvwqVaGeYHz4ghXt7TuNOI+3IwlnrwYb6LSK8a7N+TQbu2AVdFdtGtU4aT3LaOPIsM
xyOZUAso0PnLz6SV2aHRFEDBsk1vD5jXA3N4avwKQOsDD5aclqkE1milAxN5RByA1aiGGCceEMsB
DtxjOXjFEocqhvMhsMc97pWMg1lRLjRj5ui6Uiw4E2N+bzYPLUqg3OwGHpX4fWXBYYcB5Wwjwa8r
LZGhjBSgHHuzJ8NyyLTnoexT6YXxxtM1zFxhGc0FYj7zkdZj/VA6OovvKrnFHnR6lEnX9+5npyJt
Pr9araMRo6qMRhUuOmxGReWOe9Strk2gimwLecp+m+zNN3XKUgDR9k1f8aqPf/JNwmvuqEt3D9x2
mRy6sNEfbJr+ovgVcZQQ69VoHG5R/m/2eWNuXEhU/R80W0lEy9ThlHCwY/j07emyerPAKnUCFMw1
Y0svbwtDavk5wqQd0QdRi3STHK6BSL1t9CaZnGqusuEby/jLTSURJbkeBSccPSflDXR/Olcr7mXI
7pMXXyaat7gYDyssUeCclh+Ru3cGiQ3I74Y2n1F9TQPk5wZ+IOIDupPPb/BPXRLaifhh5cILengO
6YRjfHvafsWgCeMXOYBiyWwpAaOgfAXP9Aa685nEPWq4B3u2nyZOBoiLY6sEwsDBv/7qc+NgGYYf
LxlVP7BSptX5R/rQaHfb+TCJSE6jiSAV5XkYIT6A/cnxU41hF/beN51tSIW1M9FCTSduHKIZEi42
ZFj5JxGp7oGI5EmQ4FniEisbSbGmrIDnJIkHnsx93JT+nHxzM1h3Xe7ks/JQRNN8DGS2oicTOXtS
e6gZbmT6vm5la4KGQNU5ByDRrLNg1+dJd/45ETTw6ulbb88nwbolNjhahdFSTow+kkfHq9fl61T1
FBsVPcilXqEIxzefsHoabzd+5PEyAuI/f2nx7rwgeRiCXITR6eskjLjRvtCDE6et7ySG09VVZ7r8
T3jwyrSerdbUesZlaeb4pvnukRN9X0wnkgi7BvNdelUgCaETvWt/XJH3EudF6PketY7SkcpMLA4K
f4cQcVOi8dbmobbvOY0TctPJlW2Mhcl2lru6xPuKwniCMlGSKIkokR0oQG0vtJxRHJwqe72ssW/s
cNjokyL0fuK8uay9KeNnGjztLwpTU2VPyIMwFBbZMlM0u/lHWeksGrTg7nOZz4NFO7gnW8/MIfDA
yLm27k8gCg2rgy2kWz9mLyLIX3Vk02olofE3xaHF8LmFWOgn3TgN+Wxm7LJrdX7Vnf7HGewTDQww
lNNCXiOttaldqGRK2/0/Kkfly9ER8iXmufgE6oHEK9bjjO0dT39eylFGeLxaDoUKJB0cXKjZyBi/
0gc3vwXhME+5PvxNyjES/kmotnS33sTuz+WdiNO6cYRpUciHR9McrojCiBvhC6pSBBDPvriV24LR
+/M9da2AkjtAEWDCs8dCGwJjpR3aOcyxwLehBCiATMW4puxhUPuMW/AqGEFT/vyJC79Um9pHEJng
homSRxpl3kOe4a+EJDpXHPd0DMRiZehbIguyrMASg2hqTbFv42DQVq0g+ckJaewY0WJBhTtCK9Aa
rlWd92alSGgpPoCJG/USqfyOqZQw84NtDHZVwrJF/+6ZmnY1+s/W8pfiCpbSfMUsItElqj6G5+GC
+gupNdxuV3SeFJlczaG4WSoPYS65m+uH6WEDkyfPqQPJPywwbhjcGYHFvgOAzCo36SkQrGwZGJ09
5LfG+ZoDS0lAjjmWzUGb4ilK8QfQcZsjchtYnAWenqssfbBcfLvTvd7GBlJkS/R87cWDGmDOj5Wi
Ihc/2zvmUnFkSZchiytu+ype+ZtOFpOCwLxqzk2Yj4E27lsCLfV2bmhQPZVbS9u/h79kGw6gQCSA
Bz+IicMyoox+5slq77HMMnvrRaOHaU72z4AG2h5E0Jy3yLMhic7odxfpY/IED5lHR2inssHHYs6o
4Id8oWSTuYkpz2X0OeD3qg36rmqkYYu8kUoZMF1PI0zQMNYCNBJ1Tks/fIthalfrqFy/E+3Sz6fO
bd5KOHzH0Gll+RCTmw11tRr0qGie+72JOZ1Pw2qbmNCTRmEsUAvcU3Oxl5BsbdmD9nGF5Ef1hDvz
fzcaaFCBoWIR29JSCmzUZBuH8IDN3hX9AJ2hN+c1Iro71S6f9O/Rt5SvIEM40iPLqXxu58KN9nEn
qjaHSfOeMErdYDc2+U8HxscXAUzzpsr6Z7Tk4QVf4KXlA2J67IT112V58SJ7uocRJcwSzmyN0qbB
/2kb6wBqiFNXswbUCOYRFTiPUrKjXlAu/yrzgicqFC5UR7EbBDiLgGSzG7RTA52QbnJm06i35JuM
NoNvEZLNmnDJ7AYhHK/y3FPTU/qh+aGFBZwuujqoIh9IRtSsFm0TxrWWDgcblayoVD/ZhC6Z21xd
6PG7PoZ+AKQAkrUz6hcGO5M08hFvxnpkKQP9rll6KpeXaUDfRSsNFroPeVba21EzUeFnHmIHUNsz
e5ClujrGDOScpUWYXt85N6fXfZFuIRJZZehUtLuRtXNPNvwanetNan8x11qck4jtwmHsXHZ8ON98
0KIVxRkSARp06R8MH8v1xYRXCdTUxRfwd4pFBliIB0Az5ZMctFwJHBRgYWfIjul0MmSi2Oln8VtL
C5knDIypWNWLREq+bJxaJmIHd/RXlWfxZ88vHqgOU3nRvK8zV2FEC2mVfR1GYQ3Hsmxq+zZJR7qA
8MFZM217+8BRhg8NHFDayfxrMjsU6+Fn5yEI1ORV74kG1cgn+F+BuA7dJATDHY470QuAJt/C3lLT
TvaywZOEpjm6nlvWsN6+3SrpPo0T+4VmBPEpVq5CB5O5d/u/mgN4RixpI/2saFRdqe5MElLl1TLp
lVRzcNwg3105lnj8PgJ5PdjSdyfZfB7zeAOGC/x0taFxoi1Cu15EL7Qx8mI+/jxlS8k1gruFQFG2
YE6elHLzb+kwPx5XJt5q3KZ4hUdyv5JMjL1NQ7ThPBWAmGG8PZiwJ+ROyVOWr+/qpjReqG9ZeQhI
FHxOsyw70aguOfNfnk+HOMNMnP2v6giAA1j2XpgNrG1p9GziY+YbLCzEXtU/NmFGGYafERfLOZ6g
01BOL0te/JXnN9o7Z7jdPd+DMt4TTYilvI6fxAu1FoWsjnltMRf2owUH8nxm/2aIRmTqdYw669ft
b+HqaQy4MbgB6uj2UxsdjA/1yks4lXQWY4n/Wu8Q9fxb1wuukuzE00khiELbbJUxBk4PlDqpvMfE
f1oy2vO+NiW5OT5oXB28I8C4ufkOhr9S6zKd/Wg/w2J+aQ7iLEe0SoPJMSymV0ytuvRweaGSiEEr
XdJ9O4EuA76pDa00PxlOVt7ldNJdJ+ilTEXG+rGvLiqd0zh5aENKSOcBoFVhZN8njHWi7ylkOaor
euc1VpPW8i2LhhR5uHphSQXMMZToLrRMMKokLVBI1SdPphoRpbMs/yr9Vr0SehT7ou0NHSVlvcor
KheXdJ31ztwg096LF4ZhO3//LGCcUuweL9eHtq1bN5rmmocbHQNdWhZNB2J06Ve59sT1GWRq4wgF
GALmIkvTnNRF5+8RPJGfxrq1bWjduPaTH1ufi8Awgr1sDgEyHGuRs+YUs9fge5FEnD3VOkQE8ggd
oL+IjN81cgPY5Q4MCtzpRSa6R8G5GaCWfRiMZGc2M9lKW6NJgycJ59nuoEdeQjVeVtnec1jCbqBc
7LiwbvUHRjo0JIg4Pka+0vv/8ELetC65rxWFk9Xzn2ZkKLgXhXm3fGPwO9hDcfzRlzKJnz2XoMVs
P1jeMxjjAuHpro+fl1mpAlUqCouf5xRXB4LP7KUaFt7uVkAnh/RYBX+BziWB/9Z7faOC0xR61SPh
+cUn1ZsVMVL+SKYNlTO8JNrJCOmVeuxO2xdU6ZAS+RBbcXFUhkmbJYhj0lm4aAPPMld423d97E0n
v0l9cdqTehW5TeNVuXRj4fReCYdh37t+Xl0+MFOJPCdLt1w+B0XXyqpkmxM+8WsUDBHRmewwGcbA
r9EHYeVOWAfJhJmkbEoxgzhpjzDlky0tVh2PrIdVbeZE2F3MK9mbKNNuqmc8/tpGn4y82JMZuc/o
Mhu/wMy8zCuWBM/JmmIeg9V6utPZ86D/SY0pILko2TRR1sFOMYxqIBLceyeKKCAvL4FD6ovG1fne
FgBtD1a3XLXUMC1T4G9sxcLsYaGJqUBxjGBwZZaA6aVraYYw8A7LuCgLUFmX3zFb0UBX41l2BPq2
Lswodb4e20nahc1NuKttu8slFFLVSp5RiCSU98GK3CHB53gKL/X8M/9CSqJWCex538mLXkowN9l4
YSUxYBWXcastAQrIwXNsMVG+sniNhYrlJUqCegss6RqZ/O506nFVY1dZ14wm5Dv70BXzrwiDno1G
It3GhtmNRHj+Pz5MkqIUIs6SpkWTO1ZCNfDY7sL6MZXr0eAqmUMEXBhDS7KbIZdChDUmdeWGjblB
NRMfChDy96JDM49b++d2QAOwx8yQoQ6PlAdghHaFxOJM9yJVA2q5pgLh0ePtzW+t03dBewscM1Qt
S2RvpY2AOB/7D1OZveLiXZN7S/mSwjYybkTfapH0v/LMCZD9auURNlwe4HeNG+mU305kJ6eRzYHM
M/7TOFN/bHDOFkhyx06LRuUmgVfpoifjW58XVqm0pTc4tAKI7x4Q7pHGf314R7A0jhJoaa7TseM5
nHiy8AgBacDFNlKVO2IOFR0QPt8ELUBnM7qr0xQrsEIonM4FYzo7L/uAjbLps/N6Xc7YNviGduW7
h08hxiPDNeRJoXn+5PO2Ij37IOE412ULGSraekrqexu1xpY7gk8z9nr3IPExsdo7oP340CjEHcjv
FaUDGYifVoec0JvkeknrM50iMGQkk0bGoXQulN1i4TRQkfpEmReH4I4fVLbbTY9zQ2U+j64dOxBu
4La7rVbqnEb/d1IoIQuaNC/lAiV/RS+2EUl/diq735VRSsMzBwxAsI3eoeFJEKc1Fq7N3/I2HvXf
TpUQNCpVqKiTUoUbV3nPOqhppfqP1iXmfWle+N1j6EvvzvFqmvuc+cXBioish1ud9kHJ0zGUWdHW
8NaTkWKaKmxO7ge/Htex7gM3/eAagBzMAoGOjhvdR/SkmHr8Lw0qWEbdpTjH/8nvx7C7zTq2/j+H
2OKeAOOu2cq4MSRPFeqryiKfHJVR1J5dy7k5IVFTDp1YEB8LmkYmaLwrOF0yH31aFc+POqydjuIB
f9CHBFqvF6Mn2gHs4HgOwz5KibhPy2J5/PaYOyaY5AlnRRSetj6XPqaVHtHNSrySwYFB87G25si6
xZZn5Qc/ZN87HoosRP7S24okDxx6dSdEQLNjs21ALiqMVe/d2SS7sUzhQIFvJ/M0xMqGMX0LHxgf
sxu0+NoK/4eHZL5WsnSdBQOxcACBEIVfxWXemEkBtF+EUrYNidk6V3nGIGbgjWELPAO4oD6vevyo
NfNM/uibkUfHzLcVc3D3X/nyQwcLnzdC00o08z/LdzkexN9FmSGk91nL60FJbP7lZPhoQ6SCWjQU
pW2CTQDdhnzxs97Ad+IPYvzH5/btzbpPNbklZweg1XLtNcRi472STfjD00YX8LDMon75QkkKBG00
MaQgfG4fBRzuHuGG1rCje0A76BXz/KMYU0rN2C/I1nabCX9qhGZbBFRadJmY8j/nW6rbwZCsy0xL
J0BiRy+sFSgmDihrHytpG27CunBcNESCNaIJXONpGGtRm3vVi6o/b+eFP5zEqjg2b2EvuZgW58mx
9u8heN3Z0nPZLFTiqmOlqtrh5/aMuOD2acQ33GJotTvcpZy0M+AnloUdFtQZZAUz+pmLAD6XukXS
jJ/mEEYEQXl7TAkUlBvUElW3Oqyedm247XbyiNlE6bPQqRtDizpqUvfHxktO2vNFuJ5NtBA4Yusc
oDC9aA4eBkzp1UBL/3UFpe9oK55qS5R1vvspX3EsXtCD/x8w+K58QR0OmQoy2jXnFQaWmMxhTF8q
snhlgonYNG8Gt+BEqLvrZsKMt7bJp1HsopEWOlLdeo63qt8B3Hr2qTKRddEqbjoLug4o6LDMgYtW
Zh2wR/ESocRYkec71p79FBUon/Tm4BEGilF8Za5R6sMlm9yozrkNXpdNN+nXDxMSkfriQFcDc8W4
yt994zmu82SMlqXY9OlWqR7GEfPp2VKGVkrDQW8srZbuqmZtYc3yfuUys1VZNpUeYYvEMEQFLNNZ
DZWnPa1VZ+z7psZQiFkIpKVlvybFWaRUAiu4R/D/NZFZ8rl+WEItaBOdyScMxXLp3tgvcHOrbPFr
qK3ylAjAdVFZbks30RrodPee9gFbNA5xu82zYlUQ5n0GRbBXMb/YuoM3/eQlQWxGf6ZY5t1SILe/
htsMTUcz5sM50GZ0ZhfVlohIV5MvzcM2des5FriUDx8AIr60ufp7+u2puGNuD62+7Aiki3njw7TN
k91o/mDyVluRgqfYHdmEdCx1anv+tAWO9+KhdbO6HUfh6HiJ8k6wbfZiP4NkH7RIlsvecxVWJ5Lf
S2toUdyJ/J6J42Dt3JHQNF60Z9QMIG2mPnifp1H+7EIQOyY8Y8WR9y7GVu8/poEX407/U2MYVS8R
xJg1kxich65t2AjtzVuc/k3YzhKj0zz7AWNJfCTYm3eHKDKgkAgjGYnhllJwKH1J0QJb4vJDxURb
H0OMupK/lIWZ7F1rueroLERBu1aUrRpSH8cpVUatJZ6nwIkFS1B4LgTvy6otARjXjN//LbeAaByq
WWcGb5zQjmCBc3LJJF5WNoihd5h5GdxUpyCeU+rPKmE18xcCDLKODC/c6TvD36NZi9eCnYEqMZCa
+1OnI4CJIJDxnQsH5am5DMvBfSjx4QWDzhp1GCrb6pHNSLPip8V/P5e8r0TUcYEVyScN9FKirJbN
BAPVZnX961SUxGvvEq4iMFff2b+rOHj0Z3LKUvikVVUktng1yy1TCyHzQbq0l3L10ShE5gmeUMU6
AQ==
`protect end_protected
