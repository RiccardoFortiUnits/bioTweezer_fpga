`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pmt5bdFaGp0wooMXgsRur2yea4piWqe/G7fb6qoXSSqK34UcTYuwjvHU4vGnBojW
elBCOuK+KNbhQwJrzNPLbb8qEJ2T2zJFw0/g4yhrLSf3pJjM3JM05PlivFbTP8VC
hTpQm0Gjv00yKVoLVr7z8z3Y7e5BL9TAm2W/cgelUBU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2224)
wwanL1fL/PohFo1MmObCX8U5oThijLNrD/LWHD82qHyq17Eq+FXF86rBW4ifLHT6
yBDzREI9k+5DfHsb6bn2xEQ7UExC1J0dL+xD1uuaoNJ9VlFKsokdiFnvn40kmNLU
7ODE6ODrVnfiLreaAj1DGDr2XLi1WmEGfp4C32xV7IzLSqmezdJ3qqvr0FDBBETn
uZvQz3eLSA2JQSSGXPtxBcsEcaEAwE1vuKARvzu8jqbBcUtbROZFPE1eaEY6hzH1
MVfDHfBePVag9ERD7VZbGJOpnlytfWfsedohIgjhKtU38oxZedbjlQy1+TZqWZ0/
k/Un9TdmOWxyguswimP85Y8GlXfAdlWEW4xaM2gEVf4eXmMrNKtVervmWzqLLz4C
ZJJOp5oV8FTJeO7spPj8Qj9vxSPBLxHYzwNjlpfp7N+3kILlIiICMe0JDqjo143a
/nkM0FxnTCwBLIIlE7fp1SUl+8msfsz52lkTcwIibfNyJFn4jmqcDgDUMoDGuAj/
4yZsWNhujeN+Uyep26rjwuFh6zOPRisH+J/zlXOnYl7w9ZTLQsV0pf3P6dsp5FfU
ftohhT9ha7e11QYS6i/YF7zmQ4qrh8+1qXm3xauIYNT1ACksrA1uSqikKKaHe1GU
hMaii+ELccAg/b4jFhCfX9FQxMeMixEEWJbCHzBmCaZZNqu7+U0f6Bkjl9KD974o
yCEPaEBcLTsSOUWtj0eLUnHo4w2AtOaSBaSNeCNebg55J2N38rOVmm+ysWqrnU1w
hJinf5yenenYVUXBRAAq2nVp2dNPJQpR03svKFXyMeDUB5VDG0ufarTMVlgOdHfm
bFMmzxsg6PgF+ibuUYeS0e2p93bMXMa7DkRF7Z63nMPEXeV+OopraveYarXlVPQ0
IXkrKZA0ArqXnWnMAOi/xOh7R02A/LaCkbdrvdKN3gqTnw6/WsgRT4La7tbp26rF
ym/uB3Y8aDj9fZkChsCi3p34AFo0HGKMQ0rlIY3aXUUL/+zIj0jTuZ5z3kV3gewp
ZuBPTVLDwWBdS7o2E2Q+sKd83e9KrytPqK0hNTacKRgGA+Tf1Rerszh68dYZ3693
kXhQzmsoOQq4G9/ex8jPF1PxVmT1w33YGvN5AUksARHjvmmvaFijMXJwM9ZQD6HK
/DuOwgqLeLdUtjZJxcTWfHJH/2Auqu/R3JXRUVQ954lWCa1Rv38z7uoUWeZxSbNA
dE0kagQNfSvRB5rhXoUMtFwzFM7r+PvXWyHw6TCWsMeYJlXeu2zTfTEiK/LtxcN5
Qs/NLvzNkBQeSnPz7Niu9BoJVJQzve8K9q4Fz02Dr6tC6nk8QjwWM6JLgmb2WM3e
TRxYuPi8K3k/m6ZhxHrlRe0mH06dMNYQUkcgY8qTpgSRYPQmvWQLed0qyFTtaSAQ
Dg8Z/PNi5xtxYud9nG5CaoLHSEYTJATV5sF0WK8tdzcSIU3q1ac98fwGz95o+Ask
A9/AraWU4bkKzqhIMRnmMlG/5BFtll6HzG3zaTCokoH7TipksPcpGmfoAN/2jdoH
+wThtqA2nCQ3Tm0aADp7+wtoVrkqSbgCz14N8tLDHJ3K89MqxPjl60LEegnXhFy1
hEw+SzN8YTvZq4RGZtNW4DvRnNwvcSRkdHENH+BSRB++M5AXmRrDHzqYB8Gc5cTj
Fjdwkqey7eliTOogs3HrhIZCFjI3KSCDbiADyuo7eAOC3etl7m30nqFs5BAoeOrc
fHTuEgfZBsWqBZ1c07p8ZN7fQT3UkS/zlm7uJLfBLdMJAOS63AA3IuX0PXd9Bz7Y
jfFRJ7rbAdxsj2Z6uUb9LzNkF+uvtTiB712mfloNSXPUfbtZGJr49duIAQYohGRV
mrD3h+Z/isRrcGsBnb/MDEbInjk4WbdIzg/7frt3aLjk+dr/cUS9c0ooZ2T7qcIk
b1B+xPIXQ73pPuAAB+lH1Z24ESvidvzV3sIzzNCVnfNeUKInKABifX3dmPnoGvAp
tpgP+C9Gw3mu/lsu/e9p/Bc8a2dxvME7Nm6j5yAbgAqvYkIuaHJDGFbewQeVYwWM
nqsRw8WwUci7IwI3LVDt7T81VENnCbusCDuGPGZOE1K/pjNt4wg0sKIrVKit0QYz
v1ywAYvPnJNiBqE1MJTE1Y9CNFKcYZ9uFWh5gvb+QghroiVAi1D/692zCUwIR/b8
G0GYLaoRunASYgIMp9vWn37EsJzlOFouC/2QjnQPnZQFHwU0XspHKtdTkeIsxR5G
gI8Ut5k/bJAMjLiz0M/lKDFq/qOzydjCTpm1ZjER+GMwb7lCbUnknByHQ1CXqkTM
5po3x6AF5TH43wEdJnZoXJ5maOkXDjt3GMjPrmNHJ5we84bHgz5MQ0KM2XO9NUFI
wK9y4/Hflvu340p3LQgFAfeGhdk6i4Hr0X+o4j9X+kBZf+28NyFsnKbEWYTCzLxl
af04v6Us4CFq/DCVONZVHdvVlNt2MvK2f9Oj2jbNpqY6QRBUFy+XR8dyEQL1vkxC
KAD5NCST+roF1TP0Ytr7cQ3AsePu8wFLGfwvGQReIZPO+BL+7d2wOKJyRLglRlds
hW5Qe6DhyiTo0Lqz9x2WsgcD1tW2zhU4vFZO2dF2p2axNcyf1/MGiXlsmYrFg6u3
1MusWlEt9kEA+5IeYlz+c3EnATv6dgADqjlMXDcEB0RmKWAZJ0vXJQH118kz8xvM
u+H1Mvv5LfuHv943u5L1dKUxCnqQCp4AUslSaPq162EUCZiUlrylt6Su1uXoaxmi
48afA9rNG2lMhHM5TPCFZBS43A1El4reHbQi/mAV6oqtFxj3E/H1mTT390qumdBu
7iu1llMhm75q1889J7R/CRE+hOeOt2JU3y15chRM1rL1+E5288+X/nJfEhdYA8ke
ydskb+o1WO8U/NASpXhoYdi4KWq3CouHwDu45LuOKJNC9PYPCnWFBgmxbMDWiAef
6R5Udn45mxtoneokATarWA==
`pragma protect end_protected
