// i2c_alt_contr.v

// Generated using ACDS version 21.1 850

`timescale 1 ps / 1 ps
module i2c_alt_contr (
		input  wire        clk_clk,                    //                    clk.clk
		input  wire [3:0]  i2c_0_csr_address,          //              i2c_0_csr.address
		input  wire        i2c_0_csr_read,             //                       .read
		input  wire        i2c_0_csr_write,            //                       .write
		input  wire [31:0] i2c_0_csr_writedata,        //                       .writedata
		output wire [31:0] i2c_0_csr_readdata,         //                       .readdata
		input  wire        i2c_0_i2c_serial_sda_in,    //       i2c_0_i2c_serial.sda_in
		input  wire        i2c_0_i2c_serial_scl_in,    //                       .scl_in
		output wire        i2c_0_i2c_serial_sda_oe,    //                       .sda_oe
		output wire        i2c_0_i2c_serial_scl_oe,    //                       .scl_oe
		output wire        i2c_0_interrupt_sender_irq, // i2c_0_interrupt_sender.irq
		input  wire        reset_reset_n               //                  reset.reset_n
	);

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (4),
		.FIFO_DEPTH_LOG2 (2)
	) i2c_0 (
		.clk       (clk_clk),                    //            clock.clk
		.rst_n     (reset_reset_n),              //       reset_sink.reset_n
		.intr      (i2c_0_interrupt_sender_irq), // interrupt_sender.irq
		.addr      (i2c_0_csr_address),          //              csr.address
		.read      (i2c_0_csr_read),             //                 .read
		.write     (i2c_0_csr_write),            //                 .write
		.writedata (i2c_0_csr_writedata),        //                 .writedata
		.readdata  (i2c_0_csr_readdata),         //                 .readdata
		.sda_in    (i2c_0_i2c_serial_sda_in),    //       i2c_serial.sda_in
		.scl_in    (i2c_0_i2c_serial_scl_in),    //                 .scl_in
		.sda_oe    (i2c_0_i2c_serial_sda_oe),    //                 .sda_oe
		.scl_oe    (i2c_0_i2c_serial_scl_oe),    //                 .scl_oe
		.src_data  (),                           //      (terminated)
		.src_valid (),                           //      (terminated)
		.src_ready (1'b0),                       //      (terminated)
		.snk_data  (16'b0000000000000000),       //      (terminated)
		.snk_valid (1'b0),                       //      (terminated)
		.snk_ready ()                            //      (terminated)
	);

endmodule
