-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NFNdQuViHGGvw9PbNq7gwyzN9WXHA9JQHd8VvbZ2Cw04x7A/kTO3xClnHczbTXRc5TSd+YfZ/zGW
SgNw/ytxO4BkmwseJ1Ixrz9dN6zDgLARKqaLTLsovuSPORFDOSowHuNpGjfeM5sP7g60KScNO3hL
gmwdse2SVmvPLNGi4yK0/Z70EGr0KIdWkgueWvVBnnRUr+LMZ4M4dg0TV9FUXgxSkJR8cjK6ztN6
OAMXBXj4TCTDPGywT9JPOr9ewIJrV/YoQ6dwbnxfo1a2O5jtX6EEUT2Xp9QY9YrKzLR6L1E3uXmb
WgjoBmdaygQVZd+DuBF4dtTodWuzFa9g9ZNABA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114272)
`protect data_block
uhvBv3pm4FVTpapkBCJrNpAbX95OuA3Hn5XfaApdcJ0VlQkdTQ7tCkHJ3TpHAAkxnzQThN9aVKL3
Z4bF7EVP9kARvgynF3+Kohe7e6qd+u16AMs7BpF5mq6/V4XM8RubcFHBXBYdn9KY59mTXmoH3lab
sJAyNp1ZXJgKWnrcCnCjcTwEowIws2ITO2S4kMdrIX4Rktqgrf1hCQKCh9boGYN54Kj569OFSWyH
S+qFCNikpjkFK+IeLzVzKSrDlwyoZUoF5WS/0q2M5bo48mOKcFq4bhZFXyC25wKjNsNkanFn/t9i
Nru2z+qkRO1zmmV7LfKxurLCUnt0pL+wZyEjoB1429yNQfB9NVE6jM1O8NhHgpoFE0cPN98ajoe/
FpkVYQxafdiBjL2KGovLCMHl63JjYW9xSOUMDJAawvJB9T0XSJawwReHy0CEGi0mGxCV9dckNwWX
T6TUX2ZJ1bHTqUZdOnqOoMY4Md9lWCaxClW/PfXoWL3+rlUuPg9NZZHIgC4E405kqfltuT19/Iey
VtThHCnh3ZXrjTojpq0n21m/WGhhesjEksdo9Oxip4YUfYemBcYZM5XdVdSUtscITCypCAzizECH
s1z7tZOLYW5euO3T5H/kjaT2NkQLSoAz52orey9blejqt4GT71H8WAnAStSndONF/vX2/XXpeOgx
sZaTROCgK4q8f5zVz8I7vE3GtNk9MmndGcQqJQbZq16Fe5hQJQbetYAIZknt1JnhgjgXEu8IkTnk
q8hUnxfljxleGxaaA76vpkhndvf7CbggCFMM/y+jzrdVQ08EkvyuYbRRv0G4O4oNpo4H9PFpr1CP
A78Tr0Qt/xaRjQy4NJC6pEctJ2zMFHkds08jpFZfwWsDhlcu+poSTQX9eKa4wC7acWS2tP3y/wcV
HMbkEaBaw/O+QM/xc5OVEdoyV6vziQJNVIAIz2ETjuNKG+pqQysSrA5USw3pZfkq+l1kJFwDevy/
1zaT9yJF/j7TFPzoPg7aUa8Jk9lGj1uk4akpeArJlDQ0tOUxfEHqA9BAFOe5jYlJ4Rytuyb8cUox
WKlDeujohhVPtvDMp+xRcFaT9HGSwmy2U4M2AGPN4O0gmS66kHK193zLgNV/e4OhpAZ/5is2h1u8
I2wtdFx6Y4Qh9sppiFz3RuBRZIz6M7keW5msFbt3VwiLFwv4uhbKQ5ej9rLluD1IqODmUIeLZn5F
nd/YUaXY2xD8FzsRwFcFJxgGTMR/zjqdrAjy1+/uFeZ0D9Oo/DswpDXR6QGRI3vA4ibYVP1Tb6Lw
V+XkMDW83oJE/v5Uc/K8tKoVlkGUwRmti9S6bv2Q32+YR/GDNQmvSrgM3MPVw4b+kZgsmVyv9+hH
kxPPi+9XrUxUTZw80CUFq6NT9NLAIkYxAbwRxcqhXF4r0UFaIVqY41Hde+IAuXnRvSCxFnDIyp7Y
tsi9DPS0jNGzpT3be6xip4MtZtytVV7JK2ja11YXlk+JfderghEhlUcddFAOMxGUPQ/4R1KGldqz
5RHYLtxesHfUJA5lzkLLF23pl/g2Emw0qNStTDavosmJF+eQxs+TYbpQR/G/juz6W9ZRdevsa+eK
3VA2PpwvqtRjNVYHQW38aUlMfuJg0e+G9NW8HPmrzBP3PkZx6WoJsn0c72GEfFzAYcSpiImk2f71
sRUgS41Kbql8KAKOpe5hbypH0G4PZrl0FrtfOTkbSFE9ce7z85k7VnMBMUw2yb/Iu7nTUAnbSqJO
edR1am98E4gYoBFg5pswPnLMO/za46s6qNTF6zxckT5q7GvT9voC2qu5Ce4B0fOq5A2inMm1V7ZZ
+9oM05GSLjTlMOZbvY0m7riLI6aHvUv9hO/11t9zqn3nKpO3RoTqY03Ty4cZvlT5KEPyXnmrc+l1
GLkBv21vlDHfPp0r02ICpl/6805lb6HNpTdc4Nc47ScA6J/kgkKGy4n++n0f29+f2IuheGRJibZy
iutpE5rgwI1q+VwXlt2gg9A1qRsniNfR+XUYiE3hK5Mr4NtrMNpefddDXNYD0iEVKkdnf/wdFZUu
EMblrwXpNQJkM0cPq/Hb6U2crtixy5r4v7E6EDBWLwTzt06BcadlMafY9jM2g+WVuCYBOAVg62Hs
uju+MAbDHUkyZaqNBeCM0d2/K/dJFb1tcS2kI2+eF26gmmRP7QCI6hPk5EXJL6LMteyTPeZBeUMf
qC4JrRiK9Q1qQZEBWiHBMtmhXi257WQmrqalwzf4GQmbAmyPYaTO+F3ULRyxO/8H1863kg1SH70b
ZT7iT3xbXSJTJbzcm/aHuGKy8qsFiChlQH88F9XCfsXggXlgRaxKRvRw1s6IF/t754FxLTrCoMfU
dec/GfOS6ULNNFYNBjDcUoeA/eibESIofOrkuQptKuaRT52FpyxrZdDBKNrp6Y59R/NkNGcCYrBl
rxgXShIpRzSXpJGd+KH51PbGQ1txBJ+bSy7ynqINFyN84iqezNshOEsZ6do9oVHkogR05thOoGYu
RI7/fdlLINsijm/35mCKLNDBY563NVLfePYgkuL7QkU5ydvEoXZjhwF7iykwwhmaVy0ntlbmvoss
7ueepHUp2oQeOoEc10YhyylUws2OFF3dWylzSi5ibFFq6QIGZ5vmhebPvP9WK9RX1m5n6Lrx2+Bw
FhX7EPhyLPHYBvL/g4OzhyEKNTHEkafe5YTtlGGoATlQ6JXBD1uJTG5Sw7tYRey+2cDAP5LcOOxd
glXwd1HkaIk0+vvmdtNCwwjkaJLC9tajHVQ//gzz7kiNAU5hJXlLXV9TreasebLYhNOAt9xxgce7
TvJyavHuoRIyEy6f0Is7lUiCoA6Z1oRdXKWYT8sQ0m5NmoLRJtE6pl91MmKeeo0jyhJ2x69wvgJg
/Uvk31xU8jxF6VbzQUTwz4kn/oeJQ8mugLaOX339raQUnWqC6le9aVaeH7buf2wvSQZrtep9KgKA
/tin9fh01LuetI/cWjnVIHX7sg5D7v4Aou3VcefsWlXI6AI7vgBo/OPQSqjklt7TeBT8yW/E1ps+
6OOvGQ5rORsvnfWTXQtxq6iIY4O//SLNEi0MS3ge8Fjru90X44cjd3zIJbEVAkovee51VvqTPhRX
BnTWg9SeGlilOyrRbum8LKETIXr2rMkMXiLldxcK8ZsIBEOsre27tXKSM9YUqY499lLN2LHahIgf
gvAMdl5sRaYIdp5g7YBO7uH7YgNyRjvUvOS+hRibU72xG6HiV2QKmPX5FVIQ4XT1lU6DuqtSV6/u
xxrThn/RqtaItPW6x7Azb+Wad8K7aLyNaFkauF2KHLwVYm/YU6FLrMDiSLW/qlX84gKA0yFL+zxa
km4f2Fb8YqmddDkzZjqy9A3PzJOqae0/JZjQxGeJRltevTs20gQT5u7YYSpKTCEqtpZOJJXbmH5Y
7ySFGIw2adBePpgf+Eus8xw1QecXUTH9spwp0pBDa1AYhoRQbgSOMF7csPT7MuxUBUfCVtrttWEp
FZVmM6BMS7Co4uQKvhHevVZ/8YR95KrmKSIFj+q43fgesugiK4cfMDOq6An8kAL8U+3gSw01jDBu
dYBJe6ZXIKdg8jH3WO0yrpkJAQEciBnoza59ddVQQlvJQubHG1TIFRoG94m81AFdYHtJvwVkf2Ug
A2K+Tq2aYHx/xuZP8jHF4sRqlveqHhoqPAhxCgE/cZEZVEOG8aet9l2JWAAgV59nTDtuAfurVQeH
NDq0M4yLyKHomB8bct3CgZRyTIlXZxlhiywfeTAXjiBMbEy6uRzqVEQJd3ieapi0zbLbLhDmeE3Z
eL0b2TqdsxuwpXhjsneFVS6HLh07mw0L82Byc3Db5w38yTa2B99n1L55WSbVYegNjOhTQJBS+I74
6u6r5xKr78HZ7ZJIUMRrBsOIKeImKJIPfo/0xXUoIJ5/Ef/ju+E4gcj/V6WpnT+trabALnug9oQe
6jCyp63VEed55nnFrKGUzvNcqz0Pdo4RuksGrcCXlWdZ81gmT9QtYQtfIsiO9x+DbFkwdeOfZ7oC
6AB5vPjemDTJeHCoOrR8fbxWEoHs9LetFhiZdYdkAAPnVsdTm1NYF3wZaAYXtvejbQ637/hbAcE9
hQJ/NZM744XcFj+WTT918hSVbncgeaJX6sJAVpdSptih+km9OuswmuwYZAFoyay+kKkOY5o41X6s
yHPP2WZDss8vlw3dSM+anHJlBEOotwP5IProcJUQOY4Dpj+MDe3HD9RvrRZ+ILUFNlhLmULAOBsF
Tbc5v+MEetmTy5UWrMA1Q/e4Ue9li4gJcp5jT0FbS79qAr18uWIDoHKfQDTGkvpJT5dJYdWwZejX
BC9V1vqZ5KkV68SqEINnGc9nq+Z38fN3h/9UITukzcO/iGQD7y58Tv7RYhe0d+jdQ9LLAx9taN4v
mig7UnxQrkEGH9/PES1U8iCzZDhNfPaGTpOaUw4tOSxonhJMxGKGcbblmQvePSoF00lGVXvhMbEZ
VH/agXT1/Et+jMgRbEnR9ycefnmdWBo6hDyb5EYV82LI639FkA9NcnUOuno/vhBMmaV+1GcKmk5q
Bi2VZfjnA/qK1TAGWBPSt9jFtSW86b8UbDcjWXN8M04koH+AH+2gC0Dsb8Bg4l1HF534rAt3sj4i
nrM8IRAmkwaADnhBc5WJ+0jPs29nzKCW8ckqie5X/F96gEyW/1/6RutlPtUKhNBtjXy9LiKYoM/T
YBsZpjCYCb/iWWCgrhrfDt3qT2mwdZ9qkUp2vgd581gv1u2OksgWaN8GsNyz2ICKXGqwk3/RodtU
3Vh1LpZ0G4Wk5t8/SLJuO5EJ0BW+opMpxWl6EK+TilKRZoIMUId67Dr/L5QnJQU2HEZjMSvg8DWH
dCvhNxZ2ZW9xtYXhjMwbCQMgRjW2zdkL5LhGH1shz22evx+yLYP002uoX5LaTjbJ1JNcf0FCi89/
9QdKjy31PzQausygbx1+nU39kCsJksRtMCdrBank39nUrNoak6CgLzRNROvitVLZJxq7BQpBJCGy
BX5ytufyKQ5qOY15UE1y8bMJjjt4NFfnG+1ANui/yOIYgwrNc+RRRmGGYGFUk98P2EflXiQXHeoE
R9MzwDh3uW72jweyn9pjzKa6M3uclBcH3ndg2B6lAhHCadKdcwFV9zTLwUrSJy4eFP4LSTL9Dy0T
HKGo6FzZI0V8hJNaUJ5ncc75VAbNvmcFWjZ//Tr0SJ///NCaIVjnWlf3AYhCcv6DTfIimUfIuQfM
jlwKRqUG3P7M0k34vhNRVD21cO0kslCyiWpNlfJWM3n6OAAOK8tk4ZINPz4Nq63XOhTlux5g2KUl
CmGiJ4S8D2KJJVmbGMPJUood6aZ/IxqK2i0+0g2fVjgLrYelNUZiMrU/dhDX4cERW0aJjG23C6vx
0RzGb0EKSPTsBPmsR9uj31bjec8F9NJ+RzDBES+ONfDJzJlRxI0xWr2XHtbdghswKYSSNkhX/cFb
xHUgVTw0XuxdjNPiF8OvSrBEqGxKIOAwIUrxpOX3Mj5yOuz1EjlrjQGaav6ldbfGnog+7PB/9aR7
27bTG7LsiSb9S4MsAyj3C0nq43+UdgHQdS0e6m/gxz+WbheEQIdLbMDFWbjeIbwtwqQ4n1yfxjQk
Pvas3zlFh8I4slLaDmC4b5+Jr2EDIs10vcxJjVEUXOKsMSai9q+eiuU1+UT777NS7Y7Cto1EmRcB
K4frCLVzSAHacqouPYzEjAzGC4xD6av9NZYHmmfUPu+ZdR3LKr5AubcJ9uIdQZ7l6o4V7F3hI2dq
BGGl8fRBWigvdOveTBDt/t7LApuwlEhdjlNGFwS5ATPYzb9mhOSqSlhQGOC/uDpPy4LmUccdsnuZ
mbOwtBrDDOSDcr3etnd2iFsamO5+4mydCWJ5+1kIY0jEiq4T4scbKJpG4ukDkLg5bssdJk0M7tkj
1gitg919he2eUJ+EY+v9hhBZ/E8A/orzkZ0V7ihW/4IUgqmnGpmFduGhMYTwMmBnauDsXXOecDRb
XI8UA1Ed2LRl31JXx63HlCa4Cp9UpzgHQ9gUQxhRz2e1b+Tku2QFQEkBYBl3e3nhJnEcAmNiNM9t
N0Ot1VDAbPEpsKhDePU/KMsBWuWwJ/BcrRDGO3Tix2gvjd9sKI8cevSzsJ/qXLeZPfXN9zWmnLEw
dOm0fnEVhUgJfbl8RpyglR8aZ91wFXjEutj8cvBD4OZ2fIWaObii0zejX2JlQniS54N+xqWaIo1o
gza/nl9X9LywZTocr4D6ZkMmEjGnrljR20AZSalm0dAQWpQpeiWPK2I2HFf+cMPKS0t4b8nJj9bW
cXTB+EVWKzdRLRJXGp/Zn/TiWwJS/cprw/KZdi4sAW2Q4Wl366MCGAXp4ZS7E/HBhrpTKwQZ39P+
vjA4fOT6WEgac+P87o8tEsU9vUfNGtOiBzhqHS7Ef1bitpM5beSiF4WJ0CzxjKClZ/cq1YI2KP+f
3J/UkOyUtQejkeELoP9oMo9hFolAjjPRclPj1SFBaglT14gMytWjSRWhDojuUEFWxG95cNVaGL+m
w+jgTKFfKTUPI7GSn/fbNTPyj/ZQOo9wvdWM0Uasfnb32jpwh+v6HiMWTMClK0IZzjyoZYloyfc/
cLtLLhltdqczmyQSru5rwU7PpfAu8Hsway3XeCGQdoga8FW+FBbLEw9LHn7bnW7hOr8F1bm1asdg
4z9YLGDTjVJY0tS+sIKjgXlof84P1fnaNRYAqNJCD/8ZYK414Gprz/oCilem47gnYiFVGpiiIH6m
EgrEku5f5LM397+7eeDMn5meAtLsQec7N7X+JHMBhJJsOD3nmcUneWBNpf7ivym5ixPPjZARQVMq
ummADBFK78UTAobzmGz49eeHLchJcbK4qlVrbwJF8F6LDSA8+hKI975tOqxcyKVE2QNCvVmLbgOS
xwZFwBgguaLIqlF4il3Xvva/MhjzW0ZWSEiI3L9vgJi5PdQf7ipjc5/CvQfz5XyWT/8GjHG1wjQm
C0lU6iHvVFNo1lNiEWOVP/VMx/6DlEIthcjwkwmElsE+oEzZltY3TQ6MzaET+jyOs/llkt364fea
t+mIhylgYXb9GDbmVCmwSsm663ppWGKRXagYPWZwwNhsfGVwY1r8gVs/RZu7F9IrksoSJzDhY3Zg
k0Wgexc7m5zlukaWC5ey+2daGsrpAC5GlZt2IGp68DT6Yuu2UyVt6/stLhWLL8isGfy59NpmLzyO
djkqQjOTtPGGXZl1HHwpVKrcnnVD4k9VtPxp69CL4oGGaFc7Tm0BqyDDyNEOll8Y0LmRVmJ1sbss
zRGPAwJPkVAO8tjzDWbu/36OKkJ0zpsRDPgl3pzVUCXAbFbty9jiS64Bp3pKEbXnQrpBNBFXEw1m
1jBZELwGlqV+ZnGVZKeKdD7bOc0GdV3nRO+Kb8nYlrMUMLrJPx6MuaOGoa8r0Ztq0rIbeP4/tzfw
08eUBxqOikElTwWt/O3jF/Xs7N15ETi6Dvk07DBrFqGIkSqG2kjj4utsOebd6GnturPAqJdU6XyT
ST7fPMj34VVgGv0GDQsp7air8gCtK9vV4VsroG40RNkgZgAtW4qzhBuyK9pi/7S7ZRkIaoCaIOt2
xPEMj1BdldiE88IF92+eAQAUYUoxMgjk986ToY+S7qaIRtErr/NdKB41devPMEiQvbzpkEwB/N6n
9juiQc27/9KTUcNRQVFIctd07UDUMYKxjUKryJrCS0NjqY2ZCJIuxiP0PW9McO9rcvPZXMdgVK4z
4kuw4yPrS61X4dp+NR0HhcpaF03sQlR34cl6fSWpFC5OJbf4unRFSBPZbIocatQbwkpDHKC85EJk
QiYfNATQlEmeagxqRik/0+Rse0bxgzyj25pXc9AhpHxNyqCxi6YeB92aUlsoNuDNIUaiLQIYccRN
AeTRqOaWWqj96JuGjaUzUarhxoOX47f0bEWdyaCD4Ql0IQH/UnCA4M2ysar0Cph3C6qidcvJnwHm
Evv8WZ2+Sh3sUwwO1cj8CeIhPTZIcUnQWya6ehXYX0YX5wLeZ6jcba7XMcKpEFKlP0TCxOgCnuRg
Sd3k0ma+Itczbwwso2VT9xMHa9GWASW50EuuHc5vf2Qp1TbE9hKEvej8LLaviI7tBd4z4n5pefnb
FkfpkZ+ePnu8DFQsvF9ldfD3HXYYYNdEp5dwcQXEIbTlI6xYu5BnDKcVMQBMnZ3vyg+2Oi3M9HHJ
6ewHYn+uiMlHbGeO/HmtVhNNVa5c2CUOM7lntITU+qymz5XmmaHMFvGK6RzO7Jb3fAgXeitecVI+
da7HP10FbwW1bhkAlr8UqGy9xcJ/ca1CSJlBHTuOKm6QJHqd0gZg8l78LYDwpBxmHnpIiyxls3Nt
A3vX0xpKbl4DLg5u6Jb226XK9kMJg1z2gXlA/sllGVOUkn78+6Ve08rkCTb4ML4/aCT6Td3V7g4L
2vTpsDNSbTsWZ4uLEFZxmBS+jktnxEKnGYJ+n/EAsTW/LsoSYkC31imWA539HpsPZ+fdVQXE0tOC
3YXfRkVxbwfY9sdzrOthSxSto0zFSLGO85zeGG75a26R96Q/MMv5l2MtDBctwe2heSXX22urP0dj
pMHQteaGw9mtoq7LDIb8T1SYwPpDQZD3Sq5dSGRuIQ9DozwHoToMWwEit0GmrLj2cz9gOn6vpZ8F
gWVR73ls9JXtHECVqlMfnWiHxGl+02ZChXZp5hhTYc54voVu0O4C3S/JhkuF2H/Pj8PWtcjy/7M+
y66T5ktcoeg6RtgT4L/EWHLIgaaiwFrMTwsp4G03nRxdH4JBqsOP7KanfZMNMrSlQ21u85IPePF8
qHGbub0NkeWZSI7cAb0RUVjUp2NNI61bHdbm7N7pov75iJL0CPuUb/VYzCKZ9o5uSQ34P5tmfYD9
LDAOsq5pVbA0V4QPTtz1QWhLV1uiqOfIJehdJo8Mey+lYtgYv8vSroKaJsDO2fEiQwt8Tw3UARmD
ftWd8/vDxSkRSqGH54xvMCJnnzQ0fSkN8FJVvghEoyzCHr0gTDC0DyGiMO3GHRuTM0Hehos1BzDB
45Xs2Z88I600yMp6wI2YZQh/Q100wiS8IEKTnl2My6ND7MdJhrpA5GOXEZKAUkrqhX0Rj1ukkf8Z
934JGIUzX+w2KJCT/mpxoAbIxLxUxiBqf1xtfVu8UbjtnPddvhQcFrGtfVb8DTJEvT6ILgG9wAZ/
WLSVCqOjob2G9d8IDwf5vw2pn1FikUQqX9Kc86yGjMA80aRt7yaaevC0e6ZA5bs+RxJSTuTDqgHd
/vJVzkqJ3XEGfWa8Wxqo9cJ4YgpNe9+4Oh//E20QiiwWe8RmeK2VnNrwJ06hEeva+HPIZgChRqDc
8rn6gGaIAgwZFDLD013J3oNE7rh+wOECak5NiVzBRqXTc73wYcWFlaQacZCwwMQUMgPor+RgpBia
jVFwoCeLtqcUKDY35CWbSKPaDo9iEoGZQ95VeLbHwP6J7dYsx6V0/QzZmkFcVBhFbLdqAC0c/QVM
k9nB9wphq6ujQ0tMwoBB/LyQzS+Y9wyC9Ee3J5BxnjcHZiD9F96C6ZWupSV0rQfcWAw2hynoz6vn
+ChCRfiZoZKux5U5LB6dk1urVM14+RONk+D8fcy8chqC57EPW/lG/4j2cPATEAWkOTZnVMNFvZ8V
wFPcJV/zSWAxKF3XZnVsJ/IH5F8sWHk2g3jL2SM0lIBrZxE7Mx4BYA/hLYVzPHi+SfWxufdR3eGD
Rw3cjYlRPZhgTRqGa4k/i6ssDo7EhuO9GiqHy2r+epF9BhHufz94nLRLXqUEBvaHPv6iCT29ML3h
vsT9ZXHp9B/M4PjbX9zRv4cXLkMBcWA64vckuucAc9wHp660tjmMAhsUiev2tcTCSOx15RqWzWb5
zRCA8UaGrbAhJIzc3MNbqW/fMpBHhmiayLxiS5x5+GWiWiqJgdYWTNGRpxlOoqKA1vKlzjKO0voK
KbU7wS7pcsI+VO/v/8xL3nCWWPParqly7vAuWUsdSGQLZ0wLoIdivaltha+AweFirMmTjxxQ4sE+
7DWCDi9+HiBa5xuwKbUW81I3ffhix1e0AEFi5l4p5lPPG2OndPHfzT1FvR2yi2EDaBThzsIQL6in
jTkz5JJAnIIMa4p38KvMn3jWd93mi3m5EjEsf1sJqc1667y79bvi1KYcXtGJu9tvDscouDRn0wOL
rRnYYgPpLTvL3Uv6OMMPo8YeU2eSpYbvEX12tNkh3k3+Dy29j8UGVkXljs0Ef+NeCS2iJlX07cEL
Ji2+/fSHR7A5CKbn2zn/cpzPdt/bgXfbmLaxOFmT76UYxJN0ypHkuWHwD/CC30DM2KWfyJnFjdKs
lWCCIOvDCZBVWcG0I9eJUcd2bF14Ioy46j8pZqu86PNP4AY6V2wOCbwu5Am4gAYLHrqQLMyBPPVD
65OUSygVnOtE4uXRrldhjg92BtFKOgfFcR1X8nHivnW5m7NUgdwiJn5pozf8Y19JG8lCSRPvNTNg
vVBo7QVPYOyYIIYodjyNTruSxRADnuncisrMhgK5s+qf3tpdqFog+f/Wkn9B+LC4GVqPonZpg8e7
Ob2DbO2hb/yz2P01RBWCSodsRWcl0K9a3RosXjwvcatXJh78YQPYVQ+vyafJLN8+gyKlHE4qbW/u
aoseuWKAw3QBiIb4oPsKn0fgLJL2WTFG39wnzQBHNihmqfri0tW4fd/9mFbDSvIftcmFHc4XvXJP
77gOG3jqc8DOha/M/X4i1nLz565aJ0h+C2qu5abmTIGXKP2NqsMXst+8T2WOpwfsazxFOA8MZpng
D7soUcjo4t5nmc8so8/WG8vg7STMkZvl0spFKjekLxqMjOvyr4zA5dFHHsQLQZfWnuJSa6U38svW
q+BT8f+PxQkPDxVcq/4KdzP8c++kFvxAoWPyMHTOLR27/k/YCJT5NhQ8UC2z3zZyZ8qFkD0atsQw
KsNc9LrH75xaagd6atVCXoTBatOMN+ncXby/HsPJs5pVo6GuBXz6amea7/fD/lGnkOcI7yOwKS+3
xnGYEeHKY46vr6UgmGmBNnJqRVSW1UScn4HzapGi22m5p0VcKg+RutmcenxuzbEBVMeyNfa2xq57
cRFx/QHuugfAY4ulBYFs4fS9ij+0TQqhR3dtl705egsIOC6myUhIEahv8Ljyguhv1V83L2oKy9y1
FJfJYl970f9MvJ1Wvg5ePxRmphZMy+9GnkwiI6uUbA9g7ds9D366q59nU1gNMA3n92dFiPBm/Zrr
wqWVEj5VGU+jC1VbDry7Q8lPBwWleBJdAXGd6DhA2FHEgamZqyYt8OW4/yD7w3FDmnhB4huH7Zxq
Jwjm/VP8ZGw+LSxQx7RDB2izgwZHIj9QIFvO60eC8kbHtLR3r+dG8zte/sWs9kb739dnW/HKR91h
IJZmBulWOtVRmTgY2O8lkNXKQiv+ORV0OSngfz9i7U39OiAqczrpsCRbDbjRdl/tJYTQSFoijIh3
hV9/VIYTdcEnzeg00gy/JWQShH5Cd8lxTzi64vqyUwn60N/4+m6oeFdwamVVHFVAOrzvxYEkOXW4
VQum+Q0/y5JJCcSYoo+q7R7R1Hianaszx+bd8U8TMf+lyeinO7OoDw1Fx/4JywH2qS9lHKR81CZl
qlwd22P50fhrPzxrwoqkwXa6IR3JO7EbbXHjbrqOO98ZvO/HTBRSdDr1kzeLtKZX1KokZpR5+vlC
abKltJfEmLskNrhsJEYO0ddHWIwBd8nnHl5MGgXzNdJnYhppaZi5SFdSjkrPtj0lsSgjWcBKkqFg
ZZu5n8tHY5J7aT0YHOsN1d4oBfeLrIqpOGVaeF/LCD92+SPNG22hEJWV2uagQyq2G4gj4jaA8eqr
xN7jQYWlCi6haNN4Pzrr7hPQq9tNCcFinwoSWhAhHPbEWE+4oNiRxLzJnHQ+t3EXqaYyipPuYFyQ
l7TRycW80i/7QLAZi78+jb5C6OKUQzXLThXmWHuTdxED3uba/UnCQUKyYPHzWx4RFr5kQeMnBt3+
dlSPIcyN69rQ5MfL/rXdD/1dRiqgynZEZGRI9lv6gADpLUdTDdMag14agg5KiUgTpZuwtFKAxeXO
stf9yHz+w1jH4eBm/OffJQ9rZtVCwFaSPskHzCjMOL4id2wmHRoAnCCYQNt+qEIQBuK5b9KCgWat
4MjKHNb7Ul4vw1fSFus8khP09Id79Iaqnp4q+c4nVE1WU/ouRaqxgHiu1B/JEN1FbTH2G27xNbWG
A4eOjNHnCiznrnA3GR0/NYYkqaSICEbZFmpJe2WcuTyyOvZps7I6xc8q6y2Brrt6DC5OA2f4uvzL
O3hmbA8XVz485KgklZR1LlEyeFbCaV8oHh+0Nn7//5ZHiN80P9pKvKTrxHtf9BVSiTM6tu4ld6YG
V//mfxeV+Vn24Q1vG9sRD/6mLWV0hUqJlZF9rRdwTNlKr6iU9WwYp8o6q9I3OGoRc7oxHOKJaYnq
CNKEC/6iuM0406p8TKeQRAULdVE+oMc4uN90NNUZQTHpoPhDZPyc84bvuEGA4d4Mo38/at8CX0zD
/kxg+SI2HMxTyF7ZRKQUFo3vh7TBiLGdaRWm1SBv37j9lsDJy5qHX5E+OmQV7YcvI/6PE1t9pZ81
7DR+2/SomUrsu38neV7lZjdjGwZveyHR1ZwyqL3GbWUBNMapMFRKdkSxQIqU0D6GmKLGI7xbhkwO
DJ1bbAde9blHkcntdQbhdxt5RnDcsRAHi7zRewOT7mZIww/8CGlYCKmkD7EZW/vYIZpzTrzkQTHv
AECtKkVrHkRiXyi/N5DTO+H/t3HCgqLE47acXhFnF0Y/muQ09wsGm3uReH+gj76BjzrcBC02IIre
SqP9jmutAyFPkJIQbZF8K1DxHHP6iHUecyuEdM/TfgYid1oH2zApFww95ESNQjI8d3/h7dmoorwX
KxiDO3vcRMtlhsaG/aqMTtJwIIw3FnopBhj0MB2xEfP3EcuzOQixE/1YG1fbOz88GR31m4dGdJRp
XZH3frrUN5jdHlcua8kQ6vWhUzIn/53J1IQCZ49cJ4/zo7Cyc/Y6gjvDmPG3PBjSu0XZp+M4e5Ce
F0MPgu8ZzNBTppEXY9351sDJjUsyUAliAlBtjQ0L5ttIqgcssFHndJMGiXcaRp7u0tBgbacMj0DW
8V+hzLQS+cX6HZH62O42x66YMBPNPl/pcGuAzFKbXxYI8LoIXYxJozzS8Oh3Q2AwccfGSO/yaW9N
mLFCAb2SvF1XN0zIbk8y0wttunbrR4hLSiegN0vBEJuSit7kK7Iw8soSfV6xFxUwOku22UQWOMG3
jOhixf3FGA/G/U1p21hm2lZ/naM4oIxsaD46PNN/mo5pLkWQIqPYzS+CN11MRrzMyVSw3TVgFZn4
RrWEQuj5voXosdjDsftWSPQSCiZGTaqnE2ANBheDtdvMOCWFDSn6waElSSZvtg2pwyDPtTbFfT/c
FgM4JD2fAw4zBqah+S2Go3wB/ZRVoxlR+qhnRPxTddyREbRqc3b9JslRuHTR2p3Tef6m0t0pPFxD
8plzedOFi6HVVIrzUtBb3Bxl44k9ztryeB1PqoMyf3BmJ5cJEWci/lUgceliwWmiY3UpGVM1yF0v
9QOhleze9vYWwRpjtBvZ2D4YU8YG5bFtOq3OkrI4wj8o92uaLSqL8i/y7EYWgEGbea/HEdXWgRrL
nySxWopt/4nne9pFp6YfijLaOSg9w/OKR3VPSFxjHkuz5J6klk2xjW2Mp7eioEfgY4sdy3VzxP1U
YLRB+MyZKzSeCmirW/Uh13jDsBEkrKYp5Y5LNrcs/OdcOM8c5KZIq6+sly7gc2oi365aePoYmnF4
lLFMn3E+LYE2w+qZKuPqD16PGvhCe7Xxu0DZFlzRIGZ960RO6k2hxqjMQHODDLuo7zXpDXRfVFkU
BomaVjmI5ypp9yKNbsgDNPhELHeI4silShtzRNHnmX+ZP2qow4S521jZrm432JseTkhd7UTcbBIf
D8nFtkYVLAuyjsaIEOnXoD+Sfihcvv4AxwZLfKZ1HGiD1Y+sVBXyuaUTRXia5VMUhnjZtnsEtUAe
X2i3jU92JBYsPaS/Ra+00glFtdNpsDIJSG/zX3woyDveB3s35P0qT3eRMhAVi/yfbgZtnbftU/+C
o/qKQxtpCXvszlEY2O2HUUznGG9iaNF4ci/GDylh1mohmg4Tbe+gQuk81+wwVnSA5uOfn3bHkI6e
ApoB53Bei9zRzG+537ZJOXsD0f1JZfPO5CgpNeK4mPe4xhcYj6cRnT1r1j/QAod+J20UfADKgy6t
Hw/VI94KZTbkMzEycupKJC40C8U45x7AlvsuPO1k4rfHTzoNWLghrzVQJHh5OqGo8aRrETN6q/ml
Z+tRmiMPcUhoOZO0BZlW4t4XlW+dMmH7FAlmVOStp4JwBt279m2w7B5c71+atrtONR5Gn6dL3aw8
7UCtdXDculKybHcqE2wiSx9YEu39InRqhB+PmTqj8JpKPw50BP7zaV6t9ZWT4cFiEdWKVTTa/JRT
oiEElA2jE3dbr4FqpwDfx/Mw8TSZXVcExrnxZ8jO7PN0QtfgVcZTW9tm1jbOlywg0gPR9CWtJpAt
FV1/lFWe/fI68vIqrjSK4anxQNuWMo26VWj4MEpvxbi9fkxdVQZVrFKkShOP83iF9c9UAS2vdlke
plv5K1SF0Oh695iXrQZsy5hyfiQSvlHD3nFGMrnLv7gXxWkqBEP66PqouvijbChucjOpNByA2h75
AJ1lM0S/L9jPcQTy2nLzZpPoZgu6SfJS5wzjdd3kigiajRyJ8g0SdiXbzmWbHM+nAvpj9gDW8way
Nw/vNSDbcZl/V98bl2VwTEzHZ9/8biy+yLuD4/HlmRkpfqGuD+Smmm4ROljuYYstsDM6Zr/PVpMs
QVR7SzeNUeSO9yY0hDDg3iuzsJhc3ejiZCF/l5vN337YXW3PfS33f31bjGjvF60sNwBWmPp8Z0mU
N914xDDCZKO96sh17M08fen0cJQ969VX5f4l0/k6kVI8VBzKfd8PWuotq1TObnrOz2pLGSrA8b+r
2w2AtLY1e7vXBSKF1cwJviBumSE+RJGeBAe8uNzuJGF5rqz/ezuCFROzBGXsOl14621rzHlwuy6E
9Gt4SZwMJJ4k1s9wzdo/3W6h0QsHayv6ixHloKhjOMbtJdSmB8wSm5OBeILL8WHA/ezEJBgtEX5l
6XO+b92iqlR5fjP6pPPUw3ErU9lEPHMGUWhnRpUbpgkvJQPbRqzxaT9TFqNW5uyZwy4g32qSmVjm
e7nWdyeV0my9FZL+g5XEJAJqaWlOyYISFm8zRKgDvwhUUdPNr/mY7/fXMb4vvuZhFnVhthv8idoq
HEIH2n0HfodMQDDoLFs/iEPNMg/92MsCAwwNg52DIsuaaVEPSoGMBXij70RUk5uXvZHjdBM0Cj8w
GJPoFlwajCdZUVLl2J7FGU5PJ7/Yfpsx6YhvftX+vuNcn3yOuWQr0sGtzQ+FxZOVoWYic+WS2FIz
GU6fiSnGRV/pv7/TCOJ6/0jz3zYzRJJax5yuDW3+HPx72dVah31Kz8JI21ev2H0eUyLcUAU8iJwN
TD5NhgEaYcWEB3gtewH3MIHbdgw3UZ9C1hGKwVf0VRL2Mxo4OzNiXnKcBy3vSQw0L81YubOukt9w
HbMbYkiFLFMTAsTVmuQIMvZMThxVvhHOCONuY+QGjBxT6hJacyvwvmj2Zi3X9iz21JB6ZRbnf4Na
DLKl+tCdtU1aylVdS6Ei7HGv3+0s0FYaqniwd6/iyOnTCcRwqE5ga2oE3Ja3Gpuzxn2hhj2Vw8pP
HB3MnO7o/YOGNruLBG3S1tRm6uVYVHs5fIxL7Q2tvhsRq/rWwg5URtIRgPSl5tPka1bVgidBbo0q
GQ1sX7aOy82Q1cA9saxZe+abSKgXhl0gwEurj/aP+WfZzfRcXtOKpOs9ExORZj5/PiFfawrH9oV6
Xu5ski3/keTbDDab9ZAqmUW1vsUr5PYJXkiWQWr8DOOcmpTm12ksWapd3jdJrddhYd9L2RQ/uTii
0pt9I/XbSk/uNv+LhFBFfadQvIksr6+7g3RSTj1wrka+hQyGENe7e3PzJT4A2TnCGICc09YF7kY3
YfSiaETUpg1hg9Z2w5hGrLqbNO/HbF+OKz6BQ6nPiyFu7ADx1HKW35kOnmffnHu9L0m/YpdyFGR4
4TReeHTQQ2Pz95wyB1adOeJuUowjAtOh5q5IJaP26OaOp8DNLQf3wPKAJlJokRySkaZ9KkCDuLjp
gHT2tpsC3tVTo1v/wRVktBu8ufjto0QTEMCFS061MgK9dTvm511kfUifxEEzTZi5DNVSxpSYENip
Tp9c9XOraCaauUGrMU6nD5IdjXpfdU/pgxxn/iwYjF4fW7dfyVDbdV+iTwa6knIHbwRK10Wd0d8j
MHcymDZ/SeYwh6fGLY/jMMaHFe5oFJGOVeTuo6oCCaYvGwAc+Er8QSl2gH9KB6GzsvkQY7WflM1a
mO09GrpQwTPHQbnFvUiegGGwMI5sFV2ARD9uO1oRE01VW8oaw1AvorRTmOmOX7MEOdaL5dG60pro
i63FCt9TQ04qJhesnCDwEpUxc58fNzN9lWvpguRMkdYmwKaQWarmwvWqdkVxHd2FWdAJOq+RpgYH
yymijokkzrKpTGoo23aRwqkoB+nf84uZppObS7jof6X/o3sWcSOt8DtbI4XNLDsxkEZolSnAAsBd
vjmTQIqCpDBvZ5tdDsD8PMiFu2XiegPMSTe8H6mjjLOHkqM5XkT8SpaTN/ZZDANm8CBKjCZ0OXRq
un1RBWZgK0gFEXj/CNG/JipSUMURw7HxQQjPCSKa9pcvbi/eP5fccy6TVMmW0GucR2YJzXcBsvhS
OMiseuhMiW1lU8q/kb9r6jHl/x3MqhZBRofB3jIIPh2MDV9l3h10drdU6hs4VC1HZyJKfMfj+RuA
hAu2630TCzgP+RdIEwgai6Yd6OPALtmxX2x3wi/JigQDcnHyos5jSXw9WIJjdx5GeujIRO7BB6Te
7IifDryvCHyW/I0E51yonwx8blVaFsm4XQtcuiOilRaLccPq351pXZvGXWAFmDK0CCStw8y/V/Gg
y1BUb7E7LY94NW2aAuEQQyQpPnBtkerkx3c1boR34xdP7lVF7B+aYWEjGFa/Pa0uxeYTCcPNXp9u
tPDAILIXFJso/1iynIy5AwxVWteBBSwTbQkcb5CPj4O2WKKfavLUu9pIeWoCNtiXgm+tZD1745mt
Kf7A6Lfdu6mFXpNCiXNXnGIbf7EK7w1p1nmORcoA9F8WUshZ5ZlQufh/VJ5QeC3NQzjtOz3XrUuK
+blNQHVYJV0Q5K+C8XDX5QRnANxgYNb233bJNqoaN4fHKHxYlOqO4yUtxxCclcN9Urc1x+w75MM9
x9jhJJdUJ1Af4amyyAaY8Fzg5ksjNV5LHch7bA59eq21hpWLQPlg4ensSB5GtL+/Ly4gXKe4/GRc
rLujFyK4dZz6XMcmLiX4Fo8emBYuj6RIRlob6QlJkQiMvmL366Mb9n0VwxRn5SkG2Kbp1vbSBHYM
l5O+aqLFSiv/FIk+aoNfClWyor1ZFpOeUZTjO/whrnwOI/Gfu36IQkSo4DjJ5WFgmmKiEUv7SMzx
BSNIkYJMm6184y1suf7qHXJdFR/UBb4HNU2lKVgAVuvdp1aN5hfcV9Vq6BydRZUnMSpxrvocu2lk
apXkEBSfeT45nH1YP4GexDHKqCJWZpdh+v8gCMNLN6kpijFeG7NYvUB67JbQQPJA8GdmlLYi9uFN
1Zhv71o3Iw3WvKfyPhco69H9rStBgUKFri73lMNVZ23fNbpjihyCEiaEACbjAatS1ZtoIDrZoSi9
41o6rrz44ne0IX5jQldxQGeld+j2jqYnhN/xtcqQPz50u+xQ/NtxK7HX0R1CymNvvcMp7Cahe82i
i5JacPnEsEo+GEYfmGJq9zZs4Iw4f2Zo1ezqhZSaDmv3r47094C4SGG/GxnXMiPP7F8Wp8lDoA7E
5m18prICRbxaxPHwe6MNTaKhZLGjDQ/qIG9SW9UKHiu/EZ+6MmX03tU4POB+yMsMi9iRy5Jj9Qp9
tRnf31GyKwuxro6VK74XUJvym46Rc7Af6Cm6EioTWHLH5ruyPGks3LreHZ9+da0vGuq3Dit80q/9
Tn2aAoaRMftKVrT2l3+5ltNUQIHoX8mgKvWrICIZDJsxTDfxDgOAX4WY0kwJ0IvurdZVPkQ6IrH+
3Eejr8z8oMLev37zxaSAVaFrZGQSb0VPIcgkUWyx/F51WaS+xvlVEpkIgrrBflvu229TYCaUhd2+
mcvwyLtRGR+YEpRqDs7JIdA5xAHBBy9ScBGhuQNlPi6ySCNzHJGS6a/cU+TsLqniy9L20gFLzkV0
Q1AcErIUKFbJGdJbpz1yo/TCFDYIl9e5gIHFohU7b/nXKeWJ1Su85RQmbPNrcymGkkXm06IbA7wS
GaSyZ/ajUWB9f9bCiwRIRFjnKN8b+AKs794iwCNvxJA7DXpevR/DcEiIiG9RWHHX7Gwft4G3LC4S
TFaL71plkCgiTrqUR3XdqamKb1wXT0hzThn25KPYFp1DcLcaV9TZsdyZRrt6/8oUBUbSRf8lv07c
KVubZkPDRpYFswi27w27akjoNtoGCCw55Zn88q5JTgp4+FWSFVKnK6IfYv0YJg29gQZqBKg/2tTI
r9g6/QR8m2Q7Fey8s6KbQ8at1NbhgKQLwSOZTYk2IyfSxCKzW3PXV0pU5VXmxwWCN0HtcEJFWndY
WoMjmoqbbkm/g50FIEFx7C9ek770eKvUDmOluj45hgw1dUEQfx1RpemH359EDl7ZLn48YP5IjnsP
3fxU8BmU6p7gzeVRmS3ZyRSR7G37k41FYIWqucs9/iRsryhbeMyh52tLhnl6MWCYcRZRqJZWMRxW
lSBRqvyK4jLIVZOhvsffYeEDRX2g/5hv2ZaZacAv8K3OJL3Uil0+EYyRdaeunbQAfU58cdC6IO9w
1hIgjUTpPRpNPRAtpWOyPFMJLQMCYL5T6EORcTVHDrycDPl5nNKOARhQcgKOZ0i0PcvxwhvF9yZN
ncSp5qiJstznsw4qQ/VTpZ+ywbrxClwaL+BbQthl7cF+fsrrWOjGZ4DmJADu1+541y2gPKdpgJyR
Ty5QRr4WShywwRxbn59eoi9E/1rpIJC8XfZSfbDvno9AYyV4jis4anfdaatdfHWUhgaakoPCsXoD
yWSQUeBm11S5BicjRnzy/oFXzMMOJzoZP1WOezOVCpxqTW5CUNcxldy7m2RTO+KoWUoOwdsklDIZ
XbT9mwPVdeMuY96nANwdxCKZ4uh+48G7qQ4T5v/7RAT7thrKZyBvoq68pVcC0xlBKimlxp/IxItO
SqrVHN+mieF0vVNKO3edX5OeigLqLOm8vCkUneV9THb6+Bgu9gS8UGHKg3YZvFEm079C+VtU3QoV
AFguEflsLte713ofCeVLpcQQn+JFVdfuIt/SJktbPT9Wmp9dhI3GtF8/8+0G+KDy+0mPaZhIvPri
bYHQXRZ+tOO7vO6MHU8Nkz3vyNk8vPJfA85DEf3lqMKzXaAnXPdOXYGD/mWGI97F5WRUBHr//Z9i
q9PWO/d6Ud91VKOD5s6P+V4sk1QyFwFsK5c04wWvOqdO6RpSgn2qzNkcs/KMoBD8nlSxPcnTRwrw
RBWeqzyc88nAhSWhgbPNvd2viDZ6WOh5vJmfGjYX2RamQh8eFRmcbJIomdEhPlR4Y5QyJOE3RsZc
z96QUzSgF9I4jVGqHF4eiacga6gxFbCIApANqOhU1lj5EYJkMaIEEkSjvblRfiD0xeDUf5c4tN38
frHDDdK7V8TeghiJ95fpL+nhmTs41n4PZw8kqi+70snhTVbbmIB6J0R5kV+xo43dzjXW5/upHyzq
xePrglqgQP/yiRKaLzH53XRWwjZVlLnjKf9e3ehNtkXV/Ovjb5vhO8Chc01hUU8RgLRzgqILLEiV
bj96dqZU5+VCZnHFOXEgDTm5R5iBN337p509Jskt5jX5/BHiMdZqfh/wICSQmQuReAujjqweSZVk
N6G/uCik/azHZCX3sMPzxnoWOjKiOohoDcOy6D0Uj9kWyAaKBVcz+zJ1CSY0bDOYz1ipJiT6vzJu
8pEBa+CYvaCEReIsiqn5znNW6qnFokfOywsszuw7Xx2B0gPAp/b5wiup2AnmXv6MgQRsfAUR0+/2
UslPXauese9htmvN/nCyYDKWYLDSg59vW2z63OuTzdbIsRRw1Yx/5Qn/lkYuxWHzwLHvghAjXWsG
vBgyWA35F4AjOZGveYRAbtTOsNX0RwsF9ta/e6EltHdf3t/XTSHcX+6uvSgxfG/dFl/Bo2jk2two
MtYVPVi0AQ70QXWXx/F8li8JyvqowXcMgT/D0W0ZVqZve/Xshng/NKNtkLleQK2MarnjPE4FoOLw
PTy6WaSXqYFj4kbDYBto/LZ7BaSngiIqLjdbtp+g6b2ukZzy48aaUTlWeU7Vk8zpxEmJEB/Xvjun
6QsOYLxtKjbXGgYtY0w3qkmu8ldKbrnecNm3nsQpQV/ue1uKctkyr4v5cEnPzk9g9Yilum5SL1CG
DMp8Oog+Nt0xr9t2KPWpxWt4b9s2G4VhCBGsKUajMUdLbOh98OXgRGFkk6E15tA+3fejcCItJPkY
wBXIMURwXMfPtx97NQuw6QsE2Xc8zo9JzymOfo7Tl+kkuA+GiRdjdpWUnv1I17eiLiSyxdp8iWSK
bKJpTqnQJoOSVWAVsNQKKI9hc3DILG2YyLd0HEyAHzqMvhzY8pg7Cx4BIG2BvxMqiJQWdC4B2DZW
J0O/QkhKU3vruvhSPTpt1NteqMfi777zqevfiZf2sK9rw5GCjhlQj4tpY47rJ4n6qiWgx6sz+UNl
QgKg5C8GmzPR1KLde/CU5SfyIKt0dZsVYKl6f7LJpeHDpkUdpVEUzOUqQNOtRrMAXbLHkAUZNFzL
LuKD7/t5U6CLlINwtUJyOko9iu0M1mKAbreOGgeT4oT3m0kKzXOkYGFg4kdxVlhVv3gO+yxmkglk
QNCHzz52Xkiy8NJ/7xPg7pfW3KBWHHtOxfUFf6/0+06U9vDDnSJNttCTRa7oDK01KjqsdFKtRmHM
DfdiW2riOM1pVa1nMrQZWIfdBd05HXAjo/lCeC8laXBjr5P7UkvhwQOi7KaaMILF+vkIPp+Ct+c/
UjGlauexRrDqSm7EghtT5wJUD53MyL7VkDDcuKcoEB4N+wJCBIBZ0C5I7WXV66BOHT2KDJWRHsB4
WWcSOAHdcjWAls9UtjmHzC1r/KI8QW8Ntz6GEsUKnhAC5plpTMuxrOQgzsD7bZgJbQiT6yMHHLb4
cX51JoQzdrZcPl9nJWbrMmnZEx89afJGuMuBigP33Nsh9Gp2gc/QVRfnzooFInUmoDJcyU+WQN3v
bgFOutYYSrbQ5H598Z8Qz7+Qb2QWWhw2wEmo4jlnCDTvGn0pUNwEJdjX5k0g+G16yGteqRKgtCfk
LrItsharZkTFX1t/oFDlpKrtnBNyq86zWB87a3qtzX+E2pgkMsK9Dpd7MmpLGKiM9nwTLtnvFWoI
YJdXtQDemXu+jWf83xIves5JvcmFvC4ChqKf+asBKjG4LzAeIB9svStBDG8AYNo/hTdeXbgeSbYo
g199Cyn8JTSev1gMajvfTLwqaMV4XIEKcF+tS9PKWnnlCI+nqVY01nwOE5Vj8q5OgtircTs3+U8M
/SM/on0gpYmJ2fPz+2TqRRsE9nkAmxRgPENrw5tMcOuFjD5hdH86iDJxze1dY5yEEpNR4PjCLY2a
NsIzyUmPC7aA6aZgJwPtrtz+MAQE/TLMpi1SLXglKiMB9JLbjgiqWniE8iHrEEF5JUCxoWaGiAny
8Zvcdh29/nF0arU4Hro7yMlY4XwdcSH9F+bBKVs4AVJWFo6Siert3lkq/W9C3EeCZT3q6HYtLu6x
y+qD2igm2KzTYervzqg5ZI4eWup9wcWSSF19Cx+jUnyWW0pq+DP42LOhgtgCMgjViszh2nskW42z
cCVdCK3NGV0kqBepex0UpXZK9dZCYdg/tveyuXu6iWPFlIX1SYQCuY+rkzGF3K2oJehbVP34fGXK
1sdPUPQu5ri0sFlJfeuogQEmTWoSYHBl2z9TwcMzDBxsI03+qNOL2OrP9iywTertiNdh1MaBvdJ4
L1+rIbTvFUIq+9D+rouj9du73yW5BbpKfLRxne7IbRldY6ETTq1OFlf8PTmls8swW7uw08AU7BWY
RxECL3x7dEjzOloeUxbRb+CIykuRwkZVw2NoYWjHE/XsI1PnTTPNVgXrxkyL9LKp8j9oMBx1BiUt
DbX2vrsM6v1VyLm/9pbZ3kRi1s/rq2sYH+WjJDSXihl8EpajIVPkgGprunFjQqESnjB3QgAOdryi
lwJAZOZA06PpQF91o6Oe8e7SnWtBYpUNCM81TxbQCcRplidrNuofIy2mbx8I2jpWH33vVV9Llozh
S7bTvXTUO0Br0ceqkSdEyifOHcl16RsIx4VnARJbO9xHbeyZPgNQS1a8BQ03vlVYaLuxD1IPYm4G
42NfDDNRmfrPe++8bBxnADmbwafTmL6adG68qYu1/fYercVstrSsZs7TAwBFG7jAaHqdTazaFUcq
sdMYqB1CoPDv1PgLWDjoNlZswvGGtgA6KmuGwL2f0iL42xQvk8KRX/Roi+Xhq41PEs4tr5LasSEY
4XlliB0SI9++IluCzVl3Ob5zkS2lnKilv8XGKSfcuvUVGDkTUvqMMrcBEzUPwqkstDTHV4wsDtqf
wkL3mnOwhwVKvYVWmZMLvU1tDJ5V28BG/7RykKKg3ElDaEspOoUah+sR1VN3GHZ8pMMURJ/T8/2k
MdEvK4Fb61Zevu0mZugOuGuRMC9ruc5GAS6MV0HtLACWA8U0aiaG4kbUnrrA4O8sGfE5Otp7ZbX5
X53zJjj4k7RaP8Foo+QV6v8W1IbZb2aPyAvbL9ZYbVNFzwbGS8qE3iJJEyBMfXh1K7iztU7dcj1q
A4La63hOjkf0nI4tl6jNrsNE4mhPyHovZlGtSS0grTqWp75KDxBzULKZKbl9LZdm0TtVnywOER+6
elgy3y6hV+Nit9AZcVJcADapaRuyXQt+w5kl1BRO4DkmDjacg9E6lxr4lP6hoGLqEnEWMdDQDUxw
nK7hhT+QddOkm8h9ro7vlSdxaF3GNPkddTavtxkA6haeTj1whyjPosCLcMAJUBitslAL2+FzPgyX
VAyDltqLD2bvS6YJZVLNexSJJaT2tTzkGwWUYNtg372XeymOMrWvrSt+VbFYXEB81VyIre23Cu5Q
r2BwRgzGjdipwcgMlzeOegFKiafyV/m9rvGIQIFCP81nbg0VPiIZ+y6wldOaVxr96nr2qHiGWLiz
M/eJeeRkoIvq90FYvxhuy6HlkwDHsRNucbAiKA2Ht8P9MuYaQrHazsgOg//99GyABfKEGMLxLa8B
+a9QOPyCCCpHCSpqhfR3VyyyxA6tAa0vS/cy3C9z2oTLBYSycw0jvqQaFkQUTcz6jewCWWcYZSal
EmIgEFunvoVnky3n33d9Iic3PVWn3fSfmWfF4EPsgLSpbuG3Wesbp+mUyl0s4N6naNcaGQrI8LmO
WTk+sVUnYF+UKWHbcipMcx6qIhtOr6XtPEy5Fb37g4Mo1KHAlyzpgvHXrjLsYtxIO2uTl9xrCPEv
WOOcGevDZsaTmNDgIb+OyUrsl6JcYk1Z0QVTO36TtEYF4obxawPs9UzzJdMS0eZouKcPV+j0Gt7Z
ksVEUkoMgB9HsI6s/hbqiIZbfbz82XqWi/1T0H9gmXSGT1Q5djhvs9QzYAcpcXYXdqrEU3gbLdvS
s58RQeC51loRVhG+RdE1EomTjktWhSe6FNR0FgoVQJcjYxsOzhUhkGHfbpJ74tOSpwahEfr9ey1d
At9OzGPPpcyyH8+p9ehWM/EhVMYNFPHenMtQ6dKjDKYALApkZyDbSiurPaPSFazj3d98oKWXFAGz
V2lIZnkQS7a6ZcA0Y65kYNnXct5pXfgR0Q8cc0P1un7pq0KzQ1wHb7HwVk+qi/5RM6cYj9vMpGX3
h3TD1msmqb1sNPSFdsQ937gXDtj/HcGRy5G9PZ0q/BjH99V41cTb7/Dwu3fc7sriVZG/Ol7AfPy+
m6SssU3IGsVGLFuEln7rItQ9u8B0+xLoee/KXEj6ybQFHRIZtGyU/YYCq8LjrEqI4j3ounStm1ds
0kD2b/mXwnx8APeqsUhlSDi+LgFAoi2UbOdLWvbL3CqJXDZwPpNLrQdN+1eIOnAXXjz2D1qnkFEl
oYAqaKSt+MNNERl4+J3hJMOC/7MTqI4gsAJDaeAdxHf2mM4eIENkZ3bvK2mBASniaxkyXdwZ1LBx
5URq+BbICNrgfuod1GXaWX40Oie/mhZ7uOu/K3UjjEuYjb2w2PCYcTTuUJqgmVHocmrD8pEMay+f
SfQPV/eeH5VJoDijx6nhJEUe7ruaNNkszfegMvl9mXGTS/I/6SQ9J4YOekyHOqNo3etop5jlppWj
CyJrFW5YudqDqQrqF4Drr0NHUr36Gopx+rb3KmnAUousRGhdhXUpQtyjxQU3QM3bFk5YxaRsQ6MV
s1AQv3rMcalyEdt8c3QpHDWsQpcLAarY/u0Pqz7LID7Lv7Yl7nCzgVYdChMD7c7J5rj0/Obni6wW
FWXg/Nwt6ti5X8SFLh9/DHT5V+VhoNT0uLWe+PH26i6Hy1hGmOQK/T7+YUdXVLOlhZy05DEPe6Ir
HKuG7lp95FacRAMb7FqT7OtLb0yMllUMY2hdvo6DoQKfv98kuFYp63eiUPf/m9G+5h4/6hPVnb7T
9kiymujLoV8ipnJtvCn7sf1dMcABKfCfvLVLOdXsruiWTARJg1wwuz3LXvue5a8rwDobK6p5GnQ8
RTI6NKzsZs6gVKCM3OiELUMw0vRl0YbjN6OkCyFAMMkHtQOlMP1UniqzIIdoARphIJ4ZNiNIHmiq
x4dsV1ZNGUaF+bFdybDAKdLIzCGuRlcwPwi9DOvsaH5GC+w2zUpRinDkk73Jp7jteFWDjzxC6ApO
tkIDR5dfA9+SbLXi04poZIQ26sw0s2XCMbQ+NOSAkXL9JFy45Won3RvbSbqprvf4Kaj9EdKTeL8D
w3VrWKGfCmmuBSyx5n18H0Z7vZopPMfw2oKLttBH+nY5FbncxF0ewmardKtHJxr1HlobvK2tzf4S
s4/CTjvv1TATGJGXBWVLqFTnaq5q3gpcUnl3s3RoqWTLxZVKKGCvyAactsmVQCCC0NuQtxq3GRh6
htMR0755KXXkU+AoMQKyfBveoe0y4jCidD2UHZjvhKzoLrqBLXoIBAAS7GGHLP91Zs0ar9BcKhC1
5k35c5GBIhjGxGFZNRlo7h678gbGK0dEYZU/ratF5covD8r9cC0ohgP+T650uN2vtvmW53yVrhX3
dkUmmaDFQsH0kYWGuS81NnfGZZtJeg44S0E+Xve679K7e3UUS3PTPMnZigLrbGZrdda6qBMebbr8
B1rU4FFMMIUDrJElwPN4LRS0v5Y86o+VGZXQWthY13ygGyuyK909XCAyAzI41s1oImpdEUDs7WLG
J4PTTp5Vx2TIJZH6uLomGa25Rxujs+j0I02dOZKDfnlLWHTyy4ntxZ63YhTZf/Y86E2El1BvvQgw
Dcd7T5wwzVRpG75RA04GNLxGZUXblCP6blPF4XHd+n5FX8WaNA2TSdgnw9y8sNcTKqaww6b02CW5
v7wehbwYcef7gM8awaOFPzVlZzEJlo5JnL6ywoSBJVSIYMf1MdI1sn3dCC2AliHy+Knm/cuYe8Sv
DxuHIjZLUBTcKLJjs4YeHVOC9L2dpnX5uPFnzotALq8KZeCcMLtyqpn8Efni6rdCgZggnpnWBaoj
aCqfrtuEzzFeRSJ/EgXuRZ3z9SUdtVn44AAHazfT09zE7Sy0P2XS6ZnHpGI0dTh2rPparZcjqKeO
fLMLmW1WYhai5vANZnESi8aCJuCHo4e/6K09jJwD4BOChi3zWowv4gn1zl6TG8ZEhMQUv9lg0mUH
wZd4W98KuNZz30K+elyiVKY9dZwLAXj/ZdrDQUKoDWbopr19EWopwTQbDG4htJfctdvCC20dzGAz
mP8wh7Kja5e1oc30EVgIKfxw3OUYG5++gDiuIhrg3MV1iwfl9YXfori7MsUqsZsHfHkwNVyZySUR
Ji7tjKFWfhwArOQthRek/r9LrlIZ19+gRd7uDP+DQxQL9vNEBVm3Lmymrewo51/23EgFS/CCNnPH
H2qn6cBRGpgndCbEARaG9RFO7maCaI8MtOHyl1a+2jkEx4OVjP59LY5LEdZ4F/5sR6X4l7Jy5OeL
wniTG6eaQNAnA3BsZ64fXw4Ye7n4cYbRZCtFlWgW60xEQszINZVOysvKlXqOpb3QdgC4ROfcXPhe
t/DsKx+oWf42g5J2CML0Bp0zptVZqALV8EMDiSr1jBG8pynIUdDBVCvRk0dIQlZYZfGQynp4uIjT
siTImcSyPS9tCDcO4x51Ac/ZbIY6N/mBfoz5mbNLJxcDuyl+31w1SqdaEThMyX0yQsVOd5bHI40H
vG9vZXxPXUtEOTIucwbqIsNgAL5jsuWKv1D1JK0f+KSWIU2PxWmnA3j7tUykXBHjsn6CC/ofStAg
uYr6ZRTPf9L4p8dS7iCfQoigWlNDX+IyQc90CAaAOTJVcSIaskAb69GPRzf+jgw3M6qrqZqBFr1q
RP/Snnq56RimrtKVlmjZ17hU7Vq4Oh1MkAsxvJHx1AB/E12gnlMUSMUkHw2NDkl5HFm8B/BpHIUl
sORobP7jT0dJ6flZWUZ1EcS8rLGxyTe4hvdYNl0RJlSdeHpJuZt8xYsL1Av6UIYKp3DmJNwxBs0e
FufDLJ6t8vtsov/P38Wp51QXNBC3E/X5Ky49VkSPzQp1jEloKWAO1wdOq97NNZMVOu2HJN4X/IPK
mPW58YqE+ZYNgrYUT9ffzB4UBrdDbN9wlILMtpQeHCQYI1ckH8sV30QI1e+kq+LzK86a6fSU8AGG
OPmsrHedv2jze7K504lb+nDK0F/2UQLq7J3n14q4ABLtMitm5foCe/07yu2q5gSDEzphzy2RKTZU
NUvizpwPXekuz6ouq5yvPjKet5RJ6AQOTWJQ9uNNIetIGHPUwW+7zrHGby2TaKGUxiQl7lQ6ZFW4
nz2U6gP8P9mCtxEjJKbPX9ps4pnhR5n9UDOAOTjdrW+KnooyqeAsm45UOQ/AwFKW/rCnCK1mXSES
+I78FCYhruOR6ekdawnc5NOiQILrK+N0KLYS4i3LgR+hRD/aJsFho5MqJ/D37yZfVZHngwLAubBG
UgnQTiWPA4dVA5bUMUgdac9MT7euW9unri3yI+qAlPWN/pzfR9+DhvzYwTVmu2JXIr3Y8itFvXli
z65k3H2Vw3Rq0c6Wb6np7MQrKzU6MFsIOd+KaCe7+mB5zlwgTJajkR1XPbqvbmTgZ6DYwnWCJhzv
My65qQ0LjustQaHfquOM2ALAuPuKF0TzILeBn2xeASVrZCxD7D5XsosDyetTe9tASmO1E0w00xWk
mrGIX4KuuGvcXVg/QZZwU453CrFZ93n6+vjTIZdcwrgdr3eieK2/0H49awvx+ZRQUeES0E0z3Atg
AguwGCg547TpnF4SyZCNsmh1z/km+O4DLb9QwKjV4Iu8FNtjQFl8czjEkQQBXRyLC/arpOyluS8c
k9abBkjpl9/UOjJUeDWCFRWi7HiSG5nte7BvxD6XjOiSw2Bw6Iz69/UuqCunkZ2Q3Xr4EKXUX95t
1WCNUV5b+yoB6MgSxG+kBnsvaoCe7e7+A/i235HCRa2bG1eeBCagxKWUrzuxx9jlGoRlmmcyGOoy
Vs57quvZjVHzSUJeJMH88dHl+QMcbSe8JScep9zZrKM7na6RwwuHLJBhBHgfmk2XLwUmrleUKRVG
TG2zHbPZHLqryVji4TCWCicNnaZPS1Jb/A+dR+PPBcopY4ktl6d7w3aN6l8qdX4hrhjGDjpYG9wM
1k0d4ajlGb1cHkkNcIdU4rSKacjpboTdH1a0rrfviJs6tL04zZMEiwNCy3Q2lAptJ7D76IF2YLnX
MDVTltT63Vkkgh2ngbH15LAaQ7BTyOwOueMUM+RXu+L56MbgVOwRf4YbbW9s9Ap7j7btfUN5WfSW
otGQJttMckxDWv1iwZYvEtcfjqqZ6jpsHRCNCJVnZ9IjJ/bcqGzeanDxnTifyFm6H8hluVnSZhgU
N3ZU0soKfeg19GL9GbPghBHu9qHY7SO6WX0sqixjS7vFNsQmUIDxzk4GSEckqLwCxuO1/q1uKUw2
gNC63bB+Cn+avy2BTX2cM3Xbd6Y2d+wgO0XMXEDqnHDAwm4VQXIy5qRjZtv8tyS4NaXYaGU63/1F
MANrZsaLZAtlVRVhY2LC2bykRqn8uq7sjl18ET2cVGEk5ioQeIEu3rRXsdfM9oZ+JPi/df7XAFMT
RC+6CMXUJKE+M6m/3puY/n4frTUBfg28cGqEm0LCJNCFJtvkYj6AymPE56DvjDNtHuO5FGDJayDp
V+7eLWkoYk7Rg7D1KDfx2vmj3bIb/S3v1qFZo7nrODZC+8HrnRFR+cSnln0lIk1UX7Bg2VqvBYIs
bhvDrucm6nNbsm4Vb/TqIW98xVP/7zrNPLi4WwCMwWSCCDRnWSZSugh/82/R0aJCwbMgTpvlClEH
8TnSnHen/M+BXGsEbSneQI421z7RnxVVQam7nzR5OFOyGV66Di29cF/MfLKh2P2YjWrtPAnIdLfQ
AL8vyM5+b0Hslha6rPztHJ8U7nz7BSxQ2m05cGwXVly60Uf2PFFT6JbeQGlVhMUWXsBKKYjGuTne
5ogqg+cLpTB1cAPmGUx4EeDR1iWXcXFl0nVSJe2IRdoElWsWO3Jd5Xp2oNwUKzV8lWglGdK4EXGN
eHfpfoqVUeN7XOAILfLmUJ7vkIWchCtvRGLUA20UwL8ukMyEn056uNZcAvzOaSsMzOjtxFuCWGAC
das52fkGneaz3SYbbDeY9YLOkyfPlFfgtWX0DNQ7R+W8Inx6eg78gotX7gVumFGKBKILG1EM6lyW
l0oWJdB7JX95xghtQYMmgJshNT4K6Ix64H6TgA3F0I5BfCXikdDxmdKRSbiTfiadMgqKqJRHA6v2
U3t2+hiuisQ/3u1OaWurLcYe6wjYrwkwcEMcN6Y9UbVCdLmwbfIv1cAVOkiDMiI2dsp60rfa7666
w5+24PCcU1+95ZOhBsIBV4U/m2N++2TVUBkZj/+SllWbZg6I8WSr6YizEjXA5S5bQ52tcxR8f2mA
eMND4L/CvkhBbgnzYrHUcnrCPBHtJYKJbaid/8tFsBnnbKZi37gPuSU94K9/b0mQnX4iORMte8LU
SjOkTppytsmSho7P3kQ8i+Avfv6HP/L3Mf4B9XKKu5Y90+nnIXP+WIALS9kogQj2rXbhAR5xrTLi
ctgWb4fsiHz8U7kqdBxXgAw3NpsEZlGVckIi8zp/ErBLPNTMiZYJl9+1bd9dbZaGsHBU92Yo7B/7
ljXK8m7jSrfRM7jqMuodTOnBX3np2cKCuVUdnYE1TxWIoeJToFKzbIDG2pgowKF+IbTZeMInuZJo
C0SzX9J3gVLbSS0kxI44RG3DBzvHWxq5BpC5Ff0Uj/rXjVJK5jw2Se6TXTuEG5Enque8YwSJEiRs
Ua0NQIKZl3RfZYGICYXxZVW7cgNB4kaNLgvDLM4bxfUP6iIRk5afCeLs5RTjbmPGVlWe5OZL2xBd
NgoNSYUvVolqwGvvcwd+jj8jPkcS2h+FJNEZ834JP+crKJuKi1OhbPSzioA6pyXvGQDbEKGj/VFo
NMW1SaTSQip3fTHT3Rgn2vU+1sBSFLvnv6QAmna443/QE7Bdb7431iJJoLP0KHndvO3QQY06apok
R3cQ3n5EjHEuISEWv68qRtyVPwgcejpS5br2W8Cx6R1Lyo3c8RU0dI785JVBjjLTyPcuUtpyvHLZ
sWCNhILDRd1NSv2vFhYvBJB7AE/vaEDRzD9mO+v0aRCmUNuaodF4wqDvdavdDS1U/smvKkbHP0CE
1qUe3yixJ/C8jpATsfMuv4LXk9pD4haE7kdxfqxWG2fJWyMLGH5bd1cai4gx//iEtXk89zv06pfV
eM8iTlBtmtIz+Cne36r+JwJM58p3nchDmCupFw3NzkQu7NadKC6L5o+tpTwrZGQ1dP2VzYMVl5lC
b1b9j/3LpIQYZTvIAScKMHH8/cMNtj+Jv8gx6N7JtM/pOu0RDiCKejGof80TlikFXctOys2+o1YD
rlF4/2V17/LRXjTrzq+U8N7PwAPZ2zIB334zgVkUawtBz8mv2H12flC24JMG21oC5ljzXPgsIZk3
oWERNQdON7Nf/0wY3oLGEJPgvHel9VgfMkk9BrjuvZ/nOCitpX4nZe0yqtVpCSMbKk9wUqYD8Jvc
Clk4NeTR0ihmAMNyBKaGsCRrlB/ohXWwUV2+SrB5y5NIKWsu1f5GpQFiN4DqYMGLCOPoemlJUMgM
BK4iMyyLU1ztGYAWMFsl86/IMwSR5yps3tjeTFFoLEHLMvKkfm/J8YIBc8p5PPJiwUnkxrOrfc7P
Ywm4vRlBoNYeAyyT1vm9nCMDns7b7IXCsgNx4qNCsQ19Bak2bSGxbwsj/nFIwXxhS3tGRogUFpb9
KSEQWwXpK9NGRSxZUVYDl5QS0EAWRy+fQ7zO5eEr+YDAr7Ld2bTG7z4dofC37aTaFIF3WYvOU5fl
e3yMXRFwIBoSHPA3dIrkFbeBCUdtoA2/YOB83mqU6lRPDtzQcfprJ0Uhm76Qw2xP9/xypqPuWgSo
2lqB1pXuYZTPjrgRrcyVSRFYyisdd9fm+XuCJpgcjpKcU2Szpe9/VbNbg3TIEaf3twLOecM35hxc
XzO0qoP/tXBWl9IZu985gmIyt5U50a+vAT+b+YSVXnDgdhMhLW/tGx9M19W/IA8PQZTS6cyT1KPh
Cszu8oLLkre04oI8tIQPyHu9oF/f71gMc1YY1gk+jplHJmkxRMvJ6n1gSDgl+2rl+oyo+iru+3U9
BYwZsW+xC9Yb/r9NaaW/qLfZodFeZSLTtlw1jVRH0qq/vlQ0pfmmtFIFzcZq6fyzI0vPWhbrWipK
crWAJnyWieFzh83cOQk32nxc8CckSqlnxBrnYVAWLYu12IOPoXScO3bbflMkhCD/tXh9T9TA238d
ZN8QQrlhStAYf6zmWbSc/5f2vcv5gbM/ZSVD4wvFGyL49EX0tMfCsQ7cr/QNF+wyM0/rT9ySdsFc
mkaqkMD7DV7Mb3ZfHtqRBfL5h2ZqCampToMv7BvsZNdEPXbsPlv0vhisVj+pUO5ncbz1+Br+xk/c
JrVDUFmv0i6hDefGDrdvLDIRcTxIh3Y5aoawHuwtBy8tSR3khPrlT1uEU+OO/dITMUl1iIjsbtf7
khdTXHuwm0SYMmz2OgR2a21OJlQKyGuMYjGKJEfy55kKFOXGhPdlHMuDD5xF7PTZ7etej3VewHeb
48q6NQPL4Y2WYMblFFSwdVUXZ5VdxkDhYxf9omkdW2nxTlPjcfMk4zA0wlA2eR6ltSsBlpS7SxIH
5yv11Q0u5lD/ebgZTl9QHRx713TA9SWaeqHn8xaRNWRzrImB8hSvqsANLUQHTah3XE9eGfrhIKth
hMVtB6dgjVeQPvu00rQLhqflh+VVH5YWr/HrsyAvFQUBDQSIyFHBMO4Se/skPg7B/q/2fw8HYm4t
goZZ5oINZtLaiLv9P2eNK3tvO3SwLsKCig8N3IovdM6Q+N0dNNMLWmCwDunAopI8sPR3HfGkvXSW
Q1FqSdtJh3xkVVUYiEsFanpgcuLg9DhOd9AqCajIUh9tI6v+mXLi1ltBwpNJoNaWPBvC9VGFeD1l
FqNAsACLmf6+aQ0qZkDbIuv4ffiBSlzMkKeMMlHdzKn7dyO6vi18xXUKP3jRHIU0fypCAZlY8GkJ
gQQTQ3CD/2sk2u6ldlevASZidRCy+PYNowVjE+wmHd6dSRJP9mbVDxrbXFIIgwk7TpL4ktAVPCfR
w/8Aa5zlvpw+S6SUCGCVk/QBBfmzISt20shmSgRzqckjR8rZ73By/AIUcAQNh3s07WjsW4p4cSjt
WZgglTabJ7S7JcS2Ua+yxDT0y+IfR8avqoi75VHewIve8T3lyVFCtFdeH/PC3+3+jozQN6ieka5x
4qFNxhzgjEeiwdG3bW0A89QH0ADlOzpqsuSGWJcdBE/tV9ZmAPRFLFz+Hz6BoCnGDEyuitSKtZhs
p+Ft6fCjLv5Qv8t3udoBaZUipg76nr5BYZa++4O0lRNu4og2Fn2bNlS1p50l7yK99lW/1uaYRMBT
WwJFge3IBGUDsTfRCo6FfjPAl0uYEBDazz7evV/piUfIXrMf0wgW259RGxNQ9caHH7YMovJOLE7o
QBOAF/ZIE/7lvxvoL1mdllm4/0s+Zg8I+HLJKqU0mNRLEgDZGYeVy4yHa3UvywI8xjxyQdnaXGv9
f798SgP2qokARFFzKMi3NchiENDVwpXwUFyJ74x21bUaB+4zt1Il3LQLM4v4uCS/gNEuUXGeL4ek
3fYvK1qgxNIfbJtum46oj78IhcECnCuctgYaYovtRXVAhUlMY3ppjBrB2Olr4N9xp5ztozORlkQK
8Z2Iak5wBZ7tv7UQndJM1aDvnVijp5HGk5QIhFI8t6calvAySG/fyoiWiVLTUokVwIIJ4XdJEq/1
hXjFUUlZpwOOrGohQU3X3+0qwD+RU8NOPr/tHuPVLcqGxLvBc9sOwVr3GSMwNOadQWgwyDYlhJBH
K0Ls5h6b6iX0YbaKwIVhtvXjxh9o5vuIcUlKGvDPgJ5cmKCglTJtALovpgcOtZlXUsGPtOeST/4W
ZtOVe2u2yjwDxWkClAdA6smOZ3YEPl9N8W6Lt3x0QpOKLnhaJDNepVRcG/pKpRuMr9WwMENbSDpe
t0B939nYwfejiLUp1CLma3ihqUami6nDSMC4V3Z/FTVSX1npISawlacuKeISeqVq7CtBSTjbUPYF
pwxeR+2t+9MiDvyLqATm3WsDX98TUG1HPt/ksUyBvxFStKLJUyQA3q1ipmrs0J1V0u79XKMOTnoS
hoW0z5qXQpSoTXVuM14v5E1TgrNZniQb/BW9w/YLVn2GWbYCDYwSDDvw2BRbgV9PlzpmNPvPZI7t
+o33sw4/ARtaFrOIAmyz/HxFrKB8JEc2ecEbqucqa7hpIfuGeowsR3tuCwl0JbcYuZIzVgsGqYcv
UjIlMxeQaM+8cPFPUhckLbAHK4GsmO58midg5uKm1Rjb6GjWtODS2E327mFQiUuy6e+9roxcqKgu
1kox96Ulf2lRXl6/OZYqfjdGPKzIYqcQsu8GTmEXrzDAREDfmzSwuNqPqFENCHGEkE4FUh4V9EhF
I3Rp58zFOe7QrXeqdqhAqj11DZmtIc+JORF6MIDQA5OpdTG75+Qx5DH9UUcPSwIcjL2qnSs0xdL4
COTBSu995plEZJNy0CCXsxgTjNs9m35x3okzrElClnSwTjSQn2d9AuVNOhQVsZs9Jbk2bZeOHWIW
xUbo1HAaReJIR7Zef6Qrabpiavoy4ZLC8+FZaUbM9MOyQ1H11QwZDGQcF0m5O+N9RrjKCnV3UAi3
JI8Yj3E61ezusHw9Ed99SyW9cpHWFp1GD9TiB9m+jjvkWFGl3L92ddfb8sUcpfowUBaNrHYHF1A+
jjJFTdyQVf10+yTQNT53gK5fGGwzNtiEgUBZmQICBhIOd8NJ2hEYBlr2FEmJtJRT9/t75qQGIrWl
g6Tbup1l++EZqIDhmwy+KgxqapKbdiZ0XwwZAYPdU2ZNCyw7/a+aUF+pLYzfqwhWybllA7A1B5y/
vSSxaklWHfBkwMZ/lB4q+WwxZ0nJ4uEYAkq6JT4vW4dYEteeadBqgygxRfof2dhuGLXIz+EBzctu
AvIyJDQAvRPmhbkLmjJbdMrqqH8TazywT1kDVwQueyuw/SJU53NxC8pD60KlX7Sv10aZm217c1k7
GjVaEh8e9y+nNt1OhvKG0UT3LrSxf5oLXHD6l3MB1mODrRah/YGRHGzsgx4uN7tmuXLW92dWNvXN
BCIE2UEpjtmlhpMGyIpBJYp4qGwbi/P48d/h65FGj8XKTmdexCtNkAcYzB7qOsVE+kYM4O3XsPg7
JmrqautU6CJlmhRlxfr56pgzjjY1loD9cwBpUbhR7JHdU42De39HZY+S0dOBvUVzE76EErhvSdWl
qGekk5Z21lXrZQxAkJ2HGhiKPBnBG93nMXGoKiRRbFkE/E7PaYzeJYV1pEPDViKn6bMDOuH1V2u8
1jFCRuM/ejW2HZIzspGwmuPWm8RIyfvcF3xU4RaLJR7t7M2EWEmTRgZzHO2r9ZZybfj0xdOyaxdq
GNsKxXoTlfvilEHepxtGE8nPvQ3fRT5+9i6mM9oGwyPLE/eHTJhvgGHUCQWc7GSFG/NfWIb0bG8y
+DVz0rzD1gffbWpfOs1skYUivYqBk2007sq0cZ9Un94qbJ+XRo7EWRoJ7vAGrd89IJgGED0r8Pgh
ISa2bHbYx+hAv6Rc6RTGDV6HvmGTTs9yAM2Zm0QI2BiIqBLb6UqT/jSlChc3gdcFNvumSN09QTEq
jFNz2elLc7BU105+Yw36UYXS69HS6NwKxS8S8f8CDhfqQOkqilWDqprmblXDJtgL2x5dipm3Z9ac
2TtAbU1Y+AOuLROo4InRwI7IK1t5hwfMCTvRmSIt2gEmEzkoGOc8VedfV0sMGA90VNH/O48ZrLZ8
xZ2IUS+GLeJVVKr5qtOrrp2I67fG7u86QgvNUEOxPNSFa0aW/v3+s29KIUCYJbYacBXVKVJN5t+R
31P8+ZkjQszi1FL7uA2tg/tknkIkHfaKOCK4BsHSaIalj5bqX8OUsM86YQDutX5ymwImMRXohWj7
JDovLRsvMvAOdhkmEhUMoSYx7SuA8bEizbyVHb6cUQlPwBuce+PXBuTZAPaxWMwZszN1rmyWtTXs
5mO9ptnWewuGXIPYoYLgMguvtpGpicY2oKFoYSdK078ImRA4sHkEAHkuhnDQhOM/i+2dXYDQ6Q+Y
rrj8QO891RUvx/yLjyNWnwuz1jrXRqDXRuLg8LIoxXfQDb7a3ekpQ5hXFaQzjOaganZcw1ez96/f
hH0QhSClr2pzYB3F/pzt0sI6wm54tHEMWeAUMwWMOD2ZCaz2h5FXQZ54aOHjcn4+3Rqu3hGZNvz8
SqKyldKsnrkhgVY75EDF1BWqxXfF39H5jJWKxaCswpexkqtstjnDBJCdChtk8lIQRj7Mg+AklXRq
5jV2qAMKq/QKc0FSX3NtfcW5FzYbCCGPae8ucbb/g7SS92V3iYA+7DGI9W2fxc8sCEyeuGpcjlLU
PNGka/wniAzMBklCg/05q8BGUuOoMNmOp0FxJMA83LUKfTWsrLxk6aqeBfniXOqszNMmz0kp8oMg
troUsZrmhxo2THc2DbCmHRxqUwWs3Bb5Igrkj6grO0yqF0n3V3UhNa50bxfiEqETJ33wgOxmkh1b
HtHdvXEaE084oG6ThEKCzUNn1QCXpJt/CqyKNjb50TeOKBDlkgqTLn4UkpUmokRMnQ/UuTYO8rDE
wDLQ/YVx/bzbA/l697Je+Odx1Vs8w8FF3BhmNSrdcADPEcFDaiuh1o2PuUwNJ6Zy7SS8LfB1eoyw
kOo1CZiY2vobIcl6zoLRkO7MnjE/adM0wgqbrV2YjGLEz9EK/xnjAnAkFazXC5QA0+p7P82/YpW8
o7YGFVKN1h2f/npoZGf/hTWWIWSqAPuIZkxOxoj5/+Aqi8oSSU9tTLxW9r2peSlLMqa6ZMOzoDSL
kh9pO+jeWMqI0v0I5tBNr/6HRFx9BbSNBv+KG6oDonYFY6vamNVhSidRdNti4zjkKQCM+0F3qhmG
W2ayIdyPrAorqBxk2A5e4HGD1445xh8rPwxS4ppG1QzqOolnIFvK5sW80gyIy5Kch+FvCr2W8ADs
Pw0i1egd4kWp7RpJi98nI/QgyjNwQKuGYNLnk5Q1H/S8W0/HKre7fvZRV2WM8oYaSPTYaT8C+Zxn
lSQMkFwaz7YM5KnhVYPvuZQgXZ6zoVGCWqfDOek1JBh4INgYnv9eKBLRYHHDQwStg8J9sAOUV36Z
iHrYxnBIqqetD/ool3PcwDMoEA8pATd4TB1SG8vXLiqC9tS+OkPVKaCP+D3oRznsNu61UfmGEWR9
qxzjp4zhYpf1SJyEV02L5qvr/rHflIbtCB2YjRv1FCVBbNGq+iUa8AeQcbavHApBksx6Qe4Gk2S+
fEAF5erynAg9TIyzlA/U/McKBodM/swP3orHcZJa03eu0szm4hd3jGhZOdAu8C1IPL4DLOeU7EPS
5Qk2LGYB06lTFrakAIpNU7TdEB6GBXVojFniUQKD7ffOPpJRh01KNViSjZExxva4V+2icFrwk3iT
r+DX9gTEe+PnRw2ZaGPraaQWwB4C77koHYRhPIRiVfyIugmwwMFpqEMuOkUpqnBGW/fejxck4j0V
AUnjc9HDP8utav/yCQLLElBtEL8+75wSw3/yN9Q4KWRH++VxtJI9EDtn0jBGexyPMy8yI2FtuNMy
ItjL8XkQ3DQqVFBmKj76evHkAGxqts1y4KeXUW1svs6SRV57hBu4judu7OssDqkfAVyU4NknV+A2
+biVflk5vw/YT7bKYUtiA69wQvqJ2V/GWwjpxFY+t6XHthxjAuAOu0UMhKR63KnzuVMAwMrgar8X
DEJ2T47xOyWgINHrh3hS/t3OqCPFWHRqGjoKrBDS9TCHFReboy4m0Ac1nOvWMbw61RX5JU8EEUoN
onWd2l+93LIs7yi57qsy35khYLzD0bHvJHYudvF36uMD3lwLLJhxlc3rBmJyGYc8+vMb+nWw3lNN
QcXMEKCNCwJuJ2FV1aYz7kqLE3H3ULMP/sRcXFdgTWwP/XtrPks3KZvQnzPDPKPl/5gEXh8C3C+0
87qUmWDaJPRqJUH0wV72gvfN8rW2/QACx/CsoQm9z9nkfbJvj2UU9d2Xnya6gjG6haQ3SO0CYYiW
Ph43+Mujb/g3oXZxTTo9u+d4Hy3o5Xk7II+2Vwka2w5z6fkW7a8RXRDtZ0LY/Cg/NjPzOrVamx1n
pXmkY8eg0lW1O7gnCwRzplP0re+GbnBkNI73SM2ySZT4crgMGna7wgqV8nxxvFmGE12oFG/YrGnC
C1sCcAZoDMFDYa1kbXOcWcBHGfxlCLIIQSMd9nhklTABDZBFXZYroNivYUzNt6Bkk1UqhkFlXfZk
0zzknMBI5K+MpwzFKfpeG7SwQ2g2CCoEvdIP66Ae/JlRJnTFGiuaCr9eW/Iw4UPH7MCO/8jNJjWn
UF6+jsujBZWQ4cISNCQyGIdVTt2335z2DKliDU/ktjFXG5yM1cDM2sLvQtUxEFRsAxeU5vVWmB7q
of0te3RqnFn/N9G1loJQAxHLJ8p2WMm3b3p1P55Ik5XtHCEZNOcTwurgPywxmrFozk7xqrXoKgOt
CEgiXrX1zHR7QN3DPj2Fv2XJw3d2As4UtKRBSDf8kQ/OapmP0HoQmzYoqnt7pUGaBLt29WSBSt0l
0XFFy93j56m3I7aAWTXZ6E0HWuzMlnVzDZNS+UKIEyLXZN1bwCj423C5IHJ/8yK60BuN0g2sR+Sy
4OuQgq0NTggFrzSt9YGh4JGhHGktvr5uagzgo5GHo1bxxZGVinr0y7giigcLhYQtz9ijjGdw0UoT
F8OPt5VkYscrQg82NTZqsvWUBBmQa0e72lekoK/8+jVT409OAP5QXfEbTvMYxkAoREYGUTsT830S
T4lhznLtd+iPE3p/wMOl12q8e+M7hsK8qwMlDZ0CQ0wzyz1yUxB+e4V5JVYRjIKVfSP4zXRfxoL4
b9V7CTVlhmvE4589xW0yGmj/UuZAhXrNvoRKg+kwaRWgrCze5CXGQhKa9I7elAy1B8B2SXx9NhLo
819j2lwftsq9KBRHT0UDtnFGEWIZiUbvIoFDFXnDT4gG66vrggHOt5eQ51RZOERF71s0DKw1ItA5
xpcHLpti4q1DLDb946F4FSXoGk0lx+oZp2nS0QxjGAXRXYhDk6/ct/yRqf1Qmf22uDuj02Mmxs1q
JmBWTPwcKX/Glois5P7h4YfEiYPsw880ekZGyPBsO8vZr4YKZRxpldEZb9jlx/zu0wbC0Y0zMDLi
0hMzBtZeWOunSgBMzW7YGQL0taU9eDbMYls0bQqFe1kXOSPQsqarWdeDERPdjkBwwYa9X242X1yu
Bpj5fPIzdVnSZA0gk2CNrXiGx2VJuM4WL7lzHmycGha5B7mZlKZdTE5L8Yy0ugmh8QMZuYdQHkXg
qLbASHDfxdRhd/k6IPd9v+wQckEq0MSVupg2SXCLvB9Wbyu8p10/knCEZ6pCFDZc1ttOF5E5PDon
TB2Ww/pLQa64v3pNV5P4BkLKVHOF4ysr9b2oFxnZanz+x6aFpS5kj3UGc2PvDb8Rchwmrg+mG/tG
cgFIRZMiLYbMelWBu7EmMMLkjoAjmHJLGvJA6IJZ3n7GhVtZtz+5OspdDx3nXCVwKmqeoLyOAvMH
uBxnyVN9ziylKGXyHaXAR3rl8l4RD1WmdSHUlyUnaDVLArysBI2XfyF3iVc3DgcjDoyn/EJL90mW
ot1I/t/kYtaF5vozR+IOBbx0WaOskoytE0cDnAVQ3Ru+4hlGRsh8n0wqDspBjfyyN486VRT6kIzZ
xHl4DKaBapS8BE3MFTL3zjypvybaSwICFdcycGaHR/j+hN2Dm19JYMVSECW6uVpodUbsTNfgUaZZ
5Nww8sRFt2HIjElHre6SNDm2w0q+nEu+qrfGaqcDXsFHIqqEeakpcaP4NaIntqXcT7XVnetBuGXy
Q2oxYbIMUQVJUjBrpg7Rg5FF91d54riU3GoA+suMso1KJynHgiMTNxkOB9COTc2XwoyI8of0xwzJ
Z5luifrCh7dJXDsdxZyr4YHWJrZnShwwyhhOnB5t08AhZHW2vnS9hw0R8tBVuFQXN3aIGULvSmg4
M/nAf0fu5+SBxt5eVxTwrX18dpLTWn1pmDBrHmYRA5z6RxlmzZeZJ+Fv+aiRFyFFeCEgi5HpY7eK
gIBvb8gTeTqmJE2cCjixP/h5LC6UguJxgfaqpLTnN+Xuvt4nnHqCsRcWb9FAO7w+/fg80OZj3fT/
WLh3HU1IW4Z/5H3IsRwpkLIxZQyTB8u7qX8YRW8Wx7XxYhUNUoOF1TH4QW7dzN1rycrUi616wkzs
VeEZIUDJMq5Shuqnvfpog5SbdBpmv72ZGo/w5Yb/VzNE7uzOpdBboFdWwamqelEYe1U3jfvFB4Si
lwGfxMtWVN3bdUPYXGrcCO0yzDTHZpoE+lvg0O08y7/QtFVWnAi30m089qrBbtMuwL3gZZ/oIIWQ
Hr3y3pxXMAQdckGrL908YQx/FmIiKgIhA2xB792BYSddfrPLgeUVYIqzkYcLJ5S/NixsAhKZBsGh
DJoUV/OsENudQlYLadXAyw0K0Hxp+nvdipHRVdUfLRUCz5un/xk7e7lzzzKZLeRpH8jvQloTb24i
Pf0yiLLqTTgVmXV+mInDCa/7OPV2V5mq/Mt0qJUlV0Z5AWF2LNWTq0jgGgGf1Tpam0pkaV1inj3/
jSwEiu5FneUOPwFX0HVM501eeO8es7NQ2a6sTQYag1Xs028iIut1Dd14q7VIdrzlOYmrq4T10PPa
upVfddCGZfb4VhUMjOIi6cpgrJNkKXiP/tMo+kBS+NkagymdfcrGffbgWGtbd4gME+qC4nqM/XMI
15ROtH5kllVT2YZEi4ipQdvG8Eqdj/QAiNAk77uHzfDq7Qfj0ooa1KUCU9PPzn+GYdKHxaKMNjX7
7f/LZiEEwedN0lwFYllbWP6AzqAvxDsLCpm/iJiRGjn3Fj/U9UUxNW4vF4ZAroZLgL+TKtjlPwW9
vjt18uRtTsbxtYdY+3d5UQEw8VftyhEBGtL/NMrsfsPn72E0lcljdx7144QW+oMoTQfHKxbnOymS
F8yz5ntNI8O+EuSUDTeLGEIivrf8yn5tBdmHsZaWUClA82hL8kb2pwSVE+SefCKnF+YqOfunWRF2
zRd8QOT5ZXyN+7F9TkSZ1pk/g85tbzo5D/DAjvCen04gVFWtD9ba4M1h7ga+P5q9BBbpo3Z1x9ro
L57GDLZxFvc+y6y85ah6oYbzsuttaDoGjZ3DSHsWl8WhfNTgp4+bdP1lK65ncs47G+Iji9zWLX0h
Oo51tqLLsJkk2lQPAnK3C/BxxGN+/fcpHByrI4jyY+uPlnRzw166MvPOXGDSShEmGXJGwTHxJQ+Z
EALT6byD8evXG+LSmw4pZTj7vAruGbLQTylud5J8gzoKuNL2c4rjteIc39x8FSzEXRNJYM1kzs5M
L4vru8ctftpQ11TLmDyV8HAnp8L+rWM0PdMJTDT/JhnbMVouO55Y51OsElkrIi6BwvbZSlC0NJg5
7NgtSJMon+LUfi64LVYmJa3u9L4Wnfbr7wbPG4zEFWyl2WJiNdaBw6jPmN6KV+U/Sqws7+t32ga9
Qb72e2bDcDbJZdHhijphQEaretGqjsRZelly1AQcYJSvXW5curbTCYnZPjSqh0XPJezBFAiNmUTa
G7Mj2pvwAU7U/zoE2ZdNoIRDC9AXR6lxMxwjRr1GlKOQFbGDdXW9neUTESVyEDDWtupaxIcOJR9Q
hv1eqrkLH01c6uDrA36bII9AL+Nz2djHe3fs8OBhivgPCcN9J0GL7+kmw8Hbe/5RZ3s4EElC8K+A
7zrrK64T6jxQeFeoZ+vco6Y29o0P3digoOC+njyYoUjDduIVmXBMta+cVBhfKbcQakB/oBijpvUG
GG0cB9Udf3baj8MYRUJHBAc+nxqRY3p/padgMvMHKos4apjuebjvtIm0Z7T8WKlgJ/C1aX47XV0s
Cd9iwDm6wcDQmFEPvPF3L42A8ywpJlMancJUJWrn2jKCDDmbjEyQBTRWJ9ssAzsx0uMyOPt+a8J1
WLJNvz8XndlrZsO13w09CxAh5oKMCWk9uBomgoTvRccplxyjRdwn2+PBQ86iNTk+NgdwWThZeb46
uUfTX46lEfnKJD8wEWHtukhB5BryWlpC8w5gLkAVdyPT+WtalmBM3QD/wZwdutoiC6rr961Ng8z8
MMjLdBa0g/Q12lRsKyPix81eHmH91DAZVjRajD/l2Bw0ZY7Bosjb5SjHKcCgWDTQCAz1PRdjN0MK
Uc8I6wfiz0Ymh96uhQHKbg13JwFTZrXXKy9n69vg+myOny5oY+KUaLllkxpZl+xdgNA9TUuDYAWA
zRAq1dVUnBHBG8hPVilUpLWre/NtOV1x/HTvLmdEpweGe/6P9WBFWmzm1DnWA1rk6xX1wyT/OoSY
Q6mOrIsoUlrRhXSi6BGwSTWS5EKGiVIyrQ2HCGuFVgZnLUQQZZIbJM0vb4oqFYoxr7HlRPI22DNg
sFko+8OFGLXKbhNaGxxpR+/zEXSxGtdXgwMdowPHtT2hkOjt6nQ2fqBjeoLwHZWjXSC89CFMUQkM
zNjO7JOq6COIj0L0ucx3M0XWzdNls1Bkix8NS4g1uOptC9D+9ykopyby1WJpjz6VUM7muAMOQJuO
TLnB7hdtMxsOqUM0h7QVAFn51gH2JjLB8smo6VyXnAZQtMkEnz/pL7rnPhmk1kuetbXsdOSgz31O
/gW+6xD8ptDZLS4gi2uihGP35j5IqAggh6oWl8RjXFuBjbSdmGHF2ylEYcLB/7D7zsoTLWsn20dR
US6embqBtWBFtp+YPAgRiv9Boag+cP/g0UkFuqZd3Vn6DSUg8RGuV+YCIPFsEbA+k/yLWDKpZsE+
ATGh138Cu4/PPp++eMRRphQ7PMKKWdO4P093Bx7b9fffAcilUMV+rg2k0DEw8rYjLD+GKiPblx/J
XmAfxT/2EAkMDge8xjlo2NX+cFYIiFAhxVDQkqLzcY1sWUUCXmCzTlQKTGUdfa7lJkVPsobFxKu8
JIxmj/umVd3JcPn1vP4dZ+EnMT4sSp5cd0VCg7HvvBJOmRu90DDwt6kOFMSTXEuC6CPM2OCaJxiR
guatOefJ8NtNp+HURhEAji44GJ9+8T9xYy1+Wa6nWWiKSnZRtdfViBhdFVflr4jNjm6zA79rm9pL
8H7L3rnVoGWzQWGApA/YCE08tuHB9dWlRAOwOQE5zgi6a4PtX592RREG8yI5L5CTpJW+Pm9nA1kJ
uN67EeuvSkdTrONRJ/cOlgIWmiujsFNlINHoMYXBmFw/HGFxlPNa+zo+SEw30fE4R5E2QxkO7BhM
AbNjlZkJOkUbiiNIODSoCnxpPNw8Deh3core4M5FajvGoJFusU11KlBqeK+NmL/3SmVBY3FEgpmt
SYxHnq1zehGXiz4+f9zpGYfWfth7L8yHAfWecuKhlAhhq3UyvmafSFzomJmR22+eztTJbTwvj84M
gsk+sC7IciNafFVRHnu3S6GcdoXHcv8U9lLNgGAaFaiIJrShBjU0REEjtEqKqk5YrQ95/+u7OwXl
2ZC5H6LEi83FY8GdaoT/OJYCYPpUcbi7GiTBMTd70EvnDgqn2phFmhvHpDztcs0RVKFc/CQw6PVA
QyN3FIvZI+PcLt1q9IFg4ccCr/oLR/xN6/3FdqAHxpF+SYvGdzGBKuTmPVWOB5W9q5EpSqXJbXhg
QkOJ1xpAYZHjz6yZ4ORbPS6XhSBzs/aKcqEthYKxyvPqA5Vo2UfporxqyHASvCYUWg+qky2dr/SB
+DHd6NBsujSp1Iygdcpimj6SNIvrd7jzW9KnQOcNuu//W216Y4lPIemYoE+MmhH0ETVP7Rp1FaBa
FasNyFOfogv8uDIihwNI4row5Z+Xrb73dE129+/4xeeofxdNp4GO7oAa8SmhkG+dwBB8gkkvxxBn
DxoizwFCJhu35zuhvze7GENQr7U6r8jK7Q55svnQ3M/bOEpwTHMPdOJqigVzJrpKFM9qD7sl97gE
6lS0FihEL+XFG+1XH7Ouq49+vJS1XdMEmiLQ7iv8PQSjU6JOsSkq8F9b5mGyKLRtppGjG+/bhQmE
OFj30/wiGdHeCDgMKLIxsODa1jVlafaaffrJyUb4jp76pBAifYPSCNKcgzyt/aW3Y+wT3yYxrmK2
UHHtHz1LdgjNjh64SnGY3h1/PWbpKTY8BDrXOYVc86eWozRFhAtYLW0YPV1yfj7524C0OlR3ISAA
lcbV4vs4ttt5CigQZpR1hGO+YRnYMO+qWlZ+/K65YIhKIVEYzldDTE+arkYkec8iKaKgubCaWrBJ
KZGfqWVsz9RZApxY737o74SZk7Y/XZpTrRcP3q7D0VYjURbKVgFcJbWdy/c54ifsyeNRhJcJ7JY0
NpR1kuQbCfh9TwlDsfbAr7Kxq/Yz2cU5ef8F1AWlWpDQEpIg00IFx++lYYWXq+YhxIFhtFAk9HnG
45Kf28cHCXVDxGJ8/Z/JTw9tKqeJ75z4Ujj8gbC3VDbfZnrBUgZMA8eU/2jx/8v1CoE47duUn/z+
aVOTD4t3p9rtYD6UsRC9kt2fvy6PfyfgSdVEBP4Qu1+QrxUDCymxQj6/xEAMA2F+GLs+sW+5i9Ku
Pj9ezjHUaay23FLcsLgs0Ih8U/sKc09++3HwgO0x8mXqrlcsxXnbfCP7+8FlVWExN8tw+MAA9Z0H
wk2lK1ciaQzPjdLa6eq3zYPz7c2K+rCp3OfrLgKuwP9yrnZtcA/Na4XWr4zLoEgN86DOQw1oq3uU
900NFc9lCSAWJX7pqP3aNmNYE4a6I+yXGFKIzvM/1qiC9d2em1+cIYxuz2PVZdPsMTJXK4RjTXfp
vhA5pPAD0I5Zw4x1o/gC+4A3ihLW0q+1os0ESjyCP42StnRfRafiABJS2MyG+Hqzpv3vSBhpLulE
Al3SMf3jjck1ZduLlqf8piR7e0IyfD+BPM+vpPYqk+Wp/rg4/T6c8EPRWF0XphnlqNr2TbYpr4n8
GRCyn+fsbQHjg3PdEaugaJeTqEjZA+K4IfjGRUCD+ISKcr9mUGj73GbxpOACNvCTwVorFyVsDl/e
WhqYK1GjpDrSSrWhzNrjmLdRCxjCCS76gggY4upCLBWlfPV7UVdr1i2N7cjMW6amNLtFZujriIxd
+Mf+Mn8RN+QqlDMZhOxD+v0CKWzjXkK1WoXnh6kPaQ0HEh2YLpM/+Y9luG980pAeJ17n4hGOLro7
+MF+6CuNWwGdBAUOp7N6iubzzupmCfuxz58DVZEHErkQ2e9jx45Io1R6XruqXxDuntBywfCW8F4j
p6q5uVXrd27SOLWfDUx69GQCtY//lzg7KSEBWQ8fDSQINOBqS/GWUxRzdmvQMjtho0B3lCfDO+eH
YHaotnNUUfsFP2bYdzbKyecCfbI0amT1osZ1hckgaQLxmL3WzLbyzE95zfg2J5KQc11+68ZhW/dh
nElOkiDFPH556wbZitcMeGhgve23QqYdUNUg+RVM6P16WjzLuAj5daYNlp1+zY63A3ORBBvKjID3
+TfgHiTdmMSafRGZa14XS9kRwrCDLqyFQ7e3M/NGRsJxBDnRRAscSeAz6pq6CFp6GHnJRDQHUAVy
Fsc2a2A4/kQulrP3X6p6F8T+bho1MCLOWhMANVRmR3+8f/0GOvL9ZRXzRFft3owjRLQo5g7JGgS1
YAR1+Wy4SKS4PmGYhn+ha4delphxfL5x2epQ523ntQdXDslzCueGJ1zaRtXOD0xkpOy+yLFywTD+
Jh6ztJhSW6rp2shwgEhu8/ISfOcbBWrfP0Omyf7CQFkfQlitkS9tp+tGNgsN6XCExIfdEE2V83Tl
+nEd94cbVZTAzRKBwu89s3l7g74QLhcpP2AEHRYM5u7/sVSCdhkyH0mGzqIk4IMpiHx0I7ba7iHo
TyoLYQiOPNF7vZ8qEB60CtfZGcXejLdlxjv+UOqFxvSKvzoaIqfHokua5OkIlyb30mWQhzlWsdgV
90nX1GeaeGTupYaVv/oHL3r3fXfQp1ojZHg7MpxG3d9VkV0SDIqlr9AxrY/hl6qqyCKk+qzgtMJM
E5XkjtpHmW+nvCbfRjAnjqwhzPskPYmjCO/IMEgCCOHqb67vv6EggX/k628praS9VJ2yGjRYPyAq
PEj1FuZcQcOYhnubV3Ku4FveSN/n3mkFE+xHTwtkQNSVjzyXXLqmc6qzobHpydAoZO90Bx1OgRx/
PGKLbrNO1MTDbp+edAc9wg/uBlUsEKGgKqqiuDR1RCbclBCmBpZ3OQaH8XzoyF2wBghjAbdi681e
QOBg6TTUkcvNvEFi1NIeQNM3a3tkWpEvFnr4eaZV5OpSKQerlQwCGYCE13lecGs7eadH1B642g0I
CUrpI+JIVO43YJpeyK4wDKf8FjOaop/E8JtXuVGRtTccBDV6nlcLhzWjQpv7K69bSbbczVjF+R1j
9BkKtx2JJrFM8zUnZKxAW8eIWwx8qQNbTbuTF5YSJXgHaHf38Ng5DYKwc5sGq8d2XDA/RCJ7ehe0
UO0OgUAn3umO9TiLOK0JplcAKKFNQl0BzsNRr3NC9pnDCVrYFj4g3p615aQc3nmZaM6UdrAG5eBc
3w0A+AtevJ43FpSV3nuVZzp/Nca4vYrVfHudr+oRAMKZUfXY4pJjmAQ23y9lVXoEYYyXBt2iKYdZ
5GY8h6Kpm5tMcEKS9hdf2OH75B2aCdtSklDBQwICr+O/xfZw7DQdPa4rwcCau707dXP4AuF38f3r
txT2A3dhZHNCNo+m2lKbMTvDmEzHPVHM2LD/F6GvkXK5nZGQD0Mb6Zn0syrCGC4zlGcRzxNxW482
q9+oUp6n0G55OSycGkBQmDRY8IiMCpHCbJg2jamJNcTtxG8ujeP+23z+FdUYf+IjghIPYW4KlC3F
Kob8StEBg1QWqHvUKxaPrSavspNivh5S+Q7vOWPJO7e99gPYgsAaBWooRaHY136RgD5dmN4W+44T
OCjVANz+2LbW1G8XwQm/Czi6KsO3cpKXNarYmMbltwMy1+FAon7P5liZLq6EKhZlIdHhz2X3Hsnb
U30dA2zt93r9j418p9hR8uWdQD+4GbFDAWrHTQDsyRjp8X1uebpLcZcn1Afckuj9YcrxPakeZMtM
uz/xWu1elZP4iXsqL9dSdD/BVqvsdzimrIxnwua8Hppon4GS4MnTM38QSotSdOdLpJ/M8M0mkbDB
8QQ+FZo0CrCKAep7e01tUspfkcsBjzOe9IOgtXnvsS0Exyyl6jL+gqfPeokw8guYC38P4Q8A8MIr
N1o408tfrH1tDGySCiZDcrbgKcwkac+ARgppEkgHGXf4gMmsTXRQTPBzY+Zw4VNsz8L2ZJ1f1eZ5
An4Xdm8GsCUh6M324xCISPq58XqoDPxh5EMJMHLfj3WQEaGw48pFavEe+ANJdV39SIJ27iA1bDq3
88FLFK4+dWWoidHS0p4M1CRAKEuqk2El9yu78mVujjxmRJ/0EihOoJsx1jIMyIC3n99E93MhrvP6
3UeaOxzAX+aNTKcpeg7PChso2joFWl7uG4JGET7uLmctPQ+v6++QPGayFdDEDktFcHMCzYAFbuhI
gwlON4kpI0zSHaXzLNkQMezFnnxmcOqf4GzKaX/PTE3/SfjTMOUtGhwqZD4B1ayvnmytRK1DR+BJ
KV2Uc/15HGaU/cjILF4rNdgN4+530+QWP3A+Gz8dOBklLOKIqzoF35CsToHd3cgY4YVrZ+LBIplt
u3c7vdN+nb/HIQFm/RZvgBgDh1Ljud+E9Xp1wDJ9luuB9aVjsekC8OThxBI8abK2m1zyCBKrQ1lz
y0FWzdPttHB1Y3jBagKuVSFV0kl0/wcRF4FlDt46mA9C9Zjc1Vek8p9QpXz/4zWEnJLci3OKH43+
X5N73y+Zs8T/92eUIU0DxzwPADXfogtIuxJEisMBTyYnXG9OlYStLyBTTqjMgXNIk7rAQSqbQNaw
PghamjfF7ffSAOU9haiAdKnSR2LB36fAlpm/p7VpHfiaUX5iJ+9Zb4gA73ot2jJVTNz8nE/QQw8N
KmphdGRoRyq1tR1/U9zLxEN7ClVPqhCuiC2PQGM2unIHs6eThqwRiFQTNd+hqm64L0Gfn/3niX5n
Ygiqfts03FPBP70wBCBmLJbKyKv3zxMdvA90D33uqSpZurBDUGd3zO9vxJMYpBTWI2iB8ngFU4bw
a/g+9OmtLKcC6Cz+ryrxQ7UfvzESSIEhMd/NuEBFRzbk5SZQj/tIOnqc96l5JE/fw/vjYv6laPZ4
dZd6rYBZ0SUmFNU6wU2jEqvwc3Jso6MJRHYb9tTzzrNSTDVwF+jvnn28dmV8EbHt3yJY2G3/iXxd
hYQLifIllFztin978Ddu4EkOemgTw+znVMG+Bgwkdzbw5JxUHMjs4+NLUOaavALslnFeh9fjHIRw
6cc2ojPaq32aDDzLVesP6/Gk30rnNrUoFTx7V2FK4RiR8T+vcEv8y+6W+p2dkjeTD/rfiQoiLKi9
84WHmWasadeVO/HTgeakDKmQUK4ZmWdPvefMIdsE6xcHq5yF4QOr0a6TRP1k8SS3jUyjn791w303
hFH2D05uuel+xOTJH71xyzko4sy9TfH3ZUV/qsGG1edMkJfLn4y4lDB9m5TK8UdccIs8K0MOuqnF
cCOe8zX0uMYfXChzjF2qZSnQ+HzX9g9e2++EDH82ASqLNYsrNUMItmph78EkUKLrAPSjGOnd8P6Z
jiH9tmeDYjyGqtfvNrCj5LTiRVmVESc3ivPxDzMi6szpPU4KfskqgWNfYj3pvi6tBUdK0wqHfIaY
9Ly4KYTDQbzYwomxGKenTSS1qWkQ9aZxcsW7TMKlyl45zkU50Q3uqC2p7MdU790JxAEGTc/amQkx
EUydoEjZpULiq8FOzzrZDoxeckbXaVhisqXN26fDKaPmi57yIaM3aAvCEdNqTMHa9Q5cOw+/5mBU
i4oHjE8+v8o9DH5e7iwvVvW+52QB0oaNqZz2Ay+dTAue8YggN5eS91X3VleI0QLp08ZaRTefF5Lq
cRCZyN8M1Ue4tFvf0qkLGqBN1IAaCmM395i7ppBKILg6HhLj8k7nkqJxIpnWBQBbYtZU+iaK0xV3
c8cVjdg5vgPAmeiQRcQO2ciXsGrPV8neDcvPREvbOhHb6lWEUo2Ahirg8cSapopIuMn5cJ9kn3cx
fxOwhxZOKYhV3wuvuWqtqeUP7YcNvV+NoCVMqfqZpphv9VW+fJqUJYq7R23MUagYW6i5ZyuzPcMA
ciIJ/1M2Zhh2CpDZPRKs4RumtPuAPdZwwsuMm6SVOlSZ0heOEsWkMyUUYFckeEOtKDAQJGpn5RXh
8JBsDia1MMW45Z1vYXqPRBEKZdOk4fMVBDNifJTBTMGaj9/XIqeigq9DkIJuMq02NTZzj0x269UE
nzY7URX305AEJRLPPCxbI0vQwqmkhVvy8nLpE2uXNDZacHa/ZUSUZXjwbFMcx/4Osd9EVadNoWnd
B6B2WvGw8Kw/4ZFFs6cvGgVXl8YWlbFpLzgDnkbEYqc2KEI30eqD1wEb+9jDGZB0xiZXp3Tnz/hg
49bzFdbMc9GQ5bQWzVVB2QVGOf/INVaC2B1kNt33SzeSFYo45eG4Vn1cMEyRtf70tg2OuarEJAvE
wY3xwnTFQbrBt0vu9kUj1eDJI5Az3IWpIBWNiJgdG+16sWTl0XPtlSM5LFME6945KnOsiiFk811v
oE0bWhxEJPsiOksnLbkDw3PESxLG18Ab/4visPSYBLqGzTFO8JIWn89M6eQWu88jQoBf9TyRkL59
YWlQmi1KeGWHzPZ3h3agYkZKd0+7rPr2riEWd7UEvO3agvzI4Hk9q+vnbrHwdUUXtcSoYDXRcX0Y
KSsbqfPI7nBuoyqqA3Neq7T8YzfDXDJRfOfQKQ0xiJqjB9lzYi6gTto1gn01aoXvp3Hn+nUOfu3T
ZXrkaoXQO19WyoZW7O2o6uvjEWTN1Glw4zfrA1nUSIufDd72IsxrFco2HoPOZUNhFcBnI4I1Ebf9
lA3SqD20LC9hO1lw9/DWF5c4eP0MlK0jsulfJKYVq3juvVAwG4fPW7yJ/+1FZdxMgQuhyAPRFnmP
duKZcofS870NhRYPGFuhj+TtPwuoYgTLNbsk1mS6yDQU5TQNwX2mtz5vTxCJVOa3GE1LEi7cQQOJ
5YKke6idaBppB6udKKZy/0JvIzHRzAwrkWIOpVWUWRPOf3fXNXMtzZr1lerxuAl4qHy96J3UVyzF
67ioDJlGo8apESrvsQNgmdFScCgq7x4BHHqy2a/NIUW3dIl72MkuHZ/v6Jiq3DGRCIWsxtv4CJJb
V24XEvNsjOo4qNrgXuiFOB3aUJPdahtP+mnITHTAcisbuIO/OINNtQaI5FYhCR8AviLAWZSDrGUH
o9h1Ruy4U8Gd0s0FAPIkXQxoIphmqXHhu4/jZ3aGJ41dbm6K1vl3eHQ28iKZnEkYTHNJvkDXZ+6E
yfVZgpTXqlFwwhz3IeScCTd9G7EDWsAbc9RYvddvTb+LVqLsnROahkZ0nnKwBy5PUu8Ns+CiK/bU
0iXL7hs95Ow2I5gFNX7YkiWFecz1s8CPHTZKPJdHaFHNZUDeSzxXAMPy/C+Rgfr5OYe1XyxwTIlA
vG50ZDJXkUrSGvMt/6J/xfsHAmmd/j4u/WI6VJgJDOeW0Kfgt7+pQ2ISBrVEdCZusmLG2r7Q59Vq
3+ubQuVg12NASwANRPDX1RXsE/rvRuSCNg1BX9Z63TaxGehxbrh407U4iWeegTbEWPxBouT7jtp9
4UUiGNS480FnfLTsaDfQv1dM5Ia4SnXxl9XbmX/nKiPmOaFsHN9veKKtWx7wW6d8qco8bwRn1pox
J+bY0ZF2xYwkqiPooDL8xEwYuXe5msKh4DChvUWo0mYWCQPaifjJW55mms+gTzUymeaam7hJhae2
UA0Vifnr/np49OPKEBAbsVafngrpIRg8BH8i+2dC7KCW/dGLOwjeEBhbsqBxNMgVaT71pV6WLfvT
kZ+DwJrZ/cpMUPnAPhnzPVYJG88oDOSiC4NWkJ7DkgqCRfpvEyW8Lh7fO/+V57ni1wK7bZYkZMbJ
vreLiF0oKSz78YrCub4HRNKlsEjTBsYDaY2GYzan4aXBB/xv4asQ4VQLkv9OvvTIG4qPF1uGhxRE
NP6d/ix3Hpk0tluN8yc7z5Xkjeg/ayeLExe7UCMArQ4tBqxJ1RezLrcc1IceW4lcFjb7g2B2lQgj
YNb+u0x+KqkerOJfwQvE4kodzoJr821jyZojln8YQwvSDZYm4ykvq/kZxnVjGXeKG+bxu87NHQjf
XBY/hF/pSlwg3pDiUOPVhe+yRUDp6AptbOUv+1xHnRdHGqTK/krC3nqMQfoNTFkx9NLL4QuAiSct
hYJgNUpiB8NUvwX7FnWccbWnPG8F4dBLyOQk2aNl4WoZ0HJrCr22iqlrfwQIXQ1jm1/HednQbe+T
266wsFOaLw9VjUoMvSNEFpPdsqN20m0Dj3+lItmRsl/afYORNSLqSpAj12YnrFxdTuU8iB3TbuMs
Vymn1b7l2W/QpSU/S1bLLFBgJ7ssze31pag07Y087e7VWvImxfuXjlXLgy7YPr2mQJtoI2zUEWud
i4Hyt6GjExnAtocNubUeC8Kg9UUsropvVdCDDWyV1njYqs0hDDC3Doo3p6jWhhDkhyb3iivV9lSl
QgTtwoB7AJacDs884h0Rtttqv3HiEB8S0HuCh/AKLoL6foChosnZdqrAByWcEo0euwM0LxOV70tX
0zksowuTGeL/Y35dgj0DW6vwYrl1V54svu4jKoCAz1ko02ORRr5SU6UtUSFSjuDccRNsV5neK3dU
Y/qaclulwGk9Ej26LyxE86LBBypcYFFk86vjwXKaM3gsSeNI2i6fpqTdtX8M4eTmzzTLi8vavn+Y
l9KksjXSGFr2vfRNr/+e2inzcbJHQmv7oZlQYLmu/UxdBntE2DA9BGRCtmSNsCqBy7fcG1yQ65T1
xb5TMN3E3RMPlHZWTa89RLPQVzycoFBh3xbenXZhwXgzuucWhaJgv7kDjDnmVz1tiW1+yA2UOzHy
2H4BgZWMsgfTVJWfspQVUVjWjaQoBGqnxDejWvyfFB3Ys0rkyzrZJGg5P5XqIrUPvueEHseqMw5R
sy/sNQyR29BqnX7zRU5ep7XFXOeCCGXNI8Q/Q1oeNrkqbPvP5P/GVpnvWL+wtZbQPhAyoUdmMICL
Z3UDucZBQHDiL3/HmOSBBPIpzlVRvPySfm4NFm9z4iLt9S1GjHIhqMu8rGrhZh+zHLd5OvAjOFRz
twuu1zA1N0JP33fPJjDQGaCpYY0POLd/JAlv146ferruluSmQu5VtfiQELtq6GVGzB7mQ+rUywGm
5WpuicJWesZzo+zS4RrBYb8yKBfu7ShtIrnK3hjVvH/c+Ud4c1Rec0asW/4Riruie4Crhb+8ct43
yyuF32THgYjn1t2vB2zUJkPFVApyvyKcTEQZJpRR4OEUoklXTk2qTE+d4LqVR9UKfwKqHbrHnHX0
4eDxslkC0ocP4iJw85uSFfG691f94Yle3g/eOQLLl/W/y62BK10LNlV8lywQ2mt+pmnhCja3J/jB
JxyACugvdjaxXJPNEwnXbTlFoF1fo5Mj5y37xgGCVa9CKxjuY1dWzAAOQ8fWy4OiTHX65SGqNiKU
CANq8JnLHJSgfq9MLst7k8ydOAA8ilIbTL+UCLiK8y48wqGmRIx8otafm2CaVPY7pbbaKhHGukYe
593AvKySA8B3Kte1TlNDPGU/K3dwtznzRZ0rooaYkeoyK3turrCBTU26QxCf6fJQgsvO1bPS7z/f
4tKRcff/oXtgFjJ/AGJiqnnUOg+oGCB95h/HB082oFubbDZsgb7H6mYdLLeuL5XEKPpahl0uqEXC
dXcQqgLtU41j2XlXNfxOouBNadWte39Ew6wHvnOstM8WlgzWaz5kOXm8PrgRFkq7AlXRV+1L74Bh
wAxgiKIasHwnKEaCVBw+DjPyzXLoMpblyPYSNak0F3tVaLqjt1M2GF/bDCXJH/eRuitqnPSlFVWf
XkuHGjXWxFSmOMMM3QWzITinh4Mo4n3bSJcrv+EHCNrt7xEJC/R90InNoRUhso1Xbai0XVo6w8ut
WQ/G5Rhaf5bbuSvtY/QIveWeF/n1Us9PSFAqI0vcfUVPW3f1CwRjdjsDQGwuqKj5Nu+zzbcJ9XNZ
Au06QAMqrUy5Ztp1sOvfrXWF4BkU2ZFC/1QpsEv26A2EasIktA63J41Jg50wj9wWWwtRxJ24ZyDu
dkL/TO0iG/ijJEDnhQb688AbRjqoo2Z/A59XU1NjRQFt02c3J221XKPg44g5af4o7reRi1Vb+nR9
ttFgnKwwW4EwoICVBG7YkJRzPpub4zQQH0sGgvaX5X44Q6VxswLMFUDQ3knDRBrCy3LLZ9kxQ/vZ
8h33Fdc0WJ3WIMH/AIAOfA8pY3uLIjdGLISPr6AkbV57BpeoNPI4bMChq8MLVKr6enMvdTJBaA7M
uOmVMrhUDlIIJYDZ3HcTM5XS0ia0NBaQZMdwMjmrBRKUgNPMuziPwa8rav0e2mO1+7TGe6sQM5S6
P/DWjfckyo7MivksjjA9GdLtqS4GmQWy6LtS2E4Tr1zvCQNK3ehSuFXk6E5xcdQCGlJ2MUHIa2fj
+6jcrbLgVmmYCC6oNn5G4BUzTGDuzZhMp0CMSvNHFBZ+YNmPBwdvXEmKK4E45oU0jjQguNs42T4q
3S7rbQXhlSWg3D89W1GKlBSe5zF0DFolqk91p9VCH+oWnCLumevTmu8uLCjOwkQH1llEUZH+JFfC
cBvmg2t3WAOkpwqZ5c8i7uuo6XFWAmBrpdyqI8p0UZiqwUX4kmsDXBo913q4ZMxIzh/o1UMh45S3
rLAytVfkJOjHadSS8oEVxpLQatprVk/0ssRRct15FxXWNBSbYllkgujyz4IBRJQQlkzUIDkKAkE7
lXMvFhiQmPZCKtLca4Kd1e624AcVSWi+FznYvX6i6jwXZcnDBFffD1zc2mBVseoqs+sEzaEoW9Ac
ZkcryGpI+iFIXZQumNSG2pMmgajZEwbkbdFRTCmVbI73D6qClox6WNXI1VMa5CT8MvCOTBXqMCuy
81il0pcos3VzPyxpY8/cijBanCfJofZIPBXorlMjXlAjVSLszYMeAyETmUGAGFvtUR5YnGBPhoib
RBw4ZNhtGTCvlvxYdQnI/6RxOy7SW1ZOd1P/FgaKL/HSpVD0cmohVhZZZyDLdGo2VPoaB4l0f7BY
06o7jEaZgt6Zq8xaX6Dyb/bVgyPlf2Jw4ftF7A3bfSthfZLqV034ZAj6xlV3YyqMc8GAMlGQ8YwZ
c/AHr0SpkYupEA6eEaGhriU+oW942tYcCjf8sM7s0GL9vbV9D40ipZVk3qIYjPbTK1CNiu1CgzYi
sP6GsV5woVDoHInJROKXMN+sJQ0joDf0xOF/L6XWoVFyHyuKmhuibPrUF0p1ICgaGawxGjrgcJdM
g2gqgjN5I7SZ+yHDrjdl0dTVj2mk2ueWjs5Sh6vz5JtDT3PgxNkp5Lm+hYTq+Kyhr3GE4R541lkx
fVAU+FVlOwuBCs4D2UQyeqiB+IXx+5LkPQBCasrdiqz/wS83vrDG1erjNKPMPSn5vkVcNDklXIIE
WXmetp433Zr8cwOT4DEYRSXXFQ+TE5lgSmDDNSxo68xE9kRsnn4gWsbWVw0A4rXliw45t41ah7lv
TeN7uY1wD3M9833tyn18tgyONda1FRC7Au7XjQkpKUiWkOmY8JykPkv6av/R0OLy6FLJKmHboEhD
NERt56sam13373b8uEwMp/6KYlNS5SRdQDMWVEMwZuJy2AnNM1J6t+WzMbg5pdFAWP5vMLlcCLyJ
thNg/ubFuymNome/uHYUxLWEm1OujfK+Kir8k/UM0O0iYpbXoffUsP+3+uxAU/RMmY/T+PCS0chJ
qdCv2XgXP8OrSwbxxs2L72c5eZf4dIFeXZmVV8gBaZBZA6YE10QkU2i68ArzmX41Sibri5jPFc1+
ue0WvqCpSTEbyWnfHsFlheA8Ce04fAOjT8m0BhPrdJTN6KW1XxitW52tUldjd/x8mOW4qWxUyXx9
1i91EW4fA0BflqahqBa2teHvMCdgTt2yhtevb1raWCtni6cm/g6od61gwx1RJ/ErtHNnG+7UsKTH
Svj1D5Z7yKXq1HrV02AeROslLQDxw/ObzNqvd6D0Cxo+m4led2xkyI34XGZ9iR1QEOla6MyvdhPC
Oz2d4UF2r5rf/dofB4a1eCyr0gQJBKNLxIeT9pF9nHpSvkhXdHlGlULNuNHGnpyc6e+1Sx8h+G7Q
pT04xxaMNTgJF/q7UpDTkuCMK6fEVS4N6GjuRscsfu2+U7Om7CJ3tyUyJ2VoRMmPzonblkrwK/iT
PMJHZuytvMHo45QiH+rkMA0l9l4KIR4jIfsEM7MwQS6bpxsuMpf7hTGXVmIjlDj5Xm99gpVP6NE4
YRn4/cda79XDCAfIZPMhBFqohqqnkJ8TFUNc+zOs19eBLJw14+6vVGJnG0WRItlqcSvLWaZOeYvg
183lOVgUP3J4awPhVsJ4fgdJGu/GjwKpGBabrMVBBe+vYMTLekbAOvsBOjg+gCvYyeCiE6RdRV3g
znwmmLXAqXC2JcSGe5GQgmiNeEOB08jmz7J7bDFRLwGPdDZ/roukmRJ5cb15cjuVlycJHRTx+7fO
YZLQPERx9pNaGbpqsJPKDmNxYjwML5dIn1EQnPJn4fK+qZiJqEUvim6xiXwtqfNHP1hWuF1gbu0K
/x2wpWlsFNDEjN8eUtXXWJsFIf/shRa+57E85V5/zgFs8bOc1eyecFCaME3I9c1RCFxlAzXg0u33
+cXZ+AyTaLN9eeWbipZlieKu1rVlLlvdKM5l+/BnL2zwesMqby1/an+JK7las6AfAuCWODq6YU9a
vRDSuiHOhEvAITF+fzlB7DlmWetptfIBubH5w9RILPBI8Eniv2e+jpkuCydvbDH9EYODXH9t2KRB
JJr4CTm5xHY+zgN6Ugrm/XsjAgnk5wN/nH2oDs7TPCpFbkp/3QhtZZrzTkF3bnf4YYQvXv7gI1uA
hjcijhXMqC1d2L7UfibkrUmB+ROyDWFO1y2v00QqH7JpXgqKcMzzkMJS3DBVDx1a1qBcF98Wg729
Xks31Q9/QIlQKNz8+l+v5DuqvarDLMMl+1biqqFmlmmU+KhDYYWiJ8nepNJgRGU7ZmdE05ubx+WM
+bz4bOKA+VGQt5671PoKUhVZYlrvNBcZE/oyIjsrpeRexHhFZZ4+ek1XLtsUZeK3jdwKNkOqoLuL
D/JnacjSr2GcjXGiXdQcjG4cMifh+sS6xwNS/sI0glceELlRIwq+9EP+Q02AW3oMfPdPOHA4dbhb
psCRtU8xjutZG3tb9QrHzPUZSStweHPhdqkQwnIn7lg6kpu1Ug6xt9jhxT8OUr6iaQxY18HZYT07
Sj8eWlEm+CqaV+tpMf/+1tG5dLoVBcq6L4h8J2JpKmhJViqLELXjj7J8xbT3Q+gW5Kho+vDncP6Z
7co5DoJ3/PqGeVuAcyAiTJMCxUeVVvbJtCT9IYrkZzyk41NMyS4XvZbGKbmBxZ9IV/u0XqDhb+mk
zvs7TMJBa8/Oi4fQ4shyG4mxpsYI6M5k8+tnc5gDtHA89dkmWSDPqAVIPHe6ZkCOjF8nosHmIVja
ULZ/WVnDzPqLemFrNWzlUzCQw3NVtUvTgrQLODvi6oVvfodaOpewcWIDCsw1lNd3XY0R0TGCceLv
O3NCos2wUH6zVCtWIQEAburwGSApn2xu3l5d89YQdJvVaiOgzWvp5FNTgXh9zNb/AURx6HckyIPW
OpCr5p6sWfvYkPWrhX2aDZ5jiSvtTGjmC9bInf6qD3eOouexRt/HBuBSuBk0FMiMEZqMcPWey4zV
Tn/8acMV10KFoP94uTKNn9qKP5w3B2zFBPDZlWW+hq5dIC1i6mzL0LfrKp5JaZYHsVbJ7Lb/KodT
iG5NtPs9bLv17YCCP45mtLwdkX6aa3Uf0m4cOlJEVdPtit1vdN++pPsmicIzPmO55eUGe8FOUSeh
W/eNcSyJxu+jTcOdlcgKbnhWcUXlAIy7+mXw0Bn3egQ9E1QmPK8grlEmtXk0zN95yD/lKD+trsWK
vlGWHLSkhf6xexYCwJtzJMu4ijAVPHAWiTp7s05A6CSbxpDss8NkZRneA0gY6KBOM7IWaXYInZuS
yAVS9yaxL8NIcdxwn0QzxfJKDhup8B9ZdoxZ+2gpZTN+motqdel8KQtXO22kLDO2Ao+o2OEAfcau
MjkHZS0I2+joWrXE71yydIo1yU9VmXMy9fOTRviLcJXFBcvwGr6uQoo30T8Fs90ytxi6JSExt+Ar
f0cpNgfY46CI4rM7o80nNlvJj6dqAEq74CAZb845qqOaxkd4V3dKe5FjvV+DoHmNjMUmdA5BpeQc
TWAUbjEHbKWCTeHo9IN+v7qU3Psakw0wppdiGwMTN5PWoI1NahQwTPfyTGvejp+/TlQq4zN51Dpp
KKa/p3HMyC3dTgLG+h2ev8Eg9gdQNLc2aaVx73mDrBnEl3ayZ1MMJY7M9ix9H8EcKW6USTrBXrzm
GcsdxQE/ff9BhIFtCGRdWf6EgRb3yuia1KKDAvgCZ3XyN9XgxajEwnlExgn0Wmt+6hN6VqlduFcy
snb0F2poNdyZ8SX/mXNvnGYqs3wiILC9REKy91V+EFLIOx0RIiOvbde61Nuf4unAi7cyQQxXsscC
qrDk+jlRJ/B+cfw9yaYJpEuP/5PSkodkXVlrlaj4doOFqRu23CERJXq1wFSNVpDag9N8SgoVWZhi
zFDSjZ3hSNRy6UDAxJiDILh9HgoEfsgtHmnANExg3pLQOZg3dGBQJCHCzRd9jCR6/QYqQrHsg1FP
H223vVHMx1MJrMLliBnjjrM17E5EYbO5HiEzGXFc5VsZMlIkow9wd/vYcOUlZqLu0iVLABgB7hvF
4MfmkGyqCISMWSFuJabNcv19fotZPXY3dWQ7P+8ULazCYYu3XgJwk1ytNJjkjVle3QjlsnXNLvEw
fc+DUbchfxycgm42lbkJsu9j5G5v19JCFKWUTcmfZtrRHfuEwRkV6cxeH8ggOsrISkq0Boog0UT3
ES/cvAnuSy9xZ+ZMdhtC+MdAiK2ptOcdTabg6PZzggWWhXzS9UhpO+SMh5QQJU9shNftw7lCRxzl
nOdur0b2+FOMLMWqpIL6RdrrcApxdI3au/0SgzW7ifKXo4Y/fAOvAa1+1NkTLIxggu1OqvSjSbzP
8Ai0OeVw9qb2PWgWO+plS7H3qwXVi92f9TnaR2LxqLWJuSEPR9pMCX/TRBSrxa0wwykTdhHUrph+
KfNxd2gz5SZBBV7s4AHq4lbJg8Fe/MtiN2nYGXBxwLqddDkqCJuWE1jCw1VherKEVxow0sLROdji
/ZNX4pPJ4sHz6s124FZEkv7epbZfuQpuMfummR/u1BJLZ1O7FSn2VP6kxmk2ME5vvQ0x59I4H+so
4zSw5uTTZf216lv8sf57dRJkFaFnHSJTVluSNVucXGZCQnaANy2cythSPVgZtaxl4hbLQW2RKu9B
IPuMNafginSXGgTJAHVlwP3Fw37IlXGqZ6A2mWi4txlowc4MU5uxajNuUdyibXXE6Tr7qSaedEpq
EQKrknAR1p/VdTfiQ8HP3WCuWJRY5lmfOQQ+FSfHB+Am4u8k6dKKtXxqLwWL36w8tPRPeuoHxXQl
hlnL9ebMd7xM56UCkwjLIBHcgaV0DG7Jm55PTEd34gImvLkq+AfHnq+ASwI0mmLQfIv+uPsZ/EeM
1qXHXWpDtOzze7gnnlzVPzmJJLQZKQaBRUNcqJjblxiqAos9FK/uzcG7eF7puc+NHYDCzWPGS4Vy
POFMB5GzqRacEaPb5TIt8NHA2TudQhp0Xc3Sd7dnAriAXmjmcyQFFBV6cDBflrWCrfPX4rGUvEyW
iKptBYON5DQaGWQTuPiajfing4sjaiqGu6R6e5rQFTt2+hv+U9DvhBGh7xwRaO6UZWADgVhzj2lR
/eH+XAX37JvWzoyQ8c/S/lwFxyX67aOheONaiyVxuG1tPhcOuAGvi56TMq69O0sp/fWIFONsms62
W91ZTkqY7T2QG8I0+VhEwrUGL+LLCUAYQlpe/31BSkhvrkKPJ5aCxTBZnUCwtXPPtli/w2sgFmFj
O5tPlG1UyTnPHHy61GC4nUeX1Q/AGn7donqua9ASJd9r6tpZTA3xLvXvzWQXCD5K+bF8PhIAuNNh
kSrc8dicYVXexjTZtTmQMaCc4n1ZjPAZurUHyOfs6lEfzamz5l+lTFOhcuMO1w3P/rp2yGT0q0dN
YGOrGUTWYCa7t2yYSmmmBkGWltcWtMraw43kaYU7Wbxc0UhpK1bEdXGs8tK8AnDnV1qe5oqzaqMf
9sRhrNqSIwnIwMWpGtOyZfGtEwOGCAjJjz6spCAKp5m9Xjbfaoq7003dbj7P6jfecbQX4TOUaMg7
MFnzh5qO27D1B+1Kuh8f38waGeeMS83BatMHLiwx5le4GYy4MiebTx/U1hJk/Txqim5I9WkasuGu
1EFoIltdCc8v38llIPuUJAQgokoBnnFVRP6X5xaZBDeW4zxf5CSIUd3bbpCaaVDhWzPZj4KxekZ/
CJCcUDz3tiJxs6Vp98HsxCeD1fXRTQwXv0zmtsAUMRAo5h3vVLKNaaDL4Ffout7v56kdp9ZxnlMd
7G1rBqlueliwsjjRu0OTp7rlBW1iipAVIqjwqKmqIjRgpzMuuGoEY5oxw25LxLvSbiN3fkhilEqL
W9rXABYIGB7M5MCL4V7kuO/VHJC912iLPm0S2yMA7eZPeY68eeWHN5TQ7qt//5xj12zX7dgAx1ZW
haQ5nSUpDvjxwOP3SN/B1UYrmhqKeugvxWi6m7lZEgKhPJxBjc/pw4UjVTcClEPe4afoeklxWORN
rb7du9oNtRh2IZX/42VvuguPIgsof0PqDqmRrdxMIkaGPHb33PS7wRBwP6E3vxXbeArtk8RzWv5K
7NHsj7OXARLbKKJTW++j5iHTgfSjqO0HiE+83KgZ9wSZOFFBO02N1lfEIAZzD/bBQsfgMZIlc0bJ
Z56a8wT2Ev8uakfVr38UqQ4jIc/xW94wTd2gPJmJzMJE0BJd2pM09O14kMvkTEdIwMo+lxKR8A10
WH6gcRWCryuOv1udXdI1w0hsqpYGmSUMth2PLWe3BWnCVsr9s2NhSdx8A7MxKmpRDloYboi2S/1n
/e5XE1kFWDQ9iA8HdHi3SGU8s0KDABJUzRXgXUKbK71fcJ6duUIwH1wzTza3iR+nxghnp8HJL4zf
iHqd3iZ8BBJOiQGswXJjQZgamFgo7USZAXI1GALV6XOTucIyREjOI0wUD9OxSAIij2bokIxLQcoo
j0VNqLgNFLQMmWFes52r47vT1/ELmDzKoahFI5uMs+hV0rYvsQqzeYWwePolXItskuNI8+0vCpdS
5R+7q0TU65rg85Pt/2n2ZN2Y2XJwoCV5dLr4Jzhq6PAzdAIf7XDz6vvdpU+cY1qeUW+YZrHUVowZ
PabMEAJTqlS40tqpDRvbS2rno/GjFzqqHuHkjNvuAR0wMhY/V0rvHhPQT9Rm95WSQ87hFmuyPSgd
OhKlpot019CuDjCZMxtf1iq4ipgCz1LmoYWt+vyz2lGbVzWA1ktfRwqfGz+CDnwOtf7hpJBsZQuz
VYQ67a3Kw9ljNaOwyu6NH9At5cVNwwoOJSlNPaDTqxlPaLzkBhs8rqAr/GZfS8T6iw/uKaO99w9j
C8GHkdQhyvuauHcguiX27s7yq34gDUii0a1SxVZRhNUjJZpUbd7t2C8VgOJuOVJeasD07qpWPUTS
8sjMTlEr2ehqHu3qbIG58fTA8TxMzl6pH3X94XVlBmxJxsUa07W/0rTmQbSQ24EOLa0pk3B4PitA
jHdA27Zao32eKDKapzHgWvpcaAABc012dmlghMybFPlvAVgrctExrVBpeKJqlT42CMVQ8hLwCZL7
mluth9+KKqhsnh8wXCBMnepA9FT52y7RnZkwHK0lA67nYAM1T3GxArLqlzfV47tF+vxoGMyGQ4sd
pGW1Fp7JfDeBXG2OI1dLOYXi7nJRnv8sDTnFyCZdNe8hR6I9mj/Kq05R/3B0g6Mrpmy7vVL+tgoP
WJuyJf26cVHCUARagiKgtKU3SQxFrdrFv9jQDmHpLgLBXPT2HPKjMFLYrDk9JolCgZoqWkev2Nkt
MLWWA1rQweI/Gg3q5tixcSKmim2R/cB7lWMASv0IWXSpei0XfZgC4Hv84pochinpERbFwtqk4hzl
sW2Vg7BOAmPEiKDttRLVzb5weoJInLr8H6A6ks1epIxDGQPGV98QZd46zpqStwfgm9Mt+tNwlBUs
1ppzR3DTZ3ubVa7WBWJVE9PibTgaAxnL0zGGvMWhOmaMxO3teYZz4c44IlEVocCpfxVexry7XiFT
jzoVdXvEVKsi8qdvIhkigcsdZ2vHJZk15hR2oko6eKxkhM0tgOqrOUxIKBzQNvFGlSb2dJcAL5Gx
4oindTP03RMsudh8dGQlAnxomCiRzB/ugcYYichWJ6xItrVo1YOAia/CpgWKt4m7GhS3ikkWGome
zSZpFXsqAwgbaiyBSWJZErSf9gYlxjqWbw6KXmwK3l9OZOvKNw4Vy+1t3SxV8nNn8u9qm9B4KMJs
AFuw+mQoTW20FT5JM4ZAAeTtffGCV6qdAw/ozhLcjv7b7SaEORI34CqNa+ECEaLq3BzWsctZaVAq
7tipbsd96sU124DqH1zPniwb0MftLEz5G+7QKNTJPQYvXjfrddFhyeacytG8fnyDHTAQ6MC7cqT6
vKTlEyhwplPODZvxMAEeR0O8r542+7PDE3Kfh5BVPLwxdsw+Ba93g+ZL/qO9ViecaItyRcRtfsBs
PqzTjtQSZmuX2Rbd4qHekipVT9wMCdiF4CrGYZGhxsThhjA00OAiLQa0cbrSiADs9P92wtjKsgb1
StO6e6XsHc8qW+x8lyULghtxfWB4AExHUIn6lZsCTSeAderdVm+Hv7fy96j236kHN1JApg3gJMUb
2hWemZsR3OPMHVzKWtakdJWWjl7/3tbJyE4AWaPcaHuNtJ+LcvJVfX+jQyuwy6adJuNWAd+AqNgF
0JkVFwug7Co3vQmHnLQVKIV3xmqsy1OFfFFY0UHZ17ZvLa4gShAqAz2dbb9krBaXrN5b4Bcyzj5C
MNhGJcwkC+6spZCWDfE0rj3+mF3ygDryPbPgXv7lD5KdQW6XU8802avyewgIqPDo7QB3H8GBs5Lh
XEF4+8+PGXM0aXpH+Es17tggsYSPVPqsc/94j4MuqMOLPhY+rQ132Ct8heWFu6d9RXfrY7mR6rfL
aheNcbXsVUIOwdisFM1HaCOg/bMw/fQWRl2fsgj8OQUgiwIkbD81XcT+dPdGT0ezDATeoY8koY5x
YyLsCh70HrGV6AbEOD03YhbASw89Hn3HcNPfxuvJQDvZYywe/EuJZFJxtAkxzspSVTYc9+Rafb+Y
guSvCQjbsQgsFjDTeinKE3RTDsw0r53my5RBUMGTLh+ab0VdxSwXF00ihweWy1yrPSuvNrFfyJ5I
CiVqkop2NRVnxEP64XKedcdGx1WHGgJlPQGaVNxcCOcEe3C4Opsfmdkk9IbS84ed1MKVdCdSqgGE
PMlt2Ex7eWe1GmRBKXWGU8Ddg4rUoU6IywuY9byBvOse8TnwpwIW4IrNLE0aZh6ss729iAFvVThR
+ZHtIR9wRic0zyRwvXRhpECbMUHDUBjxmB8HRuYtPRJ9aleNRWTlgLGle1OQ1i4YR+oQw2jWziOh
fbp7XuGAVLEgFmZRZVr97MUVkZsdoqQOJ6zBiVjxqhS6BEF5C5r0bzBs0Du0wS6GdprNn/UExSqS
Bv0u8lOTKsLy0AM4KLKLq0qwj2kGgirXLR7YR8Nm/iwajvwkj9nHS/U9Uxfa1tqq2Dux0LUriYB2
hMODSXLhmNdgs+o54u9XLQ6h97lL3cYY7U1SuYn4tTlZAN8RKSYcdtBwwgscAE9Tq7NhLvgbfSm8
JuiswszcVbtCqcV7Gbv5JFt3JJbQFABwD7PdKdZ9QMEqOu7AOdsx4YfJaTQADvgnvJ1S+2nSe/Oz
L2hAb3A18dgF9OpC+/vnvTxabyqUWa0l5L4UBRxx7QTIpcfJVwaDSeroAnqcYs7op5q3RiWCaj4/
B9MCcB9RlNLma9luAW2Pq/nos+QoZtKWLXLeDrA026Yc8dcJSL8MJEfDODzZYWjDQrGV5oEeyT2F
wfRBPyqhvMhq/YMlofKz+Yh2WWdFiRjXxdskKHFjDnDCqMZHpfpqVEOI9aerBUYUdbKWpbcS1KQk
WUuYWNVbCf6+Frey1SXbNNFK7oLG2hfjNbJE/VpVOHxaOn39j0ogciaMGD6p7AOVMvpi7Vb1Xpq/
L6QRfOs+cdk9B3f2MdQ32nBP//jol92noYjU2o7LxnutWAl8T12+YQj16wE8d8wS5W7itYpEPttv
iSC3D+ELCrIqdVzfcprvPNjtx7tsWlxJ2UbQ9Z0fnosf2tf4jKKmfhdl94ZX99Ak20Z7I67IAqKo
ky7ZCqtdjW/Uhar6e8JgTtgvBKIXbzeTUSgblpnsK9XnB0tgwrbrVDAJKs0Oy3Y8LamK2LpxEhu5
wFpBdoxVniY2yuPxQyExr0hnlc2HGLxrcOYclFWfLQPC569lE1a0sGRHMa33OFO+6ZJMSkT2X+xA
d7xTCGuYZElY+I5rd0eWRknmBPWkx9YXs3y9YCcmHLcst/0eM0C0XneCgoDHsMQ+GHYjIJFcAEHQ
aKIBjA55M4yNYZPVWUicpikv3ZTKK0SDNt61X/+8tiLKuiRx3Q6WxElnDc/MTDCoY2oLNlg8OZNy
lIXXO2umV9BPs1uyfPPBRi+hh3MEUzVNVk6zCLzRQKHFy87V8C4ijDJykLfvJ1aA5mXTnhxZ+KVG
TuWRHUxJKr2ZTNJHnrh6HxFtBTXHq1s1HIeF/BHtX73IOUrHelNQj1+u/ZiDtKsucwnU3zIyzPVb
PAy1C9QCu9d3ZDQ0/yFa35b+u5vAlRRheq/y++z0xudDPmO6rz1dcXauLppl0ZP/JM457JeqR7NT
uUlbYuqa7LA95PvFLD5+cUTfj9K/AKIa6D2vZcmYlcbAev9O+AOzC9EWSgsbfQF9iVGo+/5BV9Ag
4GIekP3R3l+tTy4qfZ0MXqRYryZt5VCEJUw70XJDxQbR7U8tYiTnvSVqgZQYr2TmIRI6mPcng3aN
fhrTUe3l0O4oDp0/aOYVcsFN+7O2JM0q8GUZ/rvkkfLc8MChoXncpweddGC4984GSetlhjUvIXFs
s9PbIObg2pXOwcL41mPM3cO4w008Es+DmK7K99k2JSjw/L295T3r9jAH54hJUEJMC4QO0Sh/CHT0
V4QHexsEVBn3seV/1flwNwF1U8QiVZNzL1cUlqE8mxRzUvMjjwQ0Ln0uujuJHZQbaSKi3TR1zJms
l/COrQI6daer5Zeupq5S8DLHnXBaxWS80AtY1vvwGnxG9AEGx6wSKwzou6cX0ehDh+5oFmRx+/83
6VhA4sEceBM3bjSbd1Rxd15TZH2FW6Xab2e/jS4dZZplZQcnPDSq71MlifcT+yuBmrCEe+KBD98q
EPLrY5Tbi9mMZbnnWpq+eh8hB27BLMwFI/lcWy1mFhCrHUV5+7qCOpLe/dURdiTEw965DWp+Pzjz
vlj+ek9WP0VfXQVNPO/slUQRZpIjgdgWlqOf24mC5Gn64Is9ODLbKRoWR/xnBlNbukCHvojD3FuM
s+y4btDd6lixRErL0sjxYRWI4c+Fik07YDTakWeO3v3WsJqyFzwD4hgAfEf2V/TIUYQGdyvRAUSx
Qnk1mTBIjI41IlAdlGKlc9yom6BxJhSFLvpzUkYvPxiNvTXHKM22LV0jEJZ78je/GmH46Rmc+Uwn
0kVXxwu/irkvH71G6GCl39sW55zjT8Dj7//IFF6Q7IPE2wpF5eovWpdk0gAvkuOGbB8H3DA1oHll
4CFYjzFz3DrEahuECMsoLPBam5RBcNO0bujSZOGZ8UEWsgEoXspVqfCAG+SUQJAXSAWkk6bs+Y0c
yzKpQok/CjmOcU3mnH7qETXXCwRGT612BEzqrdT3DNAVMfQ1Spi2D5Dl+U1mNtCUExOfkqCcHr8f
fTToCaYY6Hn9/tOc8WAJuESE5zG5gFG2ZSnX71BkfwdVS8MeXdiQdckQ0eKaOcSdo9hKk+wmxl4S
moEKJbqYL+ouAmVbXqAvWlQ5HAVYdD4QahMCNAYKBqKr1PZQI0QfOzcrrN7Qx37BWOF/hKV82+3B
thyOtqkgZOfPsVpdb4BtToLQJmST7vVk9UNKcbJSZzZA4oZOy20zKYd0kKFCvU+V3rRYF/CJRNMu
Kt6n0zmhhDnGZUrWf6VQvy82qKq8F847+uF+hD3BqhKJXWVAdAHQNs1C3LsQuO5rGewSyiVvt9s6
sLPi4ac3974mug211lHjl1PqMZv/vjtcyo62PixBbllKjIqVUAgMW30FlsSOkvTGzSlNBkz4MO8y
FIGCzLgR/EpkmTmtxvrIg0ysHH1X6zscx4AFcU6bMMwOaI3tVYcxdr47TSInL6DS7jRn2tQhh3VG
QqwFXboa7GpGSIgDd32bFlrFn1Nm37YHz2dzhAuCMLiGaFUUnoQoZzciTcg45FmQM/sExBTJGhPI
owZkCHM5mLrd2Zni26mltISwb8QcerGWSSVJpx4gqXsr5eObgE/M3t3hxrEmkQU5l1IbPNSA3DlK
qpXJJ6So+tk7jB0hmZbOBWFukseWbBvHmU/32e6e8FqV4FnMIH7tHd7fIMwbTqUK8rL0PBSjT/fS
uXwCjPpzNgyI1TThnGz37lkLH9z4F/LStDieh1pNusIJiw+5v3Rsewmn30huLrcvL+Y6X34/TBWw
NsnTK18B9iCu8W2ytXtmZywzDILzxFP2wrGDBH/t5NEi+6fZmT/IarlphdBQfVa+6BvROctZ068Q
/Q64CQahT6SqsyAPv11K18kqvfFqVgc4GIyzaJ5KcKR/5/508e3B+v7HSW/aBSm6f9VrtdMqRrVy
2fZgjfu5P2MN/qkMTDdzkTrIsviqpte2uBxvGpscXO1m3rKWOaQbnrdQ0Pvc0d0YjWQAj3hqZva9
sDFMZIM+MkFEJNTogQKwmrfa33b4MbiIfIAGVR8HFANvJyGh5r6O3eosS42izYzaN2jnN3Y0WkIv
Nc4dATP4+27VJ8jfMZ+UdbLEwHtvsIWplixprOsjgwH01m5AcMjhaP8EvAaRdWs0RnLq7iYdpaRW
4/KvwRGXrbqIcoea/z4Sj9prYJmKwqZLH898b2sVt9Lmg7p8uivUo7tJymePgHu2+5srqIfpeqDd
8NfOvXTMOOwPignr7kdDvdS6N06fIzLWFtAccPFVDDecw2JFWz+WnPxIrSykBMpQNytQ8PgnxXJI
oZmuFZWMJ1W1EYkDMLLIj0kcP3lYr8/0ySJNjsV3fa/jdeZdqFHlwB90bOf2IQFj+NTFG8KEQpEz
9J1Rfd6UF0C7ffurd9F/PUDSj3sUqhYHZWSGlHQNTiytMCGvNRYqPn2INdfkfRtD/lYHKH1a5MXN
eVrwsJx9CGstRKqz4mQdxD/ZSleKUbvVOiXL3P0pm86zzB6UF3aTRyVHFbXzhe0JEOtISbA4IdSf
7soVSKjGXWRSTQppp0f77e2DkmCE8qt7eNU6efwR0O12N6dsTDEN6RO5YuE6MvAnAPQOe4Musq2/
CeYBi1+jsaO488JR45zWmicdf1KzOvVRGMZ8yV6S6kcayL/uQzq+gNypkQA/eX/lq54QoHKwiY8O
a/Z32Q6JzdF+51/h5bxYS8XnxXEGE3aHaTg2NzrliYKodrFC0zK2stCc4dd954ZM9bdNFdMZaaK6
/iApV5UJlRLby4EpV1/QfajLR6S2HNTOXVPgT3MYG/333o6wnV9NFSAoeeLUy6bkwO7qrj59HeqE
yorP9VL+JQ/ViD6FhlO0U/yoETDpEc8dIIg9mMHAVmKfkUogfZcDr9mh7zmWvVd4pjtIHxRsBZW5
iN7b7Jv9LfMYzM6OPIZ3XeMFRA1gw/zne5mHKLFlzvP5/c9NgY/UYjUYVI6OqCpiw7mP3e/xF8Qr
dNxq5GQNj+Rho3A5Q6dT1kd7P+cEUaAviZojRGhQIb/kogGN3aysTs8IQ2zQ2zj/6LtfQJis/T/n
3he7j0PSPG/S4274qgbWjRfQiGrgjZyrS5Rr875lcjB3b0eI7aI9i/JpB/S1TuEws3jJcasmjNLX
TvCNKi7p8lX9FFTiM0m/V/70iKQIBdXpmRb6vXdurAqDZlS0jirMKFeLBi4bU3XIxv4R2X/6aFEO
3P7KoRAmqtdFTVVj1vxZTbtFvhcXHT5yq7P1AG+ZF7trDwZuIo5ekGWsTXW/iem12s0jd0UaWoOU
8qJ/oR+egML/B7AZeZlTSrVB3qQZoXha/mb78+j1i15SRqHLypMmmkNi32S8t17Ic5Yib/kvGgB8
ZrEFGZ6879YoVvAQ1W4KqGXX2UioU3u9UTLHYYBCxxpWaWBLLRZYqS/IsWOZf0yg2k0NbI1Tl9GP
a2iOpu3KKKB4452TmAGygoVHYVPeAYy94tUyhxHCIU3/7ghPyH3v+lGN8EKauDhFPa1W+zb1tU0o
hN4xDvwAKPuV3Lji+DYybtOS3Ps7sfOAsv0vaifyPe2X16GuUHQOr4r1efIeFwGwT+Ot7Cfo/esU
rBj00fkFkHcKScJ1oQ9sTwEoKI6SQ0JG4Sc1kUoWwJ/bQeg0Ih8EDPg0FzReTpyDMwck6G0VzKQr
n3Y2nKfmyxBgRArIPXm3TT7vLm1RDTa+rJW3Qo6vHETTCiymIymrmRTdWCXFTwmYit2O8F3/XOYC
ck4xqcb7+Mdcq8zbl5eWCKndP+UVKyAYFao0UaEKSNGx2PH8eS+UNzvTlMb2q5EIn9Vik1/M0oYn
asWT8bhMtiBDQIZXJ/nuEB66q7w9F7k1f3eM4CubG2WhU78cA8aXc5uk6R215DSVo5PMatmWT90Q
r3qIEJiYN0Qd3RTyWw1SWdYgMAY8mPp7nKM4zI62LZoOoI4/RNdQAAtVHfYqCbdjDpCFDFe4rE/c
Y/KYAzoJHjJu25NtiKHA/UQX6nXE/le9LqYxWcrlXUpLHuzfdVV9fx7FvFjxexFUOBygOc4HoJAD
GyFLEWlyRrBs/2oELOh/wYfYfl+l3JGzcUxTvDKbLmJdKQqCok8v9CFGGvFGWx2656V0JgSXZ//a
P7JzOfw9GB/vdEZnZzasxtmcD5ffw2N7LSniFJgsF1xP80fm9hqk9RaAoR8gWlNS0ulsxDQT1nIh
ZXlOwQqzyoAfWvgfibkijQ75D80zf+ALt/VCs6vlc6EBt2suY+hsa8MkHRdyjTpBo+/P7c1LpKZS
U42ZvgKUwOZxhoRMhdYoB++DvpGK8IJV2pZEhrdYIyIlUD3BsM3AL9zgj3RQvoa1TlnubEF4+bUW
q5YHhNL06q/WKYd9/pGPPotCXhdyxRRiy0JgfQxOgWbcdYNI3NBlJD7AqBqh4WhhMG1h46h8hgxL
kXhUfA30BzkcBSIsOCwOIK6moLa7QOJTsC6D5kriV5bPjye2PWFrF+6aAO3RClvwiQfniZVgIloE
YxX1O5kGaqjxLuP7fgefM8sWQ0DEVZGE3mERu1CIPBOnLQQg4sYby7H97SCnfzpT5BVsW/QGod56
sz56p9JGv9kR4QeLD0XvtxaVrNzQ9ZW0v0nTF9mvgCkSRL63xJuZLjYyIubp7HDbDETjNfa3z4/G
mIGpRP9MSHbPIbJDtpU7eVPwOKeYnRZCH+frNSJRBEV0h9OzmQaUuo/yaTSDowf5QSRi6ZJXqlZ4
lEldkm92JhLbc+31jNjxDTb9Tp1rz+YYagbwxyM8KtzpMw4beiGjX2LfbBsln4V/Er90yFm453VC
yXskbi0q5fJu23kOkSEYUl0OVoLrKqIIwEo9Vz12zYhqUOxeNyhnPfNCi6IwSL/UaSsTY8uk0pNx
ZlA3jKBzsAfHxDVpHChvX9Oc04QpyeM01yqMbExDmLNUwbc606+pPD9jUUzx6Zp5Z36Ue4855AgY
A0L1cN+UCCeWugmeAcAxYLPCmeuYJzdR0L5L4LBHd3xFxqrlEkmyYpgTTN3eCZdLVJ1GA/1KuaJM
nZdgcSJZX1KJF4VkpeJ2wSwVJYUn0Twq6ct0evd8vfdxqgK5bkbVJ0gUmPB2SONv7mdRtoczxZzA
R+NPfqt04PUDNA/9afMmvrm9ISr/jROelrfKpgfCfHTcpwGsYaYJWTYI2akWDKIVEPUVkNROROub
LofafZ20Eh1VJATEeWwvbL1VTWAM2ELB0vOzKAeUVjgVWCsgk0a4qCZsjHgpN8ZECZ1n4WHYP6AV
se1bUsiP3Wanc14WIVSetYqJUODXoXfp2X2GswIoVo3KAfI/7qLtBeYo2NGvuMGnXSmbAtV3pJNM
BdqD6R3Gny7C+LrYSqoHrpeyQOerwai7V5aVwxh6PaQDGd6/pBx8+/ELVtV35F6LrDm0NWS37qUD
ETlyGpqrgrkee+fJ42pGvQsmdvA1l+OzYb1+NTxuM86jYs9dn5wsm3KK+h5yXEgohnCWaXW8eKTx
QzpKT/OtA/pvukF3NmE/OlG+7rLG1OhhnYi/7KhR3fC9J6C0sBi/d55XQEuSjvhH9xMR5OZv0tYr
Ag064g6PYhiGK49W/WlrkicZzsYlyLWLGAX+eBbTcdrdJ3TQxuLaXxJDv2yHd/8xvg5oZ7OnUiYc
TYDS5oBpy6oVmQaDla+TPLaAZqB71LimGgRqeJm9ZlVJe34p3eV0tyORJfk36XJgrKe8ymuxmvaM
/Rh2DPiP0fPsF41MnZHB2Aigs2SRXSChEbnBBDZEgNrBYb+muV4ZRrOGTVOYndwAOFdKizftsdcr
3/ET38cMt2olvTfzgTWU+QTIjuWfq1UQwUfpXUI1PWiXHv5PMfcaEeiliP4z93dLAoLL8kye9SuK
kUzcImCI6VFUSx9Q69QF5p3+fQpuuW68qdNekjjsUbhttD1s21sZ8LAuhLYydmcqWUMNpLzwe7hZ
EHlfq20P8PEqj903sbNWDxx2dExgFaQ0CzyvdVR76F4GGOPUvme8dBUdD+OscJ6DmGZ1EeFmxlQ2
+DCWUQ1Zcn0Rq9SFQInIioLS9qKQbm9wPVkIA16IbYoQiQim1VZeKPvNBbzlJVbb8LczMaHtTqKd
PkBOaNXF5AVhUNcBRRTD1+sI93Zr5ZCiJEB8HsGYiiTlKYbi5wiQX5bl2KuI0iP+fLmZ4Ph/VA36
6+5+Iv1b3V1KfULYe6QJ6KFgRBsj2zpjoqZ1zwo7G1a31pNOgi7ayYCiunq1BacHjzHllFhF03Hd
T3pOR/i35AisBbIlLZsWJdALmEHzV8Kcbh98q4nmv20qU4nL6jFeqZ3P0dTuz+3eJt/QqPimugyn
SCoZuVYQ9yjWG6lhmKP83zMRDVhqS+pArPOPIR9uAr+2tdXB1ywkpepkiG+rD6VTRSyCaFFlF6Sg
r/sSYuokz1girkem6K8EqrCJbYzvy9ymOLarj/B4PmCcwSw44K5yKKXE+DKNUOxy5WTC3E3yMt7U
noi3Yi118kl1fWcUZjooH9j6VUoXtMjlptbzp5kNp5E3R/mYf22z0ZVIJllsmoc1CaeTJA87WTEz
ShdSr5tyXIZPh+rRzLWisR0x42XwjCQGpoQRszRktz5C+k4iNAq9xKKFtJJ+Sq31Aawo0Mxy7zz/
FglhYCGJfWrZWXM+y9s5gy+ufFc66l4sRdbGYmh8Uk+U0vdf2E81kWSNqdJNJro5EfsrYJmPtqOr
7GjycODjKKXOhfkmkGkkqHKZjaV/vHSPNqWjtjeFb/I/TbxB/axOMidSNBk6YUTJUo/NrB6wlIpI
9qxubRQEAoN0n2vmC8klxtzUCf+mALmaian6gZcM7Y08YSICwguuWf/tEMDlJ8POf9jB7iFfsTpi
wwpKJ2+QsZVSbLQYijNQdeNECi2ZGjd8wvs4BxdV9y1ym14vLVVHqTTq13icJ2K9D9u9DbMfrmDU
PXiOnPsrrKuWMLSiVV6BnsThKiqO17VFX23d6mx4QI0o/eYplOMiJ0LCjAUq08UVjrZk9PM0RoAW
OVTqXNeAk31MYcNfx8+KnF4bz4nRJAB58JwFfXo1tP8U50wYnpYQf9H5GZycfIAzuuAXQHXqtYRY
1z+QHo/NAPe+PeNVKX8A75ZVfJ0GsKlg+KE3MMEOwvnZzen6jySC2PFLICpJIFpcEm7qo61qEPkb
juUsdeJ+a2i13sD3kJ30HC758LHGVZUSWErtt/4apLMQlnSxiEUGUtxDWiZG5Q5/1af/KqIgPaa9
wAFIPm+/yarizqFNnbpcdXm3D6411lAvoqAHVAz35WJvgk5yyOWMocbHg9o+4dsnyclDNwp7A4JG
BxMKU08X7CmftnL1ZFIilD7kfL4jFyfSgAomESvnOmTXZMPOghXIcyGfkpPTxPvCtyCP68YiJZNV
+CzhP+2tNeZiE/d5zlXDUWa08rSehnCXxz6WIVWZLj6now9IqYpf8QCAXaQvuSZ7JgLQwWuWq4oo
3LfZM8Cd9UPi8sCIDa3tRELaVLq5DGWLtlAdnjgMtkxEpbg4mSp3TJMib7nHbb4A1cnn0hN1hTUD
AAJ+Ctsu8CGsxNnWoD6skR/B9wGyBogOQu4F8zy5blmnDuc9U9U7b9g/tSFfeoeLlyw0WpOW65Bq
7d9MpecDT2jRyLgnnPFG31fQvtwv/f91Jb3KGC/2KPtPfaxjrHA40JMR8IXGWq4DznBToCRUBiVy
vbnW5d9deERn9HQQUd5msGlN0o2NKFhnWZNhvEMhiBIfakuO9s0Em3XjkVDM/iBT98oXD0CnqZ9S
fZ1Z+EFUGEf13WAMZXzDf2FX8aO+AsIBWCl0XIDJmVx3rJQyxS5GqYA9oFRRX4Anpx4h5tWQGw16
xLmcWmzU/S2RmCqoupJSQWGS2ltccH5KdnAfP8La3JWTzEH3Qpwyeo/phLKDMi3FSUSQBd1J3w2d
HEVCG0t+why5ugDS0U9JToOJorDy5Trpjj3P1gOBFmVXDS8tV5ZkauS46zKESe6CfKogxQspXhRz
zfA9WaDBFlVneT6Uh26e60I1caoykrMsPMUZA3H0XAzVJTjN9UTuFDry+2S8DjAwcM5TADcI1RgI
itk3J6UIku2F2cnPfcJ39AEyICg10UBReF/4D69aWtf4yfdEhYDVofKZgwfxlsRvXQKvlIckBME+
1BCC54uT73LESgVgqHkCfbg9itgZn6EiWRP1FbURhMDwZrmsea1PYEJ6FlKJAJG7IuAFU8QZ+gUb
haWIksN2rRMViuzXEIKHqPHsYOS9B62+N6Kh/SlYGQ2pfnkPzjNPUxmIlvF0zGYTnkN2NQ7yoDQ8
VcXEktn2QTCdmVYgZLP6Uv1B2BK/yWCAc/1ES+kis1wlvNQkgV2isPg8dru5etWGqAoOGxW6FZnV
b/eNpkbbWJqRe39+/QdUD9m0wBjdzzwiVUY5vKb/HslORFDbM/JyCi3v0PNpy+0+Um1UbUGRSyt3
BbRUlC7eB9PwQbaLx5XHcVd4NusILX9TKZ/Ce1fddYYvnCGdFi5d4awgyc1fwsmHlfDhWlgjZii2
CNbiX+xvVh5koo/MIUMI+H8aaiEKF27GcsBiQmNd1E9o76/0muluGRHIfOjGj2cfXWPc3F2xZpNM
1F0c5D6abjrbeAox7k1+q9qdLHa0Y+v6JPtAnCDSYdWT1pP0yzXgd7KbpdWZQIZuH3+6UGCap3HS
e6hoWsXA3YvN1cXCvbOIS9FYpQ6P8dKzLeO5BwokdsMvVy9s4DW8w1Yvg1bSM6EwkuBvPxlnMBF8
AVC2PIlJTq59HTM5jWsqd7l14kfMnNuxZghPDXliWtUOFtVBcPCNibXjl37WQ+weV2Kz+Bl7+b7G
crl3gIIN+VnUhZaO1IF+FJ+ikp5i8oEOAtQADgV3Oui3bNI8AcK6Xs6G4rI5MKJflEgdngqX1Z+r
iXV3aqn7lcciyrSFjV4RYPo8IY22+D2kH77Z0ygLitUvmsL5LYmvSNCityug3AzqUEuz3/qAq3gK
mBSs0i9MhcNk6P3IFMtwGTjSq6ixFRKdp90baX8qaP0s2PdFReVMvgh6ScuSP4SKbOmIqONjJ0wb
grWHVdpl9fEtemu+BJpgvR4XyBZx9XyXV6RZeFaTeWiQnyncUeXgb9Os3yTtELclvlWWMM7dfWAc
52aAudvNHUShtFGn0zk3hopnts2v5I2RETjWFctLT1k5uEWkD8BLl0w062Fp668pW6j3fqd++vdN
dnAL3dYRGkvvSeB3VBB6qb1pu1HWZQUBGXKZrMAndZwKuivWXct12NdfaazXGe6AhbWrwiDVNhQd
x9yzZDpJWYW1SXdvFlbQtXhS5xjhSx/FAL9321FEzRWTLtUSjVqJx0WrcsNSWcJp+iHsMf3+y2oW
JM2fA0pKXfSbvq6Xxjnam124Yx+0c7LOFKDaswcuxmaxMp3on/IiPTvZWCxyA+vIVheL/PoCabBG
v5yhpHaPEh0PFufYNDmwPnz5Q2h0tim83W34a5+WNPLLXyK6IxYpz8j5KCRwRWZOnQR3fuxZ3d7A
8UP50hQ6q47QYQqtF899IHgMbvJ0qqnac8R/NahImuF20aO1q+yVRHV3F2Zn4CLiHUhDsATn9+uq
25RO6+6Z5jVGVDqhqYlZxk+sYdRp1qv9zitRyIsNDNlKoNvr9Nd53kv1ZUzlSFjKohZwEdjWOL+O
kGifQLSzaAkbf2QKn826rytazjKl+EdMq4TKxZpD6HYUlDsRmWRrOhyyzD6N7bsiCxeZNb8UMFEt
ud+/ozXjhurLNOe2q2Ffd0dxLXYOrTZHkPHaVn1o+GudSfuvmzHyI1Gehnm0zZXlOzUU9elhX1Er
oy0cMrjdPNjQHnLQubgXbrUJF6JAXwAw3QM9SRSuszu9VsRtyuMNC53IGKVORZLXvh5Q8QIzLoQj
BTcqSg9D9mQ0aECEK9pXplkv5lB1DgCptCJklhoM1gSQRPR/01eMUFX2mUg+KWpYmwUWT3XrRfu1
zJMdG1E7LzhKjzLsBRwC6JgxWv1qlJdjXqCP5zssJK51RmtQADZW7IR5CWKTvym7Cl4+tp54fwux
EvgmpqCJV8/dXsLNuKu4pTvj1oJnXcXMSGaW3f5UEiqsLHPf3rq/JkkxC1iM/iRWc0o+BtQpqah8
/lEAQfITIxXRMcCAGGR4jWFfOZW6YVyxPvPtFaubozbk97dgqVaLE3J7ZUfUm4g3ujTZJJFglhqp
YE/exons2pNB9K2/h2uSOIKmbD0NWskVrnB9R6nFtZ8+GYgXgF/Zvw03j1WYwnxjlWDoqYqqWBwn
Ua2SWDfbJQ7lCId4c8TsdtpZ7VApijH34U32LyruRC58Ly2uzlVqbmlVegrVl0ecBHsgrCuEP2GK
Yo3h7VZfJ0G5E2yB85fPcZGPXg73MMGpD8QRhDa1TD4e1mVoA+k91H+LEJng55P5oAXxkD/N6CPu
MFGLj25rg4Y6BFkhBxVvWod2nVNhDQem5sNHEXutBICsREwbK4HBW08dp2YFLFGRfZ0eKiLpjj3E
zu12nueVdxZjEyIlIpFbLYSSW/91qhM1VMJAepAUnac3ygcE8dyOb9TTaLvXBBVGc4WsFw43uFLa
t0cp4jbWdEJXnqezsvhqNg95Hr+luoM+g0A3Kkujwom8KEZGnKE0+UTpTF/82TIfUd51EYwogwP4
Q6scwWJqG+Vm+yCK/vFpCrPvIlnIMeCe9v5V0JQQ01ubqkrGgTkr1doEK01mf29cgpmAtTdfYth6
HRditQNzpZSRZCUGpQwEhzkx3qR90Pn3fZX1OxpH0jiyk5tDIQWth6W00sPRoTGC7G85PLwS+ZjZ
ksf3fosMfEiovOTWst0KemkG2vdjvQnX4GUJnqVPK/mKp2Dc2iD1mHhOMDriM9hd9VXfv/ghifMc
h6hZ3B0M71hQMGSbA3aM2R73sObistTRE38duaA76aY4hPsYjLPOR6uQq6R26v32TVmRJ8/JnYYe
lGe6xAwJB0Hh7iwoYZng1poU3PTfCfRClmpmeHaVZK/n6eFXx9gF6w3t4u3aUwI7tF5DiaWZYhoA
A8q3xtHKq0XKeQ+ZrW5u93kN5K//6RS3G8luuGe0No/RLVq2kxqlOQYCyCStOebzSXZrmdp9RzlB
xGf58vFAasWI0Ki6o7AXTKiKD/+g+T/+rffcRGg9INwZu+KZ6b0W+HZDCVn5mHFdjNwZtX28Wp3g
Kz69E8QeoasBpz0AakO6WTxRAWV/67PODofkBMSieNQGdRzDdOirc72rVC3wBjHoTZ6UNykq2V3Z
ScttK5LeeoxA1s9RYsVVBMM8qBNEqzAbztfFfza/OF+n2vnaHGyWmlDN2ZFS8pkVGgX2W590ZO64
zLZlPGPPFc4hR+LKr1vPgZlxTXHEVez4AxE8bvZJBpGFaXSIUM7hohP9gVY2aOX7z0sgi5O4EaRx
UO2W38NEUJ3My/Xkrq1tsKysCgSn9Y2mrDBKLPQ4oi44WboV7h6u8uV8whLCoETOQSQ06J7Npt2a
7BWc8pG3sx2mvKC11Q2RDgQuJadmq/FTdQsqt/PRX7usIdu6qWxQYqnhmQyUwKAXlNuDPMDBp/7A
X+22WB6ZU9bePfVa3poa7FMfZv17UU/fXCXlc3WAQK2Q292b+If3Z/aSW/fVOTdFjPkWkWQBrdPQ
VOH566wxuXTiRpC4pB73M1t2hodumxq2AfuLZ8PDLNZBhrbVG6OH9cqUAinCu4kDMGf5kH3q/z2V
jcwKRudFsxlqqTyfLWKGul1kdqjZPsurfuyB4j0pERUfW33A0WzwLBPGBsB9qCXury16IlWzwlpo
PdeRYqz4H2CIEYP/xJGT78MHkeFgrOic8oY2GN8vmH8MINasmnWrg5L8kJuwu1SPXOBeVhit3weR
fEPgrGB5aFfg5gcbcwS+ECggU5y0Hi8i27321ZZIZK8ceyL87cN+TarjzARTTigKtgtbqt/TI+ux
puru0wfqCoGKUKjmM1W/a3w02AlVi4woRVDmQ8dSa5Gvcyh3Ier4cPapzkB8CDScapM+zF67aaJP
UxUFEP+rjUg6xBYwcVDESlc1JPd4xpzdyBwJuDDWxNeHTnNBQAMwBDuGiwIJ6UVJFTCd7x1I54VM
b9HLmpHKPeXVPzMOFfDbckxCqA29W1pYLuhff6JpSksf5pheJbCA5aKXGm43PLtjj8CrEjSZrTI3
A2i1Kxm4BfpzRHi15wGLMcHC4iB/XXg+QnoL8GLipc63jgGhoQs9sXeURzTMbf5c9xYzih+Y5BTg
vDsrq2Vr17K+I/otQmLdb7WlUt2av4fGd80UQ+5eABpdSuuXZdhzaqrPxxq7nFirVFGFBbfAXqrR
TfW7iimBUHLe3AhAVsVhyOuPe3dpGH0eGs3qBt1yIXArdesZ+jvOYNOWYORxG8fxMtV76+9iOsFj
2Gjjr1+eMf3x1HIxYDBrotrpkPz9ND6a/aSOu7B9NJnVMLzA9FihR4SYZ3fdPthcFemwG0N2a9A0
XCsVzBCbXtPNKTyfM2LaXnHqDekzuUm+Y0sRN9S2J8/hd+ez+BIIXzqOglL0I2UApmBlG3De+6RH
pHKQmq0efW78n8TCB67CpC/dj1lvf5QpbkwtD+rlrCqoWPAnTBHYJFAC/lMIxqcFyiySOPDiN4JG
LADEQCMDsX1idAxjm9DQ564Z/jQnZBJpUXPOXACr9zydiLBf02QtpeZISn5N7HYkAT7ox+aHfl3n
z9hMK1HC7BpqG0RtPQVIvFAvM4QgRCJyDx986cZ+cs+hFY4Vmr5Jny+LXjPXkLEtT7Ch619v1egH
tOJHeZnjfg8o/NwD/+lkk6WHaTmA+nyXcaBWlLAeV+kQ0YRPi06/Fqfk+9cn5p0yv6QwmLLrEIdD
LJFAXCRSW4nsvys6I/wEBI8BnZqLgPB3HhwmMwu7m/69swqMw8UOP4iWSn3+LeN8hCre+olAhYJC
WDNEn+BjpuRKrB/Mwygw/AxQfpeDqFCvo6Klm8TwH44KUyF/lwrvTSBCdfKXXdaK92mjbqPceqWs
GBMN2wgRQ+UelPqOGFyW5YURCPiJjA7vkBb4K/lUxJRjOGdsP9qEdFHU3jFzh4jYfCet/b+yGAVh
3yhilrfrHNgF3vZz8LWFHMYSNePSukH5La2HyH1hqMWLb2ijBbESjzM1tPQwVbbUYFgpn7xRnocy
UsfiEq3cZIPSxucm38ZvEDYPym/ipNIo5QUl6WSzfQjwYOAN/jIJRRBUYV1RnkF5O/wl+QiU4tD3
mXcevTR0KAI7gN9eYi0SidS9jN7mkmUkoH2g+WW9YIhCJnjVKZSO71r+tmBfFDeFd90IegZY0ILh
mWOsRZl4EyiFDKW/54+B97ncSDydNc7LFlhGpSF9SwGhty8WV2XlYWDo5wFGaQgM1qOqdmBN+TM0
+Cz1pFKhhUSN/YZ58AXQi4STzuNLDsaUWxoHR93gHOoePta61ERdFUKXp8PkbyIKwRYfvofDLLZu
oCGk8DNO7QZjsqvJA228zIu5CoktrxJeWVWiDFjUHELLaQS7ehz/NCN5ntwZ3TOSZxuupuA/R8gW
ujgpLYk9+H50609WH2BpDeUoD8fWSMiwSlrUN6oou4XYpEw+x0yhcuWlrKKYu66e5eBj0Sr91a+z
LMX+LqwfgGKAD5G0396EgKrFeSC/onf5Zphw5FNocLTalgjO05zA3S1ShST1lmsNDKcHEUcDR2a+
FH4S2EZGTO41xUfpxPaFKXAGqpWTw5I+D5R8iszXxDWNdDNOuH6IWbWTCvD7z3XLFlHsC4wl99Iv
aeXWgk7xJniJV1qcbynz4jT0VZHdxMO5g/pUABY9sNU+SIlYEkp5ozQjrte8+rrxHNqDgZ2p/2/a
HDOcjsxYgxctt103UsVvnLwF0XNtLoKFznub/DAGcL2QhyaMLe8Uq677oHsro72quUL6PVH93xnw
XDLNQ6RnLaLbov/elQm74a8oy/COmkxrINjtsRuv0WUDt/OieQLLJGm9jdj8+Abwza4EVcXceRPw
fVraqISKQxov+SLUx2pb1Cc1S2vflN0SqtagUMUASxDhVI+2BGf1vNoEtjxhRPvOxlG7rEKbq135
9vpouTvNgabiNYZL7f9sZufeO3aDhS5CKlto6KR3ZClmsWwl+rWmoHMLM08ZszBb2eRY0z6coaz4
8cTGDnbrvlrc9GIfclvz+hLZ44FloefEX/sKZkG/bewI+P5wf366VgpVELq03S+0DKR56YNIiLnW
Nw/f/VVbklLm2twqxMnkGitP0fas/YK3Ufj/OCvGbJ1VJp1P/jrs3TXUPHOx88bUHm6gZ9khQhcS
O7BwdPdHs2/JIpzld/iEFVHlXkRTKsc4YU6VbXeLhpYQdIzW+aPH31PWnbO/8O+IcxQ07raH799/
EhM2HPlYw5E8Ga/4kR7cPSUjqFVMJ/R2/1OXA7iXn4/+vXXbRnPopCmcUwcgaauR612spWyAOgYN
uKehtW0qDZpbEBlxwTcVdBOJol6BNrS3bVSoqUgQG19Nhy8bvUAp9wDo6bpO70/YBx/Fi5bBNiX5
f9Ld/SYXjODnR839SWSMxaGmZtvWdUi2a2Mn9fSYlE7v0b6WK7iDCL2UJ83qUJgkIZr0QBs/6Ly0
Hw/vyjgOc9oFy/8mrz7gfpHEwYwbvC7ZTR2pY68HMoSIdDM+EvGZFSHR5i7C+ZKidz3eK4VntcnZ
H+SsWsbXWl/4UxopXEhrqHEK1FnJ14/Lxk0ySXSL+c59HpZRqOJXHuK5qeQ7Z79qG/Lm0QqqLzJS
F6vZ6k1cjU18eXJQPViOi1Kc3JDg7jeUJDxCwaHVIkKyKymL1VUwuY3vZHDy9cBnGW2lX4mgNk1P
iYW4D1aE0ziS8CQ7+dfz4TuClFTRckPXkYQ0sDoVh9qrdnyFdgLee4UXcajpNbyksOw/HEqgnNN/
6/1mhPiXm1pLVbV7jM4kWveV7crcNBCWnM7qgzcbmuYIyDdamkX2NNWyV7TAAI5NXqIcEUR23/MT
t8EvBLC7ldKlUUpqpn8KYIpnlO0eV8fwaiAa5I+1Kjxq/wjF6oXuaR9c6kWaut/TaCh6EDRIplyV
f7mCSfrfEimdXUGViLb5fjBSi5yQzsoSqZHj3WXjGsQmQVZBahROhYLbd5EDkDFupW4wFmqkpt4Q
6vpvcFGb1J7ULfFiaXJQx69fpYrtSVyCijcNUlVxM9/3WV8J8ytokQ6TkYgVreakM8xBlb/exync
cA6+Ud0MRvFGraOIx1PRUi7n1pPCOKNsODuuT/nEoHZbykD3kmKM32jk+R9VP3UeEFUUFkNb9JvT
VEAfQH7CpBRAX7vQZl1nVvGBjieH175RwQVvf3T3EClCymfHzvnRjzx2MHw4hDhDty0XfFotEQ16
7uz955PSXjAvba5Bwu3mG0Cg73Iogh2S7ya1IIBLRisBieSd9j7dfkUyMPt00K+CQRdt9YhKxWEU
MKcCgLNLUfeFnIruECsB4+YaWlna7mJbAXrD/RjBGc2N+R6yH4FVk2OGxp1UApUbneSLQ2ViMEdt
Gt6SSy/LJegri1gFPrsOHwMO6KeFk0ndMUco7S5JQQ3J2kzPCoJL9uNO0MerAGnJF5Vwu3LWAgcj
plinAV4J/Xp0RE2aehNh2qAFG7Y0ah8ccxHtl2LGgLEeRD/F/2G8LIcx3vnwmRxs/UCbKn3epRbb
WGCSX1TbiD0ibubm4kJebFTqtIi4ax1dSXpED70mg4XhBLWYkHYIOF/+pMigEGJP/XJ4FMxHODb/
LPn63Go0B8NExj0NF3SI8kdiTi2Bb4+FLzQz7MMIjfC2BljdhS8XObxoY5m3vyS7M9W/cjGz/gaX
+eHbmbBlZw9WNMLaihgx30Kg3LKrLg5JMHR8GJwqYu4/YMdchLjUK+6jFQqF5V+C7Ez69t6titD5
DGvsnUO7rjGK1bE6nG9admDZqAYi4wnzfc/fhmkHda7evYvUisTTySHduOlOgVRK8woXv51LE2xE
1sDhWKd90qF3rksokttX764/3A2KkIovH5moRFUN/Yu50xAPORDKfXKCXAcor5zTQ1GvNK5FliMZ
4Gpe0rH5I7G7hM/+M2NS9JaCLuXn4Wz7elDEdXgxzpNX6PlDDgLEz/Pno9tT8wFEJ3qOWmSrZw+L
h6qS4WnG1eyccpwwnZMhaqz2U6RBxqhhGejQuy9QHjd0uBiLnEozx9V8rIUpHkA5FHmlbaEXOeo8
hHn4BI92LYsUdd6tcbwhDcBLZd6mXnIH2Kj2bGFh5I1pyHAs8BzwKST9WMHtI+2KKAnZCZdCfgvY
X5nXeLLDxW1LDNH+gKDWkZBw2ltETrpq7JApt63X8Sq18LayaaQdu7UF0B6vDn5unyE0urAauW9u
VZ8477moRddd+agJP2G9MR7kQ8tla4wNQEhxLxJ3OWZt4lhagul+b6lVMZFhGVEwFus/L25tvXTk
p3OiIp+bt47AYLwA4rpmzK4FaQPxHZC+GAMTV27om3liqYjzB6SCcohtxSOsb/ABGBjiH6FsyxTN
NRNXy6cz09BQIuvMUJzrR1W/QoPm58KcwNeYWgPs64CKF7oaEcgXCD0Tw2QFBOrPtC6Xh9qW8Hha
E21Ex8JV8C10hmrCnd8bQRgXFgXNUVmeTrJWut2iK6+MZxYA8sVffs15Vv6eQcFp3ZfL4s4BKujJ
auRXaymSi41Vjm56PrEuT6gSqNJOxV6eIOwgoSuFUq0zkzN4dY1fblHW8VZEeYKWBeJ4XQ8mmZ+d
dxBLM9EexvIPpN1248r2ICsj1Z7Jq6WnTNrGLu3Y74ErkRopau/wAoXF2ImDWQrJHqyFnYwxdTDB
KRN8arFaJF9BVj1KBi5Ojdj7Ne0iAmytFJbhUN55iyptJoS0WD/sCcygik5n/IrvtejiMSbLWNoX
SbxMT6K0gNGqyJG0nw+6P1tOF4iy9y9blf01xpymeJD1Ib684aRUwI5iNJY5YCIuVWivImbHhWYK
BF8DV9GRWKLan7zA9AD1R8huxE5zY6veXWgjH0P1GRgw3WK1EmEhE9P7InVrSML86Ejiim7TTe5H
SiVJD4gDlgJG9Wzmubla2hn7Iue9JrKL/iaDuqeoxF96AOGdIC9KAiyP0PC/7oa/W4pINGBzYtxu
ifUqE9hCT2Mhv6VfI7MAZLrLeZbdYVUl54FrWsVa3wzr4j6L5sx8iilBFRpBSiXleidN/sCuyIQG
q/E5ExE/CbmYLKZrDD4SAP87tSG0C6Hvanl6tRHJgrUbpz47z7KmPPMvSoR6YMXWM+Dd8s2iQOE8
kUQFU4Td2ostGLh2fhY+Wgz6sdSWWgi0wWQEFlXVTbE6g5Mf00VnMlsMk815KoVURAM7MFveqPV8
vJM+At/njIcSCCA4Sr0yMRIzSwzKB6MhcqFkqcv5S6PiWm1YPXB863+524GSW5zzis+kIIaMUyVD
jy/4jLygqbieWH9zFCepacAUhmerfCLoWVYTHMzo8/faCBJNTQ+RdtUOZ34MPb9JzDfmkuFwj7zB
giGpAUG4oVK9cSsWuECK4Lw7d4xNHf0WOjOKZBurNHaFbq+HELvrHSqXzr6qQbfn+C14oTjioPuq
HpbYJRwUnPx0IPg6d7QmlzZv7DyK5F7Occ3zCUMF/jpTTnIXJasYnm9oEFErMDUmoqwLIdj18dvg
PnSuZNiY/OnafaZYpIr1HnSH6uO2O3I+YEuZJmG4zWMRyNpxPabRLey+P7jtBKlPHMO0MleypMyQ
zjucmotb20k3+TXIiJXv6IoLrSchna6JhOtih7MOdD181heDEtbPit8+UEgrblXzg9kovlir8alp
GIw3ThUY9JqQecblNNAZlUyedGVam6j0jKEinXP8DH62g5X8HxXGWuNSdiv4x66FjHKgdljO37ct
reVr71OCaUt89FfiRN7OfJwFbVUfILfE0lEaGl9ZGo//O/3A3eJg2ZvHAr3l9kB0Ra/ICOSmu8/v
C+ALf9kH1u5trN6H+N8JzaFG7ofA+bTrdE/sjb4eQZXaENakmlNpnkg7HI2Ee3u+mSgB+ad585yR
FYIPf+4LtDCC9wjLPA3snmwuUzH/rvTw1s/IVFt6HpXOVW+Vo6C7GPadzdOVoQ3s1sPCW6E2bYFl
sle7jYRKmM+xNZ09oymQqSaleTWyAKmIg3TerfoPQgJi+AAz4TvqnExbSmK2FxUFW3DNLkzC23g/
Y+DfZR40p1i/B7fhxnU6BD6Lxma7HstHC4juYNHoiWHfSEtKZqL+x/1FJDn0rZU4JnI79jOniWpj
gridm4Z4D02NI7h2IaRN+sBMR1eFQozAax8Hwr91EzWRbI5zX9jwj759o6isikSp3+D28IsiDYgY
IHromyouCMPtrrxTbMV1fRwMXHpmODdC5yhxz8Q85Vyfri5/MJ6nhBHJqqI20iiJqILRjGo/OsQG
Xc27NYQUQbWSqK29jQw4nXEFVWWTXi2MjBqcCaYqIbxPUX1ebyd0jsMLOpZoS4cTFt/RkF1tX3Ve
HcinrWXJdCuwlZ9B2GzQ2zeHPR/azefmGoa6FnT47ImlZr7abRMi9znBw/hlvDlfXJrZv9RSz3Ud
bKHsIUozkWeCvi6RBlq9C+ogb6R1SoJfIssaqBqD2kYPQiHkR/o9SM7Mwq/JpckerN1XnwVuw9gr
0VZHS5J4OOatEyQGBDUC71e8nJToI9zwOMN9amh249dgA+4/5tuNaohV8/vX/XGMEechQ+q9GQMU
ztzqTR3ssBmPYvACJIrG/ClDYSeSBWioKIi0q5T4BymG9Dp9VFaaA4DMAZOiUy4d2o9yD/oYtP/s
eEKIRcb6c8D85tbttx2RsiHXIYS+xeJS2pbm/shs4PMAIxOUXKj8KNMoobrGd+C6PQbkr3ZDLUlv
LXuRMdMT1cKnaaGsKIHT7zk6sjr4880/TNa0vAmMBMZUEUOevGiM4EPxN4YyGwNvfkKXRdiHts+O
MaL2AarF89Ob7GxG3As7IZ8b88/hU+/Cr+3MsupowEepylF54tzicTGT+0xTIva1NLR1OLIW2Ec0
1b/caQEBkSmmICacpT7Zzjoqsxwo9cgcfBIWChM0vtg3C9k7akaYEzEfOg6vbHFk2sFKoohKzeJH
u6F8Mgq0bnUG6CCkLC2xvSeAEekOg9TIys7m5+GtI1jIUySrCUhzdYi/0YHgDEPOqG6RcJy0iTeP
Kunhyx/dVpAcfmYMQvpx/NA6ND+RIwsyexcjEOr+jAPmBdaW+f7vmEc1KAysmgSCwoB8+ZG7mIEb
PcGZBr7JMpuGImJQpGPlfypF0xfWXLFiKCbOtKjU5XRYWYctkn+DyJcmM0c3LdW34YHwA5RZrj8P
xJHVsi3gh/jNNOnrmxtabZ2CgQgt8O/zzVWTjzCtKQfqSjoH/QTzhtAKogccAGg8an2+X67ZVb1K
kHwhx8nzCihDJdZO7herGvdmOEJUDzSQT+NUiP9dCpttJ8R0JHTS4i/kwcttpx4VQ7FUvOErGdEh
N+jDB39jcpnWlJnE/SSbjedMXfvhXzise8bKFRPbZeHfh14wq5W6JmDS2/UInRyuNSe9knCNvei8
JWF+I9nuGLkWrzW4KipZghqyyi9edZNqfnk8XfLtQs7fcRWLYREPdNTBof8bsLredtqcm/kZUUZI
N+2G6ZrFJLGXd2HSYUirCGNW1TSjv9FboJkWzAqeDzhr/xHktsm/wtjEainwhOkCdiyruq8hrSc8
mzyzjrveLgd6LnwVMRZGyaUbyiXzEGh3k9L7ISO9cv/2AaDv3/0rhWRr0cvNivtHe2mdkvhjiA4g
Srtk82iCAVjB9UHq4hxCjeind3XHeJd+hhqUavCICjGgQd6laxpOi5IG8nJKIDLpvUaaXrVEqyK/
n8CcTsHUWCMLvyiO4qGrXQP6Z8mNJiDXtPVR3klnQeykzV/7Gkjx5VRPYTUJrDRZ2qndX+6cdAkI
kCQi5+D4FvQFT/z9GEzQp2fvQhHM+9KrZH8t3oyTw7oXGiLMGagCsk72YjoYOuNirfBoUi76Y0ql
ytQdqletYGRZ7T2tIAHnM9xoXkpwUwOKmzBLDDSNjDmBN+mTpT5UAxt7KJxpLDRJkrnlGSJRHN9w
EW6Coq+62ZafM62xjVKMMT/xjyE5hCRUaQHdfDb8Kbx5D6CHvB7F1yXYMZeJI/B4ZPoFU++vQcpC
CcOti1UbU0a11F5c4JO4neJ/Dg9vf0JaCLgxKXhx5z2W1bTHb1ITCkklEjmsHD3wkdhOcE/OiQT+
iHJmjK3RMW7yUztXW/BcSenVxzUriiW5EVeQlc7hC+b3jTjN76WDNQjY775L+j38Mtlk3bml2acF
2u84J1KBqGYbrrOyfMMSWu4Uv/uIrXguMIWwXbMPIU+A6pt74qeUabDeZT242r0Kp4sLpBHxUALD
C58q2RCOhR/f5+pVjizOLRWC7KpIlX+8xUmPr5LTlPq/L4NywueD7a+1dfLOIZ01E4NI7521s3p7
aj2+gNWXFs5gGBBCwS5YVt3FM5p0dku9xcUrgtqm2OesWjVMXpEgxtXvsC6L6bzFUhTxmdBQOT0Y
RKkv2ARrr0BqpbfHDTIGmE72Hhum4UE6No9RPlCUgbYL1sq5aH69Tj9KYjexYu21g3cS54CbmQlO
yfnP+qeg9Owph1dSDIgOTbAyIKZjlSeznL5Gnc4F/ZSfQkbkWdvtjUCPhgizO9jvjGekk13fZPNK
7aiZm0Zw6R52Q/2/bp4Ps9clfH99aOXc9mKIN4+hn/+W0cSnEv1R1enNTI4nbSgW/MtCMus/3qmJ
NDAfY1qZF6e5sJorf7nDdrm93y+nnmX5xa00ANYcTtbaiWXxmPXuJWxIaNGqqk7Z+USm6mJFLzpR
vPSEq7nNkmVd//WL3/6RzyG8KODNtpw+wO7UX+34c5b2pZ/H0r0kYclvFiqARhugQxd/ZYF9euMP
8LMB8yGYH4bIGRMtO7qFvqhZ2xj5c2CGMYE/uMlApUMXIyqDXkoCdKYTJSAnB4c/TvSxgRmVOML8
sO0ifwBDbjGz7JF3pBArPw3HNs4X1iQCUqiCEis1hADEEwzp8/+m+845NMylzc2dj18BqgQSNCul
kW3nE/uDZ5UsSW6aG/8wt46lzP4QTnnDKrE0L4YFtdHLpixJOoLV2gxxQ4tfgYm8VDi/nCzFJ2IC
4WbHSg1x2fnjhukC87UupTg1NZHhBdOm0DJrbB9+1TC+IUfZVmX6Sj255QI54MIxRahZnNm3vBz9
RowhPzlQw+2KL5cGMjD3JWUKM+nQEHk8wmUnBFFGuqjBv1UDco7jn8HtuGWBU6p+ZP9Zwe+HOs07
4NEEvJ4KRWkesXurKtv1y3G22zGZlofyybfSGnIdFOeMziePFy3pV+8PhegkPMmv3K7/jgLECu/e
4YjHOq8JmfJnJNV1emTDZHMDOnXel/HLaH7SxbLrDxQLBLbvxRQ6IukVshTIm3LEa0vw2hv7yMQV
6ca7ARUlQpTKC4o0vNsJNAGdVUlcsc//24M78wfS/xg5UsL2PZDD6eBcRJC4YnLYipcvWQotI8VK
p1Ca1DFWQHFzyb1Xa6EiCm4nsbZgVyW5vlyE9o6GguugLdJ7qh6S6YzuLUAofQAtDlnnzwyo8za2
iAg1JlWguAqqDHtrHk6JK1edN611GP7BXbmxUC2jubtrWUcBFmrLJX02A/SDiBHmYq+uNwbTR3HR
Jib4l03euL3s0SjajyXdxElLi9JuS0PFy7kXH4bHSLdoCxDjsQpQVcD+xNjE9SAOk/xkc4nVzSjk
nZAks+bTZI9lkn5CvF/FWMgtNtoBF8QKDPUWmTh+ZBmwfrzHH45ISeeidCKBXIgrJzul0yEF6h3+
7bpKN5nv94lPGYU93YmiBR+eh9t4CXPqm1o//O0HNOrtLrEfUnCw9yqFiQGQuMqvvzqcwknjCE1B
IHYXCSzmMgWeDUH9aj0Gr+2dQoUdN7CD/yat/dSIQnf/skG8HNgmSTl5NGf73Egqdkx+0SEZ+wR1
lyfsgskmBLdCetvI8kon3dMOBZ3bF/tTs+H0SLty9r+zNg18jzr7lVAkMpE1ILtB6US8GsFJ/Isr
s+TpgwGobDniCfyoVMctn12QnONjpvDLh++LRtoCEc2UT01uDI2rj+YmSrFWgyk2ktaWEjZ7dKEJ
tUwXtJLjJ95Ktjwgpins8xMWwv3eURqgdsv2RVicdshxe/4z40Z7I0qOmUQVDlQyMAisZYoJxBz/
y6LyDyr1vF0fH6J3UAVaUSXJ8TYImcydsCIWnkdc8bgBpLrixoaxXNwVHs1JQWAoea1GZ4JKCzP7
tIcDnhBZVfi5eU0IHx8DJJSb/5FuRGn9b6TDCbdAdqNuusyXIxwWBxx/ZA8/Ya5vGjjvciWkEx7z
gl6eocQ0mz7K+6mMHRlqxUZWBW0SveOREf0ncreTBpYejSzPEDP4LUPqiQSZi978yQLOozsWwel4
HiVzJZLpLufb3qCGrpYa0B1CcqrUeajLPochDRabUlu1FOsyI3HHGrYnD4k8K0s5iAuWcDBKEvgt
QFMct+gdvZ3KfBJhdlVB2JsueZmw8tf49RB3vE42bmFdNHijUsg/HnlkqB3RD+NDMOF593YGpEc1
dssPHaJs29rGiksJmEhwgPOG457dwR7qgzNC7r3eV2piJZSfPR34+RirpP26E1Igph17V/z8t/Jm
9xxCf0brCphX9kaPOBJgZ/ofBNOmKpEU7Kceka3tGhHZJeA5fgN0305/o6o6QeET/pYFJoO9IOgI
gaoIZrj+Q+yxAhxWeZSAxibouZgNxXdNhKd7k4FmMexNbTExNv1ylKc5vGP9Hr1OrkJWZ349bP6k
MSZtP0nlFxNIEeowgHnIpmTVyjMe2xTqjMCjQ4en6H4SLr7i6dyfoIv1/1QeEDKDNXXIiGKofFzy
Zsv5cpHxorFHo1hV5m2q3kfszB/6JmGXLfTweKiCWSW++zLGZaBytulU9DVEOuYRcY6t1FoF+8Cp
q86h4T5M0OERxtbZVPCmRQ8gqngFvlQbKcfEv3HzDwujh1lSd5gBF2GIA5MbnAwr09FZU08Dsm4Z
d+3b9BuvzQvi65DEPCPgKr+G6fpiTfJSMMToik8kDPej/jAS7PhfYQEAMrDsUvIfSj3/82Lrgd5A
sMz4T5M6vrRDKfhP+r36BLeDqWfHwvYJgfOo83dCvn16ZuCdDwOoT6ubuPA7i5JYXvsfWlLkyMQz
JDMkt+dPh9VNbR2Tg2aZrlk3kVs7ogQUDGsDCzcmj35K2Go2YhWyFL1tu8z8lO+zqXtWttqCnKsg
akvN1bDxpCu7BAVcu+yoIp4o5AXjZu0nNxAj9mLYGs9DICYlzFbv4f7duRwr1Qk+MDgK+279fQvR
+AbU71KjMS872g65ITKZcgj1XzLPvRrCI1uOdAXuYn/TuC2sWItwJG0asc7qdXiEJYgL6t6rPXJK
dWbt5aAPA/Lbs97u9lwasaHseP1+6DsjjQDobwvDVUhnOQmUr6xsH61oxe39NFkTYjnuNR8JaRVO
MOsb/6Ay+QBBXk7Znc2zjiCWh8OiOA2NbEtnssgDnjv1H5qXAR+nCtS2KyrpiY/3htmY1Otup6OY
iuJgacVsF2E52gwaetjQD0aIToZIT83kS9abSgkKFy4AWo4MRcdVH1/FLvVnbdYP5l5Amxvgno9B
zVYDrk/Y2S7n1WL+bvJmXY/5E9FkvYsjPfX1cpv/9qfFbqhfoNEXmBjGJS+y8atMvwUQLsop4dgB
7pbErvb1UCcybCxx0/ciz5RXJZzFJaO1x/8N2RIB/hNiE6+qX3Dt02SS3gAuylVzLOoj9XvmxUsA
gnL1msKeI0uJ560RzDEVb7lGmEU8ljklgJumQFXIrzR1RYSl8bMJuQBr1ZQGUrydwN26dk5zkcNL
J7FtYt1YBAMEYVL4xyoBs5GLQcmYtXo68V6rUbOUBmXHTePd9/nlbgRWYLRhszzev3QUokMQC8kl
6GYplmpb61d018hO8nfjb2UsS2RCn2oaRKW218OqhydSw1HV4YyP6E2LiPhwrVaUqDkvuX8IyHq3
XaFTybwVNaAVf4xbtogsxjl4MjOi3wGyipbXIMsRyB1MozvWAzSkS5RpiF7m7K3TldkAcywEiFf8
kE81N91ayx6iRjZnB+icAj9A7cpVeMU5KFMO48DMYHcXc8KZzHsFT+EpMYdGl3efIgvqMJ3gaTKh
nlbQ9euCvp9d8E/sYVDAnVtdGZ3HnQuf9zPbhc/3pnUULhgFMar56xI4jRQv7+md7EIEvysPBBBm
YHEKKe6REHZIqADNtW5UtWfW8cQFUiolRW507ks0R5LCGYa5PqFPhrn6KAsxujWUJUiUpBo1c9Am
uLTbpCBRGTzp0EF5NmKlYXFVRtop2WqFZgpFoMOYWY7q4wrLxFh6y8fPhbDxunbFajIPsLeuQ1qc
lNfZRrB9DtEBPR4iRrZ/Kc6Z9npy1XjEZX5dRqwR3vrmRi+8nvJH0YXy4SLkuF8WwjAXBjpoDGCG
p+DUW6zVvOWD2iWrth8pej4VvVeNiyMeiykwHGL65919VoqxhRp6/h1/JMb/8uHWZY1Gb2yIiiIZ
lLG5c/LLfwx+gjgERHDyy/IXRjRFt/60afS06YdqvWZDdYSiu76CaKRcO8EiiDy4WsoGie6byOSd
UX2khQvx/INO3qNkwvg8zlxyr/1Wu02voAPVA/hOgv/+2dLGSEX52tN2/mTXCm14a0LjdJVQSDM5
mpiLvr7RfmtQY6eKeM6rHS5Q7OYQku9nIwJxtW3V+WzlIjscVHJGkgBW0EF4FalRYLWypZwERRu+
/PEePJNKk1ex4qStZs9mC5V16SrhwuC1l2XNrF51TI89CcbCbHk2XoOvQudGh36cyaBRo15JJZxh
KUUUwX2qf7cTbiE9e+rEAuQS+g7JKLLTy1XwrUHIA+fUDtWmFNvT0ctsSyUH85zQBxktUUvYyOrb
RyR+D6AEB2KQN5ZPoWF0jnFTi+196hMk5jw/k80tEiHKPaPCi2103BJNrZBcCdyqgKSDkNle/L9w
NgoSR85+E7gCxan0jgBhnxOk8Gf3hElM6D33jBkpaFs0P7l811V0TmLDuxD6JLuQepe9rW/qXqVM
AdbhgPP6amKO9Ayf5lUZmoXndHYrwjcsbEotVKL4RPc2bOfDoiYL/S/VUk492mMfjq+cgB6LGggz
zOD9L5kSKMJgLaXMwqZwnlNSvKQpdNMaJ43AUoOpoCJswVRTAET5woprH3As5panGZOG53n4iSda
IymhFooOEQTEohBsdwVCzfEu4GRzj9CnwS6wcYFGsllQDkd2zJXOskgHRkNj9vX9VUYZH6aL1v+H
umNCZqHolSjPaQJHgfqJFRObnX6FYI/voSNV3qshnQJwE53YQrkTSdHCNkya/Akdq5sX3ooGvKBo
snIYpHiSPRyri4Cn9rftM/pCn+Glr40VpTx1pmQjR4G/GJ3S0StH1WsEDVndD4HAwgn8YLD3M3ZV
9mAEirFQbrlXXaISo0OJtViNVivzoYwC6BnjhSG+u4ucCLGI6ny5kZrXCvsQiEGo1GyM8Yg8XNsJ
7CafUuYkDNKC/j8bl8kTq9Ju62Io9uuIqujrXVquDOtYw+1f3iYuq0lioc6wwPnmUSL3Wjudene5
SDsmv+vgWOgO14HH/BODqYPjh0kWVaJT/5hxAoQrNboXXvNqaCmfjbIfJcOlgdVqPSSHZHo67/8X
94azbyLiCVi18rcr4+5F2eP/V/i+Nu5e5XOTANF+G6qB2rrklTRQccoyO6cIDf4H4eq50VuC9b/g
k3sVNFFEoImje6CFCJU7CBMAnzZ3ZncwnOCK9t4jhBtvTcs37yE8dD3A1MmnM+SWYRgfjtswF09Z
CrLbJdZGMZM7nfmb2VsAF2B+0LYqYB2OBbzjhGrHIw334AeY+kbYYQNw+dZVOeKDZ8D+AOCgoeuo
MRAP02ybqlbTohzghKRNLoBd22BcwziyfiQsxOPjeKEkUBDfNTXlS/a5VCPeA2aVA+XBRSuuYz09
1ZtivPW6YxUKWH0A3/xVuS85PMkIgFaxqIG88P3+8fuOg3bQp4VHas7WD2gO1lPE3XZYrlscoWZJ
bVMenm85qEdYKOryH+hNSzmGmUL/JXfKqg2qFjr34C2OvNpD1CelKsMBtX6+AOr8xssTj5cGJJvy
Brm/XUed+z9dnK1NXq0qpR3xgd4S4FfR28c/MnPBSdR2JQAi7wBCPbCZ4MOhQE/ka3NPih1mftQI
1UgdKO+B0KYQeJBs1+zN5adnNlygEGsUfv7wp9gTJ/ZpTXvNKnKuN5uhScs72Y6stoJOZ+fYZpVA
ep2naLUPteOruHykDQP6gvOhgtkVkdNm+Auk3p1kPMmDqq9ybgrVOxgKCuPRvMc3gjYV9m1SKzcs
qrN3YG++hXegi6AbmAHZOkFTMLTOswGdaoQCcaGo0d2fjzlC8ZktRmUcBU9JBeJO4buGOZZESiSa
+jlypOmU00wQx/ycRdMT6BySGJz+rswb0XvQkTawZsLep60dM/XDgai93RTH+lY6HFe76XQ6XH2M
RLVB8Sb9od5Wbgaok0DWO/o7Wyu/4+dwS0RQPDtzxS73KXgHWyg5W7RXLJNnp5dnRyBECzFNWp4A
NK2Mv+ZxKu3nF5YwNy6HAqwVX6+6PhOzrdNR9IXsik933+3BVIyS03L5tChD1TeZhHX+tdJcDVyw
X5mqpubQ3k01QglZRzYE9WOAZBF9fP04VT89J0uLQI0frE26MmCL/qmpBG7NqRAEP4LkAhThs7r0
rVGcwLvTAa2TGQZ9hGR4gE2T5wt8ZeaW5g8uZUlS3JQJQQYkjrPbRV/DZGqeQ5LLAbJKTO3R56Jp
UzlHUrQjWPRjbxQIEkLRQFWbkZqC2Osm8xO3lPq37iNL5c4z9IDiGKq3sMGIwokUeyxSt3qVQKO0
dx/o8NQtDPVB/x39Cxc5kRLEyZwAaNTFfjs2rC65/CMbZZC7Jp1wxmR4rWvontYD2VpuCFxwydS5
Ik8D9ADi8hgf05l9YrLf2PXOeHqrQQz/vG/PIalx/5Teiq83s7iQHmoe1bdldTiOy6NN7bus0DAw
JmMTi8CVUd0CXhy9XpaAfDsMTJWZuxcwV43DesyvMthMFek6PDXBE9weFPdhmWyAgQA2lLbeypXY
f1P8l5hIfBaRilIn8ENhuovgaZhZb5+F398Lx5rQvYvQRyCkhi1iY+VjKo9vzTcu5PKMus2xSW0c
Z6QBTAPjSuOdBBj/3cXzCXleoKqWxOY+EsPwDmHMP2aMHd90dLRTpkhSf3mGXpcKNE7n5VCJuQut
RsosKuxi2CHqOoRMfwgHvP4zErnrkzz4tA/7kr1SwoWk7joDT3YHuONWtdJaF9ba4FMx45oChuY7
rw6kcRBTumkua+GxOFFmjd4Td5994qSz3Y3JyK8HtlXoj5LCrbNZlQcwQVUYkD+Mn33fCQJE8or/
bvmRABjuOkhpPWhQ8Bx0JTl/smYpo2GarQGuj8v3lAuXLG/tHObzUNGw5LWxCj8r3plWnpBnocaO
STTCB9DZ6HoyznBCK6cuJVr/MNG1yoEHbc8uB/TEqYSAnDqQTINZbB5LP+stzn1mDyr11MndEkfI
8hPDM2WlYPtoX2z3EEnB59zcqie/o4mhp7Q9wQDANlESrEGVLSXUBufh5JcVnWUyloC0HkL5j7IP
trb5ZlKSIQ4Oy07VDPkS2wso+Z+7/rfKXC0hDuU3eFqkK1STakqoXqZ0wAmJX3co7U0RvapuM9Hm
RMyXYznvuopT9dTUsz7jbYYZnx89QCsO3XJ0oat1AXmNVfHz6MWgM8S3dO013YpoSjmtiTuUKn/2
gy4vvqregl8R+6F/1Q6OtTeho01VP9OcOt8HZcpDTdkD6esbNNb1J6HWRpJaBhVkEKIFp6hBt9+8
IIlh+Z81LYajO8z6ApjHuhXzTH735sQALynpKWEAX1k5lplKUZG1XWYe61iFsCeERuh3A5qom4TK
Q7JjQAbeTbH05C3tIz+UIOeUipcluXr96F54uy/vCM7MZ3/9+K59WGODUuCXD6GGv3sr/qms7eq8
qtNqGdhor06pir0VCEbp1dBeGh7Rg/Z2kJfwDSIIkrLRulmoRC7lbzppiZTXrRog2VYVhLOUw2Jm
4+8b7kdkHNlJw6f+jorv2V8nTXLfSBnXZdt05bKO77sKfLPBVxrSDCXul3BJKwIuJGDk/R1ihBYS
afqKCzl0gTkAobD7YrLzfK10TQ2bWi4Mjj6Ymjvw3zrD345QaR6Y5dkggCMWpoO2vi9/QAs0jWke
bFyKu/imdHYiFYGaTvmlZEMwVbpd6iL97zWfZOrkvTdxHLWWGV2BrO1hqjGZkr7QPUhNNnCyLkrl
cu6Dc06PCLsk2Aa+c9e1NdhI8Vp8ESyPldqwnFIsDzmsOfzFS+NoWvT6YCwjU2akxk6D4sTsv64w
Dzws+5+4tTb6rRlKjAlRrMfo2CJUGUnVDDvrVzzJDUx6T3tkY7G6OjK4gyjLm312xFAMTVGpaWtc
oVT+x0dhNlojqgIIVKfbA1c8bKogEfGXyDEiIwNRVZT5rLMJBI1jInUZBCH1E+pnGzec4160peoJ
Boos/vIP8lJ2Wq1KeBMNrUgmxuli4RwebEQxkaojEq4z/SKb3NvNp208jFD6nUw62NoTG9gEFpU1
f8dS8Z4gxDex+SvMNJVu8rYro0u+4CfAJCEsJRLC5ohEqzcCUEqyzpswkGdODJIbqOsOY5KyVr3r
0UZJuvlGey6fmb9I+MWTCpovrVt3uGNcOjMLZ3BzW9LRW4FFOXFjzuz2/9OGo4Jar4kfthzk7V65
3ZCeCACEO7ioSKIQPZju6F+Fr3M8qH70OT0uY3q4JEX/9WfPMgY6E06Mk4kdi1jr0aM5U8vE3X8s
wC3TGU5SpZAB1Kdk5wvTcod46i/LKLjmIo/m42923IHSY+/K9NVzgrs/NiHDePvwxNTak3FbE+65
jPRpsk571VsNaJlmpJTK24yfWxxjLXep02PB/FyC4FfoeOpNd1+JPT5Jyh8NvSybyudjvS4oK+6K
R0bcBv4aMu27agxOSZTNDCyTmSKFv3aRM5ThsstcKBWMcMW0sjSl9agwHJErSocXPGNmTLpzdw8O
arZV1WwXv/yo00uHnyQ0h/wTN3FPTEJV5hnHvr1xNFGaftZO7/iSZWS5wlQWNnFUt5/zXax9tLwh
aV3xaTiqncMpoPCpip4fAUYdMkBfAQxqGj+98FOIUzoAfPZhdL5U8qnkDfCCPOGNItLw3YUqGST+
UnFhgX4UpoH1L/WRv7I33CCgggvT4I5kBaI7hqhW6L4Js7lacwdxP+DH+H1W7/U0Q6iutxMCby17
E+9AMx5tLIpVXgonNJZc8f2OgxppF8xK6CMfWMnAS9Rr3VWyg4qnH9rrvo6N5nQIDrvq4AavoZoA
bb6UFoRV0oFoJCtsmCzHXbmNEAwpts8VwAUkZQXWvaFQ7oHviDo4Umr4Y+NlSRsw0XByN25W2qDj
m6jqIrG00t19q68660L/Hh5vgdNTh8Li8pcO0FnuWKngU56Fut3m4a6vt/BX2utS3KDKbQ0h8Ja6
h27fKRmRnqc1ssf4oENHUJcXa5uqh2kGpw1DF59lKH1CuYRPMAJe0hgPuPsHGvJU9JkrJaFsZOHX
YViY9JFVJnahndgt5ki9RDurIEsGB6azct4J94qTwX52ysKb4UGYn4TEEmcvMDKEyyf0y7eG5F2i
UAU5vWo1w+MCA7nZya9jn/73WTfns10023davVNWMMknhCM3/Sb4c3brrSkCpLrEfs9AeyggRn64
y864CYj7SrYEcClJJjNciOMIhS7tkrOSWUbx4gCHkNzke/Uvlcx8ma2RcMHZf1Gl0xBI/iqNC3Hp
zGm9AGYcYPXYnlkzfVsOiBRW+RWqJXuLElvHb+oU4Dq2GBo7OvAKU4yaGezaSp3Y5kJXgrCGxTku
oTTDXe03H9AmHbK0xq/MEdFv9nV3DFHv4Tevk8+wOzu7hC70AMe+JGfnr4UFleidlmCUzNf5bU6H
hCmMr6pbKAVfCIM8LukTc9WXj7yPUm7a0sWMrrIKRlsiL5LZwOQ91XIsSvxWbzx3fX01dfSmcAdn
Ssq70qyQJZhQP5sFdlF343nBOX4qfuS7BptYb5/4MMvLysqzonfxW7s5reBPjv3X5Hm03FzmCOzQ
qzqD1kEL9zxKgInIPAJdDeUr7v/K/PUYui4gr3YMUIFpj/1vyLrO5moJLnWX/1Rh4megmYewbBxi
j5zs3fGHHL+fZIanJUSdCLacfcZMeyy1JYrQPRqiwQf2IJ0/CupNQmWz0az4FOd44OJ0ERFIuIZx
CszE0p41ZcDRDanYGYCv1t80vaFxv2bmZY/DBNqv51A+szLfEgGt5HXDbFnAi1iWLiuR88AYLSaQ
PtN/cnu8W9XKjtSCqWlKTjMmkWfGiQgg37A2Hp8gxcFU6NryIxn+82KLY7qLYgxsMQusyM9f8eRw
Bx+fbGomGH/YNglDvIUtVcAGJHk1/xQdF9fem6EADphzSPhx91T7qmdj4nSrBnApdP6q+XprG7/y
opXcf8BzJIIdhH653zJm9sbHNISkQgd6QhBBDsZiRd0UfYOf7EQN+WsxA5N2j1R6uwj76DtU1Agq
MoQ/xPSvMifZVyY2ModleFK6ddqWr53G7H04wUo+wF9y6hjcf/L4/vxsbBPh+gbNF1dbRj0nbOFB
8wwVuEuwYRWX6f0Ml+QadynN8QyrCKvT9AvqZUdeo0aiiy0ZQhxlk9lbt0PXb3KAQCEsbJw4lTa6
GAFXG1C+ApRCvHRCXrtPM2P6Utck3ut85BQ853n4a4cF9o8YLnHe1mMjD/NJyoW/ysM2azb3N21O
GrkF0FNIXoFosN7V93zbkM+ilmVzx+oGT/Wus6VHmC4nyI/4T4GYaWtsukjWap+1xqlMK5lLbjt4
WG+81yN7uLbB4FcHu4DISVSF5OsX3d0zkelGNP8MaWwKgoszktA7hZ9lY+zIuEaSJ9J81b6jY3Pb
5q6l3ToURXj+uHtCg/+Gyi3hay3DrNKoUyAS980uMZrrZoTrG46VXOA1p145mZ7NXXBYS7s6EXze
mijS4oZa9djss+xt3l8pzx5x0s3u/ITDKoy5IhI1tKsm0QCEIfHW59or24Ryf7HUVAb/ihR/fRa0
3JrQqnbFtdC87wZKUa0tof09XF6KLnT/XVlS/hwtWUaJmFPNqDPw3/GWO2+lgJfacsgn2uiw/HeF
6bgjIoDW0vbIMjieRj8DsEOqFwkKbe8U/Oih4gJyCq8J/eGnjmhvYc4j9qndw8evvyTUhHPEgWSI
NKxkMJFOdu8KpBfp4PNLWGA1JIvwg9QHBNOfoMuH3MeT2jn7qAjafOfkLzNSbQCxVDM3Hp1qgQqe
u0FyYrWU/ekkgcIWDAryLqgE/3AUhd09j4EDrCvovS6uAnUWcO7NUWE8M/QEfy1Cs5eVsO7ML9nB
YT/EwAqeyO8KCgjH+IyVWq5pcr2U0MGqZ/KVaH468Ny6MX+uGBkaAfKxEyvoVXPAKuLUEgWwRpYf
SPGClpBLfBBGx9DEfNCp/wtQDwqe9GVBI7Jcspb9yg5S1f1Gq8fIGSAokknYN8gjwsrt2Lg4lkMZ
uG6ZjLSaghDjCz1gqBY4Tx8F4UdQwG+WxAt9NsMImRHHC5d6+rfyE+KLJE4FxKmEPAt5PP0TvUg9
1r4buifXRZihZv6K04wUxtRDF1V5hez+naTW4xgsbBXaY95R3BfLATX9PTw7lA7fr0GCDnK0BlRH
Zs4LK5HObC34UtGVEo9ZY6/SWYm1t/tORH+HvAa8jNCODk0IfaRs1JTnYY7TngxT3hpH1m/hfE5M
aIuth9g5Zpb0Rh8XUfQP0u6LrR3h3MsFLqAHRhXWbavPzmokJhgrzniRKjhwMvmhJuHiFdQmpIvb
s9dlXKEYrhI1lbXQwgVXe99uxaZeRdf74IHiIG7/70/OvGnxFxujiRrEvEtZv2h8mXJSRbdSi4Vh
HShlCSnHXEwHqk/AWosX4y7z92gDs3Mw0OQJahdnl8JCIpVcPY+lGSME9JdiEuZYkRn2P3psiTtI
6iXw2ZYRjW049m/5regE9kHJz/rRSJQK3ujL+yvCRkaNVfOm8zoiHJ3hiy18Zj6RBwkZv2ld+1pb
tgnhvlxWFf8NUbTL31t049riFXfuKIk4ccj1Szr9PAoie+ZVRJYlj9aowtkh1RwJrXHIWwuH+EYJ
ztKhlRq/I5ay1YHGaf6DC17WjTrvJY9tgvgcVdy7WGgnklsjJmsE2HUFHUDw41TaOxzcunYh80Bb
gbm/vmIW2Xn/d+760etAPIxcaaQi2hN7O6ZDPrwN8s+8oW3HM263z0v5h0k596zPnau/2cXytghk
shugsKGGv61LUdHjbyd8Hpkgi/naR1h+PGcJKcZ5SIbNLu3QOd5nHV7geb61GFRkTf8RzwoKvVPt
KPnHENWsyQz3U2M+MjUH07Fn6ama1LiiOR5HLQQ3giOjH71RBygX5GD7upJn9P+rCpX10wixD7tb
KQh221Xo53+23DENMk7XvCVHYuAB0ltgWLF9BtEPU1zyxah4qQxdJ3fxRW+JuYLWAhy+CmV4VlBK
TReSrW76pjxdt7pS382kjuDMeh5XSCIiwmjl1typUJu0LOaB1kIqq5i9zUzN0Z+WiRcKuWPwdsSf
wDSSQTod5Rl42ChF3ZpXr7xXvJ8km+u5+Zs0ty+Wk2tIckBWMvHBS2Rr6DVII76cXl6YBzFDvH2o
7eWiaP3TV2843E9Ppx5QBi0PYShaBa4QuRCY8HqIrXwVh9Qd88TODGBwCzc5xyKJycWaNYvG4HWR
XddzQNDy7dLMI07hTH2+olmOPCgSE5PDCitwrStMA9yLKXHaF1GqNfpIbseEmaPsiprI68/v0PpD
jy8w3Iqq0LYSndQOZw4XZrkyOuYTTV81oDT9Nx1EKN50xUJMuD9WfgfkYtoenAXquNdAJCBgSqBd
M9l5QSOmz+5TQEwquvhdeVfsQO9yUcMxfgBqIM4ACQRPA3hzQ0Fo90hbAPt691co6lgqp8M9uDL8
3oFH4FZAhWH8iJC/Pij6EQM1eFB+s2OjKz1PYYurvPkLFjqMcBiVP+k5A+Kwz/DFdnWXLs6VoNzJ
U67LJM8wKQR07hgVOvbu0IVN9034xJh3pDrK6/m7SV5vc19bkm9q8rnaylEUz0OagmYA43yQ6OBr
hiXY3UNJ+vEV6ILNsXE9Ab8U5gsEnYNU2Cx86vMmlROJYwnT0KMiJl1kec/rA5cdkcpPopcT26QU
WEyEkF3rstPOBjWo82Y0o/5weRkhUGAIospSV2b8N0+dFY0rAr/ueQ14nYxXVR6/szgMuKQkN4pm
RPwTRwEfCZUdKVmuxCe6WIAt+YTXzpRVYoSaVB9i9UpiboL1e32JR6JJqkdxcRmsq0CQkgjjPHZs
oa7fFIgR9R7KhLV2VgqNVGgXLyew4nsjuBvxXExcP6Sf1xPBTXkGH1EWgiZJHLyIiMFHO2ycqTXA
MY1+sIeGGovQ5vLz8SfpH5BriGDV/3kHQPq7N/gtEWyfMTpg30LPs7DRAtN6Bzar+iY36CwzTCeF
SboNwt+CFwXGytW/ne60eRdhr5zlEPs88VfWZTs/g9tI+V+OuZmZ6VuQFRo0gRyFB+1EFZSU563b
lKITtLG8LKi7NpFVS5TKNOLWeHxdjNAa49ihYW6uvhsJWi8oAy4q4ayz4pRz9okc5aRmw0bexAIV
NvSZt2x5NxJ2CfHzVfkY95NPmE6QlfsHfl2XlrR9toCoyiRhf2aM3Uwi3qzkv1dnybx7VYkiqU0l
RzDvJoBB9n++p4b1oy3zKN4BALE6fSCTzHJbNnZAu5s+olfjYOUfjn5ShnpG1QYFms08gi/ywlQZ
X2IHA5rTCP80fdZjmpgJRxg5xmJCyqlkbUbu4LacpFknfBVTa2Ujh/Gf1LjBQ1iLeA7NnZ+KBlco
Fqe0K2y88ADPmhKC/q7KcJKS99AS7N3rRedSKWg5VXRGXaI7MymGEBIMvb74KZqmAWV5Gt1gc+3T
ZTX8YJE57IswP1gq2sbkhId98ZSqOBTIejU5xeKg8WIcvI9FpZU9kTlTHIHMVdG4ExlZ2PUjgiH2
6JaR6JkSaKVWoesidx+xvfBXGnC+ltHD4w6xw+yeGCUS0WkvqYOZ7lBHEjVeVkAOq28e/0TwhOyH
LBvFHx23BbHv8/4kGZuPEZ2ugnT4uPUaAvthyrukr9ZQIQd4gCNbqmndEWwerLuiWHUcwFmNmYIK
DgT2yWz8awP/gYCmtHpnlwoYux4IaYVI5GFTgLwb6jDhMoLSEMZjLWLWW0QmCy5cPX9qj+9g/Frt
fQAkzQ7oBu1AxNm9GR12g8T+a9iAToDtMzop8usC0NqqifDm0CX0JEEOlERvtcK7gF70lX9iAClH
7K19WclZtF4XRA/Y1V3pnYdMEfW9zsy732UzyXpkpz7Xb4rdHmhvMqh4k0xICrNoUfdoUHKoJVb7
dAw72ro9G4QGAvYciyoO1nq873uzxvhEpNsNwkgC65xRVUPGlHXbH4HaoZBGWDADdFiRfeaHToau
DWxe1CNJqu6CLy7BIVhZgg4kEMg6t3AEHpntcR59bi8M7SkyO7oa4X5BdYLugMJLn15est/0/PrW
TJu5XYUp6xc0v2ZR+hnlkw9+FIHI0Wxm/D3ahcQjtSJpfO+ECSuuIWQGUzKS029HyPGWrcD7jQjv
0Ea5EdUsl8RtaoIK2rKbL2ewRvpljUxpHwrg05Seyb3IVpZTKyCYj48gG1Z16cPJYuxMSvXgJKsz
Izzw8UHRYCruxc1SeqnT+Qw+b2fxzsO8E2x3WiCIeIov5xZYI2rDj1tU1mM+6pEXNKkEAssbpjsb
aqyiPInxga5Z6ZzwZJ4VCclQQ6P0VAW3SHCc1iE/A+BRBiGuDsDJfqXXuMsGBFZZNUnmsqCf5odp
baiFRnk8OD38M7g9z9oYf/vJzcIeebXrQsj6eJydYcmccKYKfg4CMSG4EBM9nfRhPVfLu3Rp81ID
Fh4t2tAQT5Q1ApEkp7jFfWiHATmy61V7qHSUIZ6B5iKPS30M+e6zheKQh3Yms8SRJjEThPM+oefW
Ip/V1OvZtrzQaPpAyhn2jWhSeMQWP0o70hiOp7jOpW2JuBbXOFlrc70m1hr13jKuHF7Y9cjYwV+G
D77Hx78yLeHPJxQLXLj3WbpZb7v0XFGQ1o9HnOFb9czDXA0b84l/9nKd+oUEMZps3oAIHKhIMQ97
s94QMOAdAsHkiWOGjN93sy4ETxuPkx+4+nhrkjd/avJ0IiqcQPIyWkeycnQj2zhfvNv1nkqcdO60
pD7CttOCjgHKJkx5/0lH0jen1ftqRKK7UAt7q6QBBJ/zj0X0oWAX7BnYu1ISFOtJDMkVOgmNqzlk
QOCn2a1hvkEBb/U3b8Y1tVboRMjQ2DP/SjnTWEeuujGBNgY7qnjoQDjcZcCm04wkwPfWxfi6xsm1
6FgqKV4X4Dtc08GjAvRJy+grZoeQM2KYvDnFoVh0CrmDYd368Ddk110y3njrcmJqQHKSsrx5I6Wf
VpnAjTlafDpzIG6WvUgP/GTibv4U/LH7MU9NU5fzoYa9n0Oi7fx6OsOeQEwYxfIcZgMqWxfaazPD
ZE2xB1ghrKS4V0Yd2a/+QfKgr4eEfNFSeX0lzb0IG5XByEm0VFoZjSxLg7cb0/kYXlu0xPffD8sU
jg6dnpi7tPo1I8H4S7r2ILsFxZG+72NFs32IqRxiFmWmjvnZAw3bXdY2FEfye3w7pDTLZKDJs83T
GgM9upiE2p2KvMGl2UqgGCjqAFEfrwzxOZsWOjqtekb41skaslqCh5MzoDyXmPMs8SiVCF93jpOI
DV6Pe36YEJBBtlYxxJAfa8wr6cGhUVGHtuk/KD7wDweZIqrERfuFiYbse77NDKVMxQGhvOwJfAil
xuLcjjHjksJ+zW8qDzYh+L+2ReuSHGetgSj01Hr1/AXVhT4vLN3aIODwo3Cc1Ywf4BnEBYzl4kqq
PoWH5wAAfqXml/ZftasrODppfEWDm8tr1WcU5DK1lQNBMYzByCIER/jTdWk59iYoLQoOOt4TsMRn
Q/mCXY+YRI82rmg8rWtD8RiJ4h/LHQbaKaT3O+fDJ7NdJySQYITw/2/Wl+umAZJyWh4OIYMjxi/c
CrK3RGckf0z3fQ2+G2GGCCF/OCqKd53Y6Ty18lQxx6SbcpG5Wa9a+TsFpEPQXcJTxAfMxqbYA8nu
qa+ejhIykd2FAEZlB70Ryb/y0crQg+Zy1CGgVRe7TZEYLTLvri9/G2clsGYK01hCiui3Yq/jftFv
5uRp1u/p6/dfoy3NbpKehHTRZ6Nhn+kq9oaZs6IaDRgxWYg0rCmZCnK2+nvc7bwwhAirVlsJ8fgp
IOuuJZa4ZI4dIitTUmFe150OXhDfKRohcWqBVTq6eugUOe52khHTIrxrvhAaJJZlwq2+4qUbH9pn
135PiT886MiNEC6tKR5bI11Z4+FByc0OeBFuCZ43NwTPggb92k2sfwHyzWOFaCsdWHf6AuxCluRy
UINEscJXNNSivknDcdgLmkLQKcC+G6Fj2pQNS7weRfNh/Lng7oCZ5nFAEi57nrFzDYt9Tgu1hQeQ
AA7WTlavg3kH1n6OuKOhyrQC63tCrMP8Zg79Clvrh7gbE4PzHeyPjCKY8qejAfju2h1nEK1ZzL1X
2rOYZOCHhqHZepLg+zXOky1K/pQceoPLPJe7GPb8+JsQKjW9CNcc8JZLWLZ0WXsqsXprNd57ZRFg
f9ZTs+L4xbk30BJ1orEy53vbQ9Nr/ZQ/WJ9qNAzwDix06nSl7upXw9Fo/m21bUtESVsuR2iANeyk
K75CsErj77cwE+I7F2W2tr+GTgUnpX0hEkjv3U1VM2PKCLCXxwBPU0E0uT4EMahWnR07fFWC4o8h
0za0tgo405J8tHKZ7BTLh0TvJJNwX1bCRgfukY/FHMFZykzkFKzUp3b9cO2XRVjrLJ6inaKTHEbH
826ays9hb2zBuxKXV85ACV3zKoi86uPspJRGbBEJVH/c8rhjWR65boysl3ALN+XrZ+99eum/jHgQ
Zugq0kKMcPbNpCClwYvtim6Mi8kOc6w5p85DVnUbT2ovq2GwKclvEqLJarshJXIkr8tRTBiBZZj9
uWj/icSOSRdzlgtOn0E3+1EDEpRfxSD3GO3VQmcxaOqrJWHXGUvzx7IgtVYzjFih79RS9npn0QSq
Vbegod3e6+jPmaXvlurMFfeeyjTn3qPkayouSqsNmtdZ4lKYVTUoslh7m4PKPfWKEYkp4LFa57a7
+zR0eKik6gi4KV2UQCdY4YT4UfHKgc7FngFy06NsLGfejU2hyVKWWr7HUsWcMlrtozGdFxlR4XXr
+3dzSfXKSURaXaizcw+eglAfw8aoIQ2rq3C3JVFaG9e2+NEkExYghKHDT1F0SlvAJ5z5chHj7Ry9
iCp7qNnj9pQbMI//2xLb00pLoRCkNi9NtW/mmMEpTw1Ta2tnWVnirIg/RKU8MPqkCL2yOyeAnF78
DZW0bikjbwE8AoNcevewqtq87e0hgFVy2Jcr/ZU5Nur5IuIflpMX9J1pdRRDTS1s2TEVFfSs2L4k
uAS++aFOKmdIri+MSarmPOaWNcSYFK7fmxyErB78f+FKmnwVHioI5uJHtJyREBHLNx/ZpRYWWhYJ
kQ+Bqz4wFLb/auMby8uYogcUlXGhJDtOs+QTv5Ud/2pzJfX/P1T8jfOMZ06o1sXFJgrz03rScyRT
f+7f3nZwyj+W6n1QrJUMsNtYD+bfC/AQGjL6w7F0XBJ5sVR+bPxvUboFj1TTu5hj84+h0adoyp2o
4vuZLd9gPM/ZkIJ73fzOPjh6/6feOJQKBSPhw8jrFCet6kwfwMtjwKiBXCvUCWz9HgIG61PeA8+t
WMTaIgo3xMmOSWNa0K66e8i6Ed1sAYDt4gACAvOpr5rk7RFMB6zVijVTksFP8q8eIfjudJoEB20z
149bdmBShwS1/giWQfaZWds6bdsuAGKfB3nGjdGIX/YbISmqMyMnQEmVi5crneqC10xx/uxJt4Au
3U3EdamKoA8Bqb9UVVDVMjXkIq4HO9jxGf51nvc3ZEQ6GaNYTlXYkvsgzOtD9Sln5acAppz6xVr/
W+N0WIWZqxUimyWlcrMdeTXywja/bprDovEXZ8H+QFsuXxkPckkSQ894CZIOT450IuSJWc9tXCna
rzgoYpaz1+ICxYTqWMvh3jTOYfWG4w9ZktO4ksUxVQV1JxskGtwU45Pw79kWFbQyMuznifQrtRT7
9MXAMyNZA4dHuTBM0yE3xCR2ZFtfDyS8ZMyUh9SEq4vfO4wy3Vdbl3v/3IhDwDWgs5V84xNAePZe
iJQGVIgIn22607Xl1NkV6zS15GcSYJIXWK7nmmhpURgXjqWH2HL8XXJzMotmJImH2rpfNUFWc4mt
/mrK1+CHO9hyfvI8lGMODpf5GozjKYbk+OADLZGjFdjT7VsaOtC9NovjqwUMMAJaZwnHSRTL6CPN
ARo3YPgAmNBeSrMNJTy96glFyTbOGrHLamDhY3Y7VEzxEktBxIPkBjodRW97K0Zqke3jNTuIKRQ3
lzLWWd9NnkJ1PKzSJKYsCw6RT5oCny/nCHqFSPJMUvY3zHIEeyZ2s3raGUzL3RLsQ3bcfwVRojGs
/Xh/eWUlBUdvK7BAUiw0bUu8QIfboKu85447qiuBSAyW8ldIJfUiMd7raZehBO3665M0TU3jua9U
4FUuJ1fF9XG3TfUFl9ZqxrvMweyLmGJwCEyrmn68plVGa1aePQIVBvU+97rQ42g21n02jQIPQ0tS
gF7BPG7Mr58erRo57GPk2MLkIBKx6zeewONzNhr0ZvPeZK1j9LGkQw+A7R5d5s1tSVlx4syPqNH8
IA4XI4I3Oqam1XQKAmPCxfXywcsbCdT6izP62/ZeX0rqTV+Vw57xFlmOKCNX9XonqtUrnrYExYDI
zAt8xp3aDsfU+UBFjsdlNjSHH9S8wQB19m4Dn5SQGs36O2GlBs/dAUN5ZHH9VkQYRMPei7pXVUqy
ZjP+iexZR2AGl57LaEJITBOGvpNCfbijkWbRg2F0DHTo6y52ZN4BzMMlUE4GbSj8h/z5dhVx4S64
saPqjCoPHo/kGgGeDW8QJcOcS26nNrLku67Es5EkS5teXdNFXYn4ktROe8VD/Uj/g9h5p0URVoWZ
ne+2MJfddJ0JwJ5+zeMBSrSBkpkHecVX8VU5UkXpFVxi5MF0vtCChxuW1MU5ZpQ9s5EAD76+pFvT
zSaMFwiLrR3DwllXKfyc0MKlH9k3bMK6c3NXEzfQjz1WeiE7p/sRD2EX7/bu1KB091N+fj07pbvv
+Ps+GIi3Ra4hX2nafIgsx0lB1J+ZGv/Y/pVgHpezlVGe+Nl/HQcH50mBffZAFIEksFh2s90quU+d
qytYWJX1z9cE11V+SCB8JIrENIWP0HDHaMdjZ0KT6jcLY0SxQKbY03UrtFEnkf2w4hMKWIUz6tv9
qZFw/ynhUA/QTNGi2uzw6x4tSKlTDBasG/QkOpeYjAyioV6E7WpT+ouXcTqS3ID2JSt51p2w8jvz
xZyL3K72zsh9kIWZCRNuGYnuEj5n6bm/GdKRyYHPIjFRYCs4VEb5iDKDaelmZKKBYKTZPqUeH+Vr
2PQoW0gtnqtXFin0in6ShHjspSSptbou+sx3YK49xsDUyyWX4l4J/4sKXOOfg91wRFKBBOoNEJIs
IzCXm5A9rtEqtROqVAiXE1huyJ3PGnC36XxHJRmFvaHxonZKuO/KFOZuQMoaZIhGDvkVuo3ffsEQ
pZ+7in5qRXQPrqeCuJojNcMjmUE/PTyZlaRQ9WRcjlkGK34KoR5EZacKhKacBMAdtdXcOqmG/1g9
btMo+vypcUgIt+fQQPPIAw3gCy5toHnM7lIHBTyX2pdOgeCsuJY2jxVZsYMLCDUDG9YzdkXsFAdQ
xjyCUVBXIV4V32e3QhdxiCCIlvgPcPtEtQ5ndfn6SDGNn7/axt2qG2fqIcdqe0mWLiqeOiCgoPBA
YwsspCiK1MnzcC7IN8R7QaOOmn6Ga5CQ9N7aplIcCck9ixCPYHmZ0tM22llaCm5ApaXssbUYhlPq
6qpvYTZdwGyLLDLqIG8bBFS/9TwChsUFCQh4+SO9qfOMnmhuqYkUXh32wDjW5KPMIw3qGrVeKvbG
e8z6a9yvbcIhiT8E3807cfXwSkDQOcNJsDgb7Ed5tDEOG6l+vC0uQmHNqbQ7TNOgKd/zCv/YovnQ
WhMj6sdx5hcjo/pPxtheaRwWtUycKIfuTBPkL5QaBOBNVdtBmw/4i7631UPVFOxm87n4VuDyCeGA
LUGaeWG2o9xzVdpuHdbkMszq2UA/llTn5QFNMRm0HxSWdEe7ymjeTSfG5B3h3uBsidRs/OjrECQs
79aRbqt8I/H4ss15uFOKenbWd9gtRpq6yDgtrL0w+x4zjnQW63jfq2HZfrEW9Kw0fhEUOlNz3XxA
R+Ujn3jesHR5wB2JhL6xGCy9wp9ZH9bJnIirFGcgSTNmFx4QuCjlM0vQlCYw/wnL80jVkkMW4bWM
3kl/CPduBON2ze6qzwLNLAOGg6r3ISPALKX1xXtYw7tgwXAkK2vslEg9y9ojMaX3OuCKej2hlqwV
qrnahRQrHHwbvhblX9ABFDRYqVJURYxPWu4yhgz7V/72DgHitqFnlezgQgpIanEWkzB7BoxdFlX+
wm50DdpNI6MF9zNhwp3k5CCTuTQYRZVhLMrRGl6aPBZa8PFYu9OvDoS9KanoKk5J5Fcm+3zwwety
l61JPR0Ivrn2bZmk+XIdyEkuoTOeCIOyk0hCo5ZXgtfb12USyhO7hQWFhsl6/6nf/+ouhGwi9cPO
bxJ03hS9WefXPbhbz5io5MgyA6wZ1Veo6PAcw6Kn2ojTWfa0g0defY9h700LPuJsCnXPDpcS8nBa
4C/7bZFoksbdHxpWJY5KnBCDWqmez9gfOedPzrFWWg9h5V8vMUvo8LyMOwYh7TWDQ6DJoT4kifBl
W0TDbUmsGd5IoAxpjasilvqSCIlL1nJutkz5gPRBACZ71VQVM7ERPQgexhxaIJGiJSqVOxpXT+IB
VeNaHrY41G+QELTk5qf1AGrKwktQ0mVYpG5Mn7zepUvEzfze6Ql9ELcQ9WsREMewSUEexvirOmdQ
BalUf+C/GALxMmZPE+zozdnnWBNZjVt7+d54KRUVjPY8h47CRjk09Zcjn9DqcRmqlR2WDSHssO7y
umA8BYFtyYqwrvTRgnDLUw0QQKlFxeyOxLEzVHzI5ePMlfr2BaskiVvS6DcW00T0+19+1B/9JlJX
mUXijJBvbh3xjuu2m0CjY0MTCJM8LI3N3aI+FVyUOnzeQjeilFFPNkjdCScFynfeEhdroyDtKNV6
A1Zx/EQJNAQQWMMgf10pvYN2PYvJ/qDX8eAbTMf/nYWHalSWeFqLzTjAt7GdCHLVCoDewxYohGSO
o/9ll1MoF4uH3TNojA6We5mWEYS5Qx7Sw+45wrXiBpgTlEJXypT10o0gY8q9899DfAPpSh6HFhK8
AVmwLMnJsddglr2ZGVsTUImHIeNkZH0L2jm29GIawlNQHdJm5T+QMfI0dAc33raN4fFBux0200OX
uPFM+Y1LIgnXc6s7HZurDlripmBZcxKjEOE54P4+iJo1zk5h4bkmFS3JdRTq9DRfstKTHqNnyN1Q
9qyYd09KMomkKh5P80hg0faTbDkVeG4LgpV2gXy8vgI9XI5I8X32dTsTiZ6OPUQfwIxH8OvXfP7o
PQ/m41BQi5O82Xnm7rE6BYgOCiz+b6u3VeaI+sEFaytWcH/xxm6xIkKUbC/8kXW1Dqa+s1sP8ymS
5+uD+IEhbmx+vayEIOuee5Id9/7Vun3q3fZ75AEK0JhSJsyCuyLuHLoxtRA+DJlGuP6M3n+C2sQs
d0b30Re1zX+GAARxXH2ku5p7kesAaABo6htyW0Adyh0/dxGs9j1g/zQUSHJ1l/RudOJ80Tg/Dgem
NZsBnHvmUQubD8PtHoKLdHBJfOWxIMQR32hTEi8c1owNcYBG/QtKH6GFDPvT5AnAdkl3WefGVO9k
FMP2jjTpoZ+rs68APgzOuH9S+if7xMlA8t0zCB2YcEjk+S4w63IDG9z3lIk9l+YRwZYV2tah8O/N
dDi3JaqrItw9ixMNuQbb4K++AweLdMM0Dyf00BT3PIA1BefblhGPCSKkaxgU00ghNtfvNLWPVZUw
vN2y8hwOnPGlq9PR8DAFhZZatOJOU3uFYFYs9LFDPYtXup8Tz5ni8jILelmFMQv6SUbakODD5f7B
zdQrd2dW8tmaSRVWKXe01NfIL/+E1MyqXFnrfCAilycVZ/PlvZ2JL7TVvZeE8IBfaos7U8XmIDcz
c8+8/5PJfy/VLWMr6pfPsh+IulvIvs+FuQj2d1bqf0ilMdRDtiE69FkvpAUt54KM2u8hJLbnOLaL
hYpmJ1IZErwFVBWfb5NgVuJSSYXPBRFCJ2mmnOzAg/yukJSzyW8sg4YjKP8DO4mPgy1pg/lA7SgK
7jgEc26MPDhqkqeGavCCnyE/kP1lrJBGkpZz1rVp4hvjkTJINGgPAPsgxpUevfbgK5WFS0T2y5bs
1IJPoYX7kbA2mjfW+9I3pqzuC50tvD0VEoQUVuO/fjFamUD6ObxBPzo6flxYDmDooUIYW9SuF9sf
p3QOLrLuzOH7YHJcDmgEsCHFOR3MCcm8lV8L0+txoBniWLcYxVpilSLb5fHo80q9EewEbGsxqTGy
gqTln+pn3H07trQzBWPxiUVxvpYRg0N5WsP3KP2UPmRo2xq5VPZyp26qpUbpw5kDWunBa+EMl6xT
vMoEps5Sj+MktxOhM7mKWJIhG+sucu6KcsBS/gwSQLYBbOpDrUgbfgmg2aZvKq7SU7G0fPPnNtfs
/YX7qAxZ2ZNibBVBuva6lLIQVwpx3Qh3eWh+Ui+PXZ3LkWFcHuF5Dqzz3Fc1F/ObNRoILVyf5Blr
ie5hyQ1t3SVB0a0wK1e+L9HmOWOje9I5qDDogXIroww9HW6ZY4v/KY8odYGPRm6mgvg7T3XBZTE8
+Be9dtZaSvDO5SSCO5tdWxRE/v17zi8JludHKI8AL0Q+YDcK1NLFJ9ycASNzDEO2E87KAQr20B7O
g2UPSp3qWMqvmPj6b0YI6Y37ZAzeAJtiCDTLipp+uV3muunpSMjaYQy4bzDUhH6rS106sQm2Xgj7
a5mYWYdFbWy0EO6uAM4yIdoO4z3HPapC/5dscl980yq+bZ7VTHc1JN8WD71S0dB/759fSt+e5bOZ
3l1Al0zAe31RID1440689N0Jmi4oEDqCF6zrzKdWcgbonAq6rBDbM+CDuSmsC97Sg05nvBzxvQse
/DqiiOQX37DuhlM9+zqwDaTywc1PgHtIsxATW9CGi2Ry5IAjTvkaQJMdN03cQUs7ZFvLYd4Pg+Bg
pGUXRr2/wOKWxnmCVDIQhQ3sX/yeVOQPuer/vZPdFiuSAs/oe2o7AqtdxCQy+KwCoAqcGfSRk8/q
PEYpRxl/tE+4Eg8LdEZ0LS/xM29vHdyXVNCnm5VsQwPkX5AVJzS9QyCVJo7TI4KhHieD/76gw6Zi
94DEy/Ls3FdkZof7WRfIiaZaXxHJQGxmf0frqC/P4kSmvX+oOydTUrwnC7WqDffsqOZGgQ6noK8E
0r/MZorNo46szDHi//9bjUo2KDvRpWuohWQaZBGndp5Oq2KWFwDhx9nKqXsiJY5KecS0XDHXgsVW
k5SRWAv4AMULwhctIW+45jFXE2IYm+dgpHrSvIfLif1UfrLs7NB9pOD2p+lhRBP55EwcXkeSeypg
XLpuyi4BfzffmI2riDwhdAAxQMr126U6BAOE1rSD2h+QHqQ6qEvuMsBxUAAA+a5gFplAAmBU3rIo
NcUACFZ463Xa/DkuojoOj0TrbfRsx2BNwfIkeGKkDc9s0rj5/gBERxiuulGODoBrbYO084jyXoyc
NixtWMw71r4FmyiAHi3WxlblP5PTaKVv4XrEcm6s68f4z6CR39HLkCn6Uua5hk8dfBBsve25Ldqx
bgRXi7V+O5jAOH7ib69207t4cz0g/FkPbEuVtlj4Wcvwsxi6RFFyItIVa+LvD6+VclzTSUfaNzRB
JOmK5iDR2zNsHQEGOLaieKz3efm7ZNOGzEmCyIsFYK1F6FwDGmVyoy3Rh/BaShKoi4BXrKmGfUvN
Nd4Q50RzU9CqGsswKPBELzOkkzrQBE5ay9AQ63KNbSugPmiCndeqxLbvqEpSEbGZCx7/tMzliQiQ
MZHBcaJ/i2Zs9Ojha6eJPHsVmMgga8ZmUqyoDt1iQEwqvYfAoG0h1NLvsRgwZmCvvoUng/+jX9LH
xDUMZWdRohHnMXjBXjDIR4+H5H432jBTPDUMBvo5FOJ+ErWwJVBSEEfwcQCJC3fzM6EEw5z8rqo3
uMj+eJrClA4YtJOg9/8PX80rTI7PTlrEwOad1qGEPbfoUp2GqcAEOTI8xZypzVpJOA9oSikZiZXn
2h6+T3ACiSR0xUcYnlfzQMF69BQ6WHOmBPd70jJno2EVfyzTEVZN7sEJ29Yj2QIRYxSLNTHSYrOd
k+mPYih4y+ZEXPwoPNAtJkBdMXjaAbu5lzRuO0Ag9yZYv2mZv19dhdfs8uEiupnf9OzdyfxZr0qj
l68ppC/3AoCbIUve6r3+fz+BMesBFKCuJPlwJbs0Rfg1BULGlIkIW4Nsy/RC4uN7nSUxtVYgh0+9
szPdj+UcOS8WktUm3fwO+agSvx/M8c5/uw/7C4F94qUQtL5laj4fiDKpSHgi5Bt3e7N1Vlg+fYLo
zZNUrtEG9XWflC4OUqVWlDQUtJAuPNRUmWa1oyrrjThYPWCDy+D1rTC3Fz0gAvbrfdi3BBIDznoU
ao2wGvYKGd+2/EUAMCV90cIOXuZvjkwanE/LJID8zszNkBXTuvIv1CtAyS+0rK2y2M5m0uFrqnva
TVJQ8FROnHUYwMNY4tIGP6O1wZthFjAWwVrbHjtpnGfAnSKEfcWRRnf12n2cjvPD9TqcQSSchPTn
ylKdiesrzAPCnuQGHkFj0wWaIueqYTk0kFILITfeWB4luuY56C+IhPBKFgwKZcjyzk2W1HbNfb88
15vLfQvWFUdh8A+PU7UZu3eZ+SRMV3AN6lM761f/Wq6X1qyLiYwWx/Q//aOyOM3H1ErOFqhVlsah
hBQRfKrA3pgjHZUFiRoTe03O8pAJxsmHHVHc8bBniTa9gZQmJT0kL+kGJiPpOcIpj+OimX+Ge5hV
eHLsaQe/DEKeJ0QYCihJzEZPHUp5/u++cpnbdKPVJ8x2IWiLI5RPTR0m/jGtnaH2Zokz6mlnvYQJ
DsYdHCab+C3w3Dh5UUPPDNvafgkAJtBSpTHf4cLL21jBUKcYS/9pEtjCdAAmVZD2TLJ/bY8jjS4T
HDgd4EBrZWqOPi8MLp+0MKQ87NW7RaDNir+P6t1aLyebqD2eLeMO3aozelry0K7pjCH5Dz1uiKkp
ISPR4i1yB+BMIpXPohYa5/AKd4PdY/taTDeuZ7+JRwl7c/Id4DokIVFDtBzQBGJquJmHzRWi1WLN
E7xHGR4wgGmmP0uRjXhsZSDOUtud3wci5O4CpdNoKhcv5hKBkm3YG8ieb8+aZyzwsh8I7S5qvxjH
MVGb6PIeeeb148GWyPieztTLaGS3qeBugLYkkjCRrcdlpAdWHH94wH62SR3+NzfBpBbdMQ6c6/it
Ay8Qb9rVrJC617KkQHeopHYFHkmmHZu8ZbeyaEkhTXixRw7XHIKJSu20CHS+ouaHW3wytNhURYqE
hqsgJv14C/opeS0ek/FBRRuNcjTXMBKfp4TWJHhZosDabCXro0yYJ+7Xd8lrlMM+iWB7tER5MosV
lgM/+w6f35WFTZEnIvJiZbaxuX5S0yUw/+g/cmeGh1RqqFn48Pr6Ks6tAnjSpcRsFsnauW8OeICn
X1fx1uWGy2uppd4bGu+SiGdjjLGL5PQwON8Ykqv+4dWgsA/CLNd7EdxexVvcBYHOZCCsAZ+onD79
oTtafVlPZ9At+1TTKs1Yi/xYWJ8BaUCnDFcZgSoCb7wCx1slaHL7Jot9LvAbXfaEvfbLLiHM/u5B
NXVTYmNa51PbMRG91SZV8+ChMSYaHSgRxRkO3VNJZ+O5+SVqPshaaq4AnXCGvl4jJZ9FOR8HSe66
mh24rJRtVav3dcmG4OJy6MapwJWlkq0rItjFjvDJVcDZDZ/v8Gqq0cAvSpTmM7J1Ai1AucWfyMre
Yf+A7KMyZMeYF3zCAj2JiuP8g/G1iO4Ni0yEtEZSHLnMxsh1kmhdg3APaSOGzyWI34Ao1wq1HBEV
Ods8YlfCwmNzvAng341FhCTYJ7pWzmfWkg+V0HiPzKyHnq0izh1ru+pw1K6gVyeRmn7lf1Fs5eya
wFkNBxjOc0XFUcwFc19xf3JnBYr1ZHLoXcJHNkgXH0oXtaZ2AEfXmvYGdjZ/6CCGqWKnRGO1sqIH
JaFycvOJmWBCYvxHbIRsDfBCNVoosk4Tjv1JvPUDxjYFyuWygAZlkWL4A5laax4DwOmcP0/LDth1
18rlu4zGr8f5gthlZU2o3cdL/FhkNvodIrvUSqQtZY/CyvNnV1nTeavrQ0H6DafmkvkoZWCNvb9A
MF4+tV+URrAQV1Kmxky+jYpP21e8SVg3bf1y1aaOZ4P/2J3cZLNmANz3+cYTs5b9tQHCa0yot6Wb
coZIi6vxBaJtLtMh0uAHpRju33h1FIi7tsxw6viuVFLzQa82fDWzowI/NDtrvlgIZgFcxWt+FcOg
QSVjcaSX9q0sMoErVmpUQKaEgRo22CZgZkNbACwC+/UkRVAEMRAo/e1mtbjqrHYowK7UU20cgVyc
SzyV9jTt/P4sEb9yn470HnGjqY/AR1zSZjRVmY6yDohHkgIrv02BKUZa6xM/vTM4dOtpnowN39l9
Dh+aSEiYT5cJjF9jjvMP2V0KlPLPjibMEAZ0WKTQprkNddCqQfp3/glj4PGCdroNBqraxse1nj7V
Q0wSrta+VbV5t06HgqIc+kHZ+dpI8Ra4/BwL8Cs67TeIIqEvjMJT7Z2elQ2C91iFLFDERYT0qOFi
FfOZgIrHrhdtzZkFX9ARhGS53sWs0QqsD/AFr1U8hhpuCNBMNbCAT5t0DRDrSuXL8VmyRZ36fRnZ
5TSjypnSTowDp435MZ8S8+8S5+iRfX2rrJr2NKl3KEfWlMqbtTOqGVrYflUZtA1Obut5QxdIUdlX
Ci9KEFvO54NcJJsY4z3iIvbfMGbUKwi4TXYxnHhm1ck6c13mXrvFRvFiOeRNvJKwap6MzaSg5zzA
t8DH+/1b79xpfutMupqqKzjBPiR3w5t29FBq4n/JojsCWFKdRCNdCX3oirCiWFSl3NMTD6WL2UmQ
Qz1FiyfCEAIW+bTbiCgk4ANhqnpcK/i5uA6kuZq49wgTgPLtWkP/OUlKjU4aYnW8SQxCVRA3DJPP
wx1eFOQIFiHveiDESALVlwiVLUt52FH1dPOCkO6d8KqO97ONkGzp+qCUmjzW5JnT5zjvZLI+9Ut/
//ql1dxRu5LR+3+PccP86JfvgqAhxcT9iCjil1OEgU1Vutw/uptMaF66H3B9/E8IGyWulnnhh0NH
vvNcnurYOkpa/Pc6r9/gnFIBj6UfWGLi8+AwWx4u7HBTwF4ZlDfFBkS4ZJ3jbZeb7ldVSpk3J6oO
LSoSQ2Yy3VIv0pnRxuJyxceHBpvEsrKliGaANguEvWYeIRkEoGtai0WuEM6Yviz3hX/XGcnmv/Zx
dVe+iZwRdWTz0FDvfnBQtTCd+HgDisG60lcOjOiDt3WkDeL6VK/32r4utV41ztqw/DDPxnnksR9m
s+O248op2aW0oSRGuCZu8iazJAjErxWOzzKWiCp8oITQlnxoAnWBnW2ZA+0UvpxE9zdnWURaDLZA
wsWdf5aaeMeTdXjmzgYJI848u1Kr0e62Pu33f2vBC6hpRh4cJXSymX0NmQ3z48fxEIw7o81ywL/u
R940GK4fYE+q2qZDy8j4WqfFUNYV37PKOsQr5p9eOD4tExlbIzqyxiW0JdvlOs99SUUE0NFxBb14
ZMS1Qgsqdhu82ledt1cLD0NzNqkDfoSHS5X6iodFbeFblVJeb+gJNQ7MMKmPFFPw4fE0PotVTOQt
pFKqD+HSev9VcVv6noG/LcynSd8A3IInZCckHfQAzTMZgpjg1+iED+JnLRrszGlxk/ndMZWHzkMn
I3CRSziGykJaFwkmpoVgzPbvrcjk5BSrocrIAkBQirvq/u+s9UZ8Jl9Vu+YMjcQxkrOsn/MPDv6a
haXKnwms1KNF4fZ286hnkon0ZP6EHihSDyihe6pNdcz5xCUv09FGeVxqffyI1KRU0oxrGiKZWqOO
ICsyiKrnCWUptI3TpsVLhI3OfpBb6JXNOE5aZ/rMScgm0AH961bDzFknOcQMhEez0QrRN7E37bJd
H91Uhr4P868xWcEmsxS+lLhxC2ym802w01mE4M6CquMAUPr+p43uvM1HFcgxaMZOEUbY6Sbo+S46
2PD44/xg8Noye8Ye0/FZtNLs9/7GqffUoX/u1eYmAeq7MMLAwKiHKlUfmFWQOwJKUiPQ6kMH19PA
7TXgwOgh7UMxcHDWZ/gR/fnqq5H3xw52kho9wNd+4RHCvkLQ3c4lbz42xuzTMsNIjvNqRZUq1DiK
mX1vWYSIQtl9TzmKS8Fu9D1zW8LVjcsPbXILPX2xHft/VlBnM3rvd1W+hlLO6ArRZHR2KX0FRH1P
YDpb3c06YY1/Yyv8P8mVyMVtKBpbr7mvg+cyyxrNDtfeKNy55nbYElCTmF0v0hHbs0bSt1CA95w5
fdUkpNQPlf76mGfkfUj+6Hr3nKeOa3nRzjkLCCOf/9Sbq+Bu+Ggd8VepxMUeTqSdkLoQdoYqzwLn
AFRK6/VbY2IjxVA20opOEA9YUzwi6SU5ZYh0/v4KW83aVMwvDKO0eCTaKa/jWSuuE4mBgt33v8Tn
M5mcU3vPd3/nIPWg1ddZAJaUNAeSwTM1UD3wB5KToXz/7bkYjUhe4+1Ytx2J9Rrlh1k3q3jsJqDE
z7oaDUB3g37Dhgz4lDWq/aXRa5fTMf5DuIxF514BBgmIvwUplKFRTiNH3c5Z1HUHVUGmNrZI6nm2
jB19TYU2mGe3bNwtaKA9ccXA1RoYm0dvqco9pwx22AVefGbxETs2SPzat41+h/abXmKUox7hsl1T
wt3LFSiVJ1ozPSvrh7htX/CTcVd9nk7ibGsWRGknFasNRDyMlh7Ln5WsGvdI3B5GlGXFIqylDvKP
8hrJAFoDLReBOXB/fbEIw1WqNui4PjFWeoRaEcszH3XjEaZwaF8Cutg3t/YlVcnW3/LXfeb+TRrO
9o0IVNPkNOWsKIaNhOO4nT7kXAZqYcIO6PCfoj8eHy9urKdLqJFd/9G/toPujcupoexUmIkUT05E
bZwvFI61whHv/mRh+DAD6JseKmRAaYzoX4wInKZiLkEv0/olb3GgaqNn21Dihpp05rJxiMBt8UI/
PckcdpRCi4HdHRzphPDaAA/XPstKotae70ddB4xHTR4u479+9PfesiXrFiWBlPy5fpYQX551MvFb
pbyPOFmet14xxFokxO7NZF5wMHhcUSElm39vMA5E15hFf2zMe3nvELm+9Rbn7KwLYJHHcxkNNkdE
cGkvbTm9OfBe1V1T4rS9U4sEKbXee/0aJGrTDFFbW+kb1CUPxCt3VEDOjQets1P96BFmTavRXJ1l
sR/8dEi9ZgHpPsv5Czj3bvjJ3t7iuyFTNBMd7OZ9pR/CshyRLbAznMQWDheDgGMqTGYRdd+6l35U
1VGgy0E+uRP4YiKhqtLvkJQS6qwYSqJocvbF/x6Ng8lB/0J7zM/N4OR/R9TQtOG3TkexfcJzQNPe
8hN6datUT6kD4rjwboctXMhKu/bDQ08Z8Toy7OPfshE3hQKFf0nwvntOplsWZFlHYDIvxzKNA7Hx
xxwyu/w22SMXfVyn54iChTRquvZ1M18daytY+W86Bpjohla1sH6hWAtW4IvXVP93hIudw3tRAQWe
ZIAFm4ky5cCdRJkzZek7wVgqgh1NzUhnwie1wfQi2qNNOIieLQVbf5E/Rq9TEvmdL+LVRL5UjRK/
zxt1uChAbj9msqMmg0mvpTUmguD91m52K1IfydEua0raVc239XubJQZjQYiYQ6a0LA3OTalgY8TV
5jW46Osd2laZCewfrl1i9NMgVB2gmcM1nYTfrPafY6+NGpF0ZKkiqG3ejj8r/ggruF0B6IG8y1ai
351NpLYGqQgTJRuBUmtNHryth8RwXnECJnHLuu0Nt1LxCEQ4gAAeQL5EgiapOC5XYf/jshz6wGbJ
S8hWu67+BWL3FIpidSP55cjzAYI8CkdEPI4FrkIDgm7fJXw4vw4OnmKkQ7PmsCVdyndQnNAbcLlG
ofpg9MmtlioVperL3ElcCGjjYp6Sd66HEljbVpD6dT9loeKHoT1a2JRnmENCgU/KUkLBycg67PCw
WfTv5QQj/VzvxUu2hPrYL9aSM5ifC9oFxZgSIjIOexHTDP0162zee10vlZIUqCaXxrunc2WSMaI8
XFzUWlA/SxK2NJwBT4y3T15f5QBSYExRX6Ub5/yxpY+VzGsza3Q2mBnnqq/im/rQBuGr6TQJmLMZ
Noi/t4OSaeknI4kSs6e0SdvHxhkpozK1Wff1uyR7MDcXTJ9m9gKg7uuT41pfjsBp6n0aQ5oHZEpE
NqnQMh0Pqv46aLlXGvJfMPUJy4YHUEN9M9DzEzkqxU0KUUJuRKH1VU2IG1zjlev7YTYGhAZC7JE7
BUUfcdp44n3O7qb7ThLyhkuKwqDIjK6iDVr4FcX/a55jZvOANJ2VLorjH8EOYqF7M87DXNqT2oXm
3CTtpfiRu20WfuiugFE+1tBFtpfBtNZX6khoZ6LCObkm+MFaZ25KAQSJGc+zfY/xieFzZuTAjtUr
sY8lr7xYs+lqju/OHdVohHU2vsMXGtpHPYkd3XVgGCv/GKji4ZkHe/rVGTKqOVe9hfA1xixdCZj5
ARhwSc1xiz0+Q35OYoraHXz+po4ugv32e8A74toxdZLBOqRvc87dm5tN5XGHs+U8jxfUi0XcLMVS
NK1Do2+kBgnCR/35fdinPw3J4c/eTzPEl6FI97LmrIEf8CCv1RWv47xV2T7h5Vgy4hV9qt+6QYCF
HYWUKkvOFJJIq6PRlp+eEsvY/O1Dr8DXZLAiJ9jN3ziGJWBtG4cb6sJ5hw927YKf6Mdy7L2jlOOA
UXCgeysMHBdS9mm2hWodKDOuH846gp1zza75uDGYuY9u59jKKmFzRo9C2TlnA2AWNRJ/meDfx2u+
W1h1wVA+siqLYtMFS4faJ0aRwfpSSb6oO59+zc2YvvXOq3RC+hl5hrnsoMpD3y9OauC1u3hgOudV
Mp+zGgADpTCPCJ5n0E7UAJWCqaBTGI/nzscDQDTlEADS6Xu75NyHgy3LtItUQaebeSBZZ1NxbWmj
8hdy1cfILwESX4+n3obV3bU2q2y6N9GP6EK1iUXu7G1Uy80YhqF3LeO8MEfX5PAIxVbNHH10IbqU
lwOlv98Oho0S6puhMDo4/SxwNrRgYq8PJtefZrszMDEccBUeyTJgPSeWNMeFDNDBgwQpXpjOfjYJ
qE7ngQcr4HWbFw2n/X+sVDgkUPj3xVPXGmMyrtNIgkERG2q7VEg+Yn/V/+1iZMOh9VNRuo874ogP
F3rUP1088IZWccMBk5CFLiMu66cRzZY6e65JJRg9HA9GZoevH0XaRtD/jDnUpWQMAmRNoI3l2SVG
I98jUUiCNpalY7V4bJadhdn20E3aO4piWzSNTXfdOZSJ07xx2pzELE9iw2IvHf2klA9D41kZcSAF
zMnB+FKv88aRY2bjkT04nxkejta7Aouq08VFlxJsrACdlYqfF4rBAGo+3hmT/t/VB9FaVF1gHyXv
X1QJIWxshHnfg/S63v9IccM/CoRxRz5LNhkwGV3LKjUcc4N8Q5Mx3ADD1x4Dl9OdHmp5VcdEykPQ
IHb3l+2TqZNnldWNIPlKPj+63Q+G/AhBwcX6KjOtmGTNbbhvhLuKeT+IIAaV2UR5SvPEVLyTiVXH
AG8HguLi7eKmfs59tgvsZTBz8pvv90cgdQqqV08l0MZDa0ztpMT/UgT6ttsUX9jwUZ7aHdC210ip
jxYfDaB9fcT+Z1bbYw+97KCy5ahkLs65XtotUbpmDfJdA2TpjXNNpDz+4WVDHA0uwqI3JYpiXtPK
G9iF8/zhP9ZXYHl2J8oz82muOJe5IKdTzWxMdbaBuyP0XiHe1LxOI/kb3vhEQoqDU80533H/akUL
xWkZHqld7/+q2ocWwnl6raitwtKVkOeOAW4xq48g8yyfuLjl7+SoApwqviZ+fSE+TCMu/UDjSkGT
jyUQ9iSNfYvQpzkGe2IuT/IFYHLhsNcaU6LuftLPKhzFml3El2hNZXWXc0lOL6iJplBkKYTQ6iel
kmZOEjWCosnWGWmna4a/XIn6lbOBgvlBGx5X4qXQo/4jpJl16HlXmpkmQAngKbEtf9+zr1tHp9I+
NHFmroJHhLllTRMTHvgGwjiDVARd5u2KfEy7fIOmAp2RRmXzxoPMFpylAmPjMvNA9FkhdoZq3Y1N
MXAib2nMtMMn8ATIiNO9BcfwRFasMjePrSCqt7raaQGBjAGDV38R8zJuA5iVlY6qPn3Ecc9ZFekR
ZSEhfL0adoGy6NsQ2eKroFjNetkwOV/o8zUZqqvgRzHi+Bdkgl0LF9FIKkg4buItzbPD24Wqw5Ou
aMVtc2SMoIcywjjo4za9zbEFuk7KpVOun4yD7oN1a6UqWlMv33peaiod+2r/M3l9Ya1Fd+y8mwh6
Qd8S9DckDPpChpKBDA0Iay3LhCPPboURKtvuoMjofOokAJ0DmGA4E0MMLaDxGBq/vZWeX1bpM8MC
C7mwcfNf19mOn0hbf20B6UDgTpYq80QOzRza+ZYDU532sfZ+CjYGHXjwzBXHLlFKeBYbUjlflim2
IsHWkXC38rnXTIzMQMO+GmG7MTuPqIyk/mZIzlTA7f5XZNjAXhg0yfu0aOxeov+xE0eJvh6QsETi
O2/vmXf2iGa7eORkeSBxtauYFqtyLRafKvggueiIl6p/WNn8Hx+BTWteXvYFL0LxhJCXb9X2rk7F
VMJamJ+Q1TRjt0W8Bfq5WdfOrK8OyzCW1unJ/uqa4yip6noMbsVZWY9MrvVVXW3wMbrwJ/y1ao4C
IFiettmRAlK/RoTglZ1N2jX0HAxfr+CSv+561wbvmURvcgzAiV4QMllVDLhDRRWf/wGy3PvmGEzj
tp5BKv/xJ/v8HtP7CRmPWd0DLkzeIKBqFdkcv2JxpFJhLqcgA1I/01ao4DHizr1f+yl7Jq4PQMYN
yAUWfjm6kE60QD0nnMCz0s664DQa+F+wFaMLNQwJsda5CRS8IhXH45CSteF8UVpgn/eujZHc+MDO
VxVeKc+Hn4/vJeEZoQYBHLd+V+d/Buly/wkM4cSSnz2yc8ZnKeOR7FhJb5qXxhuxadl9X55kO1o0
Gj0plZSCLgyX9X6lHQ72Q6v0o+ozw2knCTh2W+P0Far7Zk6UcU27cjG0VC2Gu3PBiPf6eF4gWRkt
LVwX/h+cCMoS/CebUJNQB3kvz9umnrmi7Te0THTcve+g5rlOePyXqhytbaRQjIhpr4XICZHez2zv
IwnFpdePuEx2OqEOrBejUdePVYV5UbBBhKs/OFrzo6YcSgEkbO6Bgkh+rioixUKSvMFDuw75HwTr
BOEbvbtT/7s1dfM11VAOWeWLqn6SFiqzcEe2L36kkiBHBCm4COPYTUs8tGel8OA4AvYgbw1ilXx2
G6cYP/skcjC3ZHhADSAsa8qn+sCE1/749IKg5EyqkYftMGBjxSRq5ozqU169GvOAdLHLyjoiMxxa
F1keba0FT4Pp3woNMm0kdFk/ncdcm9s5AVcMVQwO9aF1U6gc35k9fUz7oPcz1TQcBSSyzCKx23j1
nKDJgDIcb/y3sKV2CTLBvAlz/chpOUTGdVsqI17u5nO62lRYNZOCynxm5b8cdK34MxOvc1eMhF56
O5+37thpldGMINejyuWSpPNohqVm5wRCqx+gAx98nL+9xpJXObYzj0EBhLEtdgtHOKOgmWXKJwz0
MjfAFlyFVtxr9f4ArSw17xHt+z/BTMkkhqfYBXEE9L4+UMhBT2NhuqSWUYAQQUWf5bLi66Mrm8zE
/oTHw098u5mtj5lLaHhCrGtkSQSGBLko57bMCANgMWq2+rzjdmE85OBkJ6an3D4/pewxIkOpDA2B
jZ/1yY94ewq/lc/p6F4GVrWiwqmr1DT93sivYyh9WVaH3DTVQ1WCq7vatB+8pY4tAU1I7iGzynn0
CnTNoEvXS56bqmJG0u2hvCNQwEPXC0hMJg/399kQXrYLS1nRKKtw5+1f13E0VqAr2NpOpWm+v5Dc
Am9AyyyAnE8M5Nj6myFFKuPluaxboES4NJQMP2PLQyLqhyMS4ZICT94C9yhV7M1TPd10wRWAVp3V
ICvCOSfkaXr3/wp6ZTBlLgClHYJnA8JtHNH/yPHk3F5CCtUOOU6bv/kd88EDNUlTW8Q4262bXM+D
eUZB7eBQOSKX5/zXAjKUEntyovXJNgd+kNRHYS2dn92nN7CG/vd+AAO/VJGTwyfQYEAw4N3V5Db3
kkxhWCigYWrDkcKgN+Ceg1a7T/VtJuT1zX4/LRwu3ypPqvv9MaVoFIWe9dn+DfhjNdbL/Ga0DE0z
cqNdvmjaHJsfJc+DmqRoi0Ge1YQVcUBjHIZQZ/MJ1wdwCopnsOYwf0jGMHPiABnjMktSS+cPgiwQ
yXxveWGB6DaHfYCNQ/MYEFKl3a+iM9PhjNrsnwnHb3+Kr41qcGi2lNU1ah0r1q/hvu/Z4H+/k3YT
ypoc9RIkTmROviO0S0yBASOccKTx52d5vFMApzgJ7LZG25EN/VUJOGpZkyUIh9MKzpfQ0tXtlbIh
pIzOQb74LT24NSOe9/n4DBqVZsJbEN570wroOfe8jc51Lpg0ae5ucmrxlHI9ZoaG9W0c0L35n1Of
xFZA8DLP6CefYJjRudb5FeEqeAm8h3PePgnQ7GkK1gFVNLAlr3Q/FCpJb8o1+UpZogcIWtqLy4w2
tQpLX8Z9+juJ1y6jKn2/v4nmh2zD81E6d9AyXMtzsAiZtw3GvLSKwjBUePUTTjLKDrkTkZHeofeh
ZxP9+Sh/fogKxOYu0lFCuShxoElwaHmfnCecS3m+8dmEmpIcG14QXj97jco+ronq12GqUUAc8sle
hJmcbuSpcPqaqKlNBSH7mNBdn/ufFJMQ7AgmCCKcKXOPIaW1gFymsEioYp8SBStYL1N+U8bVSAP2
OwmRBYwWBPstMm3qeS7j5DXkXKm5Rc+rm8ZGgBUT00cqEXFA3zDucLcDiMcoc+wLhqa5EVjnKq8Z
RaFvApL+0hAFcCthN2mpbo0Ffr+COFi5ltL24Ck4aUBkTaUpIfh61FWmje7WXM3sudrY305t0dCC
o6TA+mDEK8ALbzd1ive1D8+zc5kwnYyva/VF9cp2aeoBSAcrGn1z8UxE+mh8eCW9g4UF7GRdXPg+
1GKKYhxtHm4aVFt2+0ADwxkvgTZF5kmAlzmcpmYJODSfkRiCHWNkR94HxK5Xq/rS+v0gDBrNyuWM
xPg4s1z6oKn7W0NTCAvOzHhWcHnzHt/sO/R0ohhoxz9BaIFVIyFUbaWaCOk1q6ogp74rgRweBMuq
JwAHDrTIeo9+pBasKXHKr6ft6KqXUn9Uz+Mvqvxr6tb8GROth4jgFot6iMUesjg7V7F4xe6NGXf+
6fWb8RrPl4pWacBoYkdMzHhsM+6awtPi3AHHkcB1trMb79Hhv6MGC6flFhiziM9vYEnW6ZL581ae
npuuchzEZ6u4jik9B+m6SZoE91eBpLfWLfYrMXBE9ddRjDT0abzaWfstOu1xWOGWpIU/6MC3uQJc
ThnHQMioxUBHAA0CM0HG/a/V8daZPT+4rX7ST7M9R8UZbXwafbd3fESuxLqp6i68/rTD/SrYxV2/
0dQNd/dzt+zTo2DlR8kIi1JPHPibUAI5PNYwxJoOVDSco5Z+2xhmooJb5UGeInPq7OhIILjqEC4X
sgecMagSTOHsnBz25Dj9eQr+tY/SA2fAGx4ji/ng5pvBtW8+afh818tr9WG3rSJXaCgYb+arg/7h
sMcNEqq8DthvGUexab/VLJsITxqMBhPjuzEYUh8v12wFHFji0+IT21MpE5TFGCk+6JKDYQTgr65g
8tbWiwDuw46TOakntNRe/jn5jfBZMu8Ih63KSp1m0SKwPWAprsiNkSehNNSg+YETEnWZ2QlTjQWL
+qKdKjUVrn5Jzhco4JSWfs5zMs5eKFp77P9121KqpdDeS8OrAC+wBIaPlx6FA28p3GzdtSpx+3Ds
8MF2sr1oy8pnGS+fUqxx/WP3bvqoaoyoaIOmD6cp33Z/3cskT57o5UdfpPRkAGJnokNU8iUkfWbT
6MZEBvAheoI2RR7PKEpjFehD6FNLy5sA7M5bsbGNeBS0nvdbFtvDWvT7Ms03zeUNc02LU55RD3O/
NiM80m4K2G1rV6jc3oC1QBn/ZbWGPrcWJ0+WAsSNjXvCEc3pZwkEsPwH6qKsETzw0W5bm5zWVWJg
eYqA41Cl66dgPdfRsuQ9s07sZz/r0ccnR6I7OkR2lQdr4hGTy/f4gCFcyM6C35Hqd4J95dL7GwL3
sfYOJ88yw07G/VseoCsoeSb6c2OyiyDVaQnvzc/1QpMtMEcgIPAUSJwCdEMCXwX+gxPoJIz+fb4q
VlSc43sE20TK3J2UHKU2HmtsMSUn6RvnN2lnbZJsnM+EntrSMm/wl4uenC/bjNW50mZK11GXknGy
1Qpj3PzXbAAqslvJPvS73Z+LTs2pDgzBMo1/9nui5Xjnvwj+GKPYqsXIWZoTxqh2MljN/+IdP8/Q
LBk7ssyxbqsN/KIUbvTgPUafC4ydL52GOKq434TLPc2Iqg60L6TovwsNDwD9bdyUthSP8+2z8SfM
+ujItAbrAcknzr1pHhmZ9mXeBWCOJAY0dNKFrsm/UR5iLV/OCfxnsFhle42L9ALekDvNglsEZuvU
jYT5eyTqguv/RhgDkuNkTHcUV1kIQZdOrib3cj29+8ueB+K8ol6+jYe7ipa7ZiWUvqumjuRkDTmC
eZmOao6nSaF6nh1XVjcOkD7jQFocQxBcM5O0Gif8OUeC11ZUGqoRPfMyXG7LJLtm41prQe1W03S+
z4BI44Q/oitXvB6NriJiaIA+y0YIgrbGWsOl7APkEiPI4W9crWMvdqkyrnRCtK06DffBOZn3voLw
lwuPVFkgNifaTEU1Kod9k4dymg4kUDt3eYp7Ypz0FgUvMxDjKlBjib6K38YKX/oUSKQ5oNrPbMFk
VASFCS3Ku8xJP34jvnu1px2B+52MoNwzd8gq8kiA0ItQR2EFA7pxwkWsPnH9/zBkM/DrMaKTCGXV
2lN85UvoJJHzJ9LVd+2WSdgxd15Y8YtGmSy0iMIVCtM6Dd1XUc1p8vnocCvQOD6neJLkk3+c7hYS
rg+MBxIDiXzvQQRueV/YXQnGYVWSF9fZOIjRdMHL6tNsp8b2m7mzE+6f7fUs9s6z2E998BQKr8fA
U0X/bPtZ4gxNb/9/IUoY1FPm0Knj5QMQaLWHnspJ1SFVXS9MuVXUOPej9z/Lj/uj5oy0x7/r0/CI
MXYut3D6widNz9qlqOFMXMRCI7Sz3XP7AW+jP/tgNp+kVmjL87trwmhIRjH6ZDb9PO4yCZOv+/oM
8+b5XJVLaD4KNMNPBw7igup1xZ2GWD0Cbp6Bm7Cq/TZub9ijSzwegW0tck7ngeQrbt0VC6azm38b
2v3waj0B4w+P2DYxfg3kMyhSPsVU6RopwWZSEinpbpPxU0YteTVaRfphpZYh1xTz0M+ZUG3t7rub
fm5DZGzinVmTFHj1MFttwfQ/tY0QoP18uGAwsqsAV/JnLMAyUTjYWrM3EBkRzRCRmEoG0pfwpEGB
BAr2Z0lGn9vfuA+97IJgRb30tAcr/oKkaeP/Xe8NPyaPlDvYAC+ZpQFw5DFd3Wcvq6tSq/6fFwp0
E9IJ38HMPCvOWgasz78iHVgqYzwHRFbhHGLqqHw0ecdcnHC5N96I8OhxfUN338Ab3oIs8p23SwBt
ksX1yU2FklKW37xPlDpaTIvfHIIRJy/ZVdmohy6EZ0sXX33561R30qN8Y0k9XQKx+abBL84W89oa
F2B8/1HN+VQM1JDlIWNIs+f5+jV9lhzN6rzow9B/yNA7/BAP0lnln6P2sPFiXoViMBiXWCcH6O+Z
tJaCDLLt5AzzmnmGe3OJwAJZvKgHUY62hkXqZultX7g5ZAAyK3OQ0bW5x3XE2aQoKJUk+PBk6kF3
eA9NHRhUxd8gr1zWD4Nx+Hp+/0pZ2auJZJ85ESfGh+qkxacMdhqSwvT/Ong9bLOsYg+jTwKFZKOZ
8yROrgyGklqOC9p8JkKpG79fKEVXBvrCTFy9SIpH4wDssOc4lcllZir7YlJEP7mNff5f0QOpErY1
8L7wPdno4tugXv6pNW+SoNd2fqvtdZ1NVDaohKNM/4mPLWY0V23Uzidp6qNQJX6cWRil4WqNFtGU
uIz5ygXc1O0zuHvArTwFREusa1K/QbPR2t4rfYn3TiNaTjPCoZFlUwKPYQwJ/44mHTcTu5fbN1/x
mNevfYuF2ChlDlYMA+OpnvaZL7xZ6E/Z2iUEAhXcKciGXNABk0Iyo44h9G2O9cpmPCaFOjg7kYtm
9ADduwfrgsF6tD6NndkIEgHNfqAwkNidegy3mBSVcGvHCM+tjZ6qSxr2V0vVg5r3FJGVuDLHG+dJ
rF213Ziyx/n3UR6QKklhPioP9weOuN/mLdVWmu8fSly/rK63IDdltMNpYJF7w5n64GB96CVvFVEe
0ZVumyDt2Dd8Km8gtgSQg12268ymYsVUNTVxftcLzHvvHcD+AePGNsbRWC7oo1F24WvwGw7UaugP
bX7fSlFvawOoLP8OKuxi5favW+4hkJlBPpF7txzlEjkU0UbHypPUsRt4wTBH5sdKp7yGUF1BTfDs
So6ih1uBqy3IeI2D7PhLTPAQpbiXD+bQ7DsQ40x4M1Uf70XLzBYCuzdlWQBn783DFCYHLT5Bd3d/
r4cX8OYRsnAditpxEMletekF10uFYj5YjWZZDplJtkuMenERO4qLlEeyOfqy0NrfD2x8ftDY+6GB
ZWThg13b7tL4TCA5Scz2aYXe/9BFzG3YsmszyQntGxiQ9t80konImFAt+kvvusrGjBe67nYkXzFZ
ziUV94Dz/S+4q/Ny6uAnSpeX5I9AhLS7YyU66OH7exfpavYtDluuygcKURSQYKFDZ8VI1UNBN2M1
RmChosIVRJkhnrZDqbMHWzgQds+ZlxhRJthDFBubAK6Te3SNMEXIdFNuvKxxq7M39RumkcPWDEh9
/zAtEPUX7mHD7WYzczR/eDY9gvZ7YqdsfywcU4ESm2+rnsr40LsThnAPf8USPlmSHnBGnHJNTNIU
GDZNSzKOT2+Jth0nDtbHoZMk65i3dQAs8i8MkvlSCGnL0WxJRkHsl9dXjQVopCBYA4dkesuLAJay
kDj3znwsLzffPWwWtV3PlBKvYPH7vvqwMi3yU8Iln1ZxgLoTGV/BXFG7Ru0fC+KaytgEAQXSdID8
6eDi+gmdmw9o0f5KKvm2gC9nfCRps+2nsm7NVW+uj63Dbv+8eDiy2E/BXs/a8ov/4BVS17v9w69q
Qu0CPTXlGomOPiiKaEPY5feZi/OYjKjN+dlLS+UvbQ1FQbSOa3+fxAm9SoX/ZO6yrVkpAzKD6JfD
wDidxvYGODnRW5rPKS+r2O7Jgx/bA8x/TFKh5SfraG3ZVUQksPd9hGHoO3syKrvl1DDZSCPbYYx/
CRMdR4KPsFDE4FIm64Tlvc9OIT3/BJ9NFu7SK0zwhwLHXx+eAdSVH5LHRb/amqKV9Dhkt/nJSZTC
0HeY2vV9MPcAl2pRhqCclHYBRjjFmcQUMs7cZepYWj95D9eedQKM2kiUCDawHM4J003bBeV60HQr
pfH1n886jyjpxSh1XKxS6suSZvbop6YH/vsfAfb3Eo4pMQAuDKOXK2QxidAsJUMhL2Ud23JBj4fy
rcw3Lbc4v6VU1xADR7/ZveQJ0F27Oz9Gr3VbEfYfWJT6oh4piiMjnTy0h5GrRoJa8I8v4cLtXwBX
7H2zj0bBGoMn9QE4U99mmwtqmxO/fpnBksb8bWBkFh5yfmcxtYvhme2vPFMET6n414Q8yhn7cxLD
VzuTGCrOH8IVrmrHU1x6phUbsfqNtXPcqY4xLkXW6tQ5UJ4hdCd8B6NaS5C4MUZsww76Fexa5vv8
fwSZLSNBSVMKbgfT8qSV2scg7KAJXYvPMDG/NPY8YtJv2uxQeDbdpcIvvxPZclvdm1EUaVK+vB6h
708p3UKFyLA2tGg06iXNBRd2jKHcjSDXDgHAdKQ07lnLAsJtn7gqx4ygvHAp/86U2KCFHR+rbKTW
wlO4SMlHHrp3hB6qbuaDMvqVw7aXVGWRtzKn6BLEMiskpZdINlcSNl6cyBMSYpvH/dwWChSo8eA7
aq90v2QKW1K9zzK4SNXRk/GolHzp7NuWH0pAu1DRKk3wj8+6gsa3APEuUvDiZFzYPUyAy1E19g6a
fveV/XdAF7E09mLhNblZDTZHwovuAYKrkJU921T3uww+Qgm4LJdQN8nOP5a8kDI7O1tCmSoalODe
Io62J9bMQdsTpXThBUJfG3dGFWlDRtA4ESLVQggLmSD1QX0S7KoBhJWimmsXyg7d84BNwATL/7V/
NLj4nE2Zb783WNFikRIAuS2A7Frn8+oUUhiLle2+093cTG+G3u+PUNwgFlWEOE9mgM7z0NbHTtvi
YpbMxgBxwSw2ihQ760SSoCoyWzQ8fI9IzsjpeMETWWZMm7Qgu5BMHWiyRhL1OgIqBQPkOU1Hs/30
r84z8gg5ZRR6wft8gygXNARfvT/NO5V7wB5z26a4abjqZzTcrD/UEzVWnrCtYcMbzmB77tnkeWpu
vxL8pnsvgyEcTawy2/hcUTj4ViiZKPN6cjlO3ZRJUKMhayWcGAYplvw1CnSKbTGhjVI7KS/DX3Gb
q9qd+Uok9QN6tFDYqw8Ra/ZmrXhov2NyfN9ZcJfEQiHNGvlTFc14bhTBm92sUvbnVaZzEdKubeFy
ksJgPt2iJy8R6JKriqJr3o9ypp9ApeZbU9F0eU94QqSbSCN7J+5mtTiGM7LmUJd9UqXdcZqlJX62
p02DWerKu8+Ae9n30tOnwM+nvQAB5yVT88VF5d8FxqeA87Xnsgcp8RVY097r3tpkLy8QD1weh+D2
i7rcC0WFM0Q2cEnz/gwa7g9BK6yzFU5YDmN4nsXRPTaJetXCoUUiqvXXQjq2JS3Xnopuisu7yrzA
m25W85aR0eKnZTFiKHGjavt5QXR7F5K08ezWF5ok2JKP3EUJULnxkLf+sKg7W6bCKQKmmEa2BpDm
72vx2qrQMrZRdxbPoU4wBGqSXovsEABuZhYr2LBvMHt3DaZyQiMQQXLr+QPMFO6QerWWjGU6LjMz
gtaJy1cbdUBBcVh8WfS+8w/2H/df+gsWjWm8fnR8nOBnNV6BE4ZCxQ3Ecd6tDUfGBTiP9Tg4KDyw
UWfcB7dgSkT2l5dEHjo/55vnxahUPQv1w5LtFA/bPV5VLDQmesIRLkI8edetqjKUR5dX3MvjhWiW
8/0dcm0HAwX5mrtyNvbhqbiLSnGZguxDXo5VnoMUv8upV4jP6l5jB+T2wH8aixiIG8Q2XrcZT41y
64MJ3IfIshiMbNoLnk+gz+RBdM45UW2yoItU7y0XxVZ+0AMbldy9smj36H/xfD3d5Gtj0Lrz5N/L
TJDJYo5XJAm8MlKfccU3xuztw6bec9nyxMAmrgEhD4kG6y1edsIfoLyCPpLLctYRhzZlkSXVWjR4
LhhYRMdbQcaBB+vpcA8uHL4L507clf0yG4TAnxw91oOrpmFLoCbfTIJCpSxfXUJJ7L0Fw7Fd/Iun
sT3+odp5aIKjR4ROpTdEofcOtu0ddIXsuO/Awr2KeYK8/GQbuZDTfTh9J0M2135vp/AzlmzZrJqO
5OsJhvkEL7wgYf9XMqoRfdTyQczGY5zOOqv/9DUofP0Pk2ocbQBwZkNuxX1hTwwIvd56nKLOS/sm
uUAeWd7uV/9XPYE93ffEZM2uGHm0iVjOzcqIRPWXRfelHyRCu7eI9a8cCtOggO9EX2dkxPo7/67S
zOKvItK5SPWwotQzzYeXzxjuQbNT6gE0L/LuGDSjNz5WsPhezewGebz6SaaCwPSKK6sCW9WQnr/T
K9J+nr5/8aZzWOCpGwlqU7T1p5S2GFVsc01gWgb2gsnZloNHx6wgv+r/8i11ZoyaMw5b5PSsLoCK
ksmmgGF+nlz2s44La09CLusOrnGhx6jFpRYOdfXlsVukAqXcnROIIK2oyMVTtTetqdtL3An+cbOz
ZfSXocSxpwUBhUbpdvLErcrAkPdXd+qipU+dywT48tIdH9xyMPybN57RNZHJKtu7LGJYb1tv45iX
R8cLhvclsfdUWkM6KKkNeCDkmuHbplTCZuq5Pz4bQvYvWKXIJkFXtJ9/5+oYhH4wFkGrSpZvWMaT
SMOYys+IAblZtmeN7pZ+MJKVGfZp3lDFY8CnJqEm3u+/T2XDoWJWucLStqUHMkTzV0MbitvZ+yPa
x1e1itlXydeVFRQSPUQLlFijlDEdMNrDBqqvtlitA7nSlOTYj+BI+tRlULaBrbxPUu299XRz5Wmf
LCw2rtPt1QD+bUOvkfN6RSUIrbqksIGA0DUbgLtl7lhvKJ0QV08y3reTwPAS8JMN7jtTkX0BKO0Q
olmFedR8lBEhts+ohBD1Pv0zqavOb6aALrmget0rhqDtKUQbmfPlO+Irr3U7JkLOaxAR4LnZEvkX
Og4WmspIom7lfhbGpMxBxfhBfJ829vCp1mXOpLLNGZgdoV+q9QGf20X+6QcUTEPPBzM9HT92DK9p
01Vle6e+wKOxP+xKS9XRBASCd/7MWQPn4ewwo2OjD6Go6QpRlpMQ4XkYytFCRNgPmDZtbY0tb41s
TrnIWWMJPWi/3PNQifWsWC3qZnW80mGpIG7UlJ5nDLXsD0RBtHqZPn8V59JnCYRBu8uTG8EIKUkP
7N0sNKPZK92t9Bq7dXpKUsVFPNwugmmNe/7YsTPT3ec8FCpVaR6YVbLx4Ue0xEU5XQYCO4rapct+
jJKrY+qSMTaqjriDIOwY6CBpwXM/rGKCd3ogmlwV1lEsgdqqh45OZ2jFtwvqF9uDOkrd3mE6Xnzs
CTlz4kbMsh2lQnYVeXIGngZV+nGWQzzBJD0Hssw1iotk/EcoNLdcHSEpUTG6IqbEl0y3sKTfGD8E
xL/hPe/5ET84y/UZlETYxF6GlXyPMIbDmq9Bem9jWZgatR5bHrj05iT39D52zE6KiRy+8cAo0Yvb
h7YB7CWoVDl+xTJvEdqvrZqfnXuMeR+6zWpKm/a4Pmvqimq0qR5F45buNciqyYGLw7DVHSD46/Tj
Ck66sD/6NAOLRZWGHaTBM2qOnl5MM9AkktCTgr9RtNoNY+3WeRDmj6mKB/lMghSjAvrlDAJuZ1DB
MMM+nAMKDaxaUgHkc/1/IGrOkgIBVbC9mU1sIdpswBBp5cy5LkLxRXkK+Cq3y9+jwqA/HFg2Xl8M
awWPaAIRp8TLdO+M/hF+dxrVMKkQJ+zfPnla5N0KmZlTzfngrZk2MRPLuI6GjFTC12A2JDPFCBRO
y2yKRRDMZ7D1h32VL7qHvGUoS/sgC0E24WBtKAtt2jxuPLrEmI4b7NwEMKhYUwSA94nEjABD7h1t
fXp2883Z7DZoUmFuLYbpZJE0NwVWzS9qfthPGPgCCS9ABBR+8ACqmvhVnyTgO/zArYOHGq5Y5V0w
vXarTqVzQVtJeBlIUs5L63KorlUwHVRUXqBmU1Fxb0MrYsGEN6Qb6VJFZJ7rbj9AzN008ctQms2s
nRoie3qSXM0zsOb6rCF9jI155VmeZeFLsOFG2uwvijpH4mhIwGOw00+HuVHsTPo63NAtZ+nUXsQw
Qar6dwBwMXa7tIlfPp6E553Qd8WT96mGxS12xcpe0abAqASWqK4yt49+zFeVmwT3kv28oTMOg330
2Ls9guq5+U2WRLr+5tB+3wCnv0j6sRgM1FDZui1TMFs84DBspOEXuyZ5X1Txos4KJrgBEKIWbkve
2E5q5ZzzZpM1pm0myHlZzugpAcXtaw8bN4EIJH4qxZHt2lCpC6FJoldjfXnyhKLBCdKVZot0zEyV
Z3XN0dYPthq4YY8E3NbFbF7QVpaa+/jXE3c+mk+N1fFru5viqZrHkx0t5FdSZv5T15Pjra6ynMFd
eEZlW79fWDweXjVnNHDkIeFp0kElxU5cYIWUwL2IIXFXKvdFaKiVtRgE2v/d3Sh1hNC1E8WRpiFU
FAzyol7BdZFJTSk0vIWix277ldr04z+1TachfNjEHdqXYcyrN/t348TttwZIfkRdsDK4h0nbdX0G
mTSVAXQJGoqaHtUeiXLavJQhJqMcIJL35XsUAJFwOteBJsi08qIZNbGAukM91xl5wmc6CAOQuXyc
Ad6MtDVNcNN7mQuPyNODGIOcIduuT18ce1c2f2+1AQZPE6uDAWhu56vH1iqMqZ70gkTlkC9If8RN
DEi4OF4au5DEv5+T6B4B6M97XROL8WqZPlmMhEVr7mmpCgd6x+vsBDe1ehYnBxoOgeSEqEbonLvL
yVSJvdLgGbgmD4Z3xriNn2qT38+QnHNSWWmYNghHuC5Pl7XvWQuVgMYY+sb650XS0sghwrQ7Y7AP
LqnzwZmNY22M9zDmOA122KVg1toeftIduBoDwsi1MIa5Ct4y+sj/1IvuSH0hdV1DGHF4zY47awnI
TCAzE1FezheJr1UphAfYG0pm2X382BP36a58JyQ/WpJK1BoATyms5toNNY/Gb7ENqJKHtbJer/Iy
B+GBE5Nz3h3J9dphDJOFVa9uUopFqa0ufQlgKovHLy+zYG8xLLJoYs1hGrCgmeYkDJA2XVg2Tqnn
DcNMAqtfQNt+h3lrwWFqJfudlRyjb05p3CXnmgaoF7U4E9xhhiKzcHi62K/auKKBckuq2jmDYyJi
T3a5un85oaRcm4PcsaPmGsWuThuOhqqAzCssCV6HY/QBkRiIuutJ9/TjKyJDa8U3eTETzzEikVsX
UzYFOV47lmTbqBWyL5Z6+2Rpp9euqkYNVFY4ydEhTPnrp2aoxLr16kIO+RjHeaU2DY6ok8myXpuj
g0AQCQWNXSlf4nlglZmhiN/a1HVgJhsXyxW40JYmLqHUQgaOm/DggAKg4AYJCeNF1NnAysFv3BMn
pspjBHq21g6tVe+Dt5T677Hoi3ch9efIjbiC2G/GJsQ6aGXfoy+ynUVwp+FctA8nU7RjIIg44V3Y
PG0yZU7rGa8ZFkPTOL81vNbRdFchM7+d01oJKLr7AcK+XM0Q6qvjvRrxOmbhT5ONEzOpGg8ZtDaW
h43dIPtaeQoq7LBvcg61SBwYPiFH41HbdiqMYgIe/b5zglhI+BmXGZXK0wjYisr1Tcb8En15qtEP
qt5U3026W87qWV/9ytYOVLiuqV19QjKycr+kVTazP72d0vcvTttpBk4ZBLiKxwReqzp0qIjFYuaa
vhkeKSEE6q50FSFjQZFqVPluvSqxfdi9gICq50FEWjiTqzQuWa5sQjHwLg33ismg/L0XiIf7P0Zt
8C9fy+uCatHJlUEFmL5aAAxTiEGySTniIrvy3XJW57B1lNHkGL6fGDXw5jchhfpG1/Zk8b7kPbp2
XUfwKVzUzG5OGbwX/FjlRB6DAQIo3wjvIwPbrgGojmDoGYLb9/PC9NHtWd5VeiCPQmMHrhjQcmif
gxpBe84Y01UwL9k46gRJo4jPmoYkeksTrsIOUjyYmbfZv8omgr/86ke5kEd9i0AYcCvbwphdutOC
JIB7RQcQUoVjRJaCzJfpONYXlpf67RkDpa1+sybsxrlhg4rqzgmIfLbpIYojeP+8zmd/1z7DXGN2
P9WALOspg0P/R+RPaEejnCpqgtjWuV8yZyE+TfkEHK8G8sGh5nksyAcCEj9nZ8Pcmk6OXqmR8H/A
Dy8guE8lS3iQKiNcy0a0bKiHnS5o/Z/XZsYBT2iGJVCptqw79gwtnTURlUmvja5iplR5iBk9bRtC
6Qpk6S2kMXcFJjslY/S1wKDFokWsLSAOuRfJcSKUxY77jxW0zOf/QM6xP5uJc0qA9TCfwG+T5g6F
W8Pf522OESJVhlHGd4nhlV7jx3XDCXiyu5CLEhiBeaDnfY2VJVEkzqR0tQS2gJ2xPlIrSMTvWLdd
9Ra6KXt7bnyfnznUkEOKOcwywZBHsIPPrnUvEWnBJtJrFNdK5IzS8nenz//VrFv/NTD2y+rGQ9O9
NaiVRLpanE39hKv0+fM6dVSCDU4llup3DCB9tXyiPX9nCjuMkDk4PjACBJmMGlGKPovNN/sszCJL
WqerocRLuzIIQwbOsxIDcP/WTWK2Mj2EdjAlNpgIUe8TGLGD54qxe6GQG/a7mH64g6w5Shz5EzMF
RaRbQQRNZjJLdw1GX+5taViP7Fwwi8ygILBUDIIaX380fAOHWirt4irz8K5kOzL4GVe1MVepx5dV
kq442WA+WD3VXY4rXErNJkU/1PPGJrtPRw1mIEwx90Fd3OR9B/UJI0LRJmf6JIg4ZjyQrIyGgEk8
z1MsRFSkzdc4JHn1Vw2GNdRBhUxZ5iQCsH4Lwt9tPwVjuNdPhEk088E282bQbacxy+YJKcWOYob4
L1snxB7xecWC8W7xJeJAVkjg2YVsiUe9Da9kZJgRxLdJvz4LByrS/hWCz3Wo1rtmDlZaXB8rp8tI
mswAEGCNr7zCYQvDPTgrb47LiIEcAnY85HDtwk3haWb31jO7Mw5OSh4kfIaQkQEHNCfPwICdzuPN
o0zbIlzymOR8zE/77wCM9/GqkJtI4Ldwh/zfMHgn0hE7/aYqx9ac13SBbizCD+ue27ULR8qinhfM
jRs5WckRPxoRHIwla8KfVsuCzJwdU9nXkP5G4947KnLfXwZbWlxH6UXe6lMe7aakYP4u1+Mj7L/F
QLv9P0VdMN303Aa304ktv/Yyox5YqDUc21Wgxsi2Qt+oqBoDsjiW11QQuvzZeay/rOuhEK0wXBOp
Vcld2RhUyt0Un066LbUQJmSn5a1lAuuksG1Ytg4Ff2STxAIj98dAL3P8MNv1tT3H/LjRsTuqlVwu
tV4t/t+sSTkGhiKkpkLTjLAlEi4fVmSmRRDizsV5JSBhEEjGmPLhlWb44rkQ7uXpsidbxtkEocJ+
Zzlf8Ygdjbss/CnjVtzaVvcf82d3X4GUmDQsj2viSbtc/UNOERuRxkzVlRf112lIIK5rHI5xQYAk
Yn7DvbbQttk5fJANdcakysHMvB5s4SXFX7oizJJNyNKq0nFFd+PfZZBJpQdglxyh4rK3/VLumUwn
WCH5ZtKDmXnUMzOSeaPacxkN5zSXfaPXtAKkG0Fhpa7ZqjHovh35L3Mcp6dHhzS0/9Dk+c5oc2cd
PRK3lCUlpd9Y95pg7ozKs9QnefafD2mX4o2VcpFUC2dHVmV/9i9fWHVVs5zxOVNvKsSaBgN4Tia3
TpXi+q262tWCRF30pKhXtbjwOEI8Oz22T6+jrogzt8f48ozbLdTE1wY09jh+su9chy3CTNX4XPsJ
IRDC5JzFSm8oe7PsNnstvIFd9+/t8EzJgZ0hNulSqN2b8j9lm1SEO9izPsTkW58pe5Nw/ji9qBeE
os7QE6p2a8rMkuaSclr6rDQ207++MksrArY75Bc9FgaBGfBEfIHHk30SskMNHAI2bz3ItpPlICcP
HrwvuCuvG5PkzsOhDj5QZ4bY++sPTIQS+uymJKHkFhndXNmwvh6uRf7qRSJsSnkExSU4JKa1zZNF
CKCAonioZyLu2vClJH1yKn/bcFX++kJ6RuzO+N3yi7BxqGnVV76wipI4dVn8V4xV8i1+3CFVZKaZ
PwoLxGKc0tyLWRcPt3kiFUpe6cC0NCwY/Z3cPyQwhpUCPN0Nhan0dSD5rlDkFN7TxM+c9j2bGn53
52vyKpQsdfVKQbj2MpzZvJZ+/vnJ/5lIU3y+aNqcu+blJ/AONizi9HxpSvKR9kExMx4UYGiHeJUP
pONhDEjTpsHjvGEXnlzTisBxv+w2JcFmkr4fe/Fw3de3BlIwuf1I8GfG5qdvsb4fv54sUKU0ULqk
tTfU51YaR2Tgdf9JOhY2nsMyzN5d0gYGMKzWl8XaBjGwdNj/TNtRSKlKzWrUmSBik4oxeVUftXZP
PzhTMCpvYkEUBytpirLqS2bJByKMtRzJIppWXHuGl8AEuX4VcN4W6/z+2+K9IHno0ACLgXZvTm3C
tmsc796SzDG7v56GuIsKmkn8IoAh+jUTB/O5idJqzIxuQ7A5Fl6cxORMAkUb+0e5P62wI6sP2AU8
SeOPosW/4UKInpd4lgZjMhIW0cy5P2fuaHpp6mSqvs72tyeH12MlFmST657iIdy1H+1dOYx3rgJp
nNLlFrR3TOD//NTcZHPXAIE67I/dms1nJicat6WO7Tc1qRlXgsgAUC1frfzgILDU50ZoLlDbXBJu
7blCYowGcDH1Sq0167LRd/NTGRA/Dh8UjKERCRT8MoR5XO/kOmOYEZVrhzC5NnFwvFl6tt2GU9B/
igZO8FBo1BCD1DV2EodB+ix9cYh2SEHb15ID5htKAiRMReMAIv+6+lSmJhLSYHoViQx8MaPMaF28
SRzcNWuC+cvgOIQQ93/ESJfBIlqg28wba9DW8foEDIeMvOzfO/A7cBuoAgdXeugB3T6ceS9pDzE+
fvJHDnb8nTupKkbuhgouQKLXMpIpchKXBeQBSUTmlcAiyHbgctxbkbVr+1K7RsZZkdH7vwfUL4fU
JlHqikpyOJ/HnUAtvsUX9cU0KkjcveMCJvghEJwrBcdIa20SvBe0Nx2taSfUaf+wMy8oCYK/my3y
LwWiRIsIAM+2EusKmopVo2BeE8pkpZQPlG4XKQf/R+p6Gq2DSHqyRHTVGk+myoCk3mQMIOUoJiPR
EYg5mP1N/6xZKyVhxr0g5TGbTLGxRutU8Qoiw6SEMmDkdxBhJfMOOv1M4iizwPPN+fJLuJTDFCqv
j4q8vJNiYnKVdcUjS/rZBmIKqqG8JPMfIGyVzvZS3hynn6F8jjt49Bqz4+6YlmoPfELK+TUAx7gX
sD/6ALWOwd7Bds3xqX2pu4TrK6oSzyfC5pY0lBbeZ9Ny9k8r6xnKB6TzyZooeiaYkGbk4zJN9DNe
287pQfw5j33J0t9ZWdSgNCmAVz77bQNHaYf5rT68OHk+SK7ChfVA32PGcxhR0q3svlDOYa9xPJN+
H606KAbFpeHCsvbIejXTAyvbfQfH/wFbTdvzOZSW9+JyLV/W/DlaF570yw8CFO9/3iWYFQckWNUA
No5YeeHh9hZkFWfxi/Tm60ShAb57ARze1V8PnONjTXoZNQ6HTHcOhtPwKfU+QcPeHa9P7Mr/o/tE
85gq4jKBasagLeE7YUlPl7Dogl6jl2W4dnBRCt7t0Rz09eKGd4cyQkmJbx+Y1Bn86quCeR3XudPN
Zq80+3PeIwVpnZeEvotxb3j+hOLAcn5YHLSI8sdY9gU9Fe3thX5Yz5IghX79ntQ4JGmz29yEno0M
LJ7niNEPbrWHIqU99M2qyvkZancXRZlvL9LGp0nsQe+kcRSMipOpLt3P3PcjiexCI6iYcpbE8GYW
C+klxy3vnCI/l5a+al9U1XVYa6Qp2eBFirDWAscMdUV8ZNVMkAy/M7fEDc4TngKKPY5TWcH8exM8
OvAy8cgPNYfr1P6B6ODYZOtQeNathbZ4oBao261f7/VW5RHhdkEsCRGAL6HbC/KbYgTH3OUulvOT
dYEklUZNIssb1zh4xUU+gWsF9N0SK06+7xY7AgbFr6enh6EaMxaqYRa3HlLyR7nr0ciYMEziFy2c
mlcXtRKUWgkWkw7Sl2v64viOn7C3G9Hsc+61QSP0UyXPxaqcMNh6kV/QGRUJBJ7HbtmPb6ye1Nb6
evQvtVSlqZ6jQfHXmaE905OBWm0oRmMSQMWM9jR9xKbMTYwVduSsZOuMKZ2XW6FEh6X/M8GMRjC/
2z4c4G3JVYyfZNUGMLeF/sPUcWMFMEECJS8SHrCiGP+pMc3Kh5FIseKht6QuuVm3EdnZ9aGdwivc
4/kEbgJTe43iSAohgw89IEBrS4TjcxVMHP60xcrNuCfbz92VSZrQ4GnD6L9ZZFVmMVq2fihKbhJR
036n1zsGvr1R3NKNa8XK3++30dXb0uMkLCqdM5poW0vGIgWlNUILjDhLqlq6OgRyd+CDv1ACeuhm
n6K9RqmWF/IhT0Ojw06nTAfy8Ey5WgFopPOmx//C8Wl2NRJI54UZIpth4wz7/FO7L5Rlc1FNzJVR
u0Ufz6tKz3E4FiWSh2rxegjhJbRMtXxfzTpVnhX4ZD26TBewN+9HX6rlVQKTASBpK6BWcmHJIIzl
M4QZ1by58jK8VkCiCXvnx65vWZ/pFzwGfnOaixPpzhccs3KISWlnmhSvD+Y7Kcudb+7hNCs1jFI0
HlDw6OBr6t5J7tJZPlPmkT50kiwxBJGJ74Cgg2wtj8zVHCIoSUufKx24G5gP6gS0IKNHLbbNLuuI
4+Tgfl24RAlY2j0+N1v73cMFPvXU8/pZftjr9PM4VRiTyahW1oD7+zg9yNI/zOd7Wr97Ue4wJWF/
gHJXmBSjmo/+TrtLSJh0TEppEa1UkWE6tLj990MWO9eCy+jET4CFskVejS2hD5qQBpRgA/NqJZ/p
+ZX+cOyPMC2FTQsJdK2wE7Jx7hH+TCZkPDSrPIR0dTFhmKGnMswXxyX1qcDUUUZzUhEg/nXuP8T6
LdfdSxxDzZyBVZwBbuC9INqP8bwoR+Ud8GwzJkUp9D6oLlkiH2u+WT42x7O/mHmkLI24nwN/CUAc
i1aFFLyLvjzEtrm8ojeBwrs6VHHMPB/BHESmpgqvHGNXtn+H+/nK9QYovZfORApufrbb3Qwb+6i4
j+kMu2qla0VCmVwzUxXriHzvfI4jvLCg1Txdhj2rf/0TFXQSYM9lkIjxqw/OM0UNhescMqJmKPyt
abGbaEnKYY+984yqaCSI1LHHVRzyuPK4QVB9H6JcB3e/PFkTEYgN3Sc4ZOphD50IXA69w+wwwXKr
rXCAyWIIm107V0Ty6FChb3+vhFc8MWHJVifUydcqP5EPsali7elEvWVpypkRa/9CPrgWHcwMUgKh
TYkdomesLN271nTxOnNH9zNdnDQdLW8aKxGxPE+N/A4s2g/a315Nz4sl6SdW57/e+bTs2UsR96o2
hWw5TvQ4TvBfYTgMCflQ2+p+N21q+UmCD9YTYieHNST883yF/JgNLAslGyx+IFvSEYMAcR5uriDM
BcUFvWrCckpAJDF5eAAsdpX4NvZzs+rPuaHKXLsBX8DptDj4NqzRDsHDNDmST33x1611j91c02j1
NH7zkvRDyYWxNbyh+jdLH7M6UMKwZiLsYRA27r6vsdmkOB7knjwUn7upoB4aYZgDtqdQ9jTAMw0Y
GOG4d1KJ/+JBZeNPYDQFZkG3/KfKge2VOLKmCcUqJGr0iN8tHvXif8iRWAjxqf9w/d/vSxci/4Bl
tOqq6ed8BVIu2PrK7/wO+CwlcslOrPRM2g23mliyk+JuPbN2WrPGft4IqQxHd3v1Tna4Ig3H7+oB
sbk/Q4pWf0Zl84Oo2RqrNi/Jb9Ret6WjrmCZRjz+fCL6KP1EizEZHQtXf55Cwk3dsiMJsLLLh10a
cZVqvyun6HIsLgIiVpmdwzknSrtHv2vVAox2WP4GvMvB5Fq+kqYIieojkYKYGwc9kCZ10JdpsESY
JDgbMHXsMbNLp05TrTJjUE4kAvJrCrqPEiOkEwCOWPo6iGUz7kREfnNU8ybuy5s9fCpj5QYuOhax
B8ygZtxEBYnYFutP+pcqoGyULolK/nX9V61dYWIPuf0+n1feXM2ey8m7POy+EJ3CkyavOeOSMl7b
s+V24bs5qm09iCdQiMpiFqWyBgc+CC7cU/4P2Brm0iu/4yH0ukv7RQyxzHApPD3xd5JmR+5d72y9
dQWiqs1tk2qpn78MiFRBw8GzySDHut+mXmFXQQ3nJu/JPEt8hDvvBDyRumJBwm9iVUhzvTU8INz9
lUHg43peXZpxMafTCxjsFGVd1/GwD9rHwecXVqQSJK874NwMrn80wb0JbFH/IbDFGILaA+YzMd+Y
Y1hY1Bqc67tpF64cIlM8HtLMIzi79kADnWQ/Prvw9uoBDb6hSD3CoouD5u3Y9i51Kz1lPVtlR+JY
bmNUyAuOox4JiZZE0bHC58qUJyaa6T+M6loldyYcngUUOf7eyIdVLlqk2th2TbOJAn0n5ZZl+6Sr
E1xCDfjlh5mCi4JTheBsiTSTaVq2W9skD6tvINyn9ZK3ZwCg6Hunc2f5e0sU4uPJnELK7UDn+Nsz
Dc+VlhXodsUCe7L5DBPAzGNpNbzjrSJ70ZcNpNJYihqd0FzhY2uCl3kTSbGGWnjvftC2SzW/NEpJ
+QC8Mcs8tdyv0j5VKIbLgMwzdq1V4zjGCXj67okIUNZ5rvdOTqM8Z97aBq+tBxRjSkF2MNX6WMpc
1txYhnTmw0o8SqEr3aXYuSioZwtJ4PJ28YF2qcd1GxqNDJmE5HpQjrbCxA9NT6DdrbfcFHaZKcam
QUOdm541wlXmJ2RqxhI1c8ODEDh7iBzcWmj9jh8A0jlCAPHXODDv/BJNYKRzs62yVzVtbuPTMeJP
Q5RzETsT+x5IMD6ILl4Ih76TY2F2aUE5gB3Sb2Xs1i9ZQAUdq8CcbpZo82CiDSiLKRZ7saagjR1l
KbTzl8VkiBN5/4F/GczONz/GFNgIvJ3OGu5N7P4/vv0XYJkfxMv8iTV2A52a9zNXLvr7KUEzjC9q
k36Qg/Ec59yYb8yXmVdVHYWRiNOU90UV/KjWtwsUD40R6s28Fm2Xivl7X8q9smN3ODnF02pbKtwI
iT/pAi+pUd9yUVuo1DVM6plckRo62xGaiTxxfasgei3lqKY2pIZGU6ms6Wn2AqsbQHSyCewcqkbd
d3u0bHjGFKZwfcX7W+Rf0gYWYDxgT4lez454Wcmi+L0izxHI7T7bFLh5+fTl+hGCDkDFLM3bwl2U
b1ZS5RhHTnaKRWhELQws+PqUPIzJLxeKGlEOUEPvAmxfhaD5HRGnU+q/FpgBI1HSppeL4dXMGuWX
aniqZVlhmCe9tryWwohaNM2JexoTS6yEjHeePnrIyxhLK4REqMummv6JjIOAx8Q2S773uptWFFIZ
ovVQqdZjcXC0EGA5mblCCP3pzR/TzUo+yWuVcrZd2xOMb0W6XoB5YmJbuRudOmJBnFxKy7X+zs46
PJjVECJm0ZQTnVPOnyJW/PRwHuYYPzwbjei9JR7iwO4BzsnYtFOPu9i7BYHUgXbNe8+7sHAmITMN
f+Y1oG6DoAP4p04i+2YTsEHiOVc6zCE6yGxblvBFfn25ppSvpQ/6tC635XUk904wFKe+jPkoPSzG
Azvpr0c2+Wsql89JqyOG1iu+nU+3MSAgYVKCK3hJAwfCbbUtqAV+0SPo8WMw/LMZnQ29zEdS3eHi
miWkzAAw7v8M1QlCTLJU32SyLkUGom+lIrDIw4FXttmfb7179D/S2h3qFA6g9M33/TUcYKq/46t3
Z+POU3vOv+54/H+vJE5jVWSKwVCKyUrMRkpemjtVfjanRBs0Qu6KIAB7dwpnMxjzMIoaY7oJTqNg
p7qQJOHTv01Deprdbxi8YyKXv0Ugo2i2BXYF6Gm4c6pn9SuE0algVjsGo1g/bZnTts1O3hW63yEu
9wC11IimCa0y8Bsz0iMw1Xy0H9Z3bGlHrA1yIIca9QyqrgbsXoPFCKPLduzFnqm46dZMPZYkrLcd
GSPIYU9afDuce3JLjT8cv+o+3LOD/2uKEUv6UW7f7PRGqWyJNTGho7G8HCMqmxzXjErBlXXuKAgo
cGl2VnaAPcCt+K0gk8UGQ+w7sMqmiVUd/yZ2uTKPkiwfgv56eKAoXrEwcaDseNGPsILsjYw0CSSS
0RRwSymsVQaL99mGA3Qafb+l/DPXTjSP5TCaUf4Sxqa6ShFIjT81NS2b7iA5DQ1Ytuhz2Dqenp2S
MwYskmjBQnndPF70z/gQUY3czRGi3W5AKUQbC1YXo9wUBtu7qPxlQjgaYSmszABYPyyMDdVJmwDl
AK2mCytNCkhceGWLtweME+1XGZGYyu161fBD/2xuDp4D75DcahP0GxVT8ohNKN6xOu37qmk1Rid7
9+P2pX55RvFm06N3qHgu5o79RBiwmo06ywlO6rq2s5n4A3Z1D0LRTaEAXDHHzBRPh3XlOohEGpQh
fe7iWBy6xjLvSG5GR1T1hb0kWTui8PF9KND0JRjFwjYX6ScO8bSuuX8H/mQmLnqJSQ/GiwJWnWJy
HoelK2ix09lh9DpR0Cl6zFVRUigElmm6uvfU53b8c6pWJvYL2a+Hi4CwmeFMNIPd8/wu+EHF7VP+
tpkkzSA7rcZNMo1KXC5PcpIiKwU/JX3nKlkWfGvSAFA2XitKO7RHf+66w5ouyWP5QW8DfWbMrKPY
ViM2wDoXf/DUL/6Hut4BB6auoZALi1SYzPiGWNcrpoxPhznzh4+b8f1FM67hLOnmI7bEjP6GjPbR
LMHfrjrzADlnMEw8AhMilkZAqPLJxfD0MHVZSmq5eP5rigr+tynWHZcE43iCiQuemNWfpKisRWSX
4X2RmxgvorixG+VEmXvsq89HZHC4XXfYRht7x7pDkOx/o9XVF4Sqp4o4ASVdhTvcyL3+b8Ey74fx
q44QHJi7Cz7HewBD22QwFQwdC/hgbPpTJz3VT0oGnrRVFoI3wIhR9C/txEqrRPLHm/uV4guArI3z
KGJwgmhvlx8ziL3/qZ7SK6tNdTEmD0y6jocnB4WF+BpghitakqdtlFkVC7CbE6M5Ut20HY+OWJCI
ji/M85Yy2J5CciTJ0IY+29qGZJyClUCJcJie/PV3+8TRJeWcjQsQufpd8NL/TTUobhR3CgcCSKgb
Jp2o+r2CxEoAL/h8p8qmx5zbd1ipMv5YBW9hJQArDTDu3oti8cF+fAG5Us7stHgnVpBdI8OakWou
lNfaPik/hL8L5zLIP+mKe/HAi01RNz43Y6RfQlHLJWAJuIwdbfYEkxOV+vs8p34I5RlCLdCHpQw8
K5xL6G37cCWaVma85PI5C39qa9xFPv2+88LlnPrJojkLGWtSI+JBWQO1doDOJ7rvPpLUyD73G9fg
a3BwO/2SAMfHbvFhUcvArQNrwBpQXZF3qMKqGyn5y/LjAzyT/rHBWl9bLtxjGw1CQPpiJS23n3fp
ZaJocbAiSBY+/B+tlJgkeyi74dCSHor8XmJPpafdPWWBf6oFshEnq/GGHMfjDDZjaSdHU6G/vQyw
8yRc0HHlpstMJy+z9NosWBuChhqdgyEmrV84hGsxfCcHgpD1Eiuij8donSie7jtcgKFyPRwNndsa
oO2VgEW/2Ur0B7SwoKt1pl7nQAvsgcMIu3QWo4pFe+DKfWQQngXdktoQxMTVMziPxT+DlxcgQRok
vD3Wv6PPc2aQuTUCb5IWAbG0s2g+vBlW9zxSaaINBv9WcKi51aHiy72fd2WHJKLqVrQMM4mqLLv2
qbBrPiEmk7KpMPMFfTv74A7DVH+KOVWYJKIk6bCpgF3NKpyeI0vWppDopojv3xZjRwduohrv9GkD
3TFncsG57lRAOoxXeMaiYLRqRJ8/P5pOFJ0TshOcQdKgR4177aFbSlotpTcQYu0+lR/PhyZ/RD0c
HaWdcxMV3ARTc20i9lWxQsm9QVN2Z2DDtJaY3ZxHookvMlUsBnWEdQrD5HBoD6ZpZjUR7eMTMnHR
m+Zzef4TivYPbhNLuXXgl81up0BLgtYZ2SzoqrwBw9P5hG5gydvgrRqaSK9KIvPHfuibPuntKl01
ThHJJ/zOD+gqc0E0cC9BmX0GJAsKcmKXUkNpzswcKxuXsr6CLkiwVK9UjQ4SVBEA9jmTqPo2yx0F
KqVX1+0sqvWjulznkfOC5V5D5xR1xOHHRWsdm7lSerXl9e5c6f3jkKAweZPQrTUW+/ehyEYUxTf2
o6k57ihiRnuTXtlUdFKLUG6gAT74wz4+3kOxG/sz0dsA47LBBSA800Dlu7ghWVaQ5SbHWYjoeoMm
L1Po2kpNFDqnyTMndO6LwGIOne+ONF6E7Z9V7UMSZju6kUyt2l/AHIFgl6EtA0OoTXyXEjztL4t7
vT0mzDzQgysToFgVMKG+1tddMJS+zhhsNYA1S+9VZ8sG6KqSt7O3z1ZouIedHAfGVXi2GwDl5xdk
HS26PdDl/GM2cd8xUB+1MMrbnmodIG1p2dhA377bUQ1rkEGW1btqmT7EtxjbUDwESOKQ6o2CwR+z
h/L+qk0WD3A6o6wkPyO7frI6wOoEIE45UHUyYqHj3sxuCMpNc5BZpr5ViY3etoAaQaZYoPr57WtI
kJkfJW881dQO+d6mbb03rQajYrM+zo/PbJO67GyRd9QfzYGMnbtfv4+0EET9RzL3Al4vexFIYi/9
xD0UkDKQCQB6uwXjMtfS0D3CJjfyIrddeJVlOU7X1SBNuU9kRe0ENO7Rk94sGl4EKKW5pMRINvjz
7u90yL0Qvw0rasb2bb73fMkc1PS3lu9bkHfZksVrAuLdPNGABfQr+KkHrKafaB8TxODwifStJYz6
4VVv7udjVzBClChDFqOWOGeDbOCUTGf6wY+ALLzX2pi0yWsv1ywQiHVyRPJiSKvpbcm1W7FiiLMC
gJX9rtuWGGHF+dqXZV+JBUBlFUKeEga19cBzBP9Lji5jiuUKiOr6RNw60Rif7OA+UNa1ceTRg0E2
tAPP1K63+hD0JswDlu9kqtfiHscZw+ITW9ja1yPTiZOp8VnMml6pQDxSrzoZRd+A9mI85kMrQrFk
Yb82Q8T0ISJWhJSYamTCysG0Odg++lrHRdzVkp5C5gO0l2bGdaxednuPsy7eX8IMjQ2tmF5vj1AU
gBjcZB+sn8pyEN/t/NMpgVbTjZxjtfh/nco2p3VVAw2UpTunwGRDxh3mkb16ZqctnTNUWGH406nb
1+VKpt4ral+cKYrr/mlKmclWoEz3a1OyPF49HprhOg8LIpoMjwPQH8ito5WJ80xKt7/Hh6eETfEi
uNRs3+OvFI+pelFpNLiCKn5ES5e3kFJIUHwDvNyIgmsoeord3zxdUDyklJCg+PMBV3qYYclm2PDg
/l8dZIawkftbKg2vAShhrxYAxTi1mT81u7lg8gY4+PKmhrKBT45cZyjhSYPuP+jNSKxGD6kWfeHA
XsbVLTu7uGObOomqL3l3CotZ7rimNqBlAPxP36ybauqETCPq5nyDufL29XjC2c6dom3do++acYNQ
KcXWLfoG+sKG1Bau2h66XfT/aKnPfD8RQlwU6QmBpbzYXyneimUYJ7O6AG9cabgTsNyWmkxpLlPr
zSVkMLiz9goPecpxDfhqHPAlWY0mnfZUA0gZaqA/OGpTGe9I59htF4jehc/Zsvnlh1dyMpoR71MB
R7h5oP50in1Rf7Zg7gNHCD7a7ie+ZD+xRZ5MtVm+OvQYLb1K6ayXlVo6PDvLzF+rthcFAdQlqrST
Mnl9iUvtv9cZGkmWu1BWv3RAaD9AqzpXvZ9hZ9e7e99h/Dl4F4d4Cf67dbeq776+KWBeh+2RMO6+
Q4g9/+Bi1qHvSet1qmr1MAhrbOr8NusKLgw9Eb2w7MXLLLaC2i02agzBYhY5VCd9Vuzxl5ozuhup
fiYb4uJtzRDB4W7vAf8SMdIckC4tzTK5F454xX4AkL2WRwiRT0xseb60qnwywBz2i24i9K9ncFYA
T0hqs6mVocWodg28aBjy6swewj8qdmi6Hpebh/cndYUXZPewvBynqDzDLc6vW5GgxcjuV8oyla3C
68SXm8PkSYqW22G9UNLylbgbQqKPRnSuN/GGeK8yTd5bxNzu7DRepNT3qIzdogNZA83XaFmKzf/k
+fTHar56+Jis0aZpY7cFWNMGBIuR0C41cuOX2CWemQpYr8asb9wXGzexnkR2Aru6JOAJEKDIhFtH
SwSizJdl0JLZvnuQhtPAw+joH9TpI37S0egcR3SFpgZGOk+SY2BEsX1AkraE5ss2QBNpJBbsQgwl
sSaim1kmKvnxWtIvzyJM+1Q5/wW5N+PzJDH/+q1SAMvy5ZB9mHZGI7UPWuWrbkiFoFGqh10bgOWn
saqouhgR/F8Va2TtLD7y//RJpYhnj6FzSOnYCqYOvx/K5hWPjypVPEJJTrQ66EZC9aUf/3sFtcqQ
zGgTMxMoVSmT/AYOsvEwNUxaEubwg2I+awUs74L9caekKX9VYGe+yIHFIEq4mTJYgrzyOQ2weMUP
YvF93bYaI3wwj8lLM9qQ1K8D8wQt94wV3inARN7l/ZwwlfM16wAMzuYEyNCILNJJfxy1RPn1eLfc
dcmCTzvSM85XqoUjEg1WBUIOIHrEiEURbRKUS9AQTIqxceegV5YkG4UZ9hWEqLart4sUxXac5FKc
UGq3qBrRhPhvT/QEIQMiZRWK3oPoZWHhwHNRXafXTYQSCEd2XAA8zJfH71piAz52/y+CFktW3Mjh
Dps6Z9AVWsLijDKNn0kbYjUGmSPv1JUShr+4MXwCdYVfokWrZ9a4nhS8fwawVC3uIvpa/Pz5S4y1
tjvJQgf8fwtMiH+IsZzSAwy4ncjV9HpZsFi/t8YNssSIRuX/VVq/R/8TBa+hIP/00OXZTJMbBa1F
7UD+FuDSS6hZMq30tFIUdl+DaJP3ZZHILzcnwR6Z9Om4VnHviKZvaZcUH7tP7EkDn8bUAlP49YMY
xozaQGARohIhCDrJzzBOJY2XAHRMO+dkc12yLeE8XWJjYZ2bWHeDzYQ6FZbRK5bxSM+qPC0GYO48
2ia6lxGpneRG6wNSaZZ3luHS6AGSVT4F1DTQuFiw3NU6nV9vTa9pNY4LSAB1aNJ9pYFwCqCAaYba
o+E8ZydmgafK+KuKGeIBIUL9mkLosKBz+SZ9JZpZGV45v7IUTigw2HbrRpdptY9Ox8Sfc5EX73KY
oHykLBbhEcHdjuujVWiJx0a+VgzSZNwjy0CEPk1mBF0dqasSWXSxRCGBmyrcjrz7Zxdgg+pkdaQL
q0Is+I3h7OZkoSmrgpgaRzaHb3d3NbOPo4x49BO2yYWhPNv12qe9yYFvb3OnprdjLj/wvJ6P927i
OfvBD45xfQ5YRifA7pttkpNPtpVPXfcbl3psqe4SzcY5XcaW4qiX25JxKoR//iMTAyamfECq1n6z
ahRcM7Pf86DO1NaVwDl5Vs5tavOzYaDr5YWmUs+XqydZ0EQG0P/MEhbhSxYPeNmvkGKm149t3hV/
KHa3fv0jboCcVKxU3BA76p/tr8xIFQ5dsGe5N2VwTbgocKzf9oM3rFTa9hRnf1NHuBDXCWlXeRru
fPgFDfqT3CDyU5DXIb3oDT0956gINFYNF3TcungXQB/ErsgdXWf8XPO56yOYe/RlseXZbTucGxgI
3jbOmdLZlIonb8HExGWrN410HvBG+YBDY9n6W45q0ueCCKzuV/wskIRb58tNSD6L/XkXtcwYdf28
QlXLzOhK7oh5Ju1bfdgvqB2cEhTd+6kLEHFWLmTuIoSWeWFxq0Grnkm/hszPc6o9VQqK/CV7Q4in
lWAeDhGehrHdXvR3n+hFhn4lTDPChcO4Nt79ezIXdX4onBUTBzkiUpZilmnQ3IH4JoLdzxInzV+o
X2CPw6/j19sn4BLM47P5lF6+bV9AVaylWajPqzz8mvV56rztT9satudGe83+/YpKPDtwRE3cZeRS
ukSSZOPOjHsCTDU0pUVkJdCVfDkDla8PvPNRdf30e+5ccdSu+sE1AryBltuFURx8tsSqMoeI7wTQ
pYMpZ6FpG0+ySyVDz6hqOOzARP86T2LWjnpV0qZE1TXuzlvS8KqITwHeIGrPHIdHyA8Qf1tBF/iy
HQN7dNclQMnXuGP7GCR+iOT2fJzMTTKKQjnW0i8eEm/O0t/qFREc2QjHmmBPt04sYtyuvqws040v
uUqrPYWM5fKpK6XEMnQD7VxrID06KshAVE2DE7E6VSeGFXLZNJ6gN+XmXC0EppAAPpyuslJRgK4H
QJ2oSHb+4Ux+OyZfU61C05tDcEbjWZu9c466ncEvpF6CLmpZTpBklMZpT0oJfDpl7N42v013PlgR
Yg9fzmoE6G2Gkn5CS/JWel+4kiU1pYwt18aM/H0z2MfqukGIAvUGQMQp0o1wNCOVHI1gPCdMF9On
xukGxwXnxCgZhTNmxOI5hn2f8wmVqQBLMIprzEkxEpFbfsIlXVMH4AfGDyo2FAmE0R0BKoxLQ3V2
w9fb5DZWqMDsQiy3WF1E6r5FyzBJLXRQdkClHZJuWoJKUjR85OF+TVmMmvShs/dxYzR/dMFqnSXU
rIv/CXVwZ+d/T/BAhMrbfUJzdTp1T86Ad2q5hkp0J7rD+k6Sqrk/vkTCufTMKKSoDD6VFb+F6POD
mNS1s8U5+rEPH3WrtNWEVy87LMb7YDZ2HCdgOyIWGAkiAW6ZdIG0QJn0E9Cw18f4wTz5eCOX7ZkO
/mQOkjbjxsWy9KFagugOB09BaS+p30vyHAjR4yjSUMVk1ZhU/OGNAoRUkKm5gFYMpeQUy4GcOB8g
JWLnEUTUgj/6bjjTQyjZTuYAT3DZtX3MsVsNOgtbPyBxqr9ihCnHl5/qgB4HOtHEBYl+vc9YkL0H
y68vVvFTX4QOaMFB9oth9QgeYU7lrfxPc5e0X+bnj29xYpaG5sMi8sZPVWni7rGaEu0dL9wDbdnw
KWeI5pUaGtSIQNzx+2Y+V4rF0iJefT4bib2wQ7icLDwdoW9sudlK6zmOIJi456Sw3NRdVncfJxxO
Tp7mDNs/QTmLymVwQCdJRGQV+A1Gw+JBZFD3WIg/5nZqDX4BYrrx+PdhW4sqO06PpHiivhTnPcUw
Av/FkrRmYWgmZQZCQ1ekUoRkM3cLCM7iczNIxAz+WhIsL7CIpjJmn4yh7R6KRpc5MBVYanIKjZVD
c+KBt4yVasIlFX17nzN+3/aybLqPYY0E/T4KlJCg8OvRR65VHDZLwiOwcwpnXZxWACJ/izrtPPPZ
KJVeGCLRz+gl1qx/TAtJSlCxSxNJAE1arYmmq1shNB4ADUY3Bc+cqzqFW16fqaV/8X4pjKZpobiP
fephUn9UEFXc5kq4RG8lkgy9dqrXcdUZruday+mbEn4ADiFa/Uv9+8uSkFMGjO96X2mf2LmZLMq6
JbqVDmZ6lFa6vweJtrUiMc2eRAEuEHJcS8k00hlJ0GLoNilPZsatInvaI2twzzorBe+lJN2rYLv2
W8lcZlPZlG/+NBF0G5cun79nzTg5bBUTj+6o4/0vFB+Cgci+iCyGrLaWJiasGq3C3ngjibuBmcX2
w020aJjPAo9+CtpfpaDCHtPF7XsvdOTcN/N+hMmESNjSWxCkA45GwyMw+tLFQ+jchDu/ljdbKcDs
37B81Powmav8in8kz/A9CQgfWji2cYxGMeOHHv3ulO1bhLGaK6rszWJON4inGKemiIydc/v3O6lO
i574iyReN15zj9vUHl1WqwmIvvvuoGd8NNdBpOHr+b3lGUdOBeCFMok9/3rRhKt55y6O6D95m2+6
A7c+OXG+3OV/VFB2hK2pWQ7a1rr9EjkgoB/r4w8YGtYT7kPatSn47hMRtKmL3qdRN9mryUPbDfLY
uFIMgYWyqmN6NLnZ9rc+M1Dq6k067UM3wSnlo5/uXz+nhn4qXH6R8k+Bm4BEmeFH4HbOTAiDsT7i
hZcjvijY253f6oOBv1nS+fI9IbqhTmaQji5E3lmr4dVZzGJbU2u/1me9JM6oKnym6fU8vflBc8Yd
y+ghXbTkIohs08nmH2gzx1jW+y7xHoQCT42ljfHFtwFCfUW6QR5CEI5JPo/Q4hREVWLp9TDEMZJQ
9+E47DGyaxbsG39cFlNAw4D9Rmgi1zqah/X3CPnjKQkoa2FgiJoINrj+7szWa1hL6eOVk+wXPH7S
DIude2spwEJaT14TTjQ3UGVaFv5aLEMXv7fu6Ui59SWxscZitvxUv69Aao8ltuRnF5/WxAPC5UYa
cmD/VKTqnmt7o1DIZfEa+VS1eKFAIxEWw1eiwLyRMsxP/xglB3K3wEwRhrUSfWiqn5SLQtYzKIUo
nit2d4y0PCeXtlktZR4wBj9sMxPVmc9lFgtApWJC7O7qHalKwWB2WH9JuX5sSTTGBK3IO+Oh8y/+
XpV6s2nE0zXFsrvUb9xsPFXvwS4jxtr3Z+KwxA//y/2LK7edgZ7VKPr5mOclCzwB04IZ+kfpT+jt
l3+JzNYSYHbNelxldhcTe6T2X8juNeFZToJqtS1G8ZyQL8rqhIMAdozFnK2AeT63nVQEFCU9547Q
JvFoiNvdfdH9/bE5yvSI3++/wrSHfeHMVghHKzG/Sgg/RYzaLgu0fzF2zPbGHFhAvbX3FJuwosGs
2BdPgr5TtEqKLdXmA7LaMtxZa0aLbo6qYHNGJunGPj+B3YZW/6by6KFLC98tk/2E1AjbfQANpYAJ
9T1BV3Thjnwa24yOa3V5vwKrsUkUzsM+8T7s/0bkNQ90RZTDi/lFa8ZkuPLqXtrf5kt/+JOXmEdG
fkDBYdOYCZcwPcXStFvX1OejOrKTT8jrAAFih5hR3iPRUHTlBkvqfPcitll9enIc0OXMAnY9ZMEl
3juuOVplmAPhGGNZsb7NMGkN6X3HjLaMYScYbJI2ImcCpilaupFnEdCDf4NI9Rbw0CwShzKAGGsD
YptHyBhpiPwFO/CYNzRDsYuTPKDI6NukLyV0RGmK7WoBl8Kxe/eMKKquTXboWYqSLBG1pNBxXIPM
M4k4W71VSYg+HAut8Dcedq3u9MbePGd0x2FE/dZb1fB76v3v4kzko4WGevVBuOThE4svcuTdNtRG
gZn3ASlT7nzZjoQnRLnn9/Bra5wbAiZ1EmEqdArZMGl0aMsMzbkROBavL7ZTwM9Z4jvnlBPNxraN
mlj9SSU+2mIMLagTf7tMXh6aWb5YDxF2edF8Gid0Bbx/d4RE9X1wv8dVo+7qHJczxTKHqIyoW+BU
uoVvFxycwo4ai9RE+O9kMv3eAXBtUyzDzrDjJ7oCUq2JPDlHcZc7Gd1subv8ZL3aT1gVYOr+lyfK
GVCh+vM96p1nZnKoTalWVoymWyfW5cOB5rX1gs8ET+4YMfm0K3rorC/f0qCRjOhzZG4KZu3O8GxA
YFPisubZBAozYtt2fXHbWB3Z5wvotzXxwEKwwBw52skm7MIUXcho7xAzqnfqIGirRqDzb+awv0g9
4NCHv0Xg0k2T1joJMJ0LiaCpV7acjIPZFuBNqq2UGujFcN1zUyatFVVjDxFcnwU7JK98KU3LRJEY
XS6KGDGc4Lx+XbOZl1hO2/fE8HWqAc/7qtNbRWxfRyCgHP5xMnB64NW+Qt227RlqQ3IPdPxnX/vh
LZDW3PsrxNh+CszPNlLqSarM1PMwNdwOAoX0R1PsVWQu1zZfm1lvtY1jvAYy2AK8QFx5xB1+x0ed
YUnfTfBSxO1Eft4acuamq6HwqVn/5k3GGBS8NSBXb81cxjfuC/2fU2dxZV35plVmgiTX2jiXXps9
zweffR1AYNM5Hxb3BX+n2Ol2CxfoRwhwodQrG03OwiIYw32LqS7FaT1zF7p+IY87E90yEb+zCviF
/mkm3nV7Xr4yPnxAofAVWk0ayhF5Dxlut8E7N8AlqTmJxebYI9f+/on0XCMwTnDdX+O80Z2tlJoI
YMU97+PY/ey6nl2Jfj0qczzCLOq25vhehXtANGnAdhQFeMc8vesiD3Pa6q8uXLgR3ijALR+BDn4t
c5TKgDiYGrsWcDJvsIV19VeQFb/1XTwObmKKGI5YzcuxymXTeOK0SUNxTneAIMR0anN/QY324R6w
OHJennSf/w5jkhyZvuCbvYgqf8A4yCTxMdSe2u3b9M6rUvkliMlIOATxLcQq7is9BC5B3xFY7+Mo
Zhi6n/U+/9btWefTglZ7fHGPzUMeCj+5U1+HBrwcEncJ5NSciAK0sTAg0rksBDSKyNKDKhhAHJPP
IKdGmIee+kFTu1Fonmvu5acGgAZSavViHpYoYJGRJJrzAJCvCzYj3AnL/WNQp8o3gM0rjyaaTPHL
ORo/QlpkjTE9xNMP5M11y52kZOymCm17rfbvsQskcY38XMkr80hoWtyYLtXQIBVIn7uzgY2bGJ4s
Fn6na7ykUA5Fi0IQELJVrTJeFTda3alU25xt8gY2z3VUD9fArAUWC8yIzRB2pKVqWgiBTPJVZFzJ
+oJe9M/nSbfGB//Kr9DsJPP8ldDmChTXRLkJLFQ59gs/RJ5dkPn/VYYSpQFTbydaarosxjdEesCh
76GYDOTNtPEl3LpAktsBC0nvLu9sWI5baPSq5A92y2TBpQgdmmxcyQYU4zzN7bFFXKxjuNj7Idit
TFavjlTQ7RyWq5vrCpNplihn/Vv8JD5D2n8Ni0Bx4YrSg7n3Sc+glKaWvF3NyFSoM+DC2xbWpcFm
rJQij47g9xFanwLkRKKbNRYtLM+R5ftWH54+MqAa0SK/9MpuW3VKK08/3MY/n3PoUzG2oyyONMGb
BE2e+71xEvPF9WDKoTe3mBIfoClnDo9VcpEVtwwhjkIuX1JWMV8kFovEsMAJ7t9UVlaVSZZUk0F1
VnkXsXehY/kUUwDpNUZKJKXKyH2RKhtO4lNPbu374kXwQH6yQEHqIw9h3arlk5wdQKFyKKd24221
/8won4bQbLa5XB46E9jOjfM6q/rl7rkH+YvxdrY4CB0bEX+QE/E9UAyLIudUVA/3fTAdZecprSR9
dloXGbiOFJtWeutPRQ7SdB7PxLB6XLWulKK+HTp0YTJMpdjeO46A9wjJQLaqFdxFjaTqoXHk9iY+
gezTOUGwNXxOzlOZenGcnz1xgIQ0jIMpnlwv39wVy3d3X1yTOhNpZEN2xD9+bmvZDQV+8e0c1co9
FTXxKs1KlskTNzISk3jI4HK+yQFfFQxxrTWzsArU1CKcSgyNsH4R66J2K1aISCgNo4EkN0ACAxUy
Cm3Y4K2ll57He3UArjHXRmGuPiy4srcQEdDuJmD28jiuH13ZWAJJp5a2brcLIX+EAb6nBl1VGWyX
P+bKuD+dNjJvfn0p82nPhSRXOLn3VA6pcvWLipJxpnWhdu5/RVJWw3RCI/waqbH45Wjo3Sv5Iarn
F17lK2IIycZfGzSkvmyUd65dVhEoCIcxvRuQFB/yjwOpXgzoaVReuBhrOjw/aOHB0TsyxuSfywBh
K7a0VFR0c5h6RLHDBYA0rsWy+4ouheN5C2zeod+1JyZVqb5Oq9LnRJSsRxypv7l01OTebRLmyQSy
PbxtPEw2BxyFvg84KBx0NzOFNYuhxLbHJ6sovOykp2yuXnL+E1RFSEFo72tnrAf7cU7k+JuCrx5P
WVWB0HL+SEFWsz5wV/VhV+/HSGhHLB4jpTx0zOPfhuUqTDQfQ8jgchSewJgtsKAGK6hBq+/gUdji
gre463YgW+5hTfmfI8EyZ2MjrctugOOHdne7+eZE6hfkH052b5E3cTEUFC7XDV4m7kWz5VWQ3XZH
mUCVFVKkL4E/Jg+YvAbEMkzz/s1TYNdotUFj9yaSYlNrDtqBAaBxBYQiXS7e0X8Mil1Spv2YpbWK
xwfP2ogGGzE9p4fXCOeaZfruPPTCix+j1rv78xZbOgSfpsgMMsWSb/LHTtxiiPk7J2wWU8kApKPV
2zJyZzzaA++pzzA+GOoNuWd4xOHntmeaU8gYZkRR3eYY4D5I7CzDnwEdxBe1cbd685i3WcxkAmCe
8ee+q+1D1eL9DJB9hqW8Ch45+pBci7rzKa2OGVbU2ldg7uWmtpVnSomzot5S2KmCL84yWFDfKW8P
dKOjeIGRx64/3oHI1TBkW1QTsKJtL5RgW9XcCG7H//dvN70ANFZqOExNwfY5PKm/YW4jIip6q+pP
tVCeo8WCyzV4OQMZq14e3B+mKwVQYGKOXEiP70dDR3V3Awbr5jB+zFDyHyqF274psHRv39BXtgXC
3LMRM+9Ji3uxt5C23abu5GmfdoTkpga6KtGF6hrDmy9EfmJjb437OhnlnEiu9JZddtXm1gEeLkEI
2homwWhWWZnlZ0DZwmbDAzHH14vpY0ESu/BqQC9MZtGIMDBHsh529+lXnTkf8x5WjmyGe1ZWx1Y+
rlumLwPm1zJc8cMGHIcF5jMbpHJVRgmsCJhS0YQ4fPlGEt11hfbnfxjLHwi3zicFjnUS9DmTAJO7
mabj9krOiYd0tuEeisLYnONhXL759cqdF4xguXAqWJKf02z/IwwTWEfDHySIwLms63NfcHgbr3ST
HfwQlc9/iLwwlzm0H/tUuyplLK5idNwNJ7VjgleepOaOR7uHfsXM0xe1/mXBr3vCbto0Dkn612PI
B9NHQbyD1ZF7EnW1/8e7lfQnlRShbIZiM+4pn7Qdhmnf+ObJTM+r5vHTkH6FguEcFcMPtswzlFBi
lm8uLXFgTtTdpIf7ga5W+ICnoo6x0XR0M2Ek82eRdkmnEEXEjy+gdZOOUVFuRSB4hXZ2mqaxHLv3
lPDkhGBIQvuDx4OpYWW8m2gIRQIcseDjEft2A3BTlBMIE24erBtj8da4eSXRiM3E7HPmaMDrYoUM
NDJLFkg5I4eNy4VHnx1v9sEPZuUYO2I39idGmTGJA7AiKcE6E3/224rSoRe1i3ZM/B068TRvAmA6
sJdzWqKNhc7qGV8pQRHazyZcrCQ/qoK5ZKLvr/s/8eyPyRhM/V/Q6UFuSxwdsNXW2K8qrUohmKiX
kwtfdlffZKSjysOdq4Wa1343Ob2nGLNu8IBFxNLn7ehPu0qE7eY9Zkdie2E8JMXm5uUqkfCnM5KJ
3jyF4AWc6vAkLN0NDKDl8mjIiL6B0d827z6B5KPp5GuD482/MQsOiZTXDz/EYf6ajXXEJLpSUxDn
PAL1+eYduN6owQALMEE0OIfLDvGdQ+m5D4RBKDy163yw/ZPzvOwSXbCOz+gxPwOIHCGOWaUXd8Pe
UcjbrK8FIn1S6gki4T0WpeEODdBbLADcOoGdIIIRp9aTWB2McqsqwGCqJPxtYEf+zBat2GrJetqM
wd2Q71Vw3kRqg1AGIioLsEeQii9uRCq+GPjiWQNBPHvuMBfY3WWAfG1th+zJevxyWPs4yboVnS3P
2sBlITro6firYAVi3FN3/9z6kqZ8t1hCsjT4Kn8LA4zaiZaTBpe95cYSs6tmKBuMstcqR9siuzko
XJUCaINRUq9YAqRNpUHBJ9T/lOcbFJdW3oHcfO1LJyGy7qJLHLcZ1Q0mYG/hbH5Eu7P3044WeOcp
nlH9Cgeq7paZnZlPH8YMHjAi4lJUCxLfxeHAdzbO1zTuG3xmudKm5f+HNTjfmCDYWDf2uS2+PtcU
O3SyXfM0zD9O2LLAQ0xvMKVMVJNa/WmY5JXTfMds1TMw74l0yhm+D6tD6q8KLB0Kr8h3+rpZfkrJ
CIwQ7ctUs/qB11w02HKy2JKWG6ZeKTPtCmRYsCnUuKcWKejmRJjlx3PDGcLJf5i/dI1I2Fv2+LZX
UVOxFU+Su6ncEE6J80O6y3bJC19e7EjDGdCBF/W455wYUfSoMrWRGEoOlrk3iPJ0hk6eM+EH53O2
Av8Avsko0RcFxRvuf4wFP8k+3OEENDTVr5yArCmx5sVHa6f+VhbN/zRq4SzZRd6G9VMxqejcz4zR
ty+Qt31P00NhwXs8RSDa70FHO3fhwidzmiN8RgAYPkl5rvkXJDiltXDZUCgeVe0gREtwzzjJvqJH
A2bE3HEMTbXRq0GkyI1sPZp3Etk0NanDJVZyDzBQGpZs5elQf140B+lUKqdTZWcxPPxHwRg7V2dY
CMXSRqnoZ9/p9Qz+N1OY5ZaPe5XBqzbpF9zbkN41gLLOpX4dAkIpv1Ae8OhYE4xZUXo2zYWAjunr
zawiEhacsqDALkdBAH/bh/8r33VpSgzWxR53Qv1Nk+DDcGUZjrBmjVk+2r/k1YOAEWgkRQgVApZA
EE3ly9HG1hFKjeqywXRTk5QXDYkchFxELUpJeOYqnOB1omIgPj8lI4+Db4oPSVa/q0tG2eqdU15r
lXshEFRWFWaaFMVzo3eVubDhGmmiLHpjsOqarR0ccZ8hAlKcWF/WHWSaA9E6folKBCXcwGPgpo8b
F05jvoBl97/VXYBf0hZxjiCxF2khygWw07niDLkkFWTGxhUWzuRrRt8SlZPNHTRnVI0PCtqRAHP3
0X6cwQF6six+f8CJr61LD6A/lVBZDz70dvN/EexQd4OlVG4W33bLoFb0oKD6v+VAyd9Bv5aeJSpR
4GesyRt8VqzXmMcuNLVhysniICSduwpaPGZEi47W+s6/im/gRWkZ0pSNsQKGMAkdt8mMM8ABR5T7
y4UbwLNP1h+Ny5z0z29GZ636zMMFfyOgcDzXPyjbzx3XSlL3BISm2SswyyZraoVlFTWD7XNiRU+e
8/TBibRfsMRf/U7A3QtcP5sx7dKMZSqBUnhLGR3CA9NOVEYYOd6FDmsMiDpg2J9mGXxORc9eAaQn
64VbfWUjpsIh0cwbD0vlZJI9tGOHh7e+Ga11JEBX2Q6ykdBsxMUc9q7zNRXMe0v0qPRNVAr3V5dp
la7JaGjPnI7SF7WlNKelov9wjidmL75ZFsSxDco0a66hob3n+e7SbkD/Iwyf0TS1CmNu5C322MtO
n5XLRWMkyJLkMY+328hGLrACYOoYXAyzmFdOu2nUSn9r2fv5k1mcD0PlMmQHxzW4e0eeBWdTiBuW
l+cbAWdNc7sOSQksnrCzp8iZ4snKVra2tB+JifwtMqI7qIQ3k+4ajY0AWOJQGpnPIyJ/qANksIs4
z61TKPdc87AKn2gbuqgitL942Sz8Rsuq9ezADRnO7Q+NM5dcIBfG2wM06WxIqOWDivO7kX+uiLHm
8MCV+BBG5B7ChIQP+JmOoT54HnNgl/KElXnjFuK810tnj8fnSPkjx/fPEFM=
`protect end_protected
