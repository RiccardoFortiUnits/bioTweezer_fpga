`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ck1ZmGSBUd5ARbhJ1fbI3ZlVS8FWXVqSI6/EaghMo4JptHa9BbqlwxWhTSg+f9/C
D5q1Liwz1ynxzyJkQch622wg/2JRyYAyvQZxqzZSjGODpxfCLaCRYGNT5rfsstAV
d5jgUyM+8rE74aVzvDFV+t8acyfCeKrbr7NivmcJgTA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22480)
+Ul44JytZZIucbKMKoJye9+zwqX6XXJrZ+n/PQxYOTnHzLqQG9SGe6rZSmnWVkB1
F/LGVk7fl+CAjIp9ueurmXvPn3d713feA9fFmx9+8JZVgT4sHP/HJnqBBCALgVGK
iy/EgDyrcrFro0bAC4k/Ue6tD53BVT+6qCQ4jZEhFIpsgFIlsDrQw+nc2b7Pf/r6
QxToZyNhWya8/PfqXDUC7AdexSOve6loG5DU22E6o+bV7ZQVCX2twnd+TXiJTnNx
wbpZlQY6MTZPRPzbkxkpI5HziMvH2jjnjLV5WyMTSAVU2T8bz4b0epy/E2SVscZc
tQzwy9nuoaUGL+mCM9lb7PzkxFeV6hohFp2LdQz2QaA37RfSWShmdcdA8X4JcCYY
COT/XY2CoFro6yjiBJ5muB4C55hKsjRHajdJGR97+X4rj0cJcFURyC4vPMAnAyLM
f4pZquja0EeAUTWHx5zQzjymDD1br39xL82AyRTbdxM/RvJsneEMZP/HlJeFZSe/
x352pTo6vNGYp0sp8ItO1aUNl/lY7z62TG3DKv78hhdyMfE0HyH8WwtMaBUHQ1tB
xQc1zBlYrrAjw/78rE6gQ2cE3ERBefVdRBR1XZcMR0tZMYjV0bkgKKwBQb5pPEbI
w20pzBWOz+bh10zancdDfRykUwNuu15ctUSni5nbcT7Y+Tr7Rq6xecc1UsQaxkXY
a4qV04BjKjWpacddRvy2thS1pEZeLveB8N/3ICz1YCsXCivHq4j1uvhaLgE7UYAl
iqLbhDb0Ca3+4SXOG58FJ2bai/wi8RIxNu2At/RBBH9lpFiFfcV9oMVeuBCE2P7D
WQ0UOvBknXXqQa15m0nqMjb/yGWcSYGEQUHZoleFgcHI5vxmw4CV3keqbnoaRGJA
p/sQAJS/kdo9bh3RhucuXRmOu/DvS82HtZNLT1yhjZDi46Yuj6U3gbEIOseedn2/
KBqjt5h8lH8T4G1JXGY1pqs3beoFbFcOLAO4498xxh4VHunnTGEGwi0ucKNXJX0a
x7dXincnskTHUZBrPCtQJDp9i0gNhGAHfBgpJwe1CIh3fOLAzLM52EU/edGT39fo
/V0YoOD93dQuvyuPldEmmCCTaIwP97ZpYeIyj+F6u7vt4tjSdMBzQGhzzx41/Qea
RN/gxGUDN1v0ELNszkG1g23aiJXUOCp7yr9hfzm8XjFIaM2OTxNwS/zJgDsYihDg
qaZ0KEM2riNQLISSq36RyZanesrlU6JJpEW++NHYv8FZwcL9P7cOVQPDd4Hm10HH
JEc+N9vC4nfLzDH0QLxB7Ya9LabczwlwfEIz32xBsuXRXPbObfFIm3/y+GEXiZfV
P1kaCso2X6GuavFEEoyvgzIbiN6KekIXJpww6mT+CKWmpASnEkinfgjqGHCgyGwy
MnnTt726eJMW+rfl6VIHimUbCijIYzUMUveJXgUiwgIFhUMD2oqmtaLK1eP6Wz0W
Gi3ijYldeD/U0juBFSuI4PAkEKsltdYS0/8dIXJLCCSo7Mo0mdGpSQ8ukzeEWLgk
h37fdCGAufC59Um6eYDnLl/+gq0KDy4oYSK9KRfqMXkTW/vWAQafcIIVZSIL9kf6
HTWMQkcAhGePPrkHLVEM/AOenxgdfd5Ej193zX2BrvBrrDULzxYkAyQk+Ca2oQx8
QpFk+6rXB5B7d3xdSrATLHjL+Y7xh0s9VHkYCdnmyntnWZ22Q7WvKoCbOQG0BGBc
W3fHeV4hbikyudNCW+ifEKM7eFntxhwi3hZhdNfwRrmB6e3jEnr0xDMHz2ABqFEX
Dzhll95cYpeAaR7JTigotIm19mIgqmqaiBgrfxoLWHLHNzmTDDpEJtVLN5nSQa9G
I/j5Q7LQ5TuYE9gCcvt1MmjfrRtqfdGWoVNsr65MHsoZGbjszNDDsiXF5bErCeey
ehWjTTueSzKwvaavqI172Na1YvGUsnNZXTP/3sMGyOA+paxpCRCTgREL4I1E5L6a
PpF732Em5QV0vNO+L6twvAf17UQjdc/hCbZoq2F9TRdh1qaeeZ61YhjLzgnbjVUO
SAVn/4u/7n1l7QjxrZg8eMLsH2j7lf9j4qhgPBrSylB9vaIkyeq1mWvMenXXej5w
IOIe4fnP9HpNRMwEJZuP+NMC0nsBX79ygDiaJW+19c6QR0E2Pf1LmQcn2Tn9JfK9
/i6M2vygErfANNNstFd0svKX9MnTS1LPRwtG04OpIG8LBcZNz3MyN+VFo5DlRgfO
+jKbDgtd3JP5HTmqjgMfrOkfnvmKhHAbeEgi/PXeV+gL91bhyGmWU9HbxEzRUlkG
Vba+kh363fqAWy4E4whyDr5n2uB9xg9O84o1K6iWyXbfRkzAKvYgvCo/m/NlxA8D
0BCudyUbYJadPVOGvJUBySKzteD9XtwiovxBc27R6CN2UdbUa6Ege+1aPFpmsf8b
Ja2Fh4L+QdbVvp5uI2IScQ5h03ELvcQpWMP4Awi0iP5zM6jfBn7D9cBehHRdxpyF
qwVqoWrcEVdtC+y5ZH9RxtQ7EzNZw01GAWE93rnAUYPNj1e86jWQbFVc3XKEfb1B
0jJ/zMkPl6IS27PWXXTnwIYHXoLPIbnlipgZkuAtbdAim/iOL16ApVBCc+DGzZYK
fSjLx0+GmuGcPbOYVORMtnX8GeTMKCSQ7BHBOJ17JervaMxfuP4TNRakKfytr51w
iKUq+Xctg6baQg37xL0ihRxcJ4zXu2NsqGzCZ/q0rr056Aj7ck3UAGUHPzNfJDjM
VurMIx6rYuDsyPOKY/3RU3BK0+7vmfGS0c1xggrj0rMEro+4pGR7f+3yijB62Xpq
8vv1AZPzpkKUXY8QwiLGb2froig4L7AO2525JF/zUJMducmCx4ch0Igr/7LZyhiO
naMU85WMiC73fwA0ogNH37HI0nrcxo1TtgBVcNPuW3UYGbOTWitN5YC+1oHqgtRm
TgX6N/002eJFhBq9zeypO3wxhr+FbNGcu4VGoxGn/9rMxR/OQNzNCRP77LNJmrOI
wiNN7enjJvWmuKeXtFDzkViEr4UxIebGLN6FVj/PWR6ZK0wQlGicz+9UZD+lhrBG
1be4ZL+hdScDW/lsU9rRckMUf14aszovygh1POf0bbR7uTA/jaU0dhBg4efBgH0s
KhKBMfv8lQ6WFzGNWRC2FIBu2GG5Cqo8sosYCwhqpBs7VdFZHWmaewG2Vc4rfRbs
aRvuT/UNa3pmlWr3w0CdFO8JEmu2GjT+7fGQ0zT01du32+tb5I5OXULyDPTZMrPk
T0GBP8NMUAF7/HGw35uPH5wLW4vUuItPrwn5foClAxScXrQEVIqJDXGTaRXlqKgK
jRH/UTaI2nQrGcJeR26P8XGHsgZ6pVFCr0XQslmzCTClC55s7Re/lm4hP05A4cbS
QocseKImqtCEtNvSE1rUAaN4kTn0rCWVwekKYpDlFZpbiqj4f7jE6k2Ud08OiJ0E
tnsSPUTFYuyWlXhUXl+WBoXEhlfplkQGFMM9d2Vjh3aqLSRQU0yYn+wHeBVurTMs
2hXgLxPwUM9wFEQNsQhvbcKG0frGb4Rd39BkX20ad2PEOuu0mY+Bdrdyf30X1FJ6
WsgM6owO5tewTSl07IpvgDcvtPgI4Ml72ab4tClD6GbEO5SJudbGl63wFqVb1wKI
jHsDjmkS4s6e6XE8U+FojQotjJZxC0njBT5c+9gyngLuGB/vTqZy6F43gB+EYlxk
iNTmi/oC3ntWv76a8UzEwqnBlcbpLM4FjwBE0p3coLzm+uAom6dvpsaNx5fRhX9O
X2fpaT11TmTc+D0/BM9Vv9RPEfDqBKzmtDDLHwuXJU6FhG7fzPlac1i09zA6tQ7J
7i5DJCHs7A/4ztTXaD/FwzXwPfQAmdmDfYjer7iFTSePaZpCEdDGOzcA/ZCgiHz0
oYmTl+aEukCh/9AG2odHDmMiMxLGIJZcAMUvQdvQQImR7m5yyIqKUXtdvQBwEVKm
rYa++VSnyb+LI/4nmAFEF+ydwIthSifc82Fdc6DCqLh8DJA9CJ6cJiSjaOWSOhU+
d32/4UnYrnEnPERCTSjC9RCkkrhvClfr4qjczc+s4i4P2hJPAq6k6ESpSPIwEFPd
n7E5eEOPnfQoqanKSfwt22jvDfrNK6BZ5+A4G0DFI6fk43guz8O4pC627g0EhTNn
XA+8TMuwGVFD6e1xp3ks23pfNvPcKDnMfIrRkgm/3iBzBXudkxgkqvnlrMdT08lV
yMSA04F1LBMbCAzIhiqIPzTXTD69cyRAhmK9FiNmIB2X7EtO7sVK8cmnDET5IzUO
DJ7K4BrwLVmaCi0jDe0ztdoYrQFt687uLWPtmuFdiuz2ZZfpREUFTQwvT7xxC7Ny
Oirb/OI6idF5FjCd+fJ8uYiXiKV8GdGhqtZENWolZVBxpvf5lCvruToFu0jVkFi4
GhM1IauxLJn3IVckfSB6xWtWHzejMDN1kFYMqDAUSHgd/DMSaNnFeA5ZW/bZjX02
ZR24zVBQBkEXmCDY9kC/DibRfaQ4khHWRBYFZlCJioq56n4n6ZgaY5cchqzE0JIx
1vgIF8Dy1azSlvIFxj4YoMqeNBS666Dpj7t3cZvtRQ1XObGPlRbPAJPvErAjIBy2
19JKKSLbuKWuLmeqkAVgAMV/natdYECW6KiyQZAz7Pbkh4WeyieGMFlkAHFvoOxP
y77sdoUT8WX058KtpCF2AZT9S5N/4I9yQX4aJScmX6deW5UbpvthrFKzJV358UsC
KtKx8eGonZe3aY2Ury1j2PldjILN0+4991ClBWCqjCPBRXjjuC2i/qRTC6iFcw+7
K49Q2TuH+nxIkxKxTK3b9RFpVe65jebeGWyfvDfPCb6WIxRE51lBBDKAr10YVrEz
mgCXh+XEhiyYu1lT3DC/icFRxqV0xyiRFNCId8d3d5KUF8xZByVrNIOJBbTXEEoh
MMjWx8i3JLtc1e5xMSqIoWgQ8rCVbjdaB8n5+spYNTHEnS3D/vmEeHV8XZFhxpUA
pFV55DJXNhEm67nVs5Ta6aH9cOZ9CRiAm068Odu3IulsnuD3bDMNWnpkgEQhAti9
IQRhlDahTWjbzCqt0vKB8rOYLCGmzdYn5gVNkoBWxY5jk3kDU0dTekV+gI2/+VS7
jtOEKhTLtGNXe8E1MI+WjwF/kNQEAeY2aPfniNfvcH2SjYblvy5JYXZ39Vof+1mx
n1+yKardGEmAMemBkFY3KESPWr8pvA2nqfw2vVss5QGWC0t/HBmE0b232hYM8Mt7
UXVRAknvatS0q9nZBy166rhnUD6MTBpLQtqr0+YwdrE9LFcuBfsMfdPJ9A5bRwJ/
fuS31Ktz3u7sSm+HHHKq9LFJexwaAhG4EnAam0POAMBc6daLicFRUpUrdRJd/kTz
IcLbEfprZRFcN78ZtL388/6hfmm8m7XTbK9c2oc9UnLIcmlryMe5LekhBtqoPYFE
inf1dR0smIpnPX6XLSgSem9D4BliIDGBoyhZHRmV3xm6XnLqtEjWu7mw8LaCEYC3
TFLKo/IExto6JVzbl3G0aP6OB3M+Ik9VC3h9BKW1ZhuYGWRXiOId6XnoJ2YTB/xo
eglVfDuB1UBZU5T+XJ+ieZUvEqWGw4cPj7YJm5GBy+b0hAg2Czr2B6A7UNEBPzs5
LxGBu7ZGKkU8+S625A/K7WFh/Ls1jvQSoTErV1CvMhNgkuyybiUOPNY4s93X/Aof
xJig07WbSOkjiRiv1LID35KLOgG6uu2WQY/qoLWUvT6YEezp2mvC88OW1NiMhYi1
oWmo2/+DL8bPoQjy7Khxnj5v0iBNZBFyt5llYGE0deLRLR7KsiZ3lh7cyYpLtoLz
1WRRntg2gafbHnfFb95/rSVGegmtxZUDCq01B8lSPy+DVCYtDbbavVhSRm5HYWku
KLrp39LRUBNtvIJs7tWD2eXe+ZMcc7NSm+KZY9ipcAG0TgGIlf24I0HVc50kj126
luqtXN+v3Fxz9MIU2DQjto9P5FiRe76BgATobRE4EXB/QRxixzu+SoWe30/COnc/
79b1hSOSaRQln7vvJ/xer2tbDE0yYUvTej8iY7DrX1EamMywmWcnHgjUQzDcLegz
kUt56Bs+4Stg07dHv7jDgjOmH+s/mt0EIzpiO5MDmvU6FEo31B7mdTQop/6MfXte
bkimKGiTAP4C6wWp9u+I3yCGAZFX0A5NWujAYvrX2orRbVDrlz18cT6VjVit4nN4
Ixu+INfF6JavfnP8olqF0Ue/8XXnii09E0C7vrJHUov564Dkv4lV8UgLFeFTbsFl
5+bLN9Ni7vjqZ5G+7qWSw9tUSOxklmFouz3VbL6Yado4C38BpVh6NMG1J6VbeWnj
w81OMawmOSw4Gxwaw4aCGmwSHPFZCnMqcKHJfVBPhRsfbZaQZtkNFNXKhFkH5ljg
ImRXgq5zmYg+0uaLWfdSQOBKONCSkcJwOt3uUyBBTrqHq9qLX4ZjgcyFQ1s20m5C
sKvTm7bu6RLWRNR03COnesgg2BHET82aBhFwyE7NreW3QMKGhe+av+4N//p2VSmD
PgKwgqGI0TmOTOgHkg4WZLTqCC2ardBmZf0/UDWXldxerAzRqhur1dvffxvRRVlE
5PYtrPJ7sh+0zRPlXcB4jLaWOHGvAH+tbVzFlhyzXLHD6aNLIhyBkqZFNw+wTWHC
kSk7WHwX1bKbeGYlrpmc+iKfop4t4Zif1dJTEsKzjU/bg7R4EisQCurf02hnLCQ9
R1lmPh2kZbHuSQgQ4lOUoTRBUrM3qj0yF2JZ3p5LwL7M+y6AfCii3mM5UgRNtGx1
ymQHtrjcuIKcgoj46iMtgKC3wNi97LhTJPROfchHJomkdxxA3qaZnhEYRTjbHHVh
6g44jAI1WXL4Ba+dwUy/+vFs8xurk8nOUn2SkNbCa6DPBTc5QIYO8tXcC8rFovg3
0TM69g+TsiWwjFYcoR/nnq9fUopKb/fdN6RKKRO+n2k3q6LbF/Zxwbv0ji82jm/D
G4K8D84RIKuWMML/eyHKquSjfON60aL8YGHKPbFT0UDG5lgOU5iLB08UcRgr7Nu8
u/JGqGZDVxBgrqdhJwRJxd+SObLPSc/DpdUvHzOWPQteHRUjlNrp+4BG9NnJByQk
ER+LXHJEQobukDabk8LwwycN5hn3kNDwgw2Qd8BXb8MCnFBqG7Wt9HE3CVDAqFz5
nUtRQRV3FBNvTbxbomchnpnToERh5+hkemSWIJf7w0kEf++/XsnMuRftDlaQ8M0Z
CoMW2eKBJ6wJ/fUnKlGEGORi+dh7PwawNffb61G23hiSILUWmC/ZfxEE0bSEcgrp
2ByXkYOsM2NWwwhSaEHVW57DKVHlYkan3KALEy9R5SJh/WJsZ9l9J1fjatOj5nli
Y0QvjdwnvHRVKk4hHky5b4GhBvB4NG33mPdIV5TmYeA9F/EisO2E38lByDdGerPp
AS47QqWo2UCN9X38sC8drymHBq5XQ36VDougJEk15n911H5Dk2SCweXtQt44w/JT
GkIw5oUvA+bVHyP7LmvX7q7OcEgea/rJVotsOr6Vomc8LWwC+gJNtej8YHjfCJcG
/SJuXpkTJO7vrAU/BRZiS3Z5ekGgpxXJYFuKL0vTm/keltx7+MSWnx/oXvcpv8Z1
BFXd2dW1ydY8OqD8Qy9w6NAfZHQLK+YdJMb7Mtgr4VlwLMKXOt7RSocokqqVPMyI
CK+s+McBPzqWXuyXXbTzSlYtJoquQpsRXtQNUYDWb6VL3n3ZYzoar+f0X3CO60vg
bGKhjLOe+e1wYa8XinwdEnAN0e4y7n9dG/0MbtCwIywrf4Xaxfl8g5Jg/OZeHoRp
vlQmDhbE1TbThDenW9EQDC78Wh5vAjxZza0oFqyyLVWR+V6OjgAEkZpktZs8bT5l
3Y6swGgf148wxdEPHY5yXSTwU3cXMq1DIDpkpX/Ovo+Jeg1AheA3y+yVufDceq3k
Rj2iq7lN/S/1zj+9Q2FQJKzJ5+zYI1tc5rBtPaxG/sOyWXMNV55YsKLgs/ERoruD
our/UqbQ5+8KaNcZSnxcHxElywPVDLJPU+J2xFA5jeWaMclZo8jAlT/or1dfn7ju
ybFWIuNUDuK+ddo2fed1M8Zh+aw8P6pOWZunH1bOgfBfpTLn1BksDILVndMVHRW4
nEgxHqQFUq+RA1pBENZAYajDqR4wZKHgl9Hy/ykFaULKbn68sCFcYMwtTE7NO+Gg
s5tMJ5LBHSa1bRFDDCl4uoFVJoTF9w46DlAZ8BzsQ7a6CZ4kGFnjrU5C/oBPojC/
y/WeTA6HYHa76FPsys59vWFwiLh3pKwDFAjwjrE8MVNsUZnFldUupu9NCn5U49bx
z+X9JGfRFDDFWVZ910mcyIJUFbyy2E8pOwNOxQOVce9AsmxM4AgjVyuY8VTP7IUb
CF6zcpWjhOf1yd2Z1ecBI/zK47EpmYR1q6gTR2IyarP5Og0m3zCWd+yR94TKuS+h
B7AuaeOtNajngr12e8bklv2H7mcXL+j0V9eUnfEnZjuN0KVuBjJnG+WanH/dp1j5
CiAymWQcD+Vl7QrHXS4sqE2uw2+u2dgmOL/CjR/CMDLFkcfoIMKSeguECHspuk75
A/BDyPC9pGjv5YzdJ/X5XDaz4PdigeNoWeZUkW3y13//nVPw2d5uAyVB2MVc6OGW
62v/8HO4tqDG+EHDG7ETi8S0OT3a7XgUjYZjWwb4jY6lsAQS+u+j9BcDMVzBBNub
+PIDfR2WOckWi258LPI9zf7Kh2yTp0AGGX+jNAtXQY5ortx93q81o6fXSrwa+eVw
kltf+9grlr1ibNjuYq8lZamspO5TviWIaZ2vRNUKyjfB7OM9zQroM/TyXAvycBZS
oKAwSljYLuj/AKhW1autiP4Qqxi4uo+tOkOdi9AKnA/kKboR34GyxpX1j/nnhBjT
dFNdMoRUfz9InQKLvo3mOvD133tQu2olGxXl5jbauFvCN818nf2g4Va+k7xlGl7G
Mk0dT4aicLI4EmSqmDt253F7wcIsGJ0lCD3dkaSaNIMV8xujtNp+9JoyVEKNm1Av
TETD4rR6N7AMsobEZdrxK7h0uPnXVOXpVG7RntobEtFYE2r+bZlyggnHS8YBIV3S
nMhmcDod8WmeNlTsdu48F0aMKclgKl8YoiinoiSihCvYQJUYLzRqDSWEbZn/K2B5
qSzCSd4bIAo/776572KQxPQ6//BJQAeO2rbtqBtC17QTUxSP2/Q8dEao61VdccsM
EUVadaU08zeJLxixUieF59gkyqH2omLAbBCsdy1OwmQoY/JXIKZhsSdXReRGChUN
UMM/wOd2ldw3mmXuKsQnjrbaAT/hqr1JWYQ8MOlHS//Z/xoe8CgpZToQM1wQ6VQ8
tcWBpSgfLQI7OMq5rmetQbi5EaqqpPtExZ6W1B7s/2RA9AohVpY8NF6bwlmB7xnF
OLTuK160+vaUsRQ0SGUIn/AXuBcmkzk12jlZGzKKI5ggy3Ws7/aqtvYwtigyRHP8
CSgp/rEzd/TeN+n2Qyvnbkoq4z20WNeAzidKefOU+D8IASdxJZVr3/x5AsKgUu8Y
vfooDPN5od5JJfH5XnCsVxnSB0ucjZWmnmTI3y2K6irCH7GIDIBcgFrmgcUjD3ir
B9i/N6ujQmahNbSepTD9n0H05DafiFC6XTt+/+uqb1Fsq01i9r+V0zlvBTkC/5F/
2jLolH/znQluwK5GXrIrJb7gV4jWPMSaDIbwoaq7mjb3XgUS7EIUZGFMmGb8rDDt
S1W2ewDjzupGwqUgxkV28llLSVgA1aq22PuZ/7OS8sfCLw6/Zmxas9PPgFF20GZx
GraurzGtqh/9nDSz+PfPSmiie39U/JM0s39CVuVZZvQtRqVJ0BbeikBc/sVa9CPc
MMWAL8ncTA+43byk1VXfHJA9RqFzPueSEWnuyWwOdjh6qSgRxHtbhL3fPGtkvTf4
5swRblX/mz2eNwvQ9FMzWLjscAt1+n2ri6Aihhz1J875tCqfbgoqMQdL8x6rgZGt
roJ2L/v1MTCSZjB4kU0ux7tS0Hl8J2UIyur+hfgVE3+BE3zsk3q9mzO0EKHTcVmw
EmbVZqtm9nAr0tZqGWgbsRFOjRzCfga9VtD4X6noKdL1Xob4qSKsSY1SLVVvbbjY
vkxXDrOccFtE244J6DTJ9PKyigFCx9whxvzWubawXywHEO0YreijB5hDRQcvcSXW
E2/d+I4vJCejodI+asyLO/Ka85FV47vBXwCy72cFXO2JeeB1ihKt7x1XrMFOQjs8
3JCcuJBKUd35kruXWLjK3Ru2tjVMocM1AezsQucKL5FpJ42FMl2lTA1bfAl4Vqgj
0CZwlQtQ40UkiBq2h/xpB9ZMwFiookmVHxFjHIPpUutusJY18VPxqsjEf5/co8xb
FxFKKJz1wP9+4K+ymi9bFF53dtLDs06a8uwpeZykOa8qdE0lJJiMk6WBuM3Lrhbs
0SW1d+bsXA7xr43kAs59FmmO64JaTtKPIak1jUtO1QtnrM8ZBKStMU2zby0OBzqK
foNC2KeJWMu1GP/toZsgRQdBKcgJm4VK5ZERy4go4XPd9FLeDkUpq1qs/zSEmFPW
GsYlGsbhggyKfttdivCDlrYDEiyZX701xuttX5m78K7d++iC1rBHnOO8mHC8akTQ
OFby/w4xbQ80UX4Vt3iSH/Rmew+txq1cia/Z9jwSKk9hdOPC6EXv7O9fW8b/DkWO
1WQ0oStsJvx9HjQtV7tUwqY/05DOlwz9/tXEBj9Bm8FC37zU0/lPoG5hJuaTfKdD
u0CdV9eOpdQLEKcvZtLk0WaRwr0E5taPpVk65GcclCmiadUoa9fZsrUiK/Y9SbFA
q8MKZEdQbHPrA7u1ZkzDXjKVvGTTsVpxyFYjKEBiq3+OLfacMbPZRiUF1dyU9FnA
vqufPRl0LLxaTyiOxYiZ1guXbi2a2gAcCv+a4cuIC6wFj/Fl5T/6UO/E6oLLfh/5
DP7yAjRe+i77inDWUPlTwkFDhb8LGGIh8YuyLNZJSdiEc5Icmc0VAWWQMroffOOJ
TOIAAf/87JjgDbwpxywrlRrFX3Ar5xYm0onoswlTkq45ZCU4hpFv30cB7hmQancC
/gayNb8Ep+92VOpOJ1HjI+d1vhujZqXEUM8kSZs9pPZWsWB2lsysRikPYo8zWgga
SN08V/hZUNWC5TA/dPxYwergSUW/Si+Lak57muI/nrz+msBA7kABYheFOqu8jDU9
OvCdemEOP33Ty3Mk6BgdRIfjBOWuXKKgSrRRiuhW49b42uIRlOwowJvMV2LPqcBK
xxksNpKZbMRPlETGyE0OhwM+mxyPgny2WcjfHbmYoAmKa+/zipWV7sjfgoORpgNC
XIiwImyg+EdNMjHhz3Y5zPjbDU/cK44xG4rieILhueMLVUHflMRmvOz9npiazrcU
hDYCwi/t0lJz/30vt1NoMwDU6pCruHrp4L8BuBcvL7kSBqwP+TDRYJdP2Hnx1tc3
/CMrQ+BA0+/UH6/T6DbkTsZCOEWnXImi6VXuB7e9LbFyolcfgUjnhi5FHFnBgsbo
AhlTLJiqHYF/QyPyKiUtognGxEMgTXR2sh0vggo8LCONL0GR/Qx7S+ylfFl+hJzT
oUz9nWRTaNhCg53P1JIX6Fqk+0DDbujOURs7KQSYp6TluNMz3mb2mAD45YtzblUA
atLmCCxOhdGtdDZ4DkFrwIMzVmzdUiGHfQ1RYRo9LF4Xka5N37R9X4LrsaCBo0+T
8rCQ1CcviCPtFvSninC6AjbPjPbzcFT+g41MiL2sUXokH2x2MbU45U3IWkFNfzsT
Mdh38/lcBV268GpGqyCU1UYiXykDWjTmhGlxJHFjTI6LCfe5SLw2BbTVhFsyy4tV
XlQAnlZXq+97YjfN6Uds44l+5NhAQy4NPcjaEDYDsXGvWasDoTnPk1cvXNnUaysH
//Y/zJTehBc1bXRPkbcxkxKjYtsvY4e6aJmTyQuT3Bljn8g94e1oLAfRfgmTUP85
U0MEdL/62e9cS2xd8HnTNztC2f094eoFvcRqPkQZXuLwa+zj6wZcer5TfZuQALTw
rAkssltd1OlNIhMzzOK3eMWnbAc66Ub0+HefRRp0U7iWqKXx07S+Wiv5HKWsCYOc
tUsWIkUniMFOxy5rTOVjHcQNnAscH9hVhHHlbW3PUDyF8NXsWLM6W0stSLaLG29F
gDl2QHIrLPn++2EgP1IYx05K+4B3uP29BcDmcgFWBrnH2GZnt5FMqEBNZyUl0SXz
eCIO6exKsOV7hG5U5he+16dwh7eK3d2KWRusmztreopgVB+6xhIQIEQFEcAi3Zwi
fBtcvZXY8pNIhHZGohTY2CEwyGd9v1tR6KVsHh31UKqAeopf9yW5Geu8UyhViKjU
qJG+wpxssH1Yzoz4vJDzhwe1ZelZv+RnKeKSwywHIh/R8/kAjMIjrogdRzDHwfaO
VwayDnMHPzhxlQv8tmUwl3H4F4MR4evZEDGUUoxmaGMGgPxpXU4eWW/gQUrTX03j
sbxUe/1BZi6ZT5ZQF2j5aB0XDkPY/f6EF1qi0OLmClOM8PHWXoSPFGA3huwoSSvq
j+SkykCUHVDJzgEdGel+uJfrTM/F3Sh+MfUfK6q/buyObC2OOyvxQ6LSLOeljXTV
Q/REEXSGbUBO0xUK6eZcy/+zxRNJUbvjgAK4uyB4eenn+jkZmsqVZJ3bjp9vSI8L
zoWHWnISsLHhpqsOhuJ2hls9aVAwISARECZYlyVUWsKHWomv9Lbh6yZff/v+tUjz
ueiGj+MgMrolJpPey0UU293hMNU+vFOi0ZwDbvKrVxv09UvfkyluDrWycCQFeuZo
3GLAfkBZ6kQQjAOaz/jCSXHrP+SqA0FrzSQz96XxlM5MedAuFptUegTWEdRfZEm8
fJGFYnt32M/uXhV8JBPUc59gCe5X3yD8cmStiZIUq/IZtoWlHK7XL7Hv4yRKst2b
b1ZrEZ6QeTqV2JdQQKmQfS3PEFUt+KxCqnxBg5vBfFOBe4sy9vuqUHx+xbsnhRab
U4m9OsLyK5DIfbogjSBdb51CAnUkargJS13EkcdxpcuPkrDcGPj8QsJAlwiRQdUD
kk+RYMeyA17ZdId3QPb9PRkr9rlhQjQGWzLjxmaSAj7GmJqu+GvuBoLZlyICmeuX
Nb1NaqP10tpro/YMyK05b1HtrV+e6YEsJa77gcJ/WcRsFdVy49LgJZZBiado0bTY
nCgLDHMFlsku9xwx3MOjhga5F39UWN7i620Rm5hVlwakXxh3iniAfEtopogFpwGb
RRkAdhEUB64Nci6iNzBfDMdXsDihWg4hOFejVzChf6cghHto3Tdwqdjzz96nH23n
sYfkjG/vy8z/iPzF1v/odfLlOCwVOs/zGC3SaTRAnXrpt6AVzdg3UOGotGOCi1vK
QhkrpBMERM05sod48+4xV0XqeyRkNtb6905KD17kCKciBAvlSNk8f6Cc2BL9reyH
+mv6o69n39Zy7xkNmkJOiohKTqeoY5vZ4dVgAhXMUVl4yqCa6E4CcgJig3lQy0iS
R1jR2vXbuzWVo6RfUh/Drs4Q66h7hpM+LBELLP//V0vXOonk3y1mFCTe5N7XIyA3
U/pyL/kwQGGbbBjynCB+LmXsp13jfMdZkA8PvKCTbhxwULzbn9Jwt7UEsl39oZ5i
RQn58IB0igdcZYPtBvdevrtayHUlJx40wd2+uNXTZIFQS/LpLCREHmv7sH3DIxj0
MSIl2h8Nw+vlPqFZlkqW3Us9FKBb1PRfFhRasAhJ8/i1IubIMkhnA8B7qGdfhtpJ
uqQgQwP42TBV3pGr9bXpEkzRvf5137ik36odOJJlU6mWVwPyLUEx5YRcYVk/7u8/
japxupEABz9bkH61hmtFTZi0xBDFujBYE/IeQJatsRaXBYZYPsuUhjxPI1TK0NDu
aKGaU/hgUgmACV2yzj05Jeo59Q67ptnydbMhCfEhwjTRzX4gVzz9J5FUQfAfR6i5
i/3rNlTrCZK7ilzeWIvTb/VcegNvWYpUeZ4kNx7q6rz8Ooc94a3TU9rv2vkgnJvS
5c9wevCKon61pSXKlUXsG9xosGSOO/CvyoB+qFp4AhyYmyqXiA7WcWxqOuuPJPrI
aOa0dwH0BlsidsBhBE8sB27dv1eWWWVszkoSvw436eyMSoFZxwVbsUDetbThNBcK
RLFOw5QOZehwEZEyVuf8W9jJ1vkFuvGaircGMCcF7DHX/t1Mp5lHbfNhqy85q7tW
SrTWETYHKZaKDwF+gaQCa5u/+93Csahh10IbKJxCXfe4xdVKps0e2pv5F61H2JaO
rb2JxHcsIE1Si8W7rYMGlB3R8DpPLkblxjqrFizrBe2HmNOjVjz3FpckmSQFoSO/
6byhsRQAro04l4G23a9A3rDcWxNe72X+Ha315g+56bHnMchP2JnUx2OBRvZc94Oo
KKVoyQ/j7kFlUQx3vei/yMWPX74j77tLBM7yKqBCP+SVaHGNOby4J5Ne44p3D+sf
RakIy9cS08ophSGP35Jz1vjnvvZiTMKcTF2mycgYt24lNUhwoV6UVwTbu4I0CgiX
m5JEz0hK9qFvIkegmBgmwOkryxTEPtDBDZ2zZGnmYbbHo2r60qM5THki+Rm8yRbt
IQrWgQAaaUohRao/Hcs/RVLKDDk0BNg+lqbW37/KQJmhCQplUxD7GV1sqk/eA8ZQ
dEkAlcBiKLNCfC/iRKRlMhF1aw3ErPpsR2+6LHYPftuz+BrfiArLYnCZcyo8+qtK
/+VAA+bsBTnDExAwtsxKur6nosorS7WJQmCgHVIZA7OBZE2kKj9UdzReS+Tez0OX
93fCP1mjGf421WxBP4A9X4r7AazSDQk1ZFdcCJZS8gglThm8rnt7iRN6KskOB++r
xwOtSl5/5fNDxsmN6JpIBLQp54xLk01ZQFoz7UkmXT6/538tJ/DPx47exhHxJcJZ
zqf8QGlmR1cU1TXW5OlEmQYrByXwsiIHTwjIp1xB78aKz/hFrtBHZQHAYUlUOyMD
eA+55BgmpgWzJJKAjBRThiQ0soEAdqsdINT1Xc+f6TVbWED7XBtolz3DOePsekAE
NrYwq1RVv78ZlVOTPtFWj1zmxVvRbMlbYgfnqSkPBN5jCeOhE4dS10aqDg1ZJvO4
/FVWwSe0uPTicME/gfc17LqPAXr38VizWjnmNz5iXvoXgGrUJeWrVb4CeYUPsmRD
CK20elbYK8QWS5dffw+f6Wc2dDt7EzfWWZq0SKR1fPHJ7dVSi8GdVqZkDBZs0ien
wIM96ocBHMMQiKhPgtSIBGv5qEJ/8AXt49JH5KUgftRB6Cf3OvsOnMfofiLo1Aid
dzOsB+6hzlJHoumAXlPueY9lCk6ltWIzGLxRTvshfpfw1CtyRSgf5lyJTjVJ3otC
XHpqzRzEWQTboWS/tcRWv7M2teiPNn+ZQJXl3jSoLlRE/9OBEUlbLFjfTOGESLN7
bmEHKRl6pFA2eEm9ewtBKUkqXL44jzcsln+1e2eDlFpJrfC2Uiz64K7JSqezMAYX
UupdvpsrwHz55Fr6ZksJP9CcGVITz0KHaoWu86QyFbmByopWnisY2iMPICs1MLwE
f4fTAF563zA7InjdUZTnhuBZtYu4XHn6PeErl3RJB5aflL7gvixhLPLJSAP0bHmX
Lt5t6UBC4vgfEKBItyqw21yKIUC+0cNLyvZlODJUeA7JiLvvilTIKqQ3QPwpPnDJ
0xVunEiLnMVcU/71r+i8VUqdutemdgh25qfGdL6jhov57/OIns0qc6wzeJLZSgVd
/CYYKp3G00qbn8OThukEIUybrWmPnqaWCrByrj78Wbr10Hqldwlia9on6ZFlazWO
uPcKUoxDUG9ebpzuJZ/qdITWeiqzp8LEO5+XLkSpoEBAT8zKooMM/sYq+QyUVyVG
ztXa0E7NY50SqeRy7JSif0rx/4iWvbXywYAriuP/iOH9Fng3972lmzrWSmPffNcN
FP6Nksfpk3uOWOWluyR/rDZA59QVp4a2e7PcncDhOqf40nnpoab5cjQFw0vgPGKs
5yk4re6s6kV99gfKKrSKM8Qy4Ey5G9umh/2uhgP8N/BL2E8DMwswqKlUju7w19uM
8RdnN2t5JiQq0PHMM3FuUWxtwCbBWeK0UiRgYdYLjo9u59EnHvBZgjR41EDFxvB1
fz1MCyQycyFwG0Z0rpAjhtlriDMXdRu+E3Q+/iuw5osAkcy7myvH4+Wz/oh9Ta0O
QllFaJkSJmmcERj3ahLWhqXfhdWkApZ05SFdl9kEhpiL5Xlq3qzPRpvOdiT9js/F
tXmZcPAo1Vyk2zT5EcUGO//b5vp+fJ/9VdYO3yCGZgHlcLmzW7PlSdrp/6czO0A0
ezoPXAHn/qANvn1+4BXmKutjSIgl8lFchQ2UTZtT7fe4I7vOX2M2891HTWrcwhAr
7TUde+FoWYORhQwrPJebkKqpni6wjXEa8BxPy/fVA0P9BpSeSEc08b2NZaXYnJzF
M3AMNmOF84ameLKaGhf0YSn+XQDYzvm+4yJvnnhdohKU6vAAM17ZF/5RkHXny9t3
huk3lixkuyDU4gfNhW710KaVA1GR7gQOq0xmtVpO9QwHG9hTIkFp9pW6Al7FloKZ
5+3e5vhkwjmzVwdgGZ1JFF9wJQZTZgbG3/rkHDYz9yH3Ja5HniZ/bPmC9mipL+ht
LETZQtU+mItoh2mhAIpG/c2FoAFfq8GMtPxaGRUifpdEAnAYlSaV+cgDx3OXSJyC
ucx9pD8U4R9u/bahRRrsI0k1FkXnnHKkX+hdnVIZ+paC7u/mHsya/xNvJMunUsSu
7VjCnGGKxMjh0YNIbN6hfkvfeR7kDX3I/yHvJihP9z6C5wJ+QvtitWBRfdSuvZpa
7h7aWhUaaYh8o55o+atvtbbzenKvVHOS71deUCNKX8HZK62Xf04kGsb5dW7Qd4n4
+x+33GzcnxFyXaE89exJCp2VJglNIby4euT60wAcZomGLl1ndpRgQpPMtG7bdmQr
+G6A90U/VLXIdsbtwRIAA06qg8ZQHb/bByvPlN2y2dxjSFDBqUJouKuZNsbktlJI
4EDFzgeOVd8K3e8BCk6/tvNsCqJS2u2RriOhA/PWC0Fej0a9QhEoZYLVxb8bHPtI
C/jnUiJ3qL+acSDAEgm/8o3aRxYaO9fXHnEG5c1ffros3Y/gGoPpfAusC28AgUqC
UtRhNYeiah1PK0QSZzilKC3Eb3AObGYAQaOa51sTYrUSaKpkhemS3INa5T2/8kAM
KSmMmzYvGkP07zbPRVdUIn+n68hjPu68ZG/U9nswHoG7oNTWLYlgD+e10kVuYrdG
VnARvNGRYp0YGoHKhLqYLI4ezn0Q9MSw6kSI+8R78TIpHUJjqX+Qw4BpadxSsgTR
HSJVyfY3g8I/PBWptNSFgfmWNofkr5MW7zkMklWBWWlPxcDL9WLdbPVGQ44y2/gG
PCrJOZthYIzyMtJ9WFl9Yk0St533u/SAJ5/ZRxlyGzYaAuq5tJvq3GwOxkSRTTt5
BrK09efK7i3Ur5TBmT3+qS0lTd97E62L/IYUM4l0Uh7YTTAUW8y9hdOmSkA/8YUr
mI0Br14Rs5+/BWZ0EJs+g/sq1NvlMpkdhV4vwpHfGpwQMYGyjAUaH3lzmqda65TK
mFRHRERe51px64NucxS0f/TuorN3AkxEoOJ9aAWgJGumirjBoPHGPc5Kf8qwOJjV
DVsF59Oz+wCKZ7Zhx4uq5fAG5MFpDa+8qEU/oAEXvwQnm4Vb9PYmJ1h6z97+4qMM
S235Scc2lKAj7vqUyhz+QVGsvIrwxNUQ2dl/X8uZ/S86C8Cjuu9/wpGBlw45TZks
X0pnD2Pm6rmXN9iM5mU+Pa2/smEfhiemD3XnHLwkQaDPLOjkgrsRA42UfHGr04pJ
h9tDHoWyl1wJtdkb/3knmqOsyVm8R9S3ZTbRG41hxBa05p7x8pPb773+Vq6/Lkhr
DW/sl+37h8MAWHoyL3SDzBEkNcmQNhzMl1Z1RCD5kP95zEGpUODYxTJiETrRSPY1
YBGPw5eFiV/X0zv/fOUvjns40mMOqoQldPWLXnP2dHoC3ZSYXmIr6yV480auLtSq
yLzsOY4MkGcI7uu2LVV7UGzZRt4jXKxg/Ewx2niQIpUYbcMrTQ+dYHBYBEtUDN4O
zEu+JIwpjYcYK7A8iF8uus9URTWxHvymfcFU3BANgpldP0r1Y1Cf/wGkX4XM2arH
wyNuyZxy9NUisjTbrCcTyBNF0wub+DE41wA9d1KRhUjYe78MbzRLVAovSw8VpKem
X8e1l72IRAOTbhJqUMc4zGlSfwTVFIudw1YOjjcZnttOPV7ZI4ZowzGkyCZTAjUN
IfOnedo+HClUBvzqq0GRJtC4HxJWs21hVs4Fjv6DndqjQD+8AKu/Xy0Tn0HxbsLl
ispkDwQPyglhryppjIzJRSxFcJgrAXF3pcIYsAcscOgO0UpwLXk2MQyAh1WzZjTm
oIdlAnBZr5G9ziPJATja0lfzwDsr1FfZWisq+qo2jPVuTDf7mmIFRlrX/ZgqMNl3
MarJ9SllPD711rkF9WlfmI5vnZxATkqEFt5l37cUVVOAtbXRxxVPyZjn0DLVTAt9
Fcl0blUmt02xq6ksYm2ZY91aHEuZL9pYUa2WniWGuLqaaHzXZfkbBuJU/RtBN5Ls
y/LlXytPx8VgWFx1prZdlNBqbYWZBIxBW20nlyHNEfgmAPWXR+cRlnrIh6RyxmaH
zVBqc6N2ngd0aKNDAtlh80s6A7V+acJhlh8+/sM3N6z1ynygntSvhszk5pCbKAHe
qVRX4QBwJGh8q5+o/as3xF0rTHcG0Ta0eX1bpYWZwGuSJKF0VMRH3ioQVyAfI/lu
WFbCuY9yqw49NZ2x/wp2lmVnvjy+haN4pPANFn3Jda9++zqKaC9LYMWkd/gYSCOW
B1yCFwkmK3s7yf0nzR0HICybnp7mvgvQsKZtIxIsYHYD9IFfnTs45PFBf9BGS0Lq
RBzsrNBYfyq+0dcYEojd9MpbhPtZM4+tL8clN0nMlBXDJf++Z/9RWHzssmjmWMal
cm8N8lv8ZQ//U6i2wJwepLv/nNhoGq7TGMrdH/3YoRcezZ+Q9rH1YAXDTiQ1VNaz
AHVGfoU6YHIh4/SvMV7tXSqmwWZCaH9PDcMSeCgWB6w4Dvd0nbRjbgYGgXOogX0b
3HkSUVqMsnTLMElOwwcGuMBaSRh7qjUC/FOhcNudz1bXUefmS3Ld/qmxJSfQU4HX
qY1If3w/GIdolS/UWVzCNJY2uA/DiXpyeao3TaMl9sKmmRTl1DiD040roVgkAbk7
6o6aJfScDLo8AYHPPoXxGT3ekzIW73H5HfJ/Yi6woI4IZrbBfPCTrsuDKK6q1M/o
vdOqIdwl1+wt6uvIghzmzQ5rQbM3EXAhNPzIpWzV6ngfzO/dT6EuaQABqJyBFhOC
b5AfKq4X3bZmnqf+sV8eicD/A9lrrD7HMmVNDc1U7EqqvkGspfIABj626lzcxu8m
xxksDBgXD0syYFWk2c8eeZmrGZfc/C7ogSbuafb4EtdELZcyEsjkOYwr1nh2GBdI
P48G0l/7xOnDxEk3QQewWx46pd/43yZRe2XzCG5V5u1k2WiMwGe9ZLv3FUcFizZf
+IzpwuhMFAhC0QKQ+ROM13Cfi/jUWWM9nIatEXm0e3YPla3TrJvR1RtlkX7OIEDo
rbg3Ou7k6/eACS+gve6ohWGvCTrhbjkdOttR1H1NH2JWKrenaPmtt7y5LaM9B5fW
dcWkIKAF2JXpLI7VHrqDiV9mPHw2xXQdPACtdYhiLC626+bU8PN69OoWiBZ41kC8
+Z2lMPQnqxE6pCSuQYaEgMwfUTqhAaSEvd4ueEe2xmclAN+vznIKyBLQRq9R4FY3
ZH407GHjtmDyQ8CGgb28Vuke4R50DRI72NINJzhZJCEgkiFfSaaLsABofqxYLtGG
tqs5GtNw16We03uE6BDvzBkIXHtzrPIXX37R2Uw7mf86MT2zuUFDjfc/Gtey0ZFy
xfrzd5fFii6hss1e3yJRr28l6JsUGOawgYy5F8VQZTfRMcXSe96UppTYk1JxoSW6
MLzDRVpbmZ0GcAb5Mdu6y7IB+Khc2cFoZd8Ig8LWokIo8Ab8vnw5gg3a9HKtU9xg
CAl+i2Xw/1YiiASo4qK7XfiIKep0s3PC/WcuS0WbS+aAf2RXHGAP8cyGh1rom44m
DYN9b0mUE6l4Lf3Ww125wUttjkEcbzKhGD9k0ZOF055pI/6laP3V1itoJqVbj+ma
QrcNbhAkITe6eIivQcPmjkvW8odIiy07awpRLl0RroHMz76ovwSnzdu+a6oCLNRT
ZMuRRBMRtRePUzhp0ZBlXjp35bIVKcyjXFIjsQORFdZvjOWqB9uGMcVHF/QOMTlv
vmNFI5p+Qlpv3q7PNgo7eRX5eYLVjH8irk86ecniCYJda/smDv2oLw5Ua1jJOJ6N
kkanqMxVAJBzcTjwbFvmdNqenwh7RcUEF4475uVix8nz5H54Fxd6GYkmKSNYxIUk
e+9+qEXR5VqGSedFtenG5y0vd+0Ji6ilZGG3zjLP2lQ05WiV4K3yr182Hv1+z0Xz
mo0dtwoNRTze1rS9Z6Y8K/pKuTJXPzxyLlxdd5szef0x8BHdUHk3ujTNPEVbS0PA
4kjghLXtIO0LMSclsMbdlHpTRgbff6g2qbo0gc7c40WbHCfd6hBYh8Jop/Q/TY6c
kkIKXuc0i8UR5Lxozm8k+ymq30yEQ8dQYlwzCv4GpGp29vZulDfGo/aiagfZ/foW
nm8sxOBEwNcXUe+cjmQONUzDDsd28cZE4Gr0LmHdLHaiIOB7jfWxOK8auX+dq5Dq
5gmPfNBteIt3mI1rpxIQG/DeVGYUCNXSowPUUyUsSefumfHBbTt672nkNzb1uWPw
xJU6xWL/qmwPosFoeD/T1pbcmeF3I5Je1af/odATPtDbgH2t4LsEc1IScEvNhpLe
Uy8COhxpaPCfbnQnfTvGf3n+e3pn5oVcE7T3ZvApwLhM+kL/injJAx6HK/njGnNH
uSqupvxEquOUi/xV4gfpMjtMlKE4R/8OLRH8y3BiyIhObCnEOVp9rtABqjX6/EFb
Ohk+2NcAaPqvuoppGap5wxIk9tjR8g5o5wfcDPanSwvIozFxB7pgcuu3tY49csdY
z18/ZCQCGHTkWWyN93Gq4WYaju4yJA59hG1yJ/2cSIHUv2sg6RoaJdD/VjMIHjOr
lmn33ne9zUAf4paAtur5XQbQQL2zBPTssU4Lyqdb9ZnrYD+Jev/xC48eRI4tjja4
FZ7/UyTTSnA/lDByMU41UidX/UxnTKMuz7lKVgIKHAYGsvVv1BsBwuNIofsKfjZk
tc95I7NgqCCIdDChKBCUM8+DR6PBnFkFPWjIbKdvTgMg2Z3CFoRZlCnrv55STCi9
0p/lABGQ6rxIeqSA27B+/BnAaIm4E1u23WZz5VcnRpzqWF8e3I18pR8lLuBaCHRm
QpHjhDccHvN3gbvDLOqxRohyAr3PElP728/7PnnlxTzfHjeOELRfTH1uPIYunULF
MnaYPQfqmGlk5dospaxm0AHqxtZzPFJXVubaa/FXvZ7GxBzCO8IKAckuIt/l6GIF
b8eom207Yiv3DijLHEV8dLBpewdJ14ua1q6dhaI5hbwlRxj08A0qUWP8XxylbQOX
2zfpT51WmegIJuStKAQPDARY+h6EhAymjP2GMp89jGf6prEHm2LSAHoJ/zeiskHH
mV4zeIURbHy8iODTBp5iYA6r75MR6Q+LES3Bb4e5rMXuj0yV9OI1oSRnhG3yDX3o
A/oCQtbOG0r01fXWoRZFjSCboulKOS4aGihfLsV3/xt7Iem7UUp0yk3knL2zBOSi
yrf6ewEzPef0TwPyCacy/IxPue9oZiD6nq8lriRZ8VnQvfD6rJe6fQFN3L9gaYev
1jgPpHCU1/H9KTdsOeUMqVJmfT9PZa+8lO3lMc5gDJAUuJky4jbx2RK2V/sjvDpY
RRBE1d8XAnk4zZx6A78i7CtTkIb+thPqGUfIsSKuCBFcWI+C7R9hbeqdssT4XxBu
Ol2SuOTWmHCCVOgrLLkd6HfK5jV430DUJG3STzsQkJeusPo9gsXuV3k6tUXeY/42
jjVw7XDEU9QC2NOv+zn9hEJT0PHZWAZry2NNKgpzcwrp95z48h5CNeeXahFL44gC
QJdAhMw+HbIfylnOY4iWtQpt+/8va/8Hq8KhjkfrlOFWMvnStxHH8jkLzn01cQlN
rEvfnYwRzHDfVqoo4beyR7krDl6Lo5bLVNoWnRYkLXmYhAofvbIULk2s9DFTYs6p
jpXzsZkov14zKWBOeITAecM5ivKn4I4D59rPhs8IX14gtFaL99+rD750Ib/V3VTD
/GczdgjUdrXLNR76wVbI6jCh05TYAIDsu6IilrtBKdn08irz/o/gjMbrbEkHv6oa
avQ2PYd9PjYPD0Jo8IcPO/qNOfS2j8XDOrc8mLrQRXaWuBfZwlBfDnXxuSzuPwWi
vpxGqbQHkcsbPcwypOxaPltu9/UmEfkb1oE3//9HDNApo1+O5Zj5L9Y8/kcpMbxg
6LeYA8BIXPe0m3li9KNqQnGOyKbeBr+ZFChymcastAEWRNM6rPEPFUE+ESEoDXjq
x8pmp0kRaWoQkFhcOszLhjtSZ2mQ7q7GSgT4GKp7xzHYKZ7aeESyvlrgdGtNEXGb
qwX84UqXnhSx9lNgVwUYGZvDLB2aFkzqihSH7sGmVsSnf61ZCbn9ZjLNq/9QQxSc
eCdh8rGVMkMBVRCgmfHgnKCXxtJFlr4eyHdRgI2UGnHYaW1T1h4x/faLZZr1PhlD
NLug7H6926sclUWIVBHGwKofBoC8k1XLQCSGs+XObnSD9NYtXN2flofHLB7OMPgT
pgN0MIdgCIpsdyFepfLnABh4PEiIfs548x+fy/eq5jgjMh2i8s8uckgDy7W5DY+J
CihtJHp9NH7h1LFWXXqu/6rnHT/LlyyGNxrA0V6omv932qYqfGh+AyLS/lKzZ/0i
WF2sE1LI4tXE8vQvuWHhRipYpUWrOV5ONwhzftCZnLcndOYeQU/ePQefYx485Jzf
Xteo2hwoK7vp4VGhkm0YaR+9mWStS0AqeTt8nGja1bli/qgBKcjKTlXZ03uJLXCF
CmwNkamxxRKPt1EmfSb0MSAANbv9g6tioXi2RYrZkcbVMW0ukxC/ypVS/oiBdChp
jd/aH1/4cP9Q8dAK2fzpH9Nnc+olnOgzT1rCL6Bvt+MN+4LU7G/XiRmONyiyR3lx
1z4dS1mrRkeHVcFBlkkRAjo2WQL0icNEWlU73QijX2ELOhrt7ezLv20lqoraS1vV
X0NN94wxS+UIc1i5DmvBSzzjN2alxjQ1ktkXG2jUaJPA6c7IS//EN6R/9l3luqHL
Xkg+T72wFTdNgnsOg0vocXAxONC2Pb63cnVnhevxFFyuZH9pBNBy5SxovbpCSjsz
TYVtRufWkQBvAIovl+AN8L5CeFRa/unrJWSV/6KtccaUcI9ilBXw2aaSaQN06fEQ
yzhcPyc3Ag9VHAiNxQg63W+u6IAv+UrpbCbjXnTa5RHvBy9g/QExpzWdOQ0s8eLp
cyQP/vWS2Qr7XdcpliWQjZqzsKLw2je8Qws9bz9sQixlxiRHKlVgusttSGj79lg2
4JxLoYQq/IUN+AdoN6uLWDMJYBztcLDIw6BErwieVSEs5Nr8/fBNrhxmZrnMuM8b
F+3CC0jFemxObNNXIkgs0iymQQTUWiZ/uiQNku+16GYHuwMBIT0F1aJ+6IclsCBd
SlqBG4iAP3yF7yljTlR9dUaBSv+kQ57b/cHVnV5qh2yNsrxNPSBWhTHAB5alIKCV
aqs65rDZFQjKXKBgQQv7nkq0BZ/dLgCBA/QTtmRPudSukrxwKqYOXLiNPwFLbw4h
RSlJf9AfmbqJR5GwNvae/klIdGwbk+CYB99NGeN/y7QuI+RxvGLis59m/ZZaTZCP
LMZDHXj6fQnkF/Ns3FUNSTS4G3aguTEXAEFiTSgH4xq2qawz3CjYlm++v9GArTNl
7yQ07kailRXPYqStTzyBWWUv6/moZmYrxdUPSXXeGNfAXHh+CRMCWbVLHjVCNwhT
SbKkNtxE5TXGV5iJ+DaKpRFdTW5g0G4WonPe6eXSbuoU+R2OH0S1r+K1u5IMQ1ke
u8yd7dZeNqaRKAU+8d7zdhq4feKIPoxt76FnWyl2OOOWU8flLOBi2kcaLnmJzpuh
m6uZPMbtK0f0t5hByOh/0iTIndH1MJ/6yeYB9T9NjeIjB26xInvLgaynK4oDo2dE
3vPEn0vQHIvrdHKryuZ32oqpbJhK7ZH99fmNjrqdTFJZZCMpcHUBZ/KlyyJbMNTF
j29ZCjiB+GTp6l00T+i5U1hhdSxpTESSmYah+mD9IiffCPYrnLqfW7l2mgIMj7tW
FiJX5W6VkigGfuauwHn0Ab2OdAHb4wyKVYui83xlENvalEAoMSEm84pc+phoOkY+
2wxgrESXbE4nYdpfEen7Cr6PccBA4tUp5wwjtoetVzqY2bhjIEPZx37YNg/yg0qf
d1+ECiG/XRzP/MrmK8sOsOE8jWbdfE48bsDui+UYMgsrgq5amSNrWfk52uMRq1Qn
01eIT+wov9W0bA+zEY00J/aRrjU3mIWFBwrSpCrzZEJYCJhS8WWk82jyo2QpNamq
7e/nikYlTfk9HAhhWQykIP0hTVrI8IoOU70QMAClccXL5RFQZ7lIT0+D+NWiVjiI
h/peEMaxSIDE+mrOVbKLmvhP9+nLxBZEQJ9ldRW75fxVHthuAaVpYqyH2WIKjEDw
sTpV3aLawYJvLFvkw4v6vTptmu1+1qjhYP8CJ1ET+dZDhOz97PfeVNCfhq5r0EfT
j2M4yYvRd0sNKRr5obu4ZYmIZWuBkFX5inbij1TgQk1O4NppuwxwzKDRlH+ODuW5
fmEdHjfWThxlRffFjZP1YVnHt8KMosjTNJ6u4BXJoMpc/AHqveEj5MGm4XpH4bd6
fa7kKDHCCANroyqFywNd/UEFNdlWNa+sLdI+rp/JVewTtOpZgB66XFi1wysQIsdF
ikAKQ79nEbwkJ+l5T1IPqwMGzTzaHIkI1Tn6C5I5zhcCermrzb9g03bMAfnPvZAT
7AWPaTFvXvXli3NlE0dh7chjBlilnCgkcdFxhoUdKje8MlOywKwVvjl/9iEWxvpl
CboExeB3Mix/TVHdAR92L0Ej/14fnPZg3S9efIEbyJODm6pemXQmPxcL1SQ4EjyW
k2z+U9/Svg9PycnuDu67hp/qwM4L/96K7MDQAMkNMkqp6WWxrAVElcuQzU4MATpr
O6eFdB8XevvhYG1x+kdw4z79tEYo1ZvfXelY4BamIsl1xDxfYAaeE464trA1XL/s
1kMg5rWCh5/PxCgSSOBttOBaFYhPCG52PMQlDIBKpMlMogkixu6MkVQ6nxhBCigo
TfbKs/hFNBv/jWZIYtIXsSP2Sau1gV19CLz4mBPQXmaicCzXi989chMPjaYqGZuW
2G0pfbHWwkX0KI5Nlh+4fRfA+d5UtiNAKxXmshWAssP6gWQLcZmttZXC+N2746xS
0fn+o5mAiqmMCXQXRqsT4Fw9T4IqZNOXCfWi2MF0zmAC8xQHwHM0k/gzBqQn0B0H
jeJl/VrZL6n62lgM0X1sJyJkvRx9v2G94kti7pOO3w0SsAXVsFaiPoIOyZdYO8Ho
iJZhEBmT/ejkPB9BbueZiGHWgJu0CA7scxTWz2sOCiBhF++c9Hl24UHqzBG8KLEU
PdEpGdBlV0kO7Lc26O37Axb+iHTHhCIJryFDtNgnZKAoUzlx6EwgS07xV6uHXBPq
c9wn70UwmMGlPaPORi24WJgs7EvqYnZ+A6JvRRMw7jFNWZPrN3rpxSmncRK4YYyY
hDD1y3ISKr6Q+l7FqISLtSuNZq3No7RncsU1zyrBz4Qew6lfylLa5iHnB/GQ3tHk
bnWsBn2kpLPlLJBJZp/vAOXo2bc7p6Vhs0nwGbz+tADpemO8t+gahyouDGgxFMN3
+duvUmhfr99uaX+6G29Qv+Knm9KmDnlbxQoGMgWBMGW6o3cJ3INCKQRLdfe+SdpI
lKi6rxTuYJ65E0N243QJonCBbbt4bN7slH/nRRSbmNTDSI4uN1anAzcelpyckpRH
AwwzfK38UEaFpmjSNmhKBucfd0Wj+W0uJZojNjxWVpXPxdzcI7S0vm4cl7DBOsaS
R6ywPDYIV506/gRFYGYGOo0V/5jVbi6YEbGXjwK/lI1f3+lHJnAHkdD/AQp1eYsL
IiXrNecDsKgyOnqzd4JBqjT4wWqiksX6asCzdkSRxa+tYqFVA2L0O6jkO03Lyraj
B7mVUH43gLCDVbAxLe3j/LuG49H6iwnCYU1F3ceKlchidQa5mbLom4PfZsiigPp3
RBDi3b9CxraT7IUNgWiynrMY0l5Xra18w2e+vrN1i8LGbtrkZEvxhTp5MAtIchw7
kEg+ix3yOtY6Ni22XMI9WTaiSOhUp3AgNgPliB+aXPWFnt2ofmuZAzd8uzp7HDZL
ttpT7N4TCRAjqv5H7Ec8i4yRQ+VYboqLEVdpjiaT/RaRnGIcvyhMM3q2BCXxutsU
tUzFBz9yupiufGMyFAqcXpj2tm1mX69uVSxFWVm9dT1IE8LKiqlDP/+JmuRUWN/J
0HavwSK60Og0rdIJSaQWzDR7czAjEUZ7YalUJR3rO4T6RwXYLnJch+OmX89y8kPo
HN+9S6nxCFepyYMzqCkNuxjcfC9fu9gOLjMyGKmboqDGliNrfTor+SqTGvetcuDN
xIPtfoONX8P7c2ebUyiBYfRISefIQxqja5yYMkUZrxOEeEcK5dkbYEC3C8iYlTPP
z0Ky9PQVnyp3pHw6chKy0Spr0yqkl1sTRfw4BsT11wpvf37l8zK3uuVeeOrfrKDs
tF6mnW4Ek1W8eR3lA50a8vb/LIWiqrcUss3ipYfj2LbCYHjNBvyU/KZS1VrXs4N4
y9GK6EAbG7ZZZQM2/TeDzn7GsdMAw/kcTs7YuQrEHiehwMNosRCJvwfMuVOQP6Xe
Ovg0IodcIuCg3biWLe/bq13zkB0fAJWPqBabuKRGo9crOCr404BYJ/VlouxPl2Oh
IEB63UNgqUz+rgEUW7SnOR87e5fN0TmbRWXQo/X7+HqDnd/j0KsGH4RUiXQaO9YH
EMnUpgAlmsucZy8hvJVn+BBns+3tB/6u0vGZrEjTfS9nUR8RkjX0mv/opGOX+lXJ
ImytgEzTxN/pr5i3UKEFhRPkxMihzeXBqVglreKcF790s+iURmGClPl6+i/bYf1q
45OMNzqeVrvBzy2s6mrUT5srzd+7Ho5ju9KXXvw86Fz32lKefnsi2o0bYTNjlKrX
v1YjXm+V4EIlj29ZZOh00DY0Eswvu/NCRjK8ffRtzsqITGo4ORw5LEU55j8Bwk5h
IMZPisdDb1DvMmuzpBu6aDtXlU0OMz/XVZ1k4ggld0cXQVaioeEXqUV7vIadlA/K
KsY3mDjetvUDzq9lWZ9dfi0l1n/0tsIiSsPX6bImERQJ3WKGpN4e4F7L6qwbcrMw
cSSBJGJbM/aYR8gVIyOXabPjNrmMnDUD5GpNxI0cIjUPjP5HYPh4CxShdyu9wDu9
QhE1piZQ+0YY6hbC6o/ts0aNK1PCjBvFJP5fbdt73HkNj9cqLAsInGomHvr/OXV/
myQf/MtyE/7tRkQbQkNDZ3KjOYd8PUYlfp+udeSwTbiNMsc9T9WCJhZeBhwJFIp8
nzN0lFtu/GkLphjf0KLj3mfCdj8D6+J6g/ReDl2MvLeLA0KfRf3SigUGvaR3loQw
2xg4RCGcdreo7HAJUTcxaV87vr/3XCaIaeCZp0MUV5dmN5ts6baDQ1ouSX9f+ElK
ejhw2qTWmMdlIibwloybQABCbV2YPvCnskWtV3ubR3qRkN/5Qv5739j1sROkrVby
j3FDje2AldRKkLYqOYAOLatZWicHHGXfS3jVlGdDsr4K12yB3wXNVodF6vJGS3cz
WCWf0ebNrrVO4/8r8Ts+iWxtZ72mSJoc2uM6K9sQ5S72UQcXoSTEG0en1eATunh1
6rxGF8beFO3kUo5vijizZB+6Kwu9umGtN085zjXICBeCWHON1ugNRtB0vUbp77so
NVehMbBo59NC+gH+tE+WAPv5LZXG4/nSu217+hdyy3xd8TWRLSHprV8+ir14GQO6
+YVWkoP5nyp1P5/mFaaVfHI4Agpl/wkWDAPZOGHMjFNoOh140QiiHH0i4xMVXFyK
JnMvSB/F08MafmMuGMkaCeR3R3+iZLUjVQwjVwAiG/ztQVKanRaoC3ak19LE1OTY
qhO48/Ea2Rmml9sQ1xHKQmJrJjpEjdMPM+kAHZnVIVLkgFf7HwYyene4Ae+DzOxV
s94ArRn+G+MAEiCEZRqHyUkpfofF0uG8TnGtORJ4tNdD4knas9xrJreWCSjLuEZN
QS6I/aIGIpcTFglGuW9yzFaMJxEuQKjg5yzEanzLZm13W2oUvGuss76Th3qaUuGS
ptiyoDerADHIWYP7S2goBB1Cm8kteW+lDagTVe85S9kgLvSmkUNQgMMmahYTs32Q
Q7M3QcfNK8H088AEcEojCgB1qE957jNm81pj9Hj3PKtbQ+f9PN6cxHjb8bIDNU02
TKqT4Auf0NeTHEnR2Di26zUCE4UAxzipUN9fu+4P5qo9+VzGBLBgez/nyG6cNnAZ
v+odVMbcrSj7HDr5meSnzzlrF9jFI+5cIqx4wMD3eK25+1bc4ymMfkgkF9oaGswA
9898ULZhjbqCtkfgkG/eram9nOquIiEjVyx9l+0aMhfknvWLcM9KYiG7DVIr+bLb
pKDRIOFDG68PDMWM0ZmCzQMvEqWVBaP7fFH9vrK6Gy6HIijNAg/JlhR1ymlAageC
VOgTx1unisEpk7OqkuFGkD0DtUInvnXyGftzQ4Gt2YxnnkdGcFHeJwHrFRm1Gp0g
49T1mkaz5x7g0AyX4OgdhydPqlzE0cD6nrRyg93Fo7RyVSHtG6fBrVOQul/RqIMS
XwZ/BTGOdA3gem8a4MhFIHkhVfM0rttYT5mheNWGwOT1UUlFnJGTkpeLTbzZuSd7
KlplDib7xrw8Si6sratYFN0gZqLlLuAlk4e02DMC/eIjKFAGmQ7c725BNVwfD8A9
QTMWdxHnVx1B0qjGcu5Eq0y0SZ9b6o1nrpp6Vstu8seM8kLJg9Rn3VCHCdtk3xfT
9xSXVXMrb6kTbJ8jj5uLXp3qOhul1sFQvNw7ETcdd8fvE2xCYYq7SVE3yYJKLWD1
2+vNG8U7gaB61EPcG0KJE1wM0LF1AjQbOTRNSgKz171X3BYR8zldb7Rz2r9chLIV
OGNlVrzfTnIjm+T8ta5waL59aiy3BlJyB7WfyRjC1YhwaAo4TBjhzKmIg/R0Gb00
f3F4t2Z4WWmpjByfgFiDcJNnpDLLa4qe1TdudYs/gt26wy+X1eV5AGbhrmLU0nQY
UbR3lxWDLS6bsCRISRNEibqAzDuAmdsQMG0tBTYhIvpL/CYi0HIpcM44hWUZ90Ay
oWmmSjhDLdZkh7czN015A6S4rhe74y4twBkKoJ8XJv2JUoJrdOpE4WB5nke48/EK
PkafJb+FdozhDKzpVe0X+vlIpzUup8UUFL/IDpK7cih3BfAdNNi3MQu7X4SEGewG
JUTgBhQ03tlfurH2aaIQW7nYrOC0T3er05HIlach/rqvy5Z0J4AvC695FqjeJY5R
t+uFkCGAxD8eQPWOOgKxVkZN5zHD211W1GfPJcghHYT5fvvbZZp6AbwdtILlbfJW
mMJjccWw4AWGMzTkKT3uFpV471hIeoftC0zLfrREbutMuT7x1L3uJsbKBL92xMA5
5PvD0SE2hsd/y+2i7d73slUMOu5mA06dQz6HNuxaTnq4B9gZSekdgNFSnJ5dzveX
uEP8eLlz1b494a2ykoH0DEr/bOrLR3c1vSYKqzRIlz39d4meKIB9rFB2Uewxi2C2
1TRLbWPOu4122C5ExuauEQ==
`pragma protect end_protected
