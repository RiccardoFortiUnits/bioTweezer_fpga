`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oSb47FmuVJ+k9XbkMeGM9r0PyL4cIpncHXNtmHkZxqXig7Tmmf4IOMlAmYKEbYWM
bZ5p1tJG5FzE5IxIIABEhnEUSDATnLltFr7omQb43QpxB/FwIAHuxYcyZ56WdHf3
QrqfCBWKi2VGyP6yMYqHuX31/yxmJhoy4OYuQAnnuEM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2064)
AK+TWnJlbYEB2A7skTQ92MMGIAHSRXbitblfc5DTkXZeH+elWdCIP1Dp75SsRU1h
0MYGEbJCuty3s3+//MUthh1C0deL68ZCvR9cfczeBxY74NcicEoIgCck67tComrb
+W7f/nbe2vAbZkqrVkNZHI2zd55kNQmhw9GIN+JzXZ9TO09wqDczZ97SfKneW/3n
qGTJfNFZtRLXoBxzZQj7oWvOS67zurdSuUJdjDAAWN7LJdx2qhn9nyyDFgp3JTd1
GQeDVHHZDzaOB0Km6PcRDnbaw035QTRg+LOYrZnBNpelCII6Mf1Yc+L3mj4Ndob5
JRt/DxrfEPDhQapHXRB7/VBI1IKUMgIxQ+0aqhBV7dwB3gTglcHzEPs4pKXiFlR2
Unthw0mF0U9URNzNZFbnFgzoWxAodJCOWrpcAaBDVlBU9UwHqBo5esLYkFxMB6HV
aYuf2RoLETdpuHxmdGAzZSibscbRudC5qSTLXb21/gBXIaFQ4+WbOtmXpESxDNMu
z6gPHL9QyMPoP5emgTNGkv97cBzy1c6WuUV27XBTKaFxtqk6d6pHsQQIcPVNBvPx
cnGKPT9BjT8AQqgc8LTO9DckHhEOQf2qo2aW+8h1oo5Yo4YiP6QvL3qq0meLqCvh
nsWiFwCiLRD1TByUEQLG8R7xuv2/XaMjY0XXQ3870ffnXDO+G0HxwoFZkQLmMfKO
fTMsp3Gdev2PDlinel+z5APq2GMEIhaw5iZzCwZjhnaJDgNtTmE1hUpIB06yr38k
5WidOs60XfCSM+y06b3/NGIAKEJPmm+Di3Kn1O6iYkrV2lhBnQLHA8Iq4jjJ5vAh
jtqSNpyXT+KRci73arc46bHugRRYS1c8TsK2+/CPGaDhESrV/ObcyK5l5Tx9Rkfy
Jshk0Sv5jEg+RRVF4wwK6baYAZ1xVOfr0F5YaPxXI9w0+pSU6tuXZVo8uASbgAcL
FIb71gko9GarYtlDmvlk/bMSHsOnk5uFuyIPgfwpUjDhR+x1NODL5/oiSG2usLVI
w9OSAxyOGKl9Dsuei14Eps+TRKfyY6soBkioN/sj1K5rZVIcgUNsrVKGO91OvpUB
5Jn+JbNuYZ3miyOYtyl6HZ4qiUDHXK7TmjJdaupscrSQHUv/s3JFJHpKZsTs4e4w
v2soObMiFO8Us0gOBjOdvet8Sz76CyxILCgj3QNXw503NN9aXejplZlPeziBZNDw
FcQxVFDOD2lwHvLYZJ9Rc1R/DMsu6TbJHRS+ilA31wD/th9JSRnMBKfXXlR7W643
zeTAltFzN4Jgstshsi1yabuzUfoOALcc0A+Kb6eqzzW+7f/Vs2Xbw4wsojghd4cN
U8CZrbw/wgxAQBJVjbGfcLnKJNtF3on264D3ml8jSrzmr/8Lur+pSRqcLVdfVJfk
xvB1HGehFAyCp5svKyd0RAKSZbQihfdKQNahQulZsoSpTSNtaJZjQkabTd0UTQrL
HavD1icXvN70OGCNnVP7Qbchf4C7sJIaCl0ftef9Z5clO2mZnvOCrn2PxUSOFzTW
xxA2gynQ6T0bgf1k1Rra18k1n6VrxWG9NEGz6a0ioXu4+SFA2u7JzEhrBSOEjpCz
GUmXL5ergQRxOxXtcKbSSCDKq5LGCy+Yu2ujxntkgfMS6NuZiOr9srlj7ktGN0e8
9sKwX2u8adrtN51u+T81b8y5dcVmKH1i6Q0Dx2fsfypO78h57uaIU00uaNg6M84F
1JcfL9tsFsxweqrmjdYATp9sNilzSSrwhqyJmZF8EqB/llbPcQjtnuWmvvrHufK8
opJL8XQaqmJq3l72Rtcp50cIkSy1E4bVyaTatiyG986bSXamriK1KAmeF407nnRJ
y2x9Nm3JHKV086fh36faEeIKniFwAggP6QzJdccQkVfBw1/GW3g5VA4tW54SAbpQ
K8wRLrv9e+/E8JXor2Iq1ihRQxbWfrqxfpEL4fPibyS+T0dnZGjAocRhHeIwdY4d
cuQgI4XUb9Vm9nJUcqgT1QY4mjKcv7CKe3issb20K7ec5VDF7ty8x5TLoyKtSn+o
RCmyv4L6hAIW7mj54SPfMze4Iaan744q72s2hFHSTF8bZsHliNZcY97OFK1XBdnk
NoBZfX1pSVbKanoQOyw+Ay6aRYHgM+hrUQh53CWVI1waNc7M1OoIYHbzddozA8bA
6/SKtJXmzLUn8m7hKCQ8E1GAF4S8wqSCsgtp1UqLZx6qgSeq0rEb7AVnNOVxSn9Z
U+ezxxfboKrG6LnIbtQ8BZL6rzKyVyNqvbz1iy8uJqrT1apCI4tWEotb6eFhoNNL
0YOYQFymn8XhfY48LfcAaFyOb94+px82Jno01hjp/dhIqMxf+4/aSimQ+R2Da2h+
Zlz3sBRLWQ1tEZS9BWcOojar85mBu/cYtli6xN/9EdjiZ+e5q00P4vAsk+HGEyoa
P76EwFpxUQuvd1oQmkD5HYurJXeF4nnozIuCk5wOgyiD+/ybOtitaSbxUi8xROk2
tuRPTDTIVndMkU1soEms5aPG/9lguzWxKdnxAc6nnzy3wtTYjcapnDrdvqYURvL1
Ncv1Jbwg1kmVzH337SwbNaLWTwdjMaQV8Kx8sO25KySjPvhxAxWfxuoOmMa+dGpm
GJfV6iZW0Lw8+76GLhM5NnhvMqxuxC6EUniQyxh5M0AmCdBvynC8qVJKQzyLxSqk
yauydyiB1E/cog90Afuw+kvQisQG4gwJZLVUO63gujr0DASy9ZWUEw9Azk+1vG4g
`pragma protect end_protected
