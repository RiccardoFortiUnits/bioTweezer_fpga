`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TeiVI175mrzBPgeaNL+eEqRzMhi/bggaWnQ+perA5bMNCpEgqziPlyAdwAFIH23A
6/gXf4jjCCn4/wpz4I3Z4T0DFvYbfqE7E3L+77TacTY/T8II2iYzudHXiufpW7KC
J9Pff09lHwulVlpaPrWTwVZY9xA5mUZ63fUGf3vO2qY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
BRXPdHY0tNL+kO7yvmtVGi4g0y8gtuRPbnk110FqjpxD9STknwZZMg3Qgkc2bPzT
oR+PFhjDE/m74+AzOQE/ghcUrhj6HvTM43+DGVRpFBYI1797mLL/iUx9n4/9obww
dnHCkKRRv48bX02QwXS/z8D1aAWB5pcqaeAxx7+tsg465ZG05/Nlt8cP67uSA3HS
wiooMjhTvGhDVPNBKi/7zjbHWGgrJilJqTLAzKEcy2agZibzpy6nF4rfTkYz9S4U
67j+CB9MehEEDCzjMm5UpGvy/WiQXN2wHXYrTCd1OKRTacXcSnkqREPQKo5GUe4R
mxsiXfssa7j3Xpw1d9wia/HN9kMZB9VvFvr6XGEvOLAz6cds3IFvVqPVK90HPC1x
LZPs0UYenJiSN7j4LmgAX3MyeVnmh2oMj9ZVdq2ktJiFLMd505E4cW3OmjaCkQJs
SrV57RptAVV9gX9PiyhbU7y+NIifmecTKGC0bbnIkxhuSHHBjWSVM19CtakIa16X
j9SZlsphJzfuPyuNSY2IVKZxqf9quIZkMshT7VRyWZx/YkxPvEEnYexlsiaIBpQO
y4N84PeNfMP+gGYmb2yocP2d31B3gCiI1r/7Hd7ZBjRrZZhKq+ARjlayjWYUBxbR
nz2cQEILBdLeN+hBt1b95ECY6Yd88x0QNGf/J7C8y22axosG7UtX2c2kfHDS1p+i
1X+U7P1UMe6B/p2OcFD4wXLP7xj+55AEJyL6j9eAA1+iB84nB+DbB/wSDoqtXSMq
DGnBH/AWb7gg9m6BaDtasM6oEXfB8zJRt/D3Czph+aPzMZIppay3A2ZVK5TCjWkZ
Y2vlqzEnIDeJ8LaS9J9GMwWQuGq1kxz8Gl3J+eaO9Rqe98145DEbsxgUA85S+VE/
I45cN7SqBg9+kC29+LWmtdd/93+h4HkQMOVqkMB+qmQYQZCCEXsJYfrqL3AIRk5i
wY15sHO4WQZef7b65vgDPOTFYqJR+EPdciT2yNUN+RRC95gFMfH84utEH2ZL29c+
Gnree7kFa57VFuzufly0VHeXTwrdHfK4nMbZSfcNoz14Upnc2/d7IpCksOQFCefd
QGfRZ5w1Ozjj6+G/8cLjH9g2Oqeng99GbQfIRB2Ch68LWfmRGOh4kLOMjyiwo7su
YM6KnRmLo+CA1KuREmHF69bBfSryVs5FfLsLgSPd7C6YuwKjZs0D7W9+/ywaRTHC
ObvxAi8ZxL+CXdTsXWXL0m7ngCSbT595aeABBMFpZKAsDsWS6KyRHZ5LLC+1Bb8H
zNL2+qazFJsPKayY98MVOmOSa2MkfN2s9XL7nnfk0SiU4XznPmmhPWWuCK9JAo6v
wCPFTjKV3FwZxDWI1tI6D4o2KEsQkPmOqttaLlxd+hzyjHHfW7RuFEmEX0M1GC2T
s+dQSnLrNNzVfVuA5J/Ccp+6ikW9JmQsIKzOwdk9rncyW95RJzPveRMUIpfV8UUG
ACdP1+cspKDfE7a6Pg5NQAWRwkm3HIqFgpQCpg+wN3R3B4N/t4fUxfRR//0br2sg
50g/WONusCrfzuN3t2w7uSywejc1FUNcf9TqtdxswLT8lboV5HN3/tGXFhgMMasp
J/hoo5AW4aueEMZviK7dKJOmIa1vTSqrjDPP9ZH+cs7uCZERctBbm9yknGD5PtzU
pGsc6wRAR7FvS5Bx6AqlJUQwA7CjcRhv4D3XoHkdjumpynxhrr7uvjuD8Ivwaq7R
4SCb6UlsnQdPVmH8hM9d60SAtWB026YOg/C8jGGtO6RERDGjFF7nAtwtAiAn7Fw9
j3TaMuEF0WgsU9CXInqnnTFy2+JcQrudd6H/0RNnzZflXT7nwzQwa2IVcqLdZNmz
of7Abhg3dgXgcimMpdpawXh+EO3vjaLsVDRYPeZD//q+6ZTTjo+T5jwdNrugeDom
d3/SHRDjIHyAqSpNqMvnMIqaJwOytdOZSu/uvdEIKhvelMwgjcgwzjtrsFYerJS9
+EmWrUoJr0beQGhnTanQ+An6GsBzOsyYoW8t1CbJgaGpJ8jY3CkRC5Mu7OiR14AI
moJTbyVpt6SsG3EZOrcIykhfw1bkDVCQjKJ2DDVdd6xNdKD8cdZ3QPqHOnZ4bDpK
isHzSfp/CunFP3G1T+WQzv6f+fxCx0TnSiQtDw3sxu5Lw7p3QfLMwkhHuZ/sb7NN
WtvWcQOX44axmnrHPrYo/WsLUjYVP+9KfM8fJyfnwDxxcgjcvd/5IJHsEv6A0Ems
T9U/7QwpABhAT/aQ//Wx94IZ1PRgsTRiGQ+VQEA7TENfypoBJ+T3QeOCo5G4U9QX
VHmJR9LWU2uJt0oPCzskQIykHxX/4dikduErCv+qrmOY5ybUXuXuCbYB4Pl+IgSs
OmEinywhzDj+qNu7yfbfopr/Yh88KdPBQxN8AlBP1VJ5pfluU3xak3Es1MpShjmJ
YO/+4DqnV7PUPV6eEHijVXkk1znarLmvJSYE+nofVSzhQsciSThvahQKYz9ncSWa
hOOKTY3CLpf233NZfJLJY9p6NV7RUR/keBGyc3MgG/CALGkhE6DT9ZTn/VzWIuaR
HQUTb2ajE1Ek/FY5+CiKAeeq799DPdom/xw9MoxgYzl4KwqW2mjyUmndFicARlzM
0muiE+JrdnJtmxfUmo4jTrbhnZJgb+fY4Olm4rb/ZgbvRj8YzHQoHUz7+TrIxlp1
n2eOcrbzuxrOllJzIaZ4aVqvAdqg5DDXh3nckgpZ6TabYK72RqB1tEYB+iQ1Uf1U
s26S4Dn8UBzwOUr9LuTbFA0l+XDDodZtSYdunnF6dHBZ6ANPwpKExxcrzumidrmS
Ez56MRxwk9mIEpPgEL1Ii4Y9k7UrmWpWwbqHa4SkdwJMc/KZuL6rUh+GgDDKBY6y
3IlYXdNmIuBXAhuk43Yck4g3waMUPPqfRQIimgNAX44HsR6HOK0qgD0/ik33QGKf
xB3dydCERNXbDjGmcUTCugRAtLK06uAfVItzRb1p/e1xGgALk8VjkVVOmf5Vud+A
ben5YJp2dPh/hK/884lRmnCMaQSgrg0rRtD4M7GdiHeX5AadY0pUbjz6UX1RkGCf
IUacUPX0YMJ8lT0avnoXauRcydRt4tobjwqcazHKbQDfkO97voFWDPACEIfeF+Xh
tsIhLv2l9dBsyA3MPbfHQ9iDrXelplwg/rcQVASztzePTS7y0nzi9P50pcz7TSIM
6g0++mCrwkd/Cu0SVvFS8/bsAouqPzGwWn6z/3UhAd3PL+iwFz7HLcdGWBRG4+px
fcnINn825hhwDj48ciBRJdM+gm0dqqDQ6hAcnkkTfF75Oa/74/39xsU4nvDvIHlu
+CWRcntkB1N43MNjLSscY2A7puKzW9CiyiLbnF475PpUmpzCr4R5P2FVphobMJ8b
vePGwvnmu2SdvJznXAH697YJIpbif/QFHnt8MjerCdtaEEzFP8uYF3bZdDazr64S
NOqYuKG83pXegF9IHXGWzcbGgNlvkDqVIQtM4W67RsJcgkxPXoq/4GMVn4Ju5gWg
8atq12WmLgobBrlIz1tspZdOXRMEl+G/Zw9MO42il72pPWq7/AmK8NyFgt28znVH
2L1Cq8TDRY2iHqzBpy3wi5+iKzv3k2m6zUC+L48Z/Y4FOxYbfsJCNwvyype1so62
3JsDldCX/Tp8UTolE9LdIi8kUZ0mDOjixeWthUTFKEJggPZKiYLT7TGIjYPHEpHk
Czf+CfZ11Tv2t+BFfYfwQRPqnShGBstxR+MFvGgAb/Uhmbv7cG5IlTnbElXDd5rQ
jESJbmWvYRpbya6H2DIgCDtKEZYI+8gAyAvRUBD8B3M7IqXW7x0uLUvTsVblrxJK
Uxl0sDVUr5z6tRQq9X9lEZEkZOSzqedqvn3oXAKD6DVnjRUoUOuVTNazEBGK81ZI
UTrZfYLAl7/spAC+1JWk2Es6u4mrTYPBQJ1KLaYvUozTetaEXHuR6/KjjYtDWhdk
z428Ht2ChCwBPoeHamcT3rJrNLaMa6HGG+Wndri+Hd3Fb9tFI+ayltICGYB/D0Pq
DUPk9lOn5DFCmSxhzw9vZPC6AVfBLcizk8oUxG1k3kA8JuPmjYWbdFAPrSLXYv+q
Ub3qrQBSU0Fi4RbIWnrIyXllmEPWtdKMtjVB77lb9veAADgsA7GS75UsgPXAJlFe
fSCVX9jKZz1PH3UYiOE319oG7F2MG7Jt7GhLIuDdA6pA51kZ/9MG/MWv2+kbG+qD
AqTdrF/jv+4vTAdIiQVnJqFhfcZdvlBy+8vas7gh2gIr6EfZSejGFA7w7o4CvKNt
eAB8E7BvPu4EZgM7di9f9CDJHOUA4ASAJUng0p0joRDEApiUjgNpa2tOYkaZDThW
+ToW7zzaWwuBcqDm89/dViEaGG5ZSmIo5sj2YAr3qIBHSuUCVsKrG61sZwaL1IY6
dJIplKMYlu7oGFUB26/SRl6N2bsa2EJfm5zfdkJUtogXBlEBm6bfixWHqOC7QBpQ
rOUDsrswfIKUowPUGcoJIz7AIGr1FnaK9qcHGYDpL/Jv5HeGLWW6BQRVCgwbYiqz
6I5tuIGTbnAfD0uyLIMhudmtHMw0y5X3VmVcdfLdZD0zQZjYaoLJtShXWDrXDMUU
tmze8LdL83G0IF7MI7J88kHEwCaBe7kXgh2ZkM/lGfxfBraDYicHCatgW9xyGqgJ
6060TNML/e3NUwsUuulmRSnjBCLUNMZvHLvX3NFYhzZMbN4iP98s2a+GWT30lfZu
D7zyH56PZhuPLXEJy3pVNyuQx30idMZUtEd1CH1vwHTJ4d5q9ZQ+zffQyt2PEb0c
vmMv72Dr5DvK2mxfCg6hCNfS+KexDCD8fxmjAGJagf3nHRbP2+AwgnTHfUEEcmr1
//xYmcKZthFxzfOKXMqYM5C8zbsZ7RIjvyK9OlbVzsTY9mWPzDHl0y+7vX2OHbHj
klJxlu0/VRucKcdV1gfMYyVMFyPixvScrw+0wQwaHGbE4is2HkpS70PX3H65PehZ
SPH3bO2DiebsCXYh6tsqsdGUSCSzs8pZqkQDoAEoVfO4DuCE6dEssBOPI50XLtfi
RojHYFfZvP4qc9iAvWLkZCnUlfHSy2AJXTYlFaJbp8G8XjxoTZF6GA5aMqEHfql9
28EX1H1qhkuB6PIXD7eLLhYgNk7Ge2Fa3fH0d6omyQpFXTPruymLVXs8OEwkDtc+
dcUTKxHSq2BnmrGKrdnL+oNNElUtJBzb0b3MbdqHSHxv51LWsSYrEOMrXmT+9mQ0
BZ/S3uJI8tmfF/FJ83slI7eWPo0QMCwCxPoIwCyTVzHiMl8P1gNmh1XwbT1P+Gs2
1eRQV1J1vqLc/SUqMouwbWXUKMjJ3gIFBBvdlvklXnE2ravU8pe/9AM3LF9uQh1S
0LA0IITlz8NkRIAUQFYBIMssTAPkhq6eOkNUZ+p2zS5RQ+xv5fyjgXv11opgWJ6t
su97ve9T7taUnJeWshLxoMlvedMwlgqZ4uMtB5RzWUHnwlIL35rQUbg1s+WhyGwW
eU2E68OgyrXo0M0ueQBmmailNEgSr02iN6XriCJhUxHGpzy6GtJT2Qr0R237j4Nb
FXC922yR/9OKzHEkcPcximPBHcHnVFyIepjkxw/CToUzZHW0ySvz6eqH/TQATBHs
EnAM9nUkF/wrqgwCZqjh8GDMYTTWIIipRZNKPrLFFvzkT5/F/FFK7/Aw3fkE7/XB
/zVFLQ1uwgxXgr8M7RCuQnGYOh5kQESP6DVDMG8kMfSF4XEonXa5zCWe8KILGiSC
uV3PKJ+BNfgQgvwtYOnCYzLdcp4YuQ8nTLET3Tl8PPNU896D6bH2WoBMoW+gcLzo
ZyMtNrpzS50X8D6wOK+Rj9bI2FwR6gxjaL0n87mxsYgIdzZmyhiPl4kTMbxMIual
ayrdOVpxLc1J8wR/wELYRi2bG2SUZjizSBsNGIje/vzRJWtKrF4GTIU2zBwMWBio
B983il00lugsfzIyBwXz9+t8eKN9HmSAJQ4PsvOp7UFJjfYdriFV1m7WBlITfJZE
AVxM3+nQlrV8IFghVcRCioUbwrsf71PRgw/4UdFQBSJOhId3W4eQHEd4g1Uoflxw
nT19+n/qYvDX7JYg7lgsPBt3y61kmD6wJ5IufYBjLM6c98XyuV3Kxqaq+8/owHyT
Xtv4PHuPVCPY880oLQMDkWl2/DOkN5ZHug/Fvzzl5Kpc+PkBfArZz185kI5auCDl
BnR8FLGC3TPQ/+lf/QhkN3njAIcK6IDJOaYdfS9NwxB8oURywzn2EEfDmEUaupoT
1i26wPdjO5hnJeDqi/E63+poOUNFwE/DYYKyyJlonFjHHzpFwn4WAUL7H5DYZhDs
pZVMjo1obw8WvGjIArBhq9BMmhOh5+nxYzuzxQssAPwf5BEy5l0Ch/ObArSxhwp+
jYsSTAvU86/rcTNvGVvsxXosZfEIrBpx2pSD2W+DkFAqaexfaoDv4pwVBq/Fa1tN
Fz8ag4rjuqdWg8VQmb0D6Sc5JN+tYINnm0k6Qzai3uRdtFwCI5sNM/DMAANfHYVR
0UuxTxv3H0v6EPm3XtEs2hebMfre06ot5zGiQnUHe66zOueDQhDFF4eNze0pVB2t
u/WJ7PooXxTTx0DjgThkRvgcwoec5+k3ksuQEsuI9nffmG1RDmanSV8whwaty+Je
dax702q3w7OY4JwVOCOKpGQT9M8jvltKY2QKSuLXmKzE6yOWIufLTX3W/XIRC+66
b41MyYF2t58E69ieZLrXDSbk69wDECQ/YLnG0PhhsKpDWM68Dd0AKm6pJmsPLl4q
bNJtSR37XCVS8elTTIpM2RB8eXLdKS8ls6FRY8TpKB0MBt9u5LtN3gubZgPODq2n
TwhH1oUeZd6bk+8mupQb2zflqpvU6EkdKgBNYnPg5aV651Mhc9zjbAwJIrpM3HR4
E4Vme407wvylgJk6aODfpxfMq3G+uJfytMrSjJ9dUpHz+Ti1BEBVzwuGyDBib/Q+
W7LZQNnqxLLdBBW/wBh9jlJqDAke+Na/5VnreGDJRqmulFV6qOpqKxIzehZv2a13
TRx5clLJN1BT9FyX/Nlo26JMtuCRClXWScKaM6H0l2QjYai+nJ7DbZdpzF9uohJO
zEv2F8c5rY2YaEahjSdKXwmCSb5eBXByJOrWz3zeTRxXqqNgEa5Y9mCs05PQfV80
HMfhgH8d1Gj1Nh3+zVmPlHyZbXatJudQZFIceS7jrhu7y2J6TddGUg7lVHqTXXF3
HlelPOJbxnjN4tzwXus3e/A5+hG2srfD6WUiJHlQMtkAAHjUfOyrW7hVyOGhh42I
xSRdLqxZZwHpqunpBAwDDFgGAlFIx6TWH3aneLy6ziPi3Wm5IuQWrSeFwbMmRCMp
Tf2K3sd0tW02SMDe95fML1ELhmlDURmQ0zT57i6NWjOICebMlKfOjmeUY0uL0KQF
q0ICNIdbjQw2z84TM1HG0cz/JgifnNfiYPPMcXqCzsJfKTcMH8eKJpxcm9JRCb8S
iYgsfYCQcDy0x40EzbUxsq2oIzV+tdeniFwWhCyFSU2MSyK7uQiVoCZE+AhuN/7E
hnmWoFMTHGp+Uxs28939PmR/Erkw/Pr2cBAaYJaXE9TknmH0TLUxMP9hPccnAToZ
/GKdYDEfHYlnEvAIKNn9sx9Ja2wR5xyBLM1ZE8Ctu40p/lL2e3YY02zdKLsaFuYO
58LnT9/EcvGzp9jHWzT7jzO1XVvX7rI+odSbGqgopVb0ciQueSO+4PAl6plkBJA2
bS0PAs1vK1/6NDkrFkymqj6TBj1tL2m8gehQy399tJELXCi5b46tdUTPcM5ZbkYH
CIGR/KCYfvUT9zxQYjNeUcYfMWm+U7bnqs+5rDjs5lnVvFPCwuetKYtcKGw3t2B4
vy8d56/dA0PUIJJS1g+WG7RF31M9YJ1Lz/bvv8DeBbw7M1S0/iv8bEg4ESgOLhYV
S3PwKDcbAXfaCkVnMJJjVcMh/4AWKkvXPGVRd9kg3+Y2EjawPghrQDadZ0rD91Bm
opzkgh9ww77SCvPGRuCQb6ljX4JbhJZpnMJj/0SowezBfiKFzV4tkKwGJDMGbqLy
xQrZr2wbxwmncbxfzn+642yN26GuU+ti/OXhmQq9W9LprJATIpPrelchOIIW6e8r
WncvC2GD+9pCCdZ0OzXKoFOjyZZTqCaCLnvacIzXx67vbthAXJLUsiXaPcGKSkYV
6OC2oox2CZHyLw8OnKrWsIp5tdgHQxjcs3C5oXkLADBvBh5OE3n2psmzHfesYkNE
y7lUwOBexXMKzC3im5jqYpAFlvO+Yp7X50wx24lTp9LsSt5bH2/sNB3+TdwUMxAz
hvOZfLoDsc+qKP0rmw8Imu6aF9dgnzT9Jum6ITtHrk4x9ktOWCLGIvmdnyJjg08i
US1T35m9spevl7KOJyeMl58qyfe5yKA3eMjd6Qxps/Yfn2tDAJY3l0N1y79S/rL6
pUf6UNtfCfafXBlgQrlSxObzVwerQVSolPQ5Xcje3RxuZH0zV6p3ooS3sk19BI0j
MzONmdLcNhjOKqG+ksE8GkEv+aK8ybugdMBdh916IN+p/OgZrLnI50DbR4xAPtLA
wNcYdb7Lfb5fWXzDpnvGSCNUIcdNvRq25MKnHIUFhzSrqcjippYks0qxXTlmkHny
wtnk8WVs7qkzogpmTP4NwcOXKYIKalUTN2ZKpEDKFIEwaUI8w+81YtsUB3/wMiKk
HdJOqhhT//yetckebhm0P4zVN9W9bu4RjngBMuXPDA0J7GyRq/upkBiQIYu8EjAs
56gI8DfQGxmYv2FnivjbIxXI4zi9VSzQtj3UEUHZv+18Je5ZCnece8aiaVLTsQ9N
+ExJEZ+n6pJYJ1DarirbXFGwBkt5Mb57ujN4VAUeTUBJhSSSr3IwLzh9VokDk1yB
ikZQ/4vroMF4tYIy7YiDQF532yMuz1sT3TvijG3T1w95rl1VFZ7BRBVlDgwAlmH6
o+RU9OaHtbUomze2qZplIfeEjGL4NwJJt3kXMCqAYxw1WyiKI0sPUyrRQjq9xYzb
a1mMD6lnoVwgaku6AqgHFcH7EkiyGdkN/3EVg43khdl4cW1oMRipQo+bSSJSfPxr
wIZ81zFGnGm9eN6prhZh0Ou6EhOdr+N/MAIiG/FkgnpxtTPd2c6n0pNw3X6wk5hY
8csEnIj/2ObT88scRE0oOdalfuFEI6KG7lUVWI8I17BqzfQRLrjIs7TTX21Cz5xA
mrtI9YX0xy08UAoO3vYUaPDVfvM2IClJ53xHNTp/dqoPBMco8ZWJfba0b4+O/nLB
+EN8nrvVZalKTO82hy9+ZU4VgbUPGTpC1CARo93p/qRp6UwNzTHX/An0aUOnZXmT
L2EIqckUEf7OVPqTkMYYKbojdUBRKFN/LI5w+jdex5fAJQiu6rB0abQgEVWmWsi8
UnDzaSkbnpnOg/+DmaRb5sf07PcBVO3w7ItrRkaQ+rYUn3H6qo82xHGI7d8vQoqM
vTvgsGlC3pzTMDKyHTPHdZv1orwDzQQEnaQlVWYOQ4AlT+tqtJ6eb6h9iLgv6Uaf
Orm5QJu6IHP/6ErAWBX4UHxgBzHapMlwhh02GmRzTQ7ljJVNDK8E4BFK2KRtxFAM
JLdOgFugFHr+Yc1bdrLJu8EeVDDz2sjIYYob/5sYOWlFIxvM+9fCM6miDc3YgFv+
6NP2s1+sDTOQJCVrn/T9WOyUE9HwWscy0ANu68A9lv1mHFf/4zF98etJq28dqI0c
HDcxhr7BaQIIy55vMpNAwFZgMXe5jMNBJSb2AVOHiUSR+UHgKhr8uCm2gyGj5dIC
k1SSq4g9qnTE3/gT0bstI26BoVE9nwOaeUGnJJgkYpK2CYe+GN5ZpWIWN6+H07s0
qjQkJyga/07VnEO/7eZtgrsjVj8pOpIsrVYCybXS174ltGSzb5DUhvmv+sygYMQ7
OXMgQQY3g2+0E1x8QgZ0HnhvjWKegPZPERKIr3kxy1Cy/8etJf9aRoHu42vgUtM4
CQZkwRxbvEO0aaqcG/PA3y5nj+u3Ka7JgB8LfIb291GmiAZ8BJ/AEzfhDc0CZ8gc
7HQJQ/qoD82Pvt/ihS8a6Ocs/q5eGskvDv+6WpeXwHUBU7ywVgtrm5cIgE+OPfrW
umwUrABQ/KcmN8Sz/o0XW+XELBa9YkWBmxNbEowQAxcqmRB2/U28Ke4P0TM+v1KM
c3TFru84/8acWrc8B8YrUMx8XchfcYtsnlNWBbwWEv0MeXoc8Dk7m3DmCb+b4O6r
E65EnAk53rEBmxBze5rS3MXqLzJhNfQgIeGiBDtT9ohDMR/atBITUmtlE0lP0rTp
bybEZRXYr0jMK/o87++SBNriQzA+I1ZjBu9TdgBZkEOOpBUqt55h7Kt5F/Itf6z6
ReEA+gXquCNCgw86GD7kNW6LqG9pwMjyRlaangYuXApqO+/t69eCEQjZhnwXI8o3
5A8ugnlajQH7HrwEGh/mZHH+mBPSiShppSUY0iksMXKg21MW2vfHS3e5NMvFlgjx
O4Xu8Q8Phj2Dex8L9Ewf2ZD3WHfCbu4ngvrt6pFWtmnG2OFBP6N2xytcbKFtVmBy
+8BJHYKbbH3Di7r5IefZP7vJoTG3357krSCSYxlqRzNVLiFwjJCnDizhvggxWIcj
7j9JHsohMSoUHOobaai9UIuQPZE5ysNjNk/IzT6v7gvL0S7auU8mLIfjVtLiQTCx
JZi4if0dv+38joQ28/G/P9Vibqz7/BbpG81Y/Nu9gcJCoxnpT+WINCkyPET4Z/+f
OoRY7/3lyVvGZ6INiHtvD5Qir4x0mUo+qLA1r+u3Xrqd2jY0Sx7CCYP+tv7qJ3Fp
KbIYUlRBGwnc3i1EzKpm+zcQoAvw9t6Pvvuerv1H0JLY/JF6e6KmS9DLM1sD99i6
xoY74e6ShHCpQU8l/Px5e4e3Zdmrya8165ig1clpf1BW91/A0332QFtAA9XABJbA
pmiryXVKg+NZDUnWC5OK/hqNvpaQdVKX8Pnbncd0sXx9pty0ax/zVb9YPVaA5F1n
wpoWdUcOWsDmZFoZlWffzlC/2mb8j0qToYNLW23gn4LMMi+cw5Cs7JPujMiSURU6
2LYrjtRlJGxgfA15yRL2H1wakR60NhT5o3Ikjp3cHouQKUHoxsJx8DjelrZmTpdL
0uXq9B2KLR+Ghf3pEzn8LqYj2oM8uABYZ8PPHwRUWA66W5f4mLZPl9auSPZ6X5NZ
MrERvr5DzVZyoIlIBP31ZGueYLB+H3R79WXS0xW8Ey6Nklv+F6DZDQ2/Ibx+/JP3
6mk28buiDGfzArtvHndKW/DdAbvoGTpncr0oCxAt0oCKw0Js6yWfSglJeUr4Vj6X
MLK4qOAtVQpBmjPRIggNrR3TD/WYZ5ZaDt4lVyHnixnF73rncBW7n3n1TgG2MfM1
8WFEckYOPfMi4ajNGIwYRgohRFkwxYhslQ71HcJeKROloWMIbWhYWjsY7P4zdxt+
QlMTTcHn3pod56OMJEAMIWVwm68Iyu4/ydWNUW13ssUMKr36Z9iAFEjPVQ9SuZdv
E8IH8VpZflY6B/yotaUyk9lymN2qgxlOsuMCzV8+s+W4+Vzs6GCxsYP3i4ZwBeUU
bm5c4Tgk7ViLBeZZZ6bum1OCu56/4gYGbgtvSDrk3w7cZ2gt3FZPPeF6eyFFWIhx
z+UF8kTB5EKsgLHCQJtt5ZimBjVuA7GiYCSaGIBnG3UQCZytG6OrbGRTaTk7B+Ip
3NLutQbawZ2UpJk6kSA5kWzFMjkJ3Mu3AktK2lxMC/g1sdNyv5dXx/A6/jseUXC7
1ompUVsPzybpx2fZTEt394avqrHfa0n33tQRMc11f/F2Z9/KdKY91NEv0HGc0tAi
f7cPNnAkSptR+9r2DnyRH3WM4AAUl1NNczFBeMB30rzwUMaJzQ+xN+DF7w6Ew7P2
xTU1fhTNltqGe+p7MlTUkT/8FZb4UoGbfBZ2s1sQ3CQ39Z1tqbVasTvnyHiR3IPL
izPH/6DkuR1UCojGPbcEtzW4HCtR1BuwkrF9ezir8Z9hMNv1yjSaspczxP+b9Kov
abwjnqlutSPS/rIKD04sckxWqEDDa7PnQf2x/YVmsZkmHosHh5d8btsxATLdVArX
/1bKeRUsAPYTT35yFP8Amj3D16RMaZBUNOXnzl5+rW5zqBPc3qC9veZyua+RQwET
FR8sLZfuRhs7DaQs1dSD+X/YkEsRFu5jjLRCO9Uo8oWH2FwV/Rf5frMdv13X8P0l
E+mljo8uqFDOCPTzODAZZoptxRCR9Vx+zqXdF3XYX/CioGCY9EkJSkOZX3WaxPXc
bS+69Xunun+6ViQrSIDW8VujC9CdCvk89sgnPJypa6yT10x2x14rvVl9Xug48ZIl
zDIBqQbwoAyQ8RnGu79BFqQUdyxuotDU3vxQAwNPk305mr+uYbASiERJC0WEc6Ba
0AiZUQEG55nJUPkvbzpjQbM+FQZKPuwrLBQeXVUMmZRA41pcj8dUd/XYaxS99juD
nofkuDZz2iCvl0GCh9hik8XnX0GXMjhWq36BdGg8L10Lv9GmpwqCr9Df+GCggQbR
XF5Dg1MxULzePopRiJVmW4inh0DCi7oUrj39ZYxzT0Hn0fmTkI3cP1p3AP+HzRVb
BgBdm592mxR74f9iancsq1HgjGXJYqnavA61Gg3cEhEzp8QUEUJz9gAve/WkMvg1
mmbFekbk/4sYlNkjjAUB7rQtH1OiNQW81lwF4zTEkYVGqWZdrOIu0jCI/TwS5Arx
Ie2ViQPSnQoR8zfp459aep/q7LthB8np2F48iWJ8oAWIrJTydlHlqFWeK5/XjiUM
eFqo5CqVrTb4IHcMa915Q0Jm6sizpJNbhOyNfbZrU2rYrH3ElHrhTWorUgeY5MnT
i0KH5OPtglOJzTTPGBtGS+WDFyQYfW5t1M+hiZbxq1OCooLp94pKPi3Y13wBTp/d
aH8KaH4kS53Nkj5oaWxNA83SswTZz38OJHVEqh4AEd7iUHAbnkvKn9mAEoa+hPhl
VOcv2VpXAlKMs6OuLDCUEae2vfOe81nARZVdmOM/FpURwqm7wF8Q20MJ99hgFXYg
JZfpB/zf2MyOfp7/DWNZQdD6dyPyOQ84g2bA35VNgLHYjU5QAfxlOfC8svT/M93/
c9pXZtMAZIqmSBhB2bMhq0UQxsgyehbUXfgdloMZxVU2s0Rbf0QJy4WQrCrMTkop
QCTtp2koWqDCSxko4dlpsnXKTeRZN8rZ74HipyXrlhVLbDCCsvf7bf1woUyDDJmA
ae5fCxTAiCt29ZxTwPyS1x+qieVBGvjPxXt4Q0qWEIT/XFYSiyGZK+crnccBhfBi
Cfibi0BXLXqN0OfXaaaOX0C3QMQyk7Qz+FARu9Fh3QMs2OJkyUg0DUSbehhw0Lio
/6Cf5xtO11VW/5JHJszFO2nfTyOHCXBJsXX/b+v6/fYuC11gLLJrfltj0flP5F1C
FMudkyEfUFlVt89bDdHJtQ67MmveVVqJCHT6Ic3Cf3poHYZ1v7xULEDtJcAIZR4U
RM81WE6N8hhk0QxCEtorDNssY6at1fNoDAa3BWXVH15SahYbHKM+wr4cl4zQYuWG
zWOcyPElakcoVGVn+EIcxp2gmcDr+tPVxPxgEAkoTGX0El8QGhREvQK65ygAlvPi
3Dawu8JuYSdoPncRZt2S6p+JTeYcczuWbD7tiX0qv4UpZg8Zv0VEXG0uNUReDGER
advDwnUEAAh9QtWoLpQ07b/8g1UOoea3CA0K8h76bGxk6rbgukQD4MOTX8HHC6Ax
8XGROEQEnVWTfbGLJyt+XQH+syOleSwyrTIzZgWmep4xshvPVCUPd5GTdABpBPh+
msED4kKxq5/rTh3wDV+3wciFWGDxCBn2S3craFJ2UPnO+CPEfaWRMW6napyxNdzt
iUQJuZTg/b2IJ5/AtfRi55KfVRmcTGM7C2anEYoSejGi0x48A9Yn5/KTPkoDvAob
fjKz5+3V/l//yj0Nis/RuAKd55Bq+cZcu2u8s89n+H7Gk8M2HkSzwkxqRR5uwDW1
Pg63CTnNTbO9vbdz4I5KBDrfIDPtW13/ReT8AKijaStgAn0qaSgZc9y4x3AM4qGl
g06SD+xiSFvKJEE235YRDKBxL2T+zzTFRiZFdW3uvn1izTHcV9cAfwzrlbWiOWHn
xXiGR/eZkQFNfsDEFhaI3pgNpn3jpmf/nA9nE/uluDWoJUPsWwiKR0TAyzH5okw0
iv4q5VsI/ZbFwmIEAbJWajmGyCJix4GCgWl7dbb71Mav7e710j9WVAceCQgg3VHk
IvMGz7WTBQgbrM78TkVbNIh6pbxHjDUh1SWJHAlg5m2TGMlSzunB+jfow1qrY8R3
X7j4sdRSvsohU0rYHL+2RrsI2rjeasFJhGcRq9dgpodP9cwxiZwOYK00QMbsseiq
wduwqeiiUGkL84pMozCLjtnRnjTrjl+ky5xsUmmW5gsEqEIqcD0eEU9FI5ktM+fq
1RjWAE2lMTOmjozKnSr2UTEg8ePrXyyoFxXQWSF1fjlH4Z3mkIGwp4stby3ZWXRA
bqshQkfC8i+63VeNwDF6z+xs8MzIrXYAqQL9P/ZDstqZPwiUViHNl1AqWcqeQuMq
s07rjkr+wM24BkPHzkmsd668PYsYH9X3CumS4El5la22UNpOc4z+txuH51XsQkMf
vbHjjqPmJ0yqM+AYUWISJXXKA41zD7uQmlxmVeUtmM754CBG8ktrjVzUsdk9kaZG
Tp+TenPNLBzxe5sUZHX5HT1OJsSBKD+1kNsusKJtC38LauSYsWAhh16hjHmvnoP+
S2V3VLmT8DLEoYfPgG7FFQmy2LlnTAMkTxhUkHn2rDlPFDxzMK8tM4TKyqeI5VqD
84nOxsPmqFYJqBl3r9YNrxB8PmwfxHPg3F58sgK1IyqqLAucLTXTVNhXwL2NGyPv
LwhSHvHmUVGC+I0IMOr5WI7CUDGOUbcANa6IwjfmvelqYeRw5ftMxOk1m4GNd42o
Vmrh8uF+IADfmV9qKAHZfUxlgKS/ZLQAxjRlY24uR7KJ7rTq6iU/ojoHAabQdsBJ
qRLFbVj3RppUjzXEiGsI0KOY2wpMCvNGsuoxBz1M3BkiFhtp7CqIvDKNkldBP/zu
zdHg/MLzJOIFPnsfbqYQygwcq8syZ8Bpu+fmnxPu7u3EKgXPcAsBnVMczvd2i4w6
mTbvcuum690/CVg2BIsn1oo0V3uKGWExe7hdsmsn9MaxBSFM1d/RQOYnCttyahQV
50q4vEWRzdslecJoaXVzFJDZCRTbIRFJSDU39kt98Zznumoyd3w/jGByBHhF5TiX
R/VJ1itmsPjYsJHFMbQRCTAuihiNozCFs37NV1sEvDSsCR+PAos68VZypzAlY4TW
BxvzO4rwOu/QlmiH9+mhGKn/O/d/C4qZ5dXYAAt70Zd5a/GOO3jhADdDTuDsT8V/
hfUp/QaNek7DZEF/Aj4WZC/adbFj2nQyXrkV3F8gh1SALL45itPjKgDKZMdNXh6Z
KWaRD3EkIRIsqvNrCi46kAjLfvoEMBEbZD8tR/y9V5sbv1YPIxxpHwo87DAOVb09
XzLFGjV/AdnLZnAFJv7atGuVwukFH56gaf18eNJrNJ6eO6V04gFKLD4teaCBx7J8
LiDLcF3HOTgKN8YaPbBhTs8UlrMglVo2FHLfJsuHdVw5RS3NfmvR4eQH2b3327Q/
6fxyVq/28II81OCRh69zagsVahnV/UsI0odCIoOCoyyfFi4CWMP4okxPg0SN7P5b
P0GGXs2ftQvmsC3FU22kdqFfZGAAwIbpunzsG5WuNRIj562q7RZpE38qJ5/Vzi22
+ohVTQtVZIYPPB3kUxq3rOlcKTEO82caYGuHS+669zndYcUUvYdpG39d5AFSZfSs
XTfhAu09UUFPWBqQUVKxcnpTDhd0inFgKSLMFlIczFOzocz6vvRa0sbkkAPFZmxz
5uSX30ff6faviIRaJzy6f5tcl+yL24G/au37AIlPCdkyySGyxaQ328iETCXinLdh
4zfL2e0V8VayPv0URo/3iYHGQvlXuKIPO0Pf3Sn+qiZNaiFZMtS7XjsHkMvWmhUc
tJa9Q2jZ4QL2ngBRl77OJW1Dfi5vnnWe2bkU7inCLl2qzFQBFVt1cTA3m8Op+sOk
uKcfxT0fplP7Pp1WYNtC3mkZuXIQjdWSpYYclNk7uDfnFlFCixg1jtDxm+F8TbhK
N+2TuCHDmHWWAUAR3ST24Fk6rWtWaye/ZMhdLruHBGYTl/IVeyPNzCV6OjxrurnM
ndnmrXGvxJ8LgzkuhgfCEj/wuygY3Wxkh9nKpXr1T3NqFlnW6757ZWQX8Zq7EQpZ
okKkQvUBnrhIlinLy0JnnoxyInuuZ0wA5RXPwKeFHiiFtKqV1ILpFXR5l61Jt+MJ
xx9GEA8JB9EmApfNUYMjLIljOTAo7y6jubh+g9dswDu6X2uuWMCby6ACIvuAdfcz
aJMKKnw5PV9jMwi232Nmi3tU2XbfhzJodWOu9KjVVYSiDRPx6DH5iWnJVJ1Uybht
xYXbEelEoimLJRyXSQLiC/fWhl/UzIf2AeDCNmjC/sH6kn5b0Njt192PZSe8j3Cw
a2gGRsG51wDUMSJzyJHl+WxmEIIhJakdIv+mpBJZr8nu6HDRmUYKEXy17Wbcjdnh
iSHArOrOHZdEg8wA6Cc9kVigJpEapIT99Bs7fbU1umymq8xiQbAAC9fXHQeU/c8a
OuMCUBn+qUO046zoSD39q15SBsFq0Z/PkZZa2aVm4GjMN1AKbDMxyDQlhdbWOFCi
MYi5OHCfU2YFFpk1PTx0LnGoy+M17g7SLA7g+ovbeITz9nTXVkM+aoAAnlFD5Jp7
S5UdqvGXalmzVm1sOSaeaSlnAQchX0RzdY+p0GIluXZVvehql7tv8XNfLF1qeVjQ
XZYG0ZcaBBW9oJ7tDg8s8pUleG1lFe+lxSJrP/lgaufFJhez/tNyIXdtPy5gcO82
3D45fbL00SXAUXUbV81cMgqM0RdkERLQlwk3X5McCFD1dz+lIcBi+rBIrL/1YmWs
dB3KogS0yihX7yYKZ5ansIIAcwk2/ShLvJTzPO1Sjd0tAYuWj7i+KBrSH2hHTsrY
IVDzYQFQ17eqQ9+zG10PmF101jNtz7r79rk6+sY53Pe9C5WWRn1VAQ/X/VzArkoR
/7V0pS2jqocOGMVSuvtfJzBdcUANBCeCzVSB1CJUGHR1N5s8gAeqcAyyk7pe2tAk
uQAPZAHAZ0VWzFx3YTlMUbFW9XA4Dvl7eMV5h6JY8rLHbQolc9dWC/TD9hfdfYwT
fgo+SORLR17a4lPQkXtOydmZBJerfRBGqnJxqvoSsyahVQ2sN9wimiz4M6k2yM/M
lApoQ+zeWsfMz2SxyCPCoW2fa8LM0IjGiuONQXoW4ONMjafQZMGpAem9AjtPmz4J
B5QVGCi4UVrPu+E3dJmWQbyDD3yy7w6FbVjDsJ3ae9R2s+9xJIpoh9WFdHYn4wMt
tiEgKjJE/KzEt4JvWAygeMLiA6LXvtqKr6PncfvlGmHeQt+KmCqgsoYO0jKQiPWx
lYy2e2U6VW893jAwzpiIhcWLYXrLqmoaAaE9JXBDEfq+l396UsCxR8yn4iMpAi/B
/gL+cqU0xlkJqzRryJecWPIf0SrIPgMdcBVwaoecnaL80Wdj5i4wxV4+xr76Td7V
tcBnt8ocTiHRL48/DfjFeS7XTeI7Twlh3PAyZE+L+kpo2BUHFBfF8PzWYWKaqd6D
P3/ow7F4TungzdhLiSRB6AUEgxMtAA1VyZctmFEvKFkXlBKphQ+A8g2UsFQS+wF4
`pragma protect end_protected
