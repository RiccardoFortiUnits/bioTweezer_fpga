
module sweep_clk (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
