`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W14+GGRkg3FuWN+utudFyR3QyF2ZV2EqwJdWy7jfps11OLm6eDWwa2JkkPNLJ5rJ
2Npwg+8OuubsDM9WF8pSNdXjlytUdVf3UKpmJiPeZzEUHleGkU06T7basnSt0Z5+
pU4aIT6Z3pbNu7rBprWdgRT5oTKgt5xbfzXToQPD77c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125456)
3hm3vUWvnPkMqkKaeHm/Im9pt5btY3M2trYcE6CuHypEL61/qV/1TeSxtMSH33nF
RXW0Q9gcv+wVOO1LiKuko6nX50gWsGf8VhoJInx4h8jEErx8FPkC55n5UypeJKhX
dSTEmXtc+5fHW9Eh2kuwRBOX8ewokOHto6rRDUGGWjAEP9CORHpuF2+bbR2awVl/
TYWQzd0OqeaRIn5SYZD0xYhkmorY80BThYkyrtEnHlm9ZYpBKN7I6J3ICnPTusun
sgfqVUgdNvN/5OcwZD2DS61TLbe8z1wvMiXfGcNW5k1jnL31X5X36luwsTtzpuvW
DYpxCPc1m2GfKqcnK0YkffEpUy1kvYwUmt4iOfqL6lyA04biRgVtsWlbW8CGV6ah
mIhDCCrkwQVH0W2GEfJdjpfNqGbRIAd4F60f4Qfhsn24vF4heDoRZ6ON14KhftRM
vBr7swmweOjb6PfNOs31kM2T3bcn2MO+6D8k0ACuOiiE4QZwa+6PXwbobk6Cq8Z2
tUeAY59oWuq4fP+2CX+cfFRdpOFVt0ihAlkgRSU5P/bH3E/RtbSgGB8G6S1hkCey
g2f3+QPROZkmrjGCXsd0WWLqH1dGEGg554PAuTDjxVSps3kHYaN49GeJsymDHDhI
yHGvYYQEHxilW/F2C45MzngX1IE6r4ayehvtPL78UAee1o+f/ehTbg1d9w2SXmft
jLi9cH1mIcmdvpGqYazNdbyrtCBGcvTmVXdnl3/3PsRqPdysfN7fDEEg+flhacfk
McoX/2wygeA6AG1u4sSKnFSO1LsoJrMZNkYb05+rMwX/JiUHVbG5af3ZSRwFuo0G
XzPXqaF01OfjHn0PguJsWSo5e4+vytPjM1rT+NKF9yafLD8oSnCcwtOMg4jR9PcI
HAyGLNHSwGGVQR1ky9UgCIIOokRKoyhvr2AW01WYgkbLqcRvgFhZjvXEA/fVd3y9
FxGo4eRuqzynrWX3gT6ESuvO6zIkAOxU9IEEPBFjWdFtIurku3/3u7teBKF6Mez2
ymQU8Pvy69/meqDbLl5MAdVx4JBUqePMOWpvyImRErOKZCVsSs0DdMon/RjpzDHn
0G+Lb81yNTHHfM+kFV5Y1oxmOP3RgnSVY6kPgtRKhCl8hjU46dm2gYVA0pOl3AcJ
6BRZTo2EySVVyA4Xe949tbJZ8kEqldCnpa7gpFVXohVCmwdvFX8KldP9gIrOeRGn
9rt+TXO6GiYZaIvDeYLxPEbCROLh3aVEVPD753Hq1nWgSSQ1MLST+e1dsypaaJob
2Lko4qmys0OzIDpLmWtXiEEyPYkwZYzizTOy1AeYlDkwLvPJskaPLiPKiLB9zmEi
GUwvutNH5b1lkeUcH1aJQdN7NrK2eCOEeyUqV1g+37AZsjJr6teFXdAsvsEQubL7
ajT9gRW6wkgrkxJ7TWrayCetLZ+/3Z0wDegYeWdXpoILwGsYHc9M5PjACOrrNsRR
wwvqqulvafXmbPVoBbGVUxVtfF9pZvkYYNc3Kx6lSaD+fTVmEmHAup5a+ajIwFwD
e+bq4ujsFfr5qCZ9DERtDCtmL5rC4RkqCA6dAJCz2nKxJ0V65ndNbh3ocSMKKN62
EVO4h2pcqjMhgqJtyexoQzSKzigRdcX6EEX0z/GLGkMY/lrshCnwu8ac+nfZb/1a
0GNS6Qt7o0KdADJfXQzFCuRgbYjbcwSuDTm1bUusjE2nBzKbs/4qhFBVjbRBCpKV
f0gCr37tJOsdkjsgvML0DOi32EOYxZwye4tcaghWs9NI+b7QE/n4TadJc/cKyc4r
V9QMpNfECgVUBCvAwKDf+UKchablrMkNbFrRWfvu4Z+U0r0ijdxOYyPWUWRoqn1V
5jW0VqAymAGPD4czBQyE9qwmx9RTijne5OfRLiwAtwmSm9Ovu1jOimjKIy/t5dlq
judaMd0hMQuBqRmMimrvmcIpJwkocgNSWKsf1wpcBFR5qjUa8+dfrweQAsf2kpNq
nucQqzqM7D6YyAIk1O/qENt8gAbZVptXSZUcbicZbdkEI8ZAPD2jW9ZH4j4mWDAo
9yxXGTy8PU68ALTq7BqbOBZQ1wd5W1nFrsTquLKEicYLLnT02RMgPkemvfJsCyJe
7HpjmPHFAw4clT5MG7VBpsi2h2r3fIqghJSvbzjvi7ZToC2RTVvA1jloIp7/p1sI
hq4NSKJhNH/yM5gLgRQ+j/jUmFdZMpQUkYkNHxdyZH2eGblGw0zVsAHAnQoyITex
iC5x7whfUuDfFgImDlK7J23NQ40pLhX90MzK9mporZGjuhUNb4cDwNfmlFXA23eC
Ei1X70lKqtNhUnZYSzB0tVzs/FdM0zJZz5DVO9xhp/vn+hiuqPqirG2S0Eynopdu
5aIeTuOgt/xNgRVlDDcUwyV08FcYnX4CAhRECh2+Ih6osFsQQAGc8QDPgwEyJ0jM
iibI9ggCm9qMW4eiVqMMf3zCYKh9ztMPxnW+utDG7Az/SsYaFDi321/L+7wkLPbP
5eQyAjV+uxHr6J3U8Dpg/u8u126qwjMqLoKyBEYU/WOwJSRWckXewOv75jziLqvh
EHD+pfuH6qyWopQnnRGaIOzD7fTZg2cSVN0OsC1siNtwkAHd0w6rqU1iLkRrpYjq
nn4P75Ed7BvvSTAm4KvrTw3dh4mYhxF57fDqyp5UKh299gvRCnpwb7ICDFx0IGEq
2LQbW/m/1dsSOqXcwsWQeD2gCmin2wjB+7jHZKE5qqz/+ykk4I2p2ukSjbh4edU/
We5feKhU+ugQgy77L0+vdwyOyKav4vCWOs2h+aMN99sxQssKSlP6oLVMFzpA85H1
6urxEOcQ92baLKtTuzbsFDVBE8YZWF01+04C7eQM65WV9Ui9o+KXz4NOYIq1IV7a
KT805KKB1WxgDKgzOVIszsS8Hm9XxTkwMhd/dKZ9BVTgFfkbut2M42QuEpS4xyyE
Vv/Xs5NGK9adA3xqZCPkOj0fu7yv1q+xEHYOaRnx2Vh5hBoaIA3mblv7Y18svJAp
Q6Vw7lqqT7nSEO73oPBY79ABV0x2cX+WIKZwNB2K3YQSvEn3ohPnXSp7xFEBLY1r
vblm8lCiLm6N595qjm2QMIjSydsiX3KfUenvKQUNIzkjWSRYn3FFfpNypNUWLSNP
2BRMZib6ye5ILnLvCG7OnPKxys1du6IZgMW67+ACjyl0+fOY4brAXhyX0BdGlskc
FeJbzaOkAHizl+j7TEdlg8cBcuRL1y8eozZYU0X4PavkU5uBMDD7Q735DlswFf8X
3HvO/BNvhC2WTPwUuCE0a/EPRw3a1QqHYodxfA/6CsecTuRKD1KzLpvq9IAz10fT
7HU4dK1RDfeAOaYQA0oxt5suEFCaZQ01rscbdb4rj/wmcFkBpQSjaOIOs7UskYUB
wCd7is3380S40JKFEgVGGAxUYXHKszh+S4axUOmFvJF4itD+ECMUATtrTJRp7FiQ
GBxrRUh2NZXW3KXzXWD30onPvxSSGGF93pkJFEbUiOv3cRbJucGmutO9Em7NWxhR
1xFzrmnzOPc6U3pHVTQ+uUdKOnBooP3KKl65lIgVz76QnFSyAgDknueEOYXZcVoE
xxvQQaFdw+KpccRPFy3cAENw95NfHuHUNIaH7vpGURVzg1ZVn3RJ84EqdRzlFmD6
FeAecqXQf2A+QPuBSxJxJkVJJAl29Yne7CaGIvbRXz/gJvcyxc7kXA3VPV6A2rFF
nxYtTcqYrHp0IsXfbrGByzxvLt9d2ozGlJIdpYmjC3ohEd7M1qdSxIOHxELZFeuH
3hcFyrODc3OkotJ78nwUpxunNBaFZbhhCeBU2K2hLplPC/AjQ69ZmVy2OoMzFqeP
AFmbaHAFFBvslTItAFy7Ej4zGjBbkzA+NEQ0l5awD0j8mp63XyS9fK1QiW5n/wbo
DX0yT9HK8HlmVOGIZ2jorM7m8XvEuwg0tOiJ4laMlpuCjG+fHa0K7TIpXxdZ2qCT
UIq5V/QxQMH0SuE50wi/SvWF8LXE6S5fmpMHQx4CKSAcvXWkExZZyOF9e91hzYAe
utmMStIiei7HZ842H+IJcjgEuxa8fL6//hAxtEUOzFrWazbLgOqSY8+qHPaFfLEG
BGlNo9NtD0nt3lm7qhSXdSqHOcAXet9rYAwEOEb9032TCMtXcG5s7l7ZKGmdjTVz
SLsD9+TT2XNY2TeJFGpEhNfBrFYF6pUFUvktijXl3XxFbqwwO4W0Ij+ALNIlyQxe
6Si/ATyviC3JCJqzcIPH/3qaG1HikLUrSSvwFUmdPXIld5fsZcmEypq9p+UAvbhK
JGR9j843dEx5w7xFTjObqrulVHD9LPgsTI1Ex0AofLLzzcXtTTLxa+sbr9jfT3k5
nA3cEbKShPUT97z2ihUBstTtNkoK6ZaEiWgL9dkDDaREqCw+PULfbUXMyKMvXRKI
2JNVwA62iL8HlThU1wtepFM+JlhY5avZba3CSVRTzujwp2JOU0mz4GnAoKFkSSSP
nJfA4yKEmqj3JLDy4gJYwh2zwXEj97XT3lVjjflQjIxldTCaP67jPIf4ua8FBAsT
tMFjSresaunM34zp+DdPDCs1+Sbk2cYVgNb1c/DNyzkmCTAc7SKucG+nqyKkj2H2
g9HR3+zFVaVXvVl+CrnQ/QiW2ku6yUnkIkikif6tb2O2aoRUld0BguNa7S8PF0jJ
K2/6VWP4k7UPbObz9rfB/hzGRV0VSl/jMWuv4ueWzu5QLgTZ3sINkFjXI0lf0MJ/
x5i94q8SLrLcecigMRgrkOwKOMIut1blEDM0lqi2dZk12dUzkHxf7x44Ma1waTfa
ZBBNOXaAJlLGEwOih8c8JxXdVa7eDXq6NEaud1g6YR1lprs+ax53qEn2hOwPg2PN
Yud2LevRciDx8zA9RC6yyC3kqI1vlEYvBPMKsjKKN9svNDjVY2nzvR2mHOmGNlI+
w0RKXgZCUTrETyzw52R4LQ9WZ1m0DMAkh6DlgfQuUzRE3MFWSxYV37sbsjIgiv8y
qpsnehOmiIwATiIQ+It21Edvter2rzkCF24tPFVUhcwBEqVkNQ9A2vTkmgaRy54Q
p67mw+qh5vCfID7lZ1DJCuBg+ojyE6WJdjvgbTqqUbJEs/cPRZEneEv5Py4J4lLM
6tSkZgwSfk/vWSNjwfs0FzawjxFxPEtrZCWGfV9ImrmD9ULMdySk0jUQpy9UyFPW
NrLyQySWobWFX4ulnIDfyDFoVpnQlUQLNG/ldQHAQx12gkOmzwaKbDx9VAbwtmIo
G/JUoPH5vZyffkRmf99kBwpE+TpD6vems/h15dA52gGfB+943pP9v24ZmXjB34JE
ZndQoJS2CNtrYHlNSs9r53paPzbkr/QPiL4DmKq+4sz6TMeWzcwk6rEhOUa0hy2l
hw/B1YAFpsZaOjZKLiofm66aR3yrm0UzPmhNJQR5Cth8kri9yQO+Fy4ThYVcKvxd
0zfX/yY2Ye/fkyR2/tKbaXthEcVrx4AoiK/F0uAin6OKWQlWg3W0o3k70zxblJgL
/7aKvLzIY/iYDVWa+dDQcKyBTsh4lGVu9315+w/o78/biCUKRvRBN3nl+d1focLj
Khtr/AOszhSwcspLJHkAacYR4L6MRpSJ0BcOisHlShYpbP0IZIh8Xq8Pv56U+CfA
/PcDoggNlJ4ngcRxqpJPAQQugm8LisniBtg4Ma+AZkYwVXT4RCbnBkUKuB5Tqp8F
MfKu3ihnHCoD069HZ04/ruBzG9ZRIO5MIFKPnZaGt5ptaAbEgKLjUKsSCugRZW/W
OgQGy2JPIbPMoAHb+vuQBFA0fIlVuXYk/VtWyod+bcTOcwOqeLwVtjyuNygsbWA9
lJfxDtFbSgosoNE3ctH9YXjeMz/hVcvsEE/014pIxZztM52OX3vkJlsJG41Nt0Qj
qOYaxclsY9MjAluOJx6KpR46t1Q9mSNpSdRqhDXzh+ZzfzARF872UewIZMcOMMOd
IxtJCxgsj/dlT+GYxI3Y14grHxACvXYQ+dqlfRYTMgI+vS5dqfSP9u+zuJp2qzpU
/9YHmjcVVKy6X9JgoToVc9Ecp1ODY2iCx6XM5JehBGQoSBcS3ATGyQIkGCP1N4mF
xbqRd8Z6hp+MCeOJQ2Ru3No3rVy63mjX+r8UaYQqAkLVTe2+8jDE2JkXq1Ah/ekW
3FryBwlfb3IGivo9dpCC7uVWMQU7ffyq3LsF0C/y0K8LhojXgOhzxx33AXhW9oRe
YDLUE7uUovUHgDQjbT5QPI3iGzno/JIHP8qmzN5nETIDr04wioMr9o1TnKTMszMX
55sLuQjnPrStXV9/w6hW9bCxEoOOcq8US2qNAihh5TfUodGiHKQa21dkMDnAjFHh
E7qt7pa58B5YZjny7d7xVOxjXJAsQhx3yEq7bjoCSmk4ul0EI9Ufpugcmp4Y3ncx
7195NK74Y60O+n6ApGFF6eawuIa8X2I641/nzaZBbBswz1Dv4bMFNrJau1gqy/XU
hBZZVf1tzqkN29jrboIYOEW5X9dt361vJqiWPyiY6na1jL0RYhhSAGgzPMoPQKYX
8kqFZOOiEHYdQ2l/8zz7MPtN0VlJXsa22Ka2cdMv4uDF//b1/53+igYmSa5pxZrm
pigp3+a16puTFbDjiVrAjvjyiJ7GddnRuFWdOXOEZdj5pRsuMiawJaUD7UkyrHho
TOOvz0vmAi/dYzcn1jicrWdP3ywSERSuzJEVmO6ZNxVdvjqwsrsr505cWIBbNfEd
5qUNRYutiR2oVS5mSPc+2ferrcSTD8nSsEJjU7nJ16LQ0Ug+usP4lEGqeRnJILHr
lZe8i2Rcb414NtCuR5R7CgWVjoTAa67MdOV1dlLIyFRr1qzXDPDkYifDBHgbWX4K
sLAv3n7B+c+WPTBVc0e15TEFM9Dsq3GGppQ88I4V5NwiQy7GrIV0xSaP+9JfJ6Fu
vAilUdhq5Ah973RsRi7LgXQs7EUv98Wcn1p/6Utb7y5ykZOU1UBp/4W74jWmehrj
gedIFbGPYpbSaFrOTEHFM2gDXVcGeko/fdypfomulamClZ2VdHNMOZYIDI9V8fFj
qewWW5dMGE/dVZokLI6dzWjHMfV8fOwFgQ/vFQd054RUZqY0a+ElLzmd1PnaSGCG
/SskqsqlUPDTLYhUSCtlqnVGd+3BSiat818X/6V3YRp2CYZv2Rz/4sMKV2tLppPA
lg5SjXZjA3wWltdXG9p5busBBNDo2RpiFM75S//tTAM8WXYRtYZUdGYiNUYxupNv
f5bjznLIrycxWxYnfCy8X4814P974RhZpRwi1CL5xPxDEsuCdSJa923owF5s+mE1
6P/fuly6k2Ux7mvRnkdHUq6KOLFvaMtFQ4JPB/MoK/715V2hNosxPpWyhSvvt3oP
QdH2tg7qbayn0koW7twbvU/M4Pb12QJZ8N5c98+8cwTTD2eVodOwF1Sys2mMQtIT
FQub8jp3j426GzQyys6j4O06h/QrguioqYLDfhW6Fh5f/8Bb2ADu2AEz8vdJNzKc
cch9I5uSJPCccSb7aBVMtEIarTqQuSpuBDKQ6WV5GK1kg93mM62KlM2JO8M6LjTp
5HCErK5ET+eoT5UyDsDeDx0wzmzhpyJvWICmRon5eAq9o+e+fjQBG4zBH371CK7J
ewLHLBCNbWubRUrw/sXE76N6gJIAOvswvrXVWCiQ1+xA2105Pqmour//aYWNxduM
QcwQzkrnoQfQUk4LDGncvM6Kygi3aLhqatxhOAjVBd74TvkzVln11FmUSmjKPhfI
MvQkMRXC+dAxzIrx6uYzEeeHc2ApILa0mkFpXmvZQD1uCfikr43nbdjehX/Rarec
bjKf4pD55JDcSsHO1QnDbCUVyxAXX6vy6UU67FKWJ648bssAwHMkOL7BPHC0o28U
TIOg92OaojxmKnvJ/qaOJq9QdsGyobuLVCtNkj5by5hPQRk51UNOOXak5pSP1Qyy
rWssbxn6fGE7aDev04MclDQCyA9WrSAkXGAv21hvAGNs0s8hlPADaK3U7yKM8YU6
dopeCA1ZHCVIjXtAiCnICU8WqtlguvYMa6bqdHs2/4xsny/doyRJyKPX0fWSbB86
4QyRomhgN5yQRsiqWtlE6e7291ASPaY5/I5GuRcQ5rXb3V7DdhycYNb9R0rZ6Vgl
zGgQANCqdaEk0RpASnRj5QgQNN/qplzB8QL+bSj4zMbLu0DbauXgYQ+cwrDqCHkz
hT8U2/QnIe28P5nmSDBvWnT81H37zzcANFwXx3XiHAWseljkjlYq3qyOobxw4lXU
DSL3Lc11FGzzWYAw0k7uFRmaSR8Ow+7NDFODaEHTE1WFO+A7xToqkyChZ64nPrhS
cb9Z0/vbWZxJaTXRyeBkYxiG6TIq9Nes/g8Juxa4gZJMK3hFwV9tGBMmJ4Ti9nM6
jC4FcBUoVQ84HvIzRf/Lb8A//f0Kh3amS7GStQAb4FzTGc2PQlXt8Dl5OC5HI72n
pGiTuseBBmjH0P5Mp4B+imZujJwJYVGoXMRH0NXX9pgYf+9zC88KklnH4LJW54Re
C2qd9c4l8th3vfx5Nen0B8Hme1Psz6MBdOHmC32WRwjcY0R0khdw4xH+jNOLRweF
EHeJ0jt1iBiDYVX3WNbjTJvdOdsjcgQISuTZvD1w1TuY62hxFIXpcKKHgvBy2Lb+
pb4FqPlYNxyVqtpQVTZeGXhjiEym8XoQDf94SxgWT/9fheibejFTxvrGzv9GrnG8
bdQDGL4obVpC6hRGJLTwOPdxg9GxvNdK1Saj2QwRadAgRaQv0abDXrQ5rN0mnrLA
xOU4wZoeWdtO3GB/68+v5RI0RWiJfNOKDIH4xuh3ZLz5+0ZystDPsRz1tE1To15e
V4KE8X38lv1yu85qHythGhBt4OoBt6scKfvOPNujn1Jo1tuTenJJx2vOoFbSsrnk
hE4A5slpR0tkHI3j1MjN8GxVue04Zg42GmcGCojzwNDLWORYDDGgitXf99Nj4d5s
safiS4aP8BgklG2/YfGBpOtGvZne7rU9+B7cpw0TJaCXE/lW2zXM+ociqg4x2wT/
i+YFLUXefwlkThWilfa8EJJ3fS/wTFezc34EXBsG0OMG9WUyAZz/oSJtPJVcMZwc
vgIp32vY5ThFdiWXRbQvQfEpJKaU/3giXHfX2d8shFNaXGdFjn0JUs2opzk4wdPr
Nw0aRDb5zgegv73LWUbSP2qzAliuLOw7xh8PWsaJWqp2r056jUZKyYCzEMS6pAMI
z2Lo8Adv6cCxFDF3kRYGnTyn9+PpknDXiGj23JSE73EJswoKGWR1B2nKLBdwj6bl
CdCIFgz2VoitJSjcHfQCxaNaYaQ6YdRTCy/JX2fIBjJnEWQV2U/FCXvX/Y0nQBED
iPqFtqXxjn8YhChvPwRdYRFeW9+shJDh0aovrYjjF3kFhDSjEp1Pbv+RT00Jjrn+
4OA2Gdc6jhHfyEetlwwllUIkqvco9Fj0ZbHjqiBThnKmpYvJ1V0D5TZMu8npe9dy
0EpyTjcry26D+w0zizSAP1XYB1Pp4EBUfI9Jq730DgDLTsArX/e9lThcjIvQ9J3m
2Jf3SkE0gAjTc3a9oAi9Ftb+rG2g+aaOp03Ul8S5W6ekXxw+888dMg4Enck8xZtt
GAl6bItAUlfZVrgx/4V8Fr2VeTm+/69K7m1ptIErars4krLjtvzz16qehiJRk7XN
R/eZ0PR0Ql0M0/3p8AOq91Th/xfjIMJScFrGs3dzRwdQ89K0SyB4jUTw9ZRPIV2j
WSL6HMP+JGleT0NncZ/6Ry27xiuEn70gQ+p7Tji3nN28wc6o45NnbRwbQXyZp+IT
XNeKGkS1EBs1HzY3ESZdiQ4H4YgmBIAH/pXj54Sv+VPoH/SrYnQ7WrRFJDh+WjcC
lUWQ06Pu/toYcWcA+X7kOJzAuLWnj9Sa0BfthVH1IhAlhSYyj848E999m8ZETFjX
BQ2YYVqcEDqRNBZFq2zo3xKkEBVPr3ScV+vIDVsNxzWKj2AoRf8JxFWt1e/zXkb+
FAp2EaYB+Snb/B9OLZDD5hZB+joswHt7F0DfgTX/cbfKmkFigmtbQGrqrQeVKYVa
ijoxj8yXbicVtc1BaPP9zO3KCvXgI9O4XqWtUfN6haQcyGbW52vWF7sSoVfkGKST
CsspMYmz/66xFeezagrVo4E/WDiHESLWHHHCwb3I9eLjjDACB5/l2T0Patt2Qyfu
TWM6xwmnytAamL5xmrIGwa9KeRoaeHG7M6YcQABCQi0ne18mp3ZTN38PON8s9No+
TN83rISUYcLpAq+glAA9iW4+dJSsgIuhVSmaBZohoXH8hQKH3nVFaXoVm0vnRRRy
Q3L92UB8dQdHNGj7BNnNvolC5BjXlar48Awu8cwgHBom8fJouBaWGhaQSJYwK+6O
YQsvfBvcjXU2O4CZg/gymNRxys4jCR9eZrvUguK8RHzlWVphzbaDTJo+WqV53ETN
7RASjYER50l5IWKhPyeTu/jBfFGru12hAWGpFd3Y759yG/TtVxATbXkztM8Uqeqv
UvswDlT4XAQaX7bYGN7rfwThw0gzsv0NF23QEFk+rwoumyYfMAJpP5r2+kZAR4zj
eCWkKM/4Zd2PiMEtZTSD2Vp3hrYGO9rUATm7p0q8yYZmjuGy+3pb7tKySkUGgwT6
GIKSdnhs+oDa5z1VGGee6+ScKFKVLSxyuwPrjOwvic3gkPanpXLMc3uhIH8InyLl
Z4zwa2wgO+W8N0hySrzA+egx9xOwmO/KZQqcVZgQ4TjHo3Mj4tJM1qrITQaY1i0Z
6pabyaw3zPZ3bN/6mEBtIi7lpcxo3O8lmf3bx4RSmBrinyZlNMUlvdSJckzQ8U9K
Ld0+ZPO7ZqD0ZAcBMyjgkSEBEhz+MeP36D5DL81YzpdJ8WNkgXuMe1/NaOCeNaqH
bx/xUiDfPdXyy2kNzpUMCN7OHRP2CYteDkDMiNNLAW2LdzrmOxHHkR7XPXvdWztI
AmoxZOJx3qec/Z89X5vYRirOkd8DHlwFZQkKipb4cYH7eK4g3oSaVlQiHvfLzehT
jsolbQKjSDHvaEilVLuC6DowEeuxQF2kmu/53IqPRui8AFQ2asojUmqz777eDyoJ
QV8HAWQb9s05GS4iHl7EHELKJeSjooddwDTxYorei+MkD6nOZTpK45b3ObalhoMr
+kMh4WXoxCJR+44mg8LE4Tna6P7AJA6CC86TdXHk4vrHEB5plaPjVrDBTpfoX3T3
ngqa9FN+vDUqxqnaVyMtTEp7cYhJhKBzCN3LkAxcwR+TnBtK9lMrtHT9xWPPxMJ0
ZmR+zORFmwNXZRi7ou/unTMZYO3J2hOVksSfSjNsJNvTT8sXRMxd8amwTu0oPc3/
yfDnjY7ZhhVKVIjvdcTr9FaNXBt6mMIqszOh1RW/+XOBJjlyZJPOIt7E54DUlvOv
y51C0REIzmgkuzSu4qCPIbtebEwetTgT8DEeQrkKF9t90Uy4SEKxdlY/mYP3xx1K
+xrv3+y693VLcZOyzUx2z2W4kuLTe+O7o8zh1HjxxszhXks8jUV6lOO82gyhpymH
/FFP1VJkfiPm+kXFFfrm6QVBw8A3OXUIWKo+C4qugfGPB3ybEzfAn4c6merK6Z5Z
m6H+gz+MwZDfxG30FN3qUTyO23yx04BDvHpp7l1WCwL+jNiqFuOYKKuqwfJv34Mj
ZtRK5BSwhOYLZTRnBufGpVA0XttEzw1h8MO6m/Lwf666GEPK1plkvHY5YU92azVc
nl0gl2ZKuw6QL/oDuGhhjsJHdzkMt6zkmB7yvW+29qHcHh4Z6j/QjSmdfa6j5pWn
Y/3jR5+7AH17DiagNW+tIN38THhL/+MyejiJJBczrZlvs1zMlmMYBmnQMncMO+Y8
fcua611SjlAcjUECNG0qejAGAJsdrqxvBYeNbnYSQr0Vmi3JBlNkBzLaqqmiQ8st
R5gghu0eHcKzLYtLs8DeZ++lBDWgbaVsjhMpAwcPTKUZp6SYhz0RraDLxye+QZ3O
LRM6fyHqu53ff/rMLcA8uJ1Vm2EcezT2fBwGWaKXwDmBcTCSTK77/9l32FBMJGRA
vhRl1b0yVMXlu2NEEPFeXkOda92/xalKQSpGckHdb52vfIPtMN0h1FpGXDNXMNsA
0akU9cKIurb/oYF5OIyX6zO62RWe00K//ECv8xANPLrm5K6TA6dyCjfi2p3ReXC1
k61nPUNnfnK0E9u0s1Ht1t6H2qCOgEnDj9yfBmR9uujQnHSRblKp+hqMilwRrcVy
PTexMgz1oCU+uwj/hmEM5FkHRjO5dO2dZNBFLmumMbkT6D8TBHUQ5YKIXDuodMqS
QbxorER9zDmsXuCPrHAzTC3kD/RkXOPEV1yeHGlerG2eUtIlpeVw9YJ4kXvt8AG5
gSl0znAi5TS+JOb3UGUEnton0g2hnKpQjGLNIg69/xnrnqBVuS6BSstwn1C8uh3q
HZQH1QDPNNxnz0Iu8D9uvoJ+DFWaOPUiky9uXWmfdzIYI1QYCHBpffDMtdRoAtEk
p/ZflKGBxqN70hRLou3b3oRD6USpc3e9KMTpnQV5TNhkQ7F6IMPbr07PgtKNGzbv
EUyKRdBEaF7LrtkGRIKM2oqlqIui4SUrTcA5wWvrngnhGr9N8GovmPR/dD1ewUpp
TQKqpxRLsnkZT55TF1rwhqNUcGEDo7NL8RqT/EpGjpMh51NdbN7VSMtJdrFhc0Vi
ll3OQ9BQYjeqGMLjZw0Lst9GFXK1jPaPVMiZ4t57D+74uSV0DyURv5EYRlXDQRIh
GiK98B0P5ebjUU0ziDLwLzqwF7e2bypkxO9dXBGc2UmkoJgYXqcmJwKKBRiCeW/t
PiQstf12uiJfYegZ0LdV29Bo3RcPtD3/gb8V2qbBBfrD/dcl8No+ePrK/Lnaf/qy
LJ2XN02CrZFfIxjIDB+jAF529zb7K+oCKyVOH+b3GneM85ctvkZlgxexJD0nWMeV
C0IADkvNhP+sT4rPSVuweIy/nqEQiMGCBjKmXCz0ZycGNpJLC7W4WSBT4vFbZ0p2
YzvcOwwNusB8RVL66asE1sia4bz7toAdSMoIrERUKsZpyt5Rg8sztIciyzfdm64M
/Y5QLws3nl9e+KCah8ctV4vPKdcrKvLe3WHU3F1RZ++SJ/JVTt1SJk0pzE7wnBTh
VwSRY3/OlP0ImS80eLOXWOMAgkWdQ/dDy+NF4p3bvAu8u88oc5P7tRwKR8wgmYkH
8QG+Hyd8QGAfID5QJwa12vKSBkKuyGvlZ33QbYIydUkP3+sJpLZb/ZreycDqb8dr
KCDdv7dDbgaUMx/cKPgPxWD2AfI30Dee48kNgFaTAFDrNritTxeS5lClwNH2cri+
jTuF5JP9aW2JKRikGW257ZZ168UmCswYHgouIB/XVkjod3UdXvQuYZUxjSQS/5YP
UZqvqFeeuhiY8prjOb5r1R1QjHzJ1sm4LaMwY07lWuAzZhxMs/trhKqyzP8E6Hfa
nIfwDGu50kqxcXVV1USP7gf+onCW1q5it5c514+kOLGNmrGBcgAWPBb6ZjfunQjY
XppRitPcBJIGzpFJfeU/r2gBppPlVqtqqopcXxyPBD2SkkHTz57jVFlFmiqtgezr
9YcA2DGpkVWdbFypeCqgsGaWbyns72U+oVcVHN/TL5qa5KzEexJoTPrR8PXIZvTp
igYeQKGadxOgVKPqLyrWnVC/jMoq2za74WN1k0CNCxMTfG0Frrg89fApzoOtJfVA
+CT1SKEpuq6Gj2fSZ8QvUam9IG4YpBiU/ABYMbZLmMeBH2IH1JpnM/avDZjt5adN
zKoe+KY6w78YWVrmV8Ymd+3dD5xoYzrb/qaK0A7P7DXPnhtLl6J/jN9d2TxRhCHE
LaRp7348Uhk0LQmYprUKzmv5R2a1J+DgT+ddR77m+MKIn2KNo/I79vWTELB2/pg2
VzdbW6LZDr9/uAuXyemQl99qrGOQYft1M9PeksTsapsJqS/DQwzHLb7S1E2wz2gh
z1FTLlRROGshTBKD1ByPNyXPmMoy7Yo/+vOXFKjJ21wcxIhfWQmoFR5II+onP7di
qvzpHqP0zw072vDslnac+x0e8LhifebBTHWzlb2Zue4oewqNjtBBI/9wreSyEZ41
a38ZlXBqbUbqDznypOvN35D9FgVLedp32m0G8Sb1sxOPtP7OBzmElkaPX8KWT0LM
wM6HUYUMXg/cA/nov4CqvsHEis4P6Pvf5e8mxhWnwd2pzcocztjKaTOThlGRWWjD
VVIHix8H6fZfc968qos3xwrI3H9AR3xSFOpW7UlwxcOc+1T4Zcsr7UN4VwH8fSvD
C9PtoPTzHBFkv09QdAqvx+/uvpRLW9+zWjsAgLWgV590C6k7aOXbm8fUmAdTVe4O
/KdKLuDXApHql1n7R3jKPpm8SRom2t4I1KuMkgPs+v2p3N2iGOlypCPYZi/q7pJ2
eoQtt7B9IRIeppR2AlyjFr6sS9oD4BkZnPJ812aWp84c6+8W8+KfS4BG/Z3gQlW+
whFvg0R8csnseauWh41gcCNn2689IVSbewcVuUADopn8mkov4230MW6FkCER7ZEt
eJ6a1lo/VoTZl7apWREkocZTcHAqN4IMiYh990M0OPfUfEDhaNaY5g+JK4iBo93x
bst8Ov8HcEGzvkakoujkotRz+VaJwcAv4YZcDvlZKzCp59VXA1UgVClTZq/xVdiZ
Wh1NEzvE5pqdvJ5lmZe/b69Ef4+vmJaaedn37Bv+SdyfGmLqJDm0wT2P2Hc8JQT8
25nxTj0u5kEBQXPyTAmbHFZMa25ZSxOznyQXJEUybmU4qIPHnvkVRUX+GSj5OS4e
uGhBMC3CeomyQlyfR0AWMO74oo4Iqe+W9I3qAbN38kANdzlINYMwL7ELsjN9BrFV
+dTLLJr7BzUACymkYSUl/Owmt018DUnXkUPUR9eQDYkyC+NUkGMsb0UPXWzB+DSM
VZy8UT9lfFMxLF5KRP7xF4cKvstFOnl6RW/In8oEQA54/glsdAsG7kylXuw7prJ7
NozuKUukEYZFYkuNI27lUv13XANLQBCpxP9rjZDP+o2hPuoqFE9i8t1eYtjQjEtD
o/rEDgwnN6xDNf+A1GelQ6bulypFWbpWdt5ytSW8zEGYBKG13y+Zh3hgX/c+qafJ
s1ZOkuv/Dr3VCv0X67yjKJyK0NMmX+/2bXVMjBRPT+dSKtwW0cUj+j65RRHtUBtJ
68rGSRnjwXtAa6PPmxl5uV+KKBwIuSG40245HBHfbuJOO7gEbdYkGfIxgoApG/K1
vaLOet0gpi+pIOYZGWc8XVjH/66+OtY57TZtYahHwqfj5+gxmZZezvfdqK9g6FxC
DTouCx/cbXTVPX/ty/JXbnjEwMb2uiXNJ7V0+IFDKog0gnnX3o2YpLk+A4l/59YI
UwiUy62KkozJDlV1R+6xlAlJClVQ3HyYpJcaS5lzxWhxFMDa04h+kBcQmOJNhE9B
tf0Bf5qSQit+syQsg0Ro8DgxZtazbfEgQ5C5INXp/nEZ5dILkmZsUKryNb3pctxP
dXvedkRTMOYwFD+XithPs1RtTubpXPg5aYxySNsVUqSId/kdYUpVSr100opFOSqM
kq2G4s1krpuigtX3FATdxliHy6hOkeee5e3MIqLwtthQzmoPRxwalii/jZ6wvfr4
gEfRRxAzE7+UajGljOsY8SXGYWWhtB16P9HCrSbPytBIcO5Kh7x6XCyuKMIEFYAE
TxYE72gxgl+zRlaK9ZsYYYYNq6O0jUCUuiaxzF052acqoPx/dCMQBf+6KJlTIH/+
nA4/5xcRiuBoWOmVEOa7gi8VpKoBtb5wsG2BkHz6c5h8OHrk50xGuVV5V7imyaU2
DwSEde/Jv3nB6uV7rVDxtZddQ85c8qQc5g13sVm9Uznec9+BL/yHm8JRR8ivaRiU
fu3f00uDIeUkwjVOATEceizNROuOjbPTLwYFvB1ha74Wyx5ABUcDSXRcGQvr5VRz
tFHFnlqFuIHB39BHzYUf29fAWNFym+U5k9xP+Yi7atOG7BASPJ16jYs2sJ2s4k6a
VHjTuFghWzuuN45qbqBBP+QE5z42bKsCxrA0DuegYwjGMtsnTClKXEzDEBA63PXk
G3DltEJxST33QrH/9IDnjUubbjksEj+5pmBBzHgVprRVaqtqoHs2EZRD3cuiuFto
BuWtQTBOEwtrkMVJFKxyNEmrtpYZmjgZuqLTRYbukjOjXis1J6kNgfauvyKCmU7W
RXtapc5Havzr1lkVOuoXZaAMZCWyxiydn6M1gfmHQfF0GJohPRkr7nF05kWlOY01
mdciHvYqQ36Zfrh5K+fYd3Gsagm4O1fKVsij6YfLcUVKWGEFo8RYOX9LwBADumC+
jjOqxv8Kl1gFfVnzv3CzHfwuyQYFpqaTLcIJMkQivc3ZO/zVsq6nWQ07yGCXMQED
EGqM2x1miSUGtBgkIhyNW1mKBcobSVs5BO5jOpEAzY9TSe4mlgdsJw7nPVDN4q2H
42aOEMMna78DohrsMtA6deLY7mIVXOIKU/owd3pu5qy8OO2rxHgyPJqzVl6hOhjS
xBc371SA+UBs41/25x4tlLS5yMvWBmLbpTeFve0ZTRqJylebbz7Gt4hGAJcfVPWC
ZcLiVraM9TSv10IlzQmHUZnUcvZOeEIFjENKz+bAIHWnB3WROFEWIQGsXFhvkjMX
N5J3HLXXO/r/orUK1q/1s4sWUu7Fw84pPhj9rBk/I+pnOM8V9u2qu/E3fldMGVmm
ziR3TWkV+9L17Vkd0w/MzSlHysO5cGkp2d962RjdXRQyodt+yl/EcO1TCJZUih/9
CRUqQn61Kd35BHao4ve2nmCyld9Rk+n9BCIE7KPtCgYu0Gcy75HEKwb9XyRx0lEF
STEhnY2E67fKqTExSDYhPM5S10J7MYqT+2ekeqsG9xtham96I8wp0sptG1S5NcvU
tyxR6TyIcmiehe2CgvCSbf4fqJcRYsYCwQIy2BQZXJMoH3nu/C6VVr+Adjd5X6Xe
oV9qvxfx4nmBc036Tir/gRlCp2HZqX38KwHrWfOP8EiZGiZYx0u/JoON9fG3IHe5
SW7OwadvJqH91xrsiB8wSgrr8AzKkz8LD92xTsXpHDPChq9s+z2O9vA9yR3j7RLN
N8fexQ3NFwEX8LL7/v0mBIMEq+Z5BGzzGAZaZ8d5fzqRTbCErSdRc+t+aPafLjeD
sha8PW2wZiPyHCEJdc7mQvYLrAMtjouMvpU7tGaorHk3kb9atqzTBcFCUjM2yCTC
JqIRvAn5N04Fx53KMao58CIwYwZ4xmDMTRl7QOBEf6hR/f/cZGdMJIYTL2nViIx9
zHjRe1FHh/DmLggbhJCL4NRucYmB2OHvBBY6hSlH/2k06L8hDSi3X59Bh/DZgK+Z
RmWNC2Jdrtyk9c91mT8zhoUAnmAiaYEExtyQkypgMjOf4/5kkocPuyjPllACG3xA
15QIN44qZdvgP/AoKOI62Srxa1XOGFDRRqh7K3pg2PMflsHJXaUZW5a5mmd7FGwh
lKeqpdxKCtt6Nusq739re2kXkuP9fAnwh08qdOc2R3DU/76UQWjOfEhDfmSgvpy4
1xINuLiDDMxFpckT51NurjqnlnzFLKdXF51Agu53cYgojt5X0zIFvZdVKbS21Sf3
HS54wBpO4IsdLZrPII8Cd2wxcbTJMAoADR93jj2naF43B/1UXu2MI5bz8GjSWb+u
2UnW0eeypR3S3P772LySxxX2rVYFNnZoigpO+tVSZPtCp5ZWUuo7kbwv1wXtqE4T
pVZZeaxVIIzpzliu6t9ORKF/ftKbRpwP8nbOizM6200wZdK3VALvfAfX1CzYs1FT
BLpZ5889SgHNsuwI0/53YSiY4+P0L9CTiIBYmdCfFqtb/yeY/oXr0frzDJIkwNb1
xcmuKbmovisVGF1K9fC94QkUjZgiSB3wSrciUtbitG6lyJbBghkrBjIznYONHSvF
AtO/VMoICwXYYNWO5A8eKuRNvuUHW6HMAmNOJgoekUEpTxTGzHQlgCmTOs2CF3Kf
ONbPDIL7elnw8c+pxZnaA5t8PAWFlocA9193hUwlwDT/t1N4CdOHIVl5sqZspSAt
uis/Iu/eLHO7megjp9glCy4p976HqBWwATq58mTMumItK0PVyG0UUlz2lKDY7Mcp
7jIh1CBIghgISsEytK4xDTa0M9p3m5sEr+ry9/FOrj2zoCoWKMzMegeigHjd1pZ0
5XH1W9q63NswYbjwaiVScusV8mCT3kGuv8MYdTaSr1OAHg5d7Whu05ZTLT1rrx12
z89B400VxuLhdCgDhLMv4ofZMOZpAw+qfeqVc1/VcDrS40wjcx2ZW1my6DrfcHm3
wb798cxewapTrLJnW/jUH6DtsFddoPIjrR2j/MTgCc0P6W4DxO7QyfIrwFw1XV6r
LQurqPejMu2rEpNL1OCVOFrR3vpO9x355SGYIQTIrPRGlui7FuYAFGcM+APV5fRe
y85Cy79EzYJzstGZcZEeF6gp2M5QPaOvApChERFfr+Uec8q94z3LqMJYdxnde5xy
vV9yrG1HfJvog0OrrztPkmhr1ts83mNb2ALS3rLSdWJFr1llynjS397CVqsORTUd
8SmV8Kh8WlYidfSw1e9jtqvBlSaYdFd5150iFA/nC08PiKHSf42mKnWz6b4JcCXD
lBlHklpJBX/fJSMxSHY/D3xv8ClPzbXs06x0WoYqKU75Daajjtn6KquAkKiLYt17
NgVZHANCykZM+p7yTB91r8WEkW0g6GtMdKKBkQALF+1MfICZhLnooWFn87zirU1H
I+Gbn28MH7J+gNw4Xt0SG11UqxaDE64ofHLI6IwEOaKFzTh5jOj1JQFTsrvWgQM5
6YMkhRALnwRXcSfn5WTcwO5Itzw8wIUC+37VUEgaFH+2ppbe8S4QnqyBbbsGqDm2
EMD0rGLN/Ef41/G4woqF6p/oGqxFYJco5610H1psF7xI0ys5ADKYe95n5eDtaEKB
RMKrx1CZUpJb+hrtVlU+HBLSqaENaVAyHWdvLvZRUM2uhEUIAgU/KP4vlfAbfJSm
zAKYkLlPOugxFRLR/8SeTCgUaCF/m51QcxG0FMmuYX/GMA7tgdB8Owdzia5HfeG/
DSFGO3QLjAx/3JlMc3n2ijWkAQ4B8cslELIiZkFcAFshA5iX71hrIJZLCSluCkcs
TfP5n2T0i1m1xRuG/EGJDa69wlmrUC9XBY4WHL7SsW0CaYwHGLmdYarBIoLjQJy/
pqZ77Dpg+kB4MUjaG2CgzCYFIFCM269WJbE3tUwXjMFJ400y0c1rn+uPG5dff3mL
ZBU+PdQt+NGZYJU/qYq/Wyn4aOHXzp71ch8bu+Cm8VDCRd/gY5k5BpHzduqlvNLI
WtZaNwQf4DXC1760fXp17/QNFPAj0BHwmoY1fgg5bnW62mTVWjA9Sa/KWXnxHHWZ
VI9sdHqKXmsNGEK0oynxyO7guwAjUUHQueuLrSHyJSPd8fNBlVyv5JjjzWuRMNpZ
sk9b0Cii/SzedOFods4ieZ5rlENJscjhuwOHqrhYMjvKobbuK8UvuO5MUD3JkhgJ
t5p0cA0uMaBrK9AZ9atUQt6H84ieVIkzTII3YWGoN4RwFkAl/CObAdPUxGZDtz+v
3zNUdIAStCSw6EE8R+4IOdocxC124S8nW2LjHc/Tu19fpUPg8tNl1MntKvvc2rge
COiA/81EsBoIdeldjxjGavWqd0DB59BIKiWdVvrTybR139Tsn9BMLsed5S7jyl4S
mA7qUrhaPQyPrDLF3EYu03uyzOH6dF+SDlwCvEDmQ6di0IxU2u8TFShD/chM/wgE
aT8JEIYGHeBJsF3m97rzwnDBYPLA91qO8DNqlHMh7eqC/Z5ei4HagHxsTJQyY9Og
xInhFzzFB6IJuRz9e+pCLBNc39SiyESVD4J6QnpmKpNRq3SWYXKVT3lW7Qbfw7SM
ZgbXDXgKTEDPiEjlO8+WQchyXfWHnCv6SImti6ot/tkxgjoaJRNO6mdzPkMsR9I+
IG8lAr0hVDDW+c/1NaI1xYtlTjP9cmLVsmpMo2srP/5kB8hWVRGnlS+XoVcDsUEv
jpjGIIX3EOVoAo5RLxINpBiqGsgdx6LW0IfauuvduYZbFRvdM5JOJNl5SkbXDRcs
dtT/LHFlniOaz/mE4nAhk0AfTakyiLOVcIxyI6MAYiw6Se6fdrmRWoZdxvOnibrm
RcvREutxciULtrj6KrPcplWMLIWrFM59SC8Yj6FFyOcZCHTS1XcTFkcgG4jMwPTj
hyFDt6HiRdaulQtePB17436TKG5JH2cBDH4FRS53zPiTWeiLQHzdZplYopSFsOFL
kgscv7FyEe5ECVbDwvRNzLlL9dUqUg+RYmWvRqsfjwD4otNXpMDqL+D7hHIGwrHL
MN6a6Rc/SwkEwvsgqixbEAo9+thGIgc8ljA24bimqgfkm15lQpxO+aIMtrCcloFy
tFXxB8APOA9fVYpxEfZ4nRgPhz2fnTZkTzNvECQDhhg3qmID6ZUKFS7FihsckeYD
IfoCXwBqsJc+aNricHgKr8TzFiOnU2qibGoALj5plk19kEOrd5gh/Vog5TZkDmCO
SFjzCaYCIVNB1Tf1iL27RVHYtANXNwxkVd2HkFuLpzTEj7Y7FahZLJjXKlvsBVYA
UAd/hj7IZjji82L3D+YXT5SsfZVEW20Ednht18JARfGiOGgYIN3pHOQ7y3ORRT7J
n3Jd6vBEvVLX471fU3VoheTgSv3YqDMFNn/Mo8OkLzrcgw6vC+s1/Tkf/HWe1e/Y
iBM8p1V46Ic+0YFY+1hz2WRqSYIoAu80af/x8Q9xEJxUp3AZCa1doKKSGdTSYtOc
pAziReTUgz3hqDSTyvYd65zUv7epp8Q0V2Uj/M2YkrHqPTZBHYDkbrWA1d524qir
ULX4WNE5o3+2/oDw5unpDv/lP1TIhTXWjJR0GJzgf/cUS4oo3MAxeFqYK+UywOlf
bLy4uxFaZGBiLw4bZ6QCniAZ6TH2yOHswWSx7gehP70bqUtvDpxFU8rgTjqv+DIA
x4iohph9DKsFZj/vzIitkpAmpd4qDr5WTF0evfkSumh/EMjUzkWrp6A9aUgVvvcj
gsClwrT7AmvjKEaUq8jAm3R+rH7ANj+4RSWK9PTZyq6NfbRVeYXuwhLx/MDAlTK/
QyAPNtCX7BhRo3JW49S71o6bjQJeG24pqqa4CziKuIj6EuVp4aDyLzEy9hYJZSUU
JV6vWzQ1h17XddjVTxGq8cJciTDeF0E+QLVEeSqdeBBjSDvOxhbevsrC46Mz78cP
WK6Lfy5sFxUHJSKbAPFQy3He7FoYmfN/PcB86syUU4rIQH72J1un2xOcnz6ayjfl
+ufz0ciz3NcNpvxobKlwbn4fbuz1xCUhfgjoV8QzGutFJO3DBsZm5LnqX2MKU7d2
q2PpH6DoV6pqkhb2pb5RWu0a4RHtHP4Oxfidsf2CHR3MapZYw+MnQ+i55P2O3s/Z
CCdyEtul/G6VFs6hSI/aNU0cTll7l5n0djp9UmzZZqxbo6V6wfgsOIvFnescpyqN
km3TYngUKIv3XMPyw00enrjXbA9ge6TeKpTBhHmCv/hqiYsEP5uRgQRqTIH7nWNz
DCZmv8zJzf+2DsAYEGtlf5qgVxDZdgpV06l/1+ozipOZZRlXga9+d/dzdAVDcWMC
lMeDxgrax8LlMqjQQ18gsaPGHvUYc8KxcF8gfKBMULI3Hr2AgZqnNZnWZDFp9oYn
C64a6OjCW7WVoodNxLd++Cc4ckAbjeuL2gPUchOGmRBw5j7N0HNFN72DAc22sPEW
ui/bq4Fwk57VxLDMEbZwUYm9FAbT9+AM7/hMssULaH3h8yH2pP3VEyh6TcWv8dei
F+72B077gg3ofdlIMOSZGFKqQ1WXvCQHO5p+6Ne18uysgB9JzcX83G+syS/GWveN
ZG48SMz8cZN49x6lL2NoQIjy6VHwJDFHdNsmyIzqdkyAHPMybci2sBrmumrb38Do
OOZVfsWWs35sqoCKFRQUc4kfoKu6nYIGYm5vPtppZYXnHPnidVcptXggWI9/crsS
lVlLZeUOD2O56axUVQ40nu+qV5nMsUxXEAsatDpNW5rBy8uE3uLZDj4soV+umlsb
7Y3zVhI/VpMkrladgHpPmgfXE26b7AAAZaDMoThGlS0T+6OqTKQ0qfRB4rBbZA6A
0bK1e/3abzmYkdxU0PCKUUUuR34npLlzmsChVy2Zbgbp9nA/y841HY0PIQkmYGxS
gMYRRnTZRs+Crc7RQVkPwbUCWUer3U6VRDgfIjphCkxswrZlhK2xRPvN1u9s3bye
11UFc/5Pn1Z7FDae/El2yKl3gau/PCgkjlkI5fWuyuoU0hwTHGbCecwG4JOyrqzG
EyAiFr7LoT+o5z3p+93yJxxvQhUr/3Aylk+PIV/ikEL0gmUuK7TbL79bPzCz2pc0
A1TCa8++/8SUmkHijxjTJ9HepEyjwxlT6JCLKvX9cr9wp1pMOKtKTqPye0ir0Vof
YrewTXVHf7NLB+fTv+uObjKQFc21dRcOsishFug/gv2Lg8VyShYrMl4ufWzSJb5n
fckMg1yeuUE+L+7bSZBF+48/u/aKKCxvf9baQks+Lnh8Pcw48VJ2mYkUHxSlK6QW
6QoM3KeZm/EVckCOwlx9IarR8Qz8LZsoNos128WMNxthRR+lRUvkrwktiXrDu03W
toP0y60TfLn/8FvALUMzyDgnSiHzEAImGMuaVXxhE7sqCm1gbPgGgzTPAwRKWcol
wPGKFNNKQaV68+IGQgqN9ckcFRa8Jk9Vqs/7UkWZ+2gHlyObdHSO3QEb4qCFpT6E
1rLMzcROkCKyClErLa9lrqIklusssjcHjeNiXBoX2Ceuu3nGdHK3k0ti09UIXMYd
E06mqdzIwSFLnWlJJqemD90zJBBza9/xdEzmXNoRAjodTYUTjLNr9L7ULXiIX/qE
KGu+IobcM7s18D327QEBFrnBqGz93kOFVwzrxLJeGD+UQMqo+CdFN++Sj6W2JZs1
aEXscyG+8aKih1Q6uYWtSfYQfJNNcAi8JYozvaEsTlJcq+4CE+wM0iq4wIaQIzMW
mgea/5BMg2P4FDkVkZ56dYOS5eMTGQW8yv6WBCEbC1YxEnbNQRU4iLGNkxwmKtrh
MDsjjZLQkmsovdohaLR4VdFx5MqW27CvK3NxdcrZe/fjHpP/qY0IrxcGHTIiHX/Q
kPfyu0aCIHiuJHdBmJczJg0u0pMyRLx8iAsWIQS/czpW0ou9TfS/7XM+BqN+uvZ2
IsuMO6R5Vl/3kJ4Jz9u3ZcDkPudE9G0p1KBucdIdIhh8zryWsoTJWAqLrqTyJi+O
iMHuHJCkGQ0FbYbvwGFKU2Zuyvwl1Jn2ac20jxoPqHaEhbOmyUD0IF+38CSuTD7z
DsqkzASTf+IYwSF5rhT78j+4f1RpMsNPe1MXiC47l2/kNwptfZxOQATL21rYxMLN
ACrIYhJqfbYfGEN/R/ZYIhMGIgVjSPJR58bSxCaHHtw0f5850gtRyt6uMZ4z8Hir
rLXNHoSG1BIyFgu3V/qCw81PcpBJk0fpaCrmH5CR2dCeWjdngmxX4AdZiewd5l2Y
rd6k7n9mwZvhfESFRC9wduJXEq8s4JYgGagRyk9clbaGS8clOY+fr8fqDPnQ5Oaw
YYPmlLGrOb+KAreYj/QvZbC3oossVm/mLCLxSN5M5041DHnTxh6vhb4P16tUNCpB
r6QLfrjAV+IC/FJl0okI1gw7qrTLOhe+83H8D2KTl6xvCx2hKe55EIZpjjavmLqo
E1wLv+hAh4NvaTis+aC+SmSO8XRmG3rNmr6kJMsNKruLN+liwde+/jq3MeS9ldQ9
D+ZIFAEdkuDy+SUTVfiCOPMTGJcT1uIjodw21wIIS7T5XeyW7Ld2suW3TevqIQkg
NvTbM1ptJx1EpBF182wEkQ3X82pw6hLsnRtwOOjSyOlE8rbvDiP0ypJS8v335db4
EACo0fx7eqoWnx/T7v+Rai2zCwMOGsFgLuNL/nj2CCEq4x8Ycva83ZSIgCFyIEOD
vXRJzYJCRWBkRVtdQml7Lywb0Tp5D0SL20qWG6UMuYLAmpg5P/mjXUqaqxMvPPWr
lQ8kGptVGlxgWXU97Q71PHmG4X76a5vdmTgPcLjUWtDOSNnnus54DOmEcd0sOrv9
uVeuRkonYo49pmdzNo+/Gtx7dzSh6G60HG46AeL+cjzhoZ56wnR/40+e0XJQZ/jH
5afMDhAF8SomnyMiiBryG3DwBpbiL6tdGWz0FvQobU4mllxnQchyhPXw9+OGi0FI
Ngb9+OJy9+YU4rDlq0rdjzBMab6DIQP80lbtRFT2IKZuTIlE1ywEG4e/gT/nZ/3C
WhThltL8wsgfteqGM7kh67hUTYfsue37QPZA5YqZQFep4HepEOS1lANySZXkoQZr
DA74pVRjbGvx7MzyuWFVUvBjAwkmKKEP9EFM5Yz7TfrssN2D0bluL2MCmnchHuRw
MUcTBPeQo74S5wuRCan7vjIvvDuoEqPT3k/pM/Yo0lny2qBt985A4sKOYMtjq3IH
aL44c1NhdYG2sjVtpU+r11J33vHQXa4V19hlX901xcBQCUrhv3ULZY7XY8nYXHOu
EZ1ny0nslKGN6CLkiPtTQP4devHyvR0rYaIaEidHkm2Q9JN0sOuFkJJw326g5hyz
fS6MllXRbmKfEQ2lU/BAWw5HQrkXTXjsoHF/5l+dU+cOKwHUbCQEbm0ta/0gGejL
0OYwaPAfdxZRu37KFY8ZFZZQsMmKMQgUYJNoqDSPHNL0cg4tpZLFc5gM0h1+AL4P
GdzpIRajCR6vTh/LNXmDhZvbsNoYUk0TMky842MSBbCmkD7Y9pUOLSvh9jQwFKWi
fp3QMc4kdX4EaVU7L3BheX3yNItNtIUp4YVWoefOTdDbmwwRG8rlSeZSRKOTugNS
GzvaVp77ExkI+3z6UgcndyZpLJaRQRgx8iMSP/mzbMX2Tm5Ix9cKq+0CmsHxyP5b
XhEIzO6KwsgC5cDME8mp16LMaUpxn0a8BRG++O1hiqOiRpRr+y0sY6ecu7c6gItj
GePUY5L+sNDZ53yBnHHsBrIjW5NFwPH/tRHUpscgbRobt8CV+/kcJtqeJ10vypG9
hZJgpcp+0cKunrK+HOTzXgvrNGwxi4JvAneCf0zRiMAXUvGKN6hxUVRyaSNn385C
tR3Ier0tk+QAvpe/CPQLeg9GcC+f3wva9BMwEeSyM+T7F/6gbz4wgFgo7zA7Ya26
6y+0moenl+zDneM677iy3gow5jCPCWjxwUzLDisgb6G8O+GmSLBbsplfmlyzn8lZ
8BVlCjNoMLLsbnzAqkn98570gczUh/k9ZwgRI1PHPqpfdXj7SDJ91JIPd2L+GmQj
jytPYaI9OlSEm9f79fTOPk9W/7SD8XtFlbFaO+Ni6XmIZXDouRoEYwDbIgwtdL9w
vKi7xpje4SFF53x/dPb2KiCY4aGwGtb2xd3YKbVS+5hLRWU5ausI53YwMs+RozSo
jD0L3xvqqg9W80AUUuLLR5jVUBEZyBc7ZAh197DlRdmB5xcFAV0/wjdsRCXT3Ifb
ZJPDlbLM1mifHyDlnG2Jc3/dSMXW8NWhTd+apurHlFf7f5oQ7FiTGIfaRUwpOuYR
kqkJrmpaUI5XNNu+FaSwxc6xfDQxu15ERJOv8dSOAP4eSmSKkQCNpjBB9of3n1qq
qrQ8R9u81pUHCBEfSpNmrpD8AXZ2o5+iLjA+wMyba2kGiaVXReov1v7dyzked3vO
WnlQ5E5ZNrLX7w9en3IgZ62qG+SsblTvdeQy+f+izPBXbNSt2QJhps4+D5kv4VuG
6kpFijOYxGmtpdb3bYkGukM/VBozHgnTrfNH1KRb5JVZJs+X2bYH5Bwz5JHvPy8/
iOZFJuH1cremiq5lYEv4HrnqpDAk6NFFY+j1O/3puVYGMQ1Y44M8Rm9xSpgMScBv
8WQpKTCa0IgiXquqHjPWeAaJrgiYBUNzAaUOf+5lBmXqJ5Tn/2oR8u6/f61xhU+P
R0fQ7QoDg1tIMynhDJOnNZHfwqNbUmvyTyAu4OBxB0pHiBBqvLowOpMOgk/K54T/
4LYGkGTyT7844J2B0tZMyc3n7Xrp8Um+9DnlJG/b3g4VXoB09ZEwm3jfxL1MKzCE
V0PF+ILTgA6DdLXbyrw0ANTW1FDh8dI2CUDsrUypJ6hfyuObfueI/ETRfi7ijde2
3bEVGRO6gCKewxfAuUkrTxtn5ni6LFlXGHhST55hu331MaseoyQgaZuxH4yN2+fu
Am8IJK4ZEvBHBTPoEX5I405WBK5EidlcNJD6Z8WgCYDs/tlRQHX9fmYTkisgPEhI
N2AZOLh3hSGL6ws2XUABschzhcowMFiW5/Chyd5LJA45yZ6d61AHczDEos3fu6I+
99ugUVwcCVd22O8rAX2kuDQDhHgAft53nKj3SkLYC+RpQN9S1zWOJ8IL1SaEK5cN
6ooRW81EQe+15avNYdDJbIYl24uENe+KVROfmaIgArxEp4zXX+7ScrrleRG9zCYD
so19OWOQ4yG7oY7/AJt9CD6d5txhOYjBIG7IOm63N9KxX57iKdGwNgpRqGutTG5i
cYcmMY5x2y77ofSHrn3ZnSgU8EIC76yDnj9iYgoz0ceVbmWF+XgMRT42VczjpWQ2
MzQhimShvMcDYPy8ia7vLGL6MJJE5thVgxgyvI+3qnJOuJktB8PNVoT1zL2gMZJk
Rk3iUIkQa6u1KAVpatJEXoIs3J2cgQwsbf82ceuIKvvHtyFpHHgCvdEzGQhNBBeg
KVLLftjGWYTdv2lF1mtF+jQ0en/K/AImA0OZH9SmjKNpSAryWMNdtlGm7DUG3hde
17y5emMddMRCqDYRYf03wUiJ0oKuA8N8h7DE7PYou72W8aI8vQ8F6bjsgv0zQgec
cmW543TLAlXI9efPIfg8dKDlCBUs/tYKhltKKssQakEqUAlXiBj4Vmg+6opXa+Ou
PUovA9G3fADj5ATzVJXaiUWZs4lmQGxOBA80MWpvsyTuueLsvzjrJj/7ngWXw7vI
rHE2o1pacoTqIRESZFLrvENseWRbd+YrFKr33bhJge4cmmX38Hbp9r+RnWNdYk5w
VYok2FkL6gV3fvT2k7PX695PfbpY1TwlZrfncI5cv+MnyYDpkTqvoLMJk/H3yw1F
WR9jCjzWal7teBEV3RN7STKXTgXRAfFapQfSKwV6ZkUWhE5kkjxUbZD4WKl2F5OT
xDJfhoHPHviLkoi5mGCkSK43wnr5fbiuwTua5BZCcd/PGTixiqOtjaOc1fyS6J9S
6/Kfaro1nfxMN2bsUfBJfQ8cwXBlKEdeodDaiYXC366GojoICdRbKJT+RP2mjoNj
34qsg438QN4wjZuXSajo7ucnIycR7g5r6t9pgHpv4eQPV3b4ZYzOatIaBFcbiBOd
0CKm/Nn+17vSOmn8jxZlLaCv+oAFDieB6VFvJZBmkPKfZONczkK+7SbPCxmCnnBU
wG9zUpQaYZstc542w55J8jVBvPQOy+OwWGRRHns4NBye9hBF72KG5+Y3UyXhQi/N
Fjm/7cbUk/aKBn3EZE79cA1gc117Ge+WNMX76BgXgy40hHUwa10NZthif4HRmniB
YEascAL6tKIchZA3tYLoNdPTk7dy72c6N/hmbMAnfk2Sl8uKt9Vj7jzRfWvOzNnq
PbHb/eCdZ/4OhJFro0RxUB7At4RH5JBVsrhsZsSjjiPEnR080d/EZ6YUhIxTk5la
fHnWOQd4KiNwmyhBZhzYVzgEKJllJqdnV8i4WcP3hpsadAu8wRVMWl0KlSuTTj2w
iPgmcRigK/3FzO0xBryBMC9jXaiffaS1hLgPw8YN4AxKo2jSwA5IApb090KnuRAf
rdmYeSxGxDjNPDDVyx6aKsPuktsGWjqFgfk/wQI8v2K1iIr0Epq7X0JwvIh0r+IZ
TLGx8FTR9FDpaC8YzaAmLW6zNx4neXkceCvoVQczImmHPI+7SWKgRFbgtgKAs1lj
g/jz+OOZshKiLb9YKJ457+/+AyEguULdSiErC1YKxqGlXK2vpMxtfK6y/59nQkL0
qLAnxZ2vzqZ2OwUvUxWtc1P1JjkqOBZp7vlWlEidReqy/LbuOHyHMGx3OasCGJN4
fUJ/Ixcg7sn7pkwSIkyYlDg6ARz5RNWHelKxEZnhLKeNRVjcXu+rVAPqE/UHle7n
YjiUCeu9+xrfrscuQz7nyfXCmWS2/KAdwW2TXoNr4zHtn1ZVfUbW3fikhkHq58HS
lf3l2Ouvskmaz+UGRKIxrlq5qVReorop+pbzdW5zjAKLBFJHQV68vG0gAV7DppF0
6n7lhaacNlDEya5uBz9Os96ruuOs39A5Bu+TX7Q1xK9BgWVXOcK5liwsKCavBeGx
wip8StOS7pcRIg8+nLCng39fQAQYs5qqAzZuPkIHII0UMV9fZZypujgu5IBu0q9+
aV3+JSPchRZVHrctfbjLH+RLvHxhPUWsDWspmBDLddCzhAMS1XI+Fa9PYOSJjbQu
gSwRMOCwV2PSLwjVQQ8VUVrNVN5QTYdTQVdTYI02b8xUqKDCoBUaQbfg7YvXS4v9
T3oowXwN8oPOQUcwL9B+t7U2DwY5N2+oAyxKWmUDreAD15P53LnCY9Cs+lQBr/M8
0v6cEPxLvl2YvXVbvmPfbYiyb6MsQwpZ4c5QV0MgIrkVS87hppJ93+hP6Q45JcEn
s5TGvVZ2U/a5BPEoMc2T5hBW6qRYkZMOPMtc6wAiQlUCJ9LqZBLKeCQs1I/Ti0p9
qDzQat0vqcJIHioKEmTSpPDrzO/hfeXSwdviuwVZ8G9qH0xykQkn3EDg9a+akxrW
bLpA4N9q644tQiv1rnrx/A5j8Nz8VWinQKS/O3JCAfxx/k/9avsZRGvPUzqNRg+A
q5hZ3bbFvF94i1Y7eXbN9w1HU37ZocFJe0dn5QlpVd2lr1w9MVgmUOttGqvFMJjh
JtsIMKH47euWwdwXPmuoLXSYvTJgojHrecry3C+xbIb4jmYtRvGOheLeO02N6f56
OIfTKcXvfkZcYawSrU5nG1onM+eQqohF1kJz/Pm0dqcEHEBqcSjlXY8XQCPKY4DW
2i3ZpotIOgiBmqJ+m9wJ2J1CFPIeLRxCNPJRXw4YdnwfCfILYUN8vRPAwwDo0C2E
Y42MsRMuBbHQ1BntnLB12/SNrHCFFPeWeFFWThRfMCPyqETLhcJMKsteiwjFcy2N
yJ9iArJ8Xwtw6rlC2GfhcgWMmbO8xxBshnFu3e0sui2t7GbzIFEmd4XVBV3/7Di0
QHQYrLBM64lYn4to+aYriQXB/Pz7vj6Fh2SQ8oRVplX4ZnbcmfeX1Cx7qB4Q1XXQ
8z7vx56Q4elOTy6GSltnaqW0Wqpz2TbBOJHlBDtrjDbP41ftvpgQ1uTEfD8g2i3N
0C5/UDUUG8S2L0teBQ/9KefB/1FUVodH582tV80UZNVE0hTuWN49KhLNrN/OLtGb
MvndISXY7UABravLHFyBepthaV1I/HGpeRPa+7j0X6DSzi7SQP3BmNEAEwOkjE5L
+S2zYmKpIygHXQQ0igOna34M2zKfnwAqNp0cwUPSDqOQiBaatlNicQTRSrbx1ffq
VkqJVj1v+YN4f0Ha6RKA1kzIkrrPjRainfBrH5xF/tmbH6E6ew2ByP0jFruuLVID
9PnEnehiGeiTASmdF/5Yugik9t454rZySQMP30yLFvsGxcNJ3RiSgMA2tl6r6xlv
fveyemxnf+FupbIe/v+Vo6/45ja+vXlDzhIW7Waq7yL4WJ/A3KHhiuuADXIM+Lch
+kt0fweIvdjMkUYkQPraY1LhheAwY9PXYoSMZgd+w0gsJFIe5qeJHjnvf4tZbQka
nCAGk2BuqfRwGa0SoQIo3QM78YxpCS7BV4Gjx/UhBmkVYJQy5Wi8RYyWp9UmIpEO
NhTGjhwws+t+Ncbx692L2NteFbMh2rc3lTHi8I89QenO5AhdfF2Ff4nH5A0E8Gzd
rng1xUtDQ3JzM7CS5GGG5xZ8ttbo/OfhzqhqmsBt+Vp63mmmFQCMnIl+787y0Yn/
F40KTTQFryJsr1eljn8Ju2S6l4vHnwWtgdjIOlK5rOeZSmStej/MxXUxUFzp2SMv
gTEG/EJZb1lgxxhoUWRnPH8DWBAC+IujZJlLM/o++1w2lF1+ztExQMgbjX5BZsFe
1b6D865iKb6MCG2co/ymuNMhwKai08FS05a3piKh3ZBD9yRwwbpNyO9sQU2NggyB
t/Lm6oWp6CXs8fcwDtKKyjscL//nOvphrfLrx5qgXJtStFdjz8RuPEiOG9LNkygB
gWxtiHoAT7JaVmONIZOtl2Y9u2v0FCod7wYJu4YIfjQEjOrzcfLOiTgjZzS2+nFP
ERIhWBJtR4B1/Vc4u909u1rTE1v0XadBKnjmbgw+BKZy45JCmKqVo6ZU2pTttxAL
i7sSAEcev0FbjU1UsSMaKlON7nTYV5IQ0wBsxodOthaJ2z7bM0oUDryOzJQL/B9q
f+UAK8mz1o2HVlMLtjuHMnBx/NHrXTFJFTCov2qrgsxCcSvnXLmM4Nw0UFBv+RxB
ARsNGUVqS37nB1JGehlRdCHDQ3zBFZAfg9oDDfRSsROPlltW8N7715y3bj+7pSAD
BLiAUVMYBjA43jl0oltfEqQHpb0BzcdXr9n2ByIFhKXEDMOrsv5F0mZug0uMcQjf
l6ETvKjxxmX8vgiuI18GS5IIFyDpZ+rpYdnhzp0ZSVNT3aF2D2V6AtDU4rcwLm02
PB2qI1xwNwqFyFDkB8akPIrFiRMuxKXiQ6Tdoh37bbeZhUMygyVpznlGgfU9xqvR
2xfoIHSxpQwcjaoKyT+co3TuZxRc+EkIaQw6MGWVhEDRLk7lRnjMSxfssXzEJk8k
WY1XFfeC3c+4cvMD/aaJtrnd3TahJ61BP1JHvsod4Wb6t6U5ZPVQk4Dt3+8aXDEI
szLUP0RFUHh8ItfCgC2xcBwbte5aSBcubVqMCIE85IUui+wwELPpwqUVCXvhf4Zr
FyXpXdsoPgdVV6/WD/VIeULB6/3+1nqEtY5ziQtCgerR5hil+txvtS50SUwenTLa
GW/OMAG6eDtVWnlOqSURoAU2Y8Z7N7eiho7YDMTnNHww9mbElz09ZfR7iyJdi4d+
NylwaEXUSuMxRKM27OvvTV9gPSuTwV35IwpNvpJ4xR3+GNlnvCVwuFLdTLG68yzo
W4MEaOkrmGCinJZhHbGSB8wf+BR9HY1S7XSX8otoozSRd1WKN3NUhnBDH0DIj6i2
D0WTXSPmT+5ppMb9gx8uV/tbx/KUhegwhsfbQB/BcIMG22i+pq4E5Y2Vr9D7QLik
VG3N/+OMRIMG2Iby0KaP+1/u0xYIvfw/0MgWxO12ggXA8UrKRhO9b/+5HFzVt5em
MYQaUkAEtA5oS8nFc+Bt4Ny7uxtpBNPthdLWzs0IB0/Ey/dIkl9iLRH8wSGJEMlH
R1zBNwnYa4UYvYzaHA3AvjuH81S7AkfDVrA3s6EBd2sjy8+xEMIW2sNMpYEehozM
KI6sLzUNapfa+7ygXNzMvUZO2pD58we4tdLlzUol00zs7JQ3f2TmcNdJdxPkZi3G
FzY+LPkxh1Rpi2cKAqtMwef2BXi7zhThuIkBd95bee3h9AEhXjk8pF12z+d1WnJX
PHSWzdwqcigMyE/O83NTGw7UP3q5ciStaccv9Hx+Ht5V+t0BS6BYnO7y1e52pqVE
l2TUGGS7XMRDwlnrOAd8NzvHjkERipFqoC2oAKD3fOZC22EBQSmd3w/j4ZgvgGo3
KL8HuYGuJDrTcpAorAsax7iKAgJorpNIP6XRTb/v926Bnmk0sZJLMiD7Htwq93y1
D18jYyxuoi9mG/clv9bk+vVOYlddZ+IXAo1Jn8R684oFB0wjy4U8sCRHrYhJ0JgG
CzKDfcNaOm5F5ccFpwUsrHcZyWURmLZUy7Rxs46hcnXHgVPevLY9sidZMmNCOCqO
Rg6NzgSbzGBkkiCY5inE+uBxBGptHkkz2SrQ42d7JHKn29gq3qro+QivO4Llu8KL
HM7tS6TgJxP0i/Og53xauS6E3asXBqfaxyyzaka4a8j5RNPp/++ixvQXr0Z5WWj7
hA0CIHMc8nqJ6SwY/WVvIpmjflWwq/YRlIAk8hN//dZbfllB4LeUArPYXSJVNeKO
U4hKl6/PFVyH3RV0WeblvdCkfxo134cFpyc/Cq5V01uGtpRcYdbv2KT+qYoagp0k
m0YLgPM8G6wzGcaAkIk7HONkMdCrlTUZVb43jvdqIsom5/eNus7Om3W/HrBs2yuR
prv+FrhWVUwOomvEknhDMbInk9unO3AeAixc1z03w0OF26FJxzB2sWW6PNsKokyK
WApqWsJn5JMkHHT/vLmsFjtn802UfoY3C76D/ONzqX3iapDhE/mcu+MafPPyXOE1
zU0MBVlpiNqnVN/IBCluXDnSiJsKHVI0EB7vRalyEdO58m8JYWOZvmjA0wd/AUam
ZcPFo1YFACPqD4xneZUJAs89+XlVe5jKSzTtyT5y3cSqThueTmwi3d2lWzZpdj2+
9hLZRDvF1t1ZVa3HeW9Wf3oFAHHWBhM+o2AS62pJW7bYVVkVKV04IjHWlqSkW/JB
ARIpWgf8kwrtNTohXpe7bX7n789bkmjz8clsTD+GkAPiNMpo3d0IzydBrdUd4xB9
+GtRHOCuXPsOIXlQ3cL4lawv2V41m/TPtRJhDq+icGMtTvLW2v8ZWNLLdTOyIwYZ
Xskzic2/izALsQmkNtmZFTVVD3xVWnYfiFW/XeH1mSuSoqVNxDot074xvweFxsgr
jYMoJ8ziNpoTL4JOxCBJGTOfyk9S2pWLVtSRKi7oTMrPbVmGvG4oYKzVc838/0+D
1WzcPm/usToCh5r6h/CR4xviikOT6eysJQNJ7begPv97J6kVMHhDfNKtXdsNTeq4
yDbE1qAajU9IJq6VuI5lwCIkreJ8Vwuza+v4+LBg8Ycqg4KcmuD093thM5PNP2ae
eXE61paNPVeMjHHvGFJREmqpZjBhHNF/C4MfdSOsz9Pgb6WvtRGjQv+Xn+ZnHJyB
E3dZn0DCpZTqcLr/XZCWKmQqd8+1NowbHKQzTfh8L46+hYp5KiEOra+UHsZCKFsC
HS999vEuvMeKrWyN2oRoLTet/+GnYQIkytpLuJZ6w7WHeUnIsCCbga4Ya2/Hfj/Y
ZfOHj9FgIkxcqiSY2WQLWQR+wwFTrrlWT5BSE5Xz7vRLxmbIc40GgCJQiVGzjf8g
voTvJzFqUpTzNEGANEQksQheEEq3aNgUHXp5L1TYSrqahjArX0S0HWb22prlbeSA
MiNc5RiLSqGoM/uVs6MLYw/0EXlvKfQka3G0Y0M+txLLLA5/sHxRDMijZ3oOJ0sT
xU8BgWMaTqVl/KWkedm5y/CbFB3R1mNr4wK1rWJV4ZCB1KX8ycotaBwbocjtRR3G
PpACpIHqMsdA3V1iSEIiCVqL0wM1gg6VVmy04FEfBkqtOdvgR4WSuGSeauoUNDCC
l5SqVj2EsnWReV+PPnn67FX7IjWDHUeA2wezxn+4YNS8I+s/5btwFacqNCuJOZGo
Phwt+Pic3n+CQIBqh4toQ7ZpWtXD0IH8Dm5W8BfkzBry9Rrpdd8dFHWjCyuZ4mzO
pHKxx8qSP4eycSaYLE6GketSS5WVlatmE7lI2rDFEam2YgNdoykz/lfaC8aRX+Ss
4Z3KnMyzXHou68Ip7moYp0L+tmzJaUz9XD8xQlasowh9IK7JaZtujV8eLsL4dzoo
OCSPPRAe7PfBqT2mzI1snBlwszbJpIlHBnkpd5gEZE15aoI8rYdXtZrLWV9RkrCb
dbxmvBon0r1mgZ8ncf5nxAxbKW48u6UHU5sII/ZvFxBbCOpl+eYIz1djf4EpLwCt
mmYzFZTpIxOzlGkl+FQ6odvqrHF0K5DE/qBLaCUnJrq8O2ojSMovwNoI5IDNyZsj
0uxqlGwozf5dUcdcfLq6/T9pF23w56c0EUOHMlYg29v/2Q90luvnNHqxfLiDxYfg
9LkYxpnkXjwtV6SNRAt792Mr6FyGZRqAOaa41VxIRwgejODFrYnrduMvxHEcempK
TB2E0tGVvcJvCfvJCNVyRCXSILWbgDAr7auHmycg6RzqhMt4CVoYWIYlDxtRFe7i
hI08OQ2xpXeHsOn64NFeJnWvdUbZJ7cX4mkiObqyMUajOQE8/d3ijnM4KvVluWlZ
dtDrqyajXpITboo5VxG+9kV7hJhqMFfo4slCarOTORkqh418Pk7DWOOSKHF3A9xR
e7G/c7oYmP8Yuw9LT8YIjp8+3NcOBKa2i+t0Qt1WD3I2dj+BJIn+8CAUHkJneE+f
H6kN8BtaaXVST88557dzbHWA/eZTmq5ELXDq3PXjBIJ2Y86hmzt/7Q6lBvh52NoK
bCz/vAe3K54VBHDhYpLvkqioLpTzCLbc4t8THasH9mpmcA79SPO0JHdD9mVfb1Cg
LNZgutE24h/HcRNNoStw1mgM23xiuDsPeSFLzMX3uqp4nVBnFdptfzP/5mXFAmKs
u5XVnaJFUu5rtxywyivugsjSd/6MjKYPGBGmdKcG1jDihmOmMuyJkMijnYztyr5K
w2eRliojBDKqiS5Wih8pHe6p//2SQgAtMWrYsobkrX+ayAgj2LJJxGb3d1ycsdrs
fl0XDs3n2RnFIkAW13ZwxW/mBUj77NlY4Az/vaNQK5FqsbXbH3JdN0MunxUPOLUy
lCxjhIpD723Ra2bQCMcBh68FRjSZxWumF5n9jnLlnFCiZed3t9b5osm1d4IoLd+v
MRcuthap9zwr8tCYXgIYmjpb/sPANK5bKWZzoTrSNsqWIBuZYR26TQKaCn5LRiNU
2wPyegGB4Rmdi0hWND1a7TV/c3c1CBdAzzwOs3r2lMNm8JCrmB0YTmQeFl8SclVK
zN2XzB9cOU+QHvp9+7BnA8aXAZp8KXS9RG+R4gBEoViGOAKiObD5wYetBfFA4J1P
qMu+UHpBwpy2O3OvTmC57SHfd1jUFA/sdA1+TysDJMVVQW6VvQeZvX3EaYkQRKa3
aJ7vgAw9lxDbsv6jsSl9vC1WuVbIvm6qJAmr6QaTIMhweaBUg4Wx8XIdH3TL7YHd
cCgFd67NZ6Rz2wHrHK46B4PXDe5MUBTCuBasdATmxZ2XUznWhEjx4aQ77k2/5Hka
TgLKwARdQnoTGrCLo9oSrBmgQUazdi4K5Q/7M2ewDfz9gta+oGHueLtQ7Vd0qffb
NbVEG0aPp/Ib/qUGYnGTSyE6BjI74q9cSDDHmt0+y39Bj58VCr1srCoDaAClN2op
eGtZZDC/8fIxq0Hlp2kI9dEuGj6y+rBZn0zbkUJGhnb6bkNIu7fLdhLsIMkhywTs
8DunwB+y0TAmCfoPa+HVUiLkt5FC+YUFrOEX2NCbKfBJUdb7ukt83zXRvoFgECJF
nKudbluUAY6wA5A66s+KB4ZuMHyWO1Cd67TJNrsccTVJCA0JWu4Vu1ZuhlZRvS6n
HCO2qTJJUme/9uUdmkYZKiq4vJo+xMlhjwAGQR85b56YnY0BzR+n6dY/HHGhnhEd
13aA9QTLjcokws+eEot+m2DKLdzPAV88virg4p4RR5X6VtfuzldUd12E6pOoLFJV
llwuHstvnrxqDeUYshCDxDV9Kg2+TOg3vQoOHfEcGOF8QdE5xWMCA28ZzFIjG4pu
dm4g0sX+C8nbv+uzbA3aGib5zCIOeHn9hNgj3RNUZmNzcOMMem9orKnD5N10xdAH
SOLG2jalLG2iXy9MUz4CF9fvDhWAR+lTn3mbq7MKc37oxkaauR5ZGzbPz4vCuUfs
9vyA1QPPgcp9ETMUwTS0jclyrGfF4qyG7hmcM5rNNgOedrZR53shhjzkk8tClSwI
3AZphza9X2wR90+WJt6mnrpouhTYgEfZuzgDPMq9au/XlbC8mAzHG3Yl78fBSSkT
x6OJypc9IYmh62C2HoZBzLCTQQ5keyb6R+fKh8eCeUsQ6shizfd6KDcHsj+18Ks6
mvTwQ6Mg3DlMb5S7K4nAgyvg9dNCrZrsySlEDFeuCc198TiB+HNjlES2fCeSy2rn
G2K5vBP2J1bSMaz2kt9sqYIz1pfe07ohq5C8QrRezsm5UWVRbTI9tDsmb8sQgtLX
r/loLf2/n8U6kwTcthqMTt6I+zDyTBASfHN8BQNnE/druHIhVndndgEFQVt9vvoE
BmMx8VFOpX0X42+pMJGwtMuqdzIBYfFYvWlBkxkGKr2pqCi38Fbsi17oKJmFjsnF
9VQpO05qWii/LzttcThp2+6nbJTUFYjoCZ7sVFIEnsAC1QL6oF81gkC+FBUdfwal
zXpokyXj4reKiqCZf6oCVrOMVZ7Lm3TFpO31dTHzt/uCO/xMBE1xe7vocIo3mh7F
pZoUqcTc78MFvzs0H1r1dFqs8xK8hZoODrn1NuJnIDr70ULthX3by0CRrI2VnA9J
/sTze4PjIbp5Y/3YaAvVXnbihqKIqJxhBwYde7tABFe8E8ed4sMJ+Q8NXj4M20dA
29l2uz/baWMfFsRUoNelCz3vmddk14jr/Ntn+eBaZoLFviU73eYl1E+aoy2sfuqB
ut2552R6fVpnVvweKAdzoBYcoX9nFB/3wDLiNPX0eIJWwpofM7IXnLQ+KtUnvNWX
18+t4NY8xjypeG8/ykLCQmcqboDJM/FdcURhbh6Dhylp+njHMQ8P7u9/nwwPXjUE
YXJddFLd1ExF69zMBQqyGVZ8P2FuPP7YYpvNmLNFXJuZDj/LSp4TPhfAIpbyZ4Kp
kSOP2TNkbRWHLDSSQ11LzfL/Asf5acdPfeqrpnEZuUR6Hy+jXfI2pdNBE6TDHENF
ZBaZ97Je0te1HoIELYZ+P2Y8n4zp0glLQQWitW7X2Vi5X3eLqaQ6x9+pvAnCBNRc
sSZwsn3GnlIPK62UqC/2Snwg6PRmw95FXNv3XBUZc3mVLDWtOf/zdoXJCfuNupCy
3erCw/QDiOZyDg5Q7IVJkBHXFp9EWd1kB66XotYRxxoRJw7Q8zYJctpdITVm+etT
f37uocC5uZ+VijsZ0Nha83oSmPEjCerxG8Vv83lfnO4B6MYKOuSNJDxHImHah50u
2wPDrTTGjtP5iNpK+9Uj59mZO5VbD1Mr0+NQImxiC/nX18aVmbRXSWn9Z7XMT2tW
VliS4MWZ+BDJ5KoNpnHSn+8vMx6A8k33frLq6rCHBPFJTFE7XRXLZEfydCXKoHnV
o9DdU3qG9wK9i0wLK/5NITJnQZ8+w2tGTRtUPfxFkmj4RQaS6PbdmK1mHK/6bIuO
c+AcKwgmPTfY4bUEbPsDeBnXZaAG8kx7WCvOBp/wHZnvri+7+NSarWuj6kU5CKAC
A8jgH9IFMCfyG4MPV6x3GNgfms1jah+Oq4uDQ1skQ/8RTILP2jpspBSm12nagF8l
3uB7tF6fH4X6wD8Uhl+yncvWQ7xYJFAquAtqcbYYKNW8KXdznxx3v9upKfOvO+i1
NDUOf3uPMaLvNhI+7c8ZbridBcA2vhLExU2shJ+T8R3BRtFQBTSlYtpY0aJ2kq0U
BMeD5ymTPUDXnJ7Pi9Q4Sr+jzI7Zv8q87f5vGBtep3NtAsCydmFPmJobWKHoZEOU
+VfFXLtEz7BuAIH53zQW8KqAyHINaPWBSQV48YWb/OyrWxSuaZs05heHdiFP8hs+
OqwILodV9zabchBv6g5hsPbScW0dfrLUSHG370dl9Q0AyKxTpSIZI8ddFab55L+B
YJ4/zZnoGowXUTZo2HtZBQ3b7jsievIoOcmx5jr6lvcbb4ZymRYqC79shJ6y5KWO
+EtlsFFe6fMhmNVM/e9N78coEIQzLrVlqTZKhey1Fh4HaPQyjeJLHlmE1nwiNT9W
dNSAHmmR9bYAnSALP5R21Lv/g6GK5ufIpxbbZRDO/hMCXKUo3QCvumXZeMGDR19w
J36e+1SHMLAsVc0NqW/OOChkRcpD2MdFTzKS1/etSkOuI0SXga0nkvB2lpDuO0xi
+yXA3DUb5K+rkAmddS9X4tMbgx+BW9Pw9ID5uQM43noCBzhgsuIfsxjCwuTkWqYA
S2gQeEezt1j65NkSxLCzSW69E+0t9Y9BMqbv58m/uUQRreLiak3tirDQSuCqZ/Yt
HCcLltFjVZKmwslyDuRj1pb2gELgrAUXF4yARqS/9vV1dIy+lA6ibPR8AwvPiQ0c
fM2LIYQKYALrhHjLw4ji3BkmzF/mn+Q1JUZQ6ahxbCRn7f521C6F2QdfZicofkye
nkfnmeKDSwahhM3pmAzXSg283gEPPoH4+xHKGoaEoaLDz1+1LzVVe6HcFuncgN06
5ZVeJgXEo1wtjdVY4n19GGy9E5JyYkumrKS0AizpGtHy1ql/gcaJ1jemF4v1+djG
jm5GjShjx57BCnst/X0/m81YiGtoGoif+q1VuF5VHUl7QR71E1w5Y1xtGckAfIOL
CnfDPajHIxzbyv/PZFTxLHSrHv4EJSJEbuV2W20pEzv5GNryO+NLyXMrYnoDKg4v
KJMHUAN0bDsAaAlvXp2bMnqisra8V6CuzA+JONphKAjqGL9bziMfrdacQt7Qi74I
tUAFwgUkTTcxfOnK5W1nIhV6Z3M2J2A5I8X/MMLakPH4JSuUta1vvHhgJC4yJCZx
DMwLAzbvGnc1uo0ce9yxclDL4NO+ahKpfLJGH165HKPZyjSwYngjRZqMG7f5Oi4D
2873tFGgnT+wOQC7e/ShOi6TvPdLVIg2+n0J7DC1C7A7+nEVFr/jJDkzLX0/cZH2
QtvbrC7nq8i3zrDR2hGYImU/ysJCFhaFlryyft2mgPZB3BqLh7V2gJEbsUvFunav
SMTu/1Tq/LgQK/YBCplzYEZS6UjB2E7jBzhJCrFh2PeBMZRUTuk+ZJOmhaDKbNUW
n/MSmy06WfC+LmdYJ74aNYwBpxjpZ56KRvc+JBUnDw0+q+5Nmzrl7P0GRaUUY7pp
n+xZnQgIk8qzxPVE1WsJ0obu/K8wLuysZ81PsvCk9XCmHJT1Mwl56c13nKxPcLB+
uDIvLGfOnRgCkmRlhygzJB/ULviQ5pnN0AmfMo8sRErsvP/CfvixwM3C+Q8oiv9J
g7MEBhtd4iZpfwRfueX6xjqO5PeRri1troqQED04xmr1xVMoSrpXTgEyWZ0wZ50g
zRvPL1j0FsvfpoiQinvFirXk/YjLvGjGQzF9rtCkrpPEYDxW5my59cZn0TKYTFDt
QroiiCkqWeNt79rnaljf+ONKaUv27opDguVLnB/d/78E5mllreALHJiRvgkpmu2s
fXEFTza20kG932T3yoctEtHkawzNfLT0dd94D3FsR4aDqJphIsuOczCHTKJTF7+a
Hk/xqQDDXkUWQLQk/hLWT+CT7dhAxBeQdk5Jf5hfvEY/hxfi3H87e00PTMtD+QaL
XH9oZBMkkvL0zH99nrG1eEP67vZYz9dASgMTiivAh6gXmp1poY3EY5tepMCGka1F
tkJolVTFCqFaqNjcmQxEZlBpecCXyIHTxCVwBvwTfi0GgpdDfVxx+vaY4i2UH2mM
YBlapILdIkymx5XqmPEcyyWdgr7ytRSv/8Gqk2Ha3X4LnaKcqLLfCLg3ghZMq3Ee
+/ARTvhDwpInzys2bi6jEjJ0DUAuWGsx4nIWpmivcqHwe+dI5N8ncGr7KOiZctYP
J+21jMgAyxflnI6KnGD2gNBAtpI5RTf1aYXunAwvyPdaANxaRh1lv7LLRsyaP27E
Fa0rNGK+h7Iz8Afj+MpmdqsCduA9KIh8VtGutQE3BxmCjHTLLFix8F9TmtKgvaZd
C5UkBFw5jUVsoStJZJnAawJ2SMiLwlfxU4YByH9/Pam+Ub69fOtye0qZ6DloO4hx
OVmPgtGDYEohC6Udr/JKZLaqj3inO/pBum4GvFGiR5Bd4ynEQKIypfCq6vqu0PIb
Vuzt14baTzI7Wcfxo0EuyJxylFCEQ6ye9Lnz8TWT+uXxvrj99Bf6TOa9u2lKuHl7
iVCOZ36BRC/4BbaGLrZ7KwJFTJ9709QiYT5Vig9GqYoMYh2lISzfpZ03I+lhJbqJ
qaayVotvga0SrOngwG6mny6pZ+qBXSwI9DgjXUL2ZmLMsF935TRrEX6Ox+WxyBHe
6+f98i+GWBusSnlHL8IX2P8U6JKBOzdmdUYLS51Ah8Y1gn0tmhsdQBeciUGBxiHL
GwMQD7Bgey0HQr8SCCsNyytdMgcFF80CsPxk4koE3FR4D45wAxZCmMu85pFAAa3n
1xngIBIbfDY0EUm2HxRzF7XEeC3GJtNPfPOMsYtoKvY8qU4MZFKMvPdDSPVtzNTW
TJ4FCH/47jLeJNGZntDW+P44ST3GK6RsGXpU/1igGH5voxjVr/JwAmUHw14nmJd5
11zDJX9azHhg9p9qk6N5bM404oimdKkQP71IbvbkDve+QQIDYeexJzgxWo2CwGit
im0R53OgHJCgyxhbBhXoVE2VtbZ4ofSUch9m9FbkGE8VsNjBTJDwSXqFaN0WnwdT
7ChjnduOVNSxSp9rPcrPr14uEk+22FuQOfYnZplv0/HJK5kNkwVi7hxQmkxALYw5
64w98wuWtFf2KshTC+9fu7CBJB8GOtOQkqgIu1moGpXDNEnpjEHe7jkZIec7owRo
uRZfwLd1AJdhHQEQr8pRV/Nc9pNhbMiViFnJJvM8+KqoIJPVNqeGdTGmOZO+3zbE
bQujBPTgVUVeVI3VL3jUJz3oGLbi9jW0bT68xUVpirar25JEdbw7Ku+TRwtaZNiD
i4IG0VmYppCwBQgj0UgM9yvef3zzCzsE4VC8mjH6/56a0GMV/KIs5lr7uK+qMM/6
EBAPjRyyYqbsHiJLecIvW5DAZg0z2gKQCszeTGd1kYK+erfydcjJIln4yaq1Zmw8
dPaHeObsw/j0bO/kFmDxwQWLJ9VVU5sQqZIP1FYBCG9WHrDH1Imk+66H4N+/CFOj
XM9KwBlutdBk0+n3u3UNgijQPrG1/wN+mmReSaWBn6qlb5hM4B4yGB3n4aoAnTmm
m1P0L33a6Fe/RT4dSe04Pi/z9lcHV2okuKBPRCPtse+yiOjkSIXH/3PZ0r7LFTR8
iDuPrqA6pL5fol8pOvLYYa/C1usFgVyNK1yf6AYlLTeDS26rD0LRF5vD0KGjLvMT
pPVbRHYUXvkzDx5S4UbnmMfgFbie5aq61LI0DWKXn7KBr5J690Z5u+9/Gi9CFicC
j7znVuRqhbBrnh7vqyof4SOTQHcA5IebQyx+5rsNwwIV92o1q5LCjwP3zVxamz0h
KkuGs/FBMG26kmbSBRJ+A6D1DQvxwDiuTtHsHfR3DqKlWh8wue2v/ETOA+GXKPKS
3Fh5lvnlAZ1ApC8ZyjFaf8BCxQmeh1jWUh7EKKrCx5LG5vwJ3DDfLU0w5i/tecI6
MpNYOLYghDiQLUAYHa7Zk3nD0sKnHYUBhaPQfjGXc1DiCsLRzmQACxSUZ5+1qQMP
lCIJBbTTOEsrThhoPF/KxbSioNLcuROM9FxXK2OyRKyxCHTRbetA3dmb5h+eaIPP
2CDA2YQoLjNR5/Vx8EiU9CMIZW1JRPpKSfs1lNOZTg0WOFMAPUEB5fGPWBsoySrs
GJcC6VbSmPIDzKYztQawWFamx+CbLVVozoO9upW4x1zlhtOftsh9ZxlAO6TFFNBD
YHmmknbM4jLnjArj6DrKheOAvWf+3AwQx7MjpWVRRo9wAN5tJYbjpLTfMTf7YkPW
qGOTxvc6/A7NQDb3kFw19bhNqPGm0Xd1mQnM9sYm9zfB09BBwrNoUVbvlhInYQhq
cNYlQrZ3ufrhWEO8BTW607EGZPuEzT2t6qDnZprgcYhTJNPZMdDI0W1Md0lHW5Fn
ume8SfjuiGWJk3tHp9i0VmZbeN702XCY88ssN209FNkb/IhoZ6t6vqWy17Lo0/ei
t1s9KqPwLLOdk2SBTkzmvzKzDu0aSP0oDTtjBYT6iheG1Zv+azBIEo2BIGm+jY5Q
Ec2i4m8gSS4tY0oz99IzO06oE5HEAj6RAB+8H3GH7bZOPAEiJLTOV/uob4JYO7JB
GRxKb+kdrDZFFGpi4S2ir8fTdXEOC76POW+39fatWJUx4ycSs2wuRVR9M3XKsr8z
E2DHNH2MxrklUMTo2Q7F+HrqYrOguLTKhYZsEKk2CnwsI+/KWN2qLbmnuWqbu99l
IjHXWIDYuEXOADAde/UjB2XAnttWhBX5tc/AUasdbCRMs0ODF9zaCnwaIsmn6ZSn
6OWMCugTK2MTR4eYiUIQwCZ1VlvpscgKMoX+C3DWcwfoUToxZkAvhifxdjOZqGhO
qszCK7aWRE0+J4RKECY1a9pWk+Hqpw+1tYhOQ699Hj9PWzHLKJNE5iN1B/tKVt84
qvqcNGiYA8kWEaWtx8guFDMtZOoYk8bi1U19fuUWH2Vws5y3sUaoV/KsB2rLeFhQ
hnUKTLDEfE7mwp4j5mX7xJoNRoiV4UusMVWLMzHHK3HYygBUwvQehYgr45M6tKeh
JL1XD5r18gleBJv4ctKaHraMMRnwY/ZCujV4zmXRB8HICbW2x/BKRwB5tQVMKfCt
8FsERWYAyxyFwcZh9KBIf2SQS7FBrbbbgAoLOAAeDXyHu8TaJ7kt3w2EaXXZ+fKx
rO2Qki1fHHs9Zfk/S0y5VhwkGulzya4cL00tliX27WSDOa94l9rVjAlOikFENBD9
ioW+kPxkvoPEfvXk0svCmTQPtn8PFS5CjJB+C/qL1PGt823t+tw/cisP8TTToRD2
5cUEVLN31Rv7euYPntdvl05x8898CMoWYSvX2P2FIprkLvYkNj1j2Ijz1lAqZEXt
Xuqy1Lqz2Qz04ViyTgaqCUuqZJ/qMyj+bt0N/oYSKYfjd4aCe/UCYrRikjlFgs5R
cFJ+jvatU6r33OwqQtyRa9QJlEzwVIUhsS2gIf7yzRv88r8Lu8jsqAw+9LJipw0d
NR4jhXAiV5y95+//P7ZhY3mK0KDcwYP35phVNtGPKr64wE3kVhnir2VJfYg2RHJF
0D9HiwXbwokwCCx232TZGdsyPZdorBlKLNEjsF16JC5+uma8MJCp3Jn29VA4cVXa
9SNU3VkfwquxIxy4D7KSim0ACU6Hk6GBplmFbYaGMBMa5L+VM0oMHqlHEGNVWWf/
GAhI8Duqyh8pOJgplhcDgBHARswPUMgXAcfRkINoJZmlsMWVBOqHPROHsMCT+n/q
Z6lHJ3UWN4OsxbYmxaNyKFkMuFZPTiHz1I2h2PzLxkR66zeCM4fexHbuQVyaLs27
8Wdi/c5oVjuiGvqsxIbQbg/zm95AVk0FaD5cLxybZVAKXO4Ur/hBSCRKPFiVXgdX
+CSSFHwlDWdYrHMygo0mLnmKNJPD1HKM7DVllrbS3Dlb7w2WwX3JQJKPCWjaugZR
E15uTdVFZXkf7hryr0OvdBiV+RCv4HmFeei2IwM8lgkan6agBRGNTESRvIzKsUC6
p/BK98CASiz0R5SMZznfPIzO7enM+YQaDqBbKgBQJy/RTkpCe6zGENCWYnxLZuZ0
/8OhvSA0LAf8hQY4MhYGO4LzC5/yLa1KB5I/F6pR2kV8eJ/S07nymOyBNhMTJDiw
l/l4z8lVZOUYErAVoQ63paqosIslfxsExFcFcQ82m47JTxDSV8ZpSXqRSFb10/5O
qgVphIuvoW9TQ1XXeOoa2xCguEqJlbiaPoCqP1raeoebJVo0hveYT8fLsEUeDwqC
yjuzt2e6L8OlFk1lqOLrH23CTVyCvYGRol9o26eYe3edsRrK+U00+NNY9pGuiIFN
qLU8FyOZ60jcNnuux/RZ4OTc6N6ogoUePgyu/LACAV7/y9jx3lKpCZPVse74oWPi
SFXwR+PCjqDr8iGf5Dbvq5xWLoxgjYpeJgks6dZJ3RPCJ3dTjMXd/sDi1wpGs6EK
n93h8cVjfYWI1lx/xz2vp3hLxPiv5KL6LNX4hDDz+CaozsUXVXWEJtb3PNs565Th
s6YhHQFNHxwS5ri3AURk9vfbKNdo5V0HMsmoXrHZi7Ryc7Z3J6XeunY3jz6vszS4
qQ6IqqU863hbhlIAqw5SpoxLAvRJVrDZViWbdNOQJ/b9Ojm752SMCUuFHFsaSZt9
1tjWTflZuIhrZkCnmrS1HowPcnlIRyjcm3zoO4H0nbQccP+Bc65RHwlsTXQ6L2Ks
m3X1TAWXY+S8YHZ00MuwXeI+awvXbYK/mzie9/qNFd67l/LTAVApoN4auHMo17W0
zXY4fA5D1ILlpbZROwFO8r7gcrDVlkTgO9UWbWcCAcmu4/dX+O6fAV2HEYA0S+0i
P9B1ZiDtXEB5HPOrBMI5hOiX5pdmXWj9v9bkLqhic0G5HjufbyWeLcSACEp6ZwgE
8IaNpZW6GpdXlgtBPijYfnZSA82FC7qVPV9OK3g/FfOjrvUCAKk2D/PHz/9WdCZV
itTtvNFlItmtU8G5u4F7d4jVUG21eMirVZboJ+CVFsGXFpVbZw95j8fX9gxK9ajQ
qYTzai3dk0QFvdnvXw9nczEjNc5SoeJ3t3rIpGmvzqddl/ivDt8LQgmeM2kM+7Ed
5L0Xvyi9lMA0sN1EKKjDUyNkEWoSAo+H1gnbejspKZXQFdZZQOe0XfTEmfYQdCTp
+qyniNd+/4sUhydl/LrlpgEr+R02/KrpLNaMJDKTvb6ad/fsA+loDHikJxeY2C1M
0eNYwXOsoWM9rQupKgszlle5JJ9vYY3kFRR4PCwE+ibJaDC0yqamJZc6YIYoXH+D
jOwSnVn3dmaRv24vuJ9prJKTUMzataTw7fGbSkMyv94I6qfOB7wgxh+QCnWrWn45
RBF4KDgtpdjd8Z7M/AI2NEIf5DJBOvyBJRod9KH2XowfqEPx+sD3hPFyNz5Un2RO
OKcapmvRQjz3tsVC85krMp0McVG4qfpRAvDsrmE2pAzgegmwNycQSdKQJjrPRQIE
FQ0aAka6VWn1uyo5jm+l+oJsfecBhJIQc0/Xyfh2ggYnGqJIm42xdhza5hVYVZcX
9YXj72wDqg6S1SWMaoMmKow54NgEB0kAr8E45kDeCEMz7JkUmC3fnDjPXIZNXEGq
uoKqSjdfcTvBOkPydJk3rs6G5C/CcuaA/8XJadasgMJz1r5bpSf38pmsOmLT2phR
CEdAmvPJEpqDhkYMmnAX6BDIgO1YFPhVT4r2iZDVZQbMwSk3x9NcuafBc7YcvqLG
2DstvGxGZ+5VXTo6OKNuJLTMHY5MSku3fh4PcKZ9Ufuj+PRJFuwQJcRlHpEWAOWN
KWGmf+ezoUQesfCHVu2AXKgEEPZespoc6dHwB6TBmV16SEb6AuDyi7wWVAu9Sb3h
h6QZTAaemGjG8PkWmH7Cg06ZvlVK4DFummkExdvQkQS60fDsoCqkBNPhXPxhx4L0
TB0JnMgHzSSYyonJNE/o6mSdUwL82hcFgNRSGCczw+Vig87gfkdF8nGLlR03B5M4
PJJZyYRjPzw61hDzki+/dgJSoGVVVdNYPkgE+efxsegjae3Ui4vyY7bOvx2QiaYB
08A59iZ/VjQh9nPsieEbUwz9SpvRp+SrTKnfWEUZv8KVs8QCLwxrFuhhEpAp0TSm
T00sRz3j2SdQbQUhCpiAT8Cs5FcZBHwDV067remC98lmbDsedo5pEhAnMJYfU24v
3yEqXeyiT6gyrlTvpdv6BiMaAO2fpzZTfIYr28kMe0Fd7JpWIUlKt+R1nhANi8Ra
KhwlrcQmEgsZPp65q1jMWDcEAU06npZOHNq6628u88xYPGgkB0A6nJOUxqyW4y9o
qnuS1vxPxJsl8g4vQJgpJgI0VkTwlAfpunRqBk3L1u/40jtJCzMneVr2aINP9Btb
gUwOCAgNnfnXslFk12Wkg4nFuITQCoeDK9wMdIG6BEm0H3egMx13UQ9hzrt2s48O
9yiveP+5ADjgiNp1G68wDaQRN3T9j4pTDLzwrEx23SS28VeYFNwPJ+eg4xSyOK4I
hqnZXMEXj7x83AGdi0FtP2DFDuD/8EE9CrJaxUOG43s0slhaEu2/pYxmIwqv5tRU
D3nShZzN/QW8DL6mdcJ8fgrDPTjpeoF4Mo8Z56T7dUYYkSDYpeLVPaIrxYfCFiiq
dP6jl77YfaMQklqvEfRQ3lBxBDEFEENmNtoSb9zmLW9tMWyJR6dETyh3wkP7PVyR
hfyNpUa1tZKN6m5qNIG0dWM+tlM6cyGYd8MUBRBsJsd5ypg1FxbNF4A327xVLsD/
w7UxrjbZqg0JTig6YBTyVO/JxwcoIATFqR530OLR98U9m5Wgar2We3FE8cmZeIhn
mwKl2Ss5Xnq4tPRSSQO8O6isAwhGxndTk1H6FUIPCDQ5sLk2d+zO0sIx/Be0EFnA
UAlXu5RDvvR1/Kn9arn+V8AqTlmwEerVQGqL+tRG8hFt/KwEUB7iFriX82xBhWat
BHFcTnMx4GzW/JbX0KjnGi1Jv6yU8JH316EdXDpAoPnarJ6Nte/cGqR0pjbZzeI1
R84MAhey01M1ecpWDxQq3NZ3p+QMItUP7cvRm/xXlx3TvdCODWzKfpC9v6tNLDGl
/PdcB9f+7g8Fu3nCRT3+rx6uoughkrD1bnSIj+bvAIJpITdQOPv/NHKZOFdaaJRy
1HFKyXkV5YG4dsV1QdlfVmalN/LagaFuKUVv67airhsqxaMYtR3iA7wSzvq9iTT9
NqC7gp8Bv1oiYCcU9AynSjNby9lPqPPH5PsWQCIfu62lDz06iWdFkwS+pvx/ZxKm
lT3D3UTsEoH7uytEfNAqEFHXslnHlm679j7c3ipNxg/ed4GhIbIYFTPD3hD0aHUt
olAf6az4ma2FIZCn2spShSmuSRmM83B//FyA6d1enS7yKOwPnpgOnzbAV5l4Xvqa
W/tqg6xgsWS8mgjLq/sDw7iOsXr0AQv/nnWRFUXpayGhUM3PDEX2CksziPMFg7gb
o+5e89T0Mw8fldj//SAZ8/5TfUKd51+RybRM4Ep2cwv5zinF6h4wFsRJWVgr/Gq4
TK+cVXr8yUdV5Xslnpp7MHgdEv9ilSRwdqr78ma9zJK5VT2k8uUavG7Z2/QekNvu
q5Kt3SrUVQXRI3YQDCaMc0LjiV3HP/umMcEkSFQvncvReLGsbTlx1utg6YjBu11n
IgXDkb2bpSfVjlJktkWvw4byzuq+fUHVKR4eHNu7jKTzvoeT/UUXOgjpnkTbIWFS
9ZJEq9XxBOxfuVnQm8Gjo/0q73JuO5Jv9BuiB7YzeiXMycsddXDM+DL2ZSbs/fnH
YH2mZDwNP/x5hSmFET4c9mlWZtZyWf2lnmZth/MEcU/YBn5N6ogrkJfA2NrOVlGp
n9YJViUCmjb7kJ+mIR6zulpaWGSzN5MxZ11zt+3BcBvJTNTgESKdBwh/hCZpgB93
YLbCe2vURKEteMp3zL5U+1l5gYdCWoyaJaKGzoT48uURDlIDKfTzlItUshKur21R
D01CIJ8zSVIQFNiKMle31l1iaVIfZSZ3agdQ4DCME9HoZ4QMbhU3nj9Pk9xSPD9p
WI+CqbS1dqhACBAirjYDKkFw7Zs3tAX97XOBQI0OyY6Xhoyz6Thbg4jgPwNt0mQU
Zquzbo+nJSM53w/QkJGLjfHbu4aXNLM/Hv+WI8FnICT4m9bucaWmHM1PDQLBhlxL
Oa0lVFwFcSuMrsWuZrj1S8XjmYi2+D3GxVaXxSKcwM0jOURDQGZSmjQDa0I0Z1mf
JqNiEZcn66cQ/QmtFTWsSyaVn+O4SlysgiplTAgvj3Fz1rYQnypHYYeN5BpAcVi4
IH9L+yZh5MQhXaV/2jmr+Sydh1Ns1N9SHL8AcYNQRN5q+uEGLH0Fkx4Hf70iv/6Z
kodvln91wMYw/G3MHoJuKyPxG77AJ/r2cvFpl6pdjMVwEDyZY/Wz9kckr+lgQBhF
bTw4YvpWj2+VUQYQ1bwrNqOUqXR76OI3dAPtHEevYS3tRn/4Ub88m/6Bf6zSkREa
kcZI2hzAZZ1iGStUgVXh4ivx9xnpRE3+zHpj8IFtAWBOBQy1O/PLylwN7XHFqlOO
J7BlPVTFhcbbuuYUFAWp1B2zjpOPwcN5lKqD+eOxqz6aK/IveS0g8dckP0rt9LE/
ima0l9ejLD03266FmTJ74F8keZMaZl/Y5gliEGscN2hFmm2l3tBDrNot6dk4LY+s
0669KWurG33T11KDut2265ueG6kqcUtexDu9PAN92LS5TwV9Q7KUNgKuo5XpM3AU
TnM3xB3S6YE7whhPNII5jL/taKT258HHRpaRM1sWa3NQ3na0l3+5qNlRJt/s11S8
yhaBPcKk4QQXOuIZON+k+s/9VWNAPYRf9etyS6Mv6HfpT3B7UfyoBUqapHXtKRU6
jQ3pPM46FvQfm+ybOPzigAMwbsrTdaC0HdzkDUmZNBDzVK6eD02U0I4RQxocyyBN
NP3zXgjKBZFGa8Z6M2GNLrHsVKfxysQC4UM3+h0w+wiY0TRB7vaI92ajhiwczYyT
7D/jFa8k77J23BOqvO8d2cZshutq2YpT8vQNonXRpJ5BSflg6hOiZC7S4OwUuqkk
owOJ0Hc9K3hhLfUX2LiwSVd91+ftetJJlg9XiIAJHUnmrSQxt5w3CF9VjQZmPgPO
MF+3dpW/fCOCH9lAukRF/X+rqnVZEoUeiv+PiXvfFvkOCYpWig81eJPAhGw6m6sh
HLDHpYqamXn+xrme22DiPHy1i+3SFQpXVaZqR+aORo9lYt6N1sbzNkSjkkpKsjgI
4Yy6+iL7dpK8kMa2MTHlSAL7EpmJoMJDHhWwlBXbdA4tLwNKG7txXTi9E5xRTydl
uVrqrU2DwYF9d587MmdR2dFEjuBEf8wVNHtZgbUlSSPmqm/LkX5ZIpzwtvOkklVe
qUc1zdVALAVAjQVhhncu8L7vvlwY3wtUj4e8u+Q/tEk9PVUpzn7rE6fxa1AXP6bL
xlVX4s8AVCwUp3LYC80MnMIzqnFap8sS7gW0meTg2U1Wb5VTAXQbMKAMfKyWrvov
m9Q2s8GwERTF58Ikqynz+xVc1Do21nfVn7N/XgQxzAK36MkZ76JDmYoKTu9IlGVW
RZoAHSiiBMli2R7mpCL2CGyII18n0o5hKciDpMQvHU0RLlZnZ23Y2fFSOmtKBLTp
MztrCEdu5RQ84cxV522OpFCrf3SY4gCeh/iBsLvD5O0UN62c/GrST5djfJ1bXcNb
9G2Y5XzbByLn0vjxe3D83aQ81GR3i1uHUHW24hXvjOn/nZXtmGQNwobb77kSmEaM
2NmxZQWa9gU4u0X+IFOq0FI5qZ53JGJKm38G6ugO9gyY/uRd3H0jPpgs5APrycwz
ecrV9Kx29bmtD8YCJhFNIlYEE6c8TfkSiT6hlIQQ1d6h7az1JnY3WmJrFtCFXfJ4
YuXcbQ/s+UzKmwdWKJiikeCkqL3T+Wg2mSebzeTLO+cJxW7bw4Sj9jbKPrpqRVem
rr9keYh7wzwNWxyJArKfjogLJfoJujdpHbsAj+GP20Ia8e3aUCPtUybx8bXDe/Dd
jjjcpVZH5NFaSrrykRWCmm2x1T/fwyM3DwndkH/S0BvlGV4Dx+qDRQ0RmSUlivIs
BFWbQJCq30Eb/tAMumfO33zJ5zJhqUB7Hfwt+XObPYzeps7CbH6b6+NdavEDSy9E
1fdSpmPW84V9B0fi1bHW++VJpwXhM8mJ8XYwF600Px1fpec2Oy1B5q/N2Sp9v/3a
qqXA5D2wRPx91pGI0l89NNjE03qZOlXaYBtCdDcRrhGjPHhdqE1+V8Kdt8zyzCOU
+WT2RWiLn/cYGz7d1SO5/X+MuLpJd4bFLmEXlpiCgc/Il8FrOvKzcvwuDK0l3oz+
oizmPNFtdGzCT80g/77wTZmE7kC2CjQ/EYIJ+jIyLBK1ppS4+X0E2fkz25wJPWSf
2/6pIHBv1+/qjo3fkbj/JJ5Ikz1Fo9VXUM2H2m6Or1WBy5M7Kz0sEFiUDb+K57FQ
OEmUCToa4nenIgwzPDiLr3cZyfCtmxRAnW2VO4CjtMzm2mN4IrHA8WSKruO8NLo6
yFmW9nuPsiYLFdkaoMX6MaSHSO2YzZKqBwGauGeLGeylDvHMQYTVlr2snnGbAUT3
Ai4esGrCneVrYsK+97aZ1PJkrlG61g+ETVb1OCbWvzRwQBn9fRmgF2f6ISqZOKcU
hLhKWq6yKRz4NYpX8lRsw3rsK3LT1bbYcdO3bMOEnSTVjlBsk1X9RRRJy13QGTK1
DuVD0B56sfoc685GfrbSB7pXsGLlU57DgfUW7sP6oLWbvI5mSGj7voAAbCFA7jqj
1WhzVaBhFhjGkB+An6FrRjkyN3V6y+R0/LXEnBd4GsfsnrAXnvV71T7NrTzEt+Wq
XDDB9Trz/D29vArHg76HjueUQ1liPLE2TstLPR3v17bcoBz3phjxq5Mla+u4n59e
T66HyV5uashPGni6IMyQydSSSNHS9mMea42knudNl7R+qRAghtjUdCq85jrpF1Hh
gXG/EovLzCwjOQQxrIcapd+xG0oY4nP+HCIblXdnpG/k0vV/quMpcTynZ+9+sz04
VXIRJWUCUQs2gZIKLKWgMx5xEohpDM38CY9W5wWbJ4Lu9wjuFfDGVZIQlQZbS98P
Tn8XrvrrNtvzZvMzEW023hal7nytPztbfwXXykiqVlDCIW1Ne1I3bbLXiDcNoxUl
+ERPEPyNC9wLgnE77MSs7TveTCIi7IdhUkxINQwnPF6QwvgeRbQi4/cyPLGPEC09
cBZnHy6z7/cUu6zetkYv2mxi6H3qWsp7JIvCIPVSigrBsZdhhHcifU81bljUUfq7
O2o0ZuWC5p/6244WWdhOp5Xg4R6Onk7gsc1Y7CvAGpaBGwmmX7l6RY53Q32Jw8eF
tdfhuVheisyJgS9A9or/+sHDwiPwrfEYXM+IJ7rOw8qcVoTKLYPuxw21Jn1L4auN
BwoSZOcYd0tHkVHJuc9SDh9h226o3rvCYmoF+e3aIS8MPDZVYT3vQoNsPab0igw/
OzdxaTBMACd9J0gyDdXKAxRKv1oIoV5+5tkY9KINeRegwnEAibETLLAC+DkhmUuQ
0iic12g5I8BH8mjEI/bJWL2FeE2UbYIk95DJLyw+jAMMob9j2PXHONDT9uj+c7qC
74sZP25w8Ev1UhN7vNLBslahqlLZDXGRh9SFUQJvHsPL4GDMXcT82dgU+uIijtQV
QLnsX5WMzIsWX2rzL1u7dpXYOjVznQm2MCK9NmDNMTGuGdKT5r7GWzz/we/0bXr2
8gkbeyX2IDmTPtsVozEROa1+G1SdFLLQBVWt3Sm1WkSd6pOkY8xLnmPiS/YEfF1G
iqNVwEiHnqcmI7OxwdmJDGsCxAWPQ7MVn64H3whR9Tu+wY9ckgm8cY/T46lrp7qH
0bHFv3QdqmlFfExJTA0+YvX/3r2GLFEkMRxh/p6AmbT9OorYJZPpO2W6gzBCT8gO
ib9sjgqL4LAgw4G3bnygA2fq/Hu/TenVSYucjptIE8nQP+SMUyk8rMXsJBpQUu4D
kcxd/doCZydZzhvWYf33tRVRvvfhfpDgMpQWVNew2V3mjKW0i4AcRQipObgaT4YW
q3BKYZCfCvW7HD7Oo71Lml044EuDiwMBIk7fXlddn3TBJphmlhYJT7q7W22noeeo
RhT8kLxCkdYfNm5tb3gJHc4cgAu1sZR87daQs0bFjuDfzPhToqvtcsqyVgjQHf/8
fr33o1yBcKMdus4dd63HybLx1bM6nlKSw2zcc2RO4+p4kv86OCpTjD7NPF5ADdch
9uUI6pxj581CQgWk96cs3C591epPVyDmZ2Aos4PhTfyJ4iG6or6BfQsNYiFIv3UD
DO36sCzi3iuhQkTJ6c2tcM/Hf4I4r65m52SyU32/CWx7l7s6s74+wlbyIlGQah+U
kqHj8eV/bJfzhZVfBSuHJxshmylrlSjrl1+snFC96Dh8F0oARW3fnLgmVqQzXFpr
OfGzbr3E2bTMhbExZibHCdpshzMDRfTU89Oo/SEr9/pyGtuIka8FflWJuSLJousD
SbZ8v2V5AXPzFmwzly/UiBlQ0XVlqdqnYqT3+s85dlpx0iwu71+4Z05vcTsbHD/G
DTQEXQl++WewXOHd617mG8neWrpEmHZrb0YwZ9tZXI1lKRgKblF62qJeDy+me9bw
RjxCgFfAbOkjbJKwko7vF+TPiE3vwmXXFFL4IbCOm0blJy8S68LKizTs5WU87rbN
IB6O+WtYyWGedlmz6nU9nqNceRHD4pYObCtmSOUBJMvIbouLM9lPZ21MjWXevJa6
YpNrSRN589Qcns6zv8ZYWwPhWh6LPb/9A3GsnYKK+hnsAgXRMDUI2h5RaVp39EkZ
pwaHIUvB6BiJiR/Dcy5StUUa3GotjlWcEomQ3pQEXVmK08agbDIpAXg9I7kXotDr
UT7OqJEL6Gda2CYV4QuLuPUkSPyNgtkIBk6S9TR5USFXQB7MLov7Y73Sivbtq3f/
4n6wmkhrC8pXpaINkIegCjWMEHDWPtmf5BeoN4xOcflQlEe7rWukn7w0LgIS79a7
QiZQCN7IwVOi0tBYKxlQO0fIPzPfG04lzeHNBo/4VeQ0aiiLD12B75P7C7x3pXno
wZyhXN3dGzYLk6g6cauqfUhYMcr+xc5xfPxj4B1qneMmzR/PYoD+QGHJg5D4JV2d
0TxKlqo1VXVUKdl2dtVH2GBtqLj1ojtCa40BYEP931l3OQ0GGBRIKRfJB2R+hC9t
GFOhycgq1TYLyDmuc+1Rwp4vs8GgUzZMW+KZEslor8I34JfjRqakiEIQcLCE0oQf
UWx8UzX6IYHhdwMBKe3gZGEP0LDhcoXse2MuPJKJ8wmpqx1fsYTLrDxPcWMEHDL0
FU4ho5Bou4PyBOSSp5YWsQoOMWNLrUkS74JleDndmLeDZE94IR59HywfskkhoiTm
RgjkpiqXej2mtgRf+27PVkzZj8TVT+XCD4KFsynVCG3Ek32VmDZrqDAD+QTCRjku
p+NKmjgMg3SZTLnCnRpnP1P1BjAt0d53ag3D5Gz5F3kOsZc79MfazEYpMTHrU0zT
+SJ5j22z25CktWWnhu3Rl1uduwCTyUnV0eRt00KQid0b+GB7Q63Sk3K4e7LsZqqQ
552KrsuoaQiMMwOy/D4R/1nM4Fzj6R+AKLkSmfj2yDSoSsDuSpdtG2/ITvEoH05E
LsBc+Ndw5W8tQCS+HQnAAxuuT7gicY+Vwnoh3YPprjKR1fWQBftWAJIYJ5NjykBJ
DB/1Dikz+y+0TAIfIL/Ib3hbLb6x8pvc+gggvdt/LjvkHhNBs/crYaNibeqJ/ifY
M3NmosZvInsmAT4yTis1MMLObC3/at7WHCr6O1Xrh2bxOWm0avhfZZbaj5XhwMbo
zJpJ1Dw0727OUtDrOulMXYVLzX9Z2dhXs6Q5TvrZ0BCzUYEzQVKlIx+/GTJPoeOo
Jf4FRbxmOpYA3G4pjCCL57JorDivY5hfrlc/H7CuZJnf+/vgWaLkyLhNDwG8M49G
tOi4AtqV2of+iJn1bbpGgDpbM0gbNPK9MEkpcDOj9Kiut13coCnOQWk8kquzS2ZE
vFhGTw5izlu43k81ehqiXMAOAC6At4DBhO6hBGCpdwB4yCfYZJ6fRBFPHXG7aoKb
s5JLAi3Q2HaykisaiGGqXKY656F95NNNnxFE8pZbFyMxZ+cXOD2/WXAXZYjNoVeb
GGqxLvYID3XFfehaR2v6yU5ROpzAmg5zoUzIUW8i4ZEVz18b7jTWbcP4tiIeCjgz
N2+ZbI3Tv80P64V8lN9ph4HYqjAuJMko+LIkRB0R7Pv0HemtS7W537UCINgorRPY
m7I0Vg78o7FI39ySwBs6fKCf/sNtDC5gd4lox9ZKuJEG0fjhYnogezFk279ki8yo
Vv//tarTzT8Vye8hGkQlpZ+P7CXS7h0MO96/xdgcUgtcQgz/zuvRmZ5QC+CImwd9
w+Gd22ZCb1lJ/J6JT57aZvMUJ+K/fM7YQfgdzoXdj22i+lR/WEcGagzT/ItzoRcF
66XU0hfLpwHoxoPx4iFyOGcFVYZsunFvY/uD7pYI7JO5yY0bTyFKeYNZzFaU0Ts9
W3gytBlRFu5KDjIBHJAN7Uju6lruXrNCSeeLWhMTkCH9N71EAXd8rbgov+6hfV1y
s8+JbntHeKmir8ncsHV2AcrKrkCqUUYQoBLq7OepBGkBQAz8tsQn/BLEFTf2utp/
DOVWH2zmzr8cW3QAsuGNlVmvH558OsbE26217R4QdItJMLlbLZqJiVwhAzlmIvPA
VQM+plvyIrufINqEf7V2dbhPhkzsmNVedbaX4mafhJSNwREXCq43L1GhB6l+MEii
mJUOg8tMjAJ16gAKScgl3rVNMLv+CDMuL6JZi61xjyZBwFiP60/bWkUaJPktIytQ
xluWVzZzNIijIIXcwnfHO8PSHDnqYqv1HY0JS8T0z9ygHVENh83hujyzmDo7MW0c
GbdU0y+HIJwtjnmXo1tIOXe9sUHfB/39lUMnTEjBxi5Oty63MzlcnNrM1uZsF0tA
vzsgPs7aV/wZ3S4eghiAuYqIpCNbuYy6spiRvbUo4qY6Z4vPLNdbQUoo7zQEeaDP
gsXvzKtPe6xlUU3tOXIfP7UvHpbmJdGdFIFIEYCpSvbxLINljA0mZdNrMD/wZ516
TrX8unuD7tlRpY5FViPAjKvu4yaUapo4AE5qM/YDDiZRV/aWMZfgcZ7CBoyzQXfm
abXqkmr/RM0TN5FEQlcijruNryNmu74KN81xXRnggRMcXzJeM9UbxKLdhX155ssC
QTArRQqi4Q1Kzgk0LbLH8WjtXiYBq7blBT4nMLVsmY8AvisP/YBG0sfz1AT1rNde
nsEQLsCM43QMg0OQ3nR3OIy6+Emm81/fn+xP/ruZqvC68fQKaCKjd2D3Uf7jFz3w
5+9o4hp7km14cOsVGveBOmf4vjKN+Ysu0uIb30jn+0XzPJ7FvdI090aX1tzXAQFq
cYXNqO8Qb2e6ChMqVcDGiICm+JO1KFEvTrMYjDmf3KRoB6nM8wgiPgghHtjeGHyq
35Phzg7/H+CO7N+Ckaq7lNXDJPoHNeOjsa+9D39GIF52U/PHAZpACwpaYAmSdkka
iX6gr2QZvf4LI71/oaMdzHe1IbavOkIG+IrdldYRPAKSHM0zyc+ekxd3e0PE7wGw
+dKvqafABpNZDQuh7AjoAS908vVxo20Mz66IX5rCaMT/n2tuJWTj4J29C+4DHU/C
8t45ATQDdo/agwMEZ30coQBhGZwOwebRty/1AlLmfAthAU7IXbpDkyptu6eNSMh+
fmGmtM5agarcbV/IWNAiHjsbWnMLuhgpqGh7m+bJMC8GOC1U8VBrwXaEMhHCm0Ux
uYHHdJ8GkerC1odCzJ7eb/pjs3jjJRM0MbS9iPfN9+Q6aqnIj2rmWeSWCAENt0/H
gipX+Inipfr2nQ6ZRbs7yowdQ7WiBUnWR/l1L6UqpPByeXcTKXBmA3PHEkY+17Cm
gv3qvhhJorAWtMyoYdgEB8iQept+CgFGqBxUxwNeYQT9coVlZh2jqwQtVkxLRRhF
yErFijEXfyXty0BEyhaqk6yweuPKWDF1wxWH41PgU5eCkjJocbG2fQdl858UJPa4
G6PuJaZgDZbOSq9+zfisKSd3XUMq2x5xRNluPp+H2NM1+7bpk6WDOfFj2XXoqtPs
vitbc8eRMNbDRhCGcoMwkdQhEzhFuj4VatmByGCHzXZESG6X9X50AXvMyDo6Vo8f
fgx6pGqrIC+ZFNhExCGLv+GTLAdtrIDGy1uGKFbxVFR42OG7gWcF4eR8Kf5N3tb/
6b0yP5F4Z1hJ7T3gTi+cvFsaNUsnPsut9hLjr1FPz2lQ7ljzBhOnj30YT8Nja0f4
PsV+ub5SnsWJ0UUE/c99fWYlhhchpIj63xDW34psqfXDihYYgWYKgcEDUItz323w
x97qt3yC540SRKMuk1N0YV+EfYPXiOKS9rlE2rThIOTEHd3YUD9sCoidE1Py34w1
tAUmplK4sO/WwUjoJg3wf7sXSpDIW2sTd0u6mMF1QUVPFdVA3YYumlM9MdJddIBP
i6ZHeFLDSXyYcgEiwU2YcqwhtwsOCJFnqE2g5wFj6w8UyUulAQ9/3ApuPZzWBrV4
rs40j8GEY6wbHDQmodaw2wIRws5DP+85tOdyTn2NfKD8JksO52a416VV1wGXSpqw
ZmXjVjodrZ1Ee1y7y/7osDNr7JhrpF0qXBwCPjxspAdJUeoQjMVc3T5zXW7mzTE/
rVXbsb1gxsJuf4lAa9EeuiC8SCpf1JVG6uTJIEViobr1Z9CBKRfQvb+OUgoPVYKA
GNdLJequuVRUSHiMztwxkmspQblYr6W314s4E9KzKHTPjvRwFducHknW9DBVXyUM
Vz64o6JSuRN8Fm7cjxgoLfjbDrb1Anl2IDywPlNZt47fsSdkNhv6+N/b6KxV3ssE
R8jaLy05YEp9JLKDusR1aFByjp4796v8ZInNqdTg2YtQZsKPNEabqQ66jj394aP5
nlsQ5wSmOqieWySvuPyn2Np4+P15ylagK39fsg52jJwNFhOFcN38w934lEXINSvs
Tw/l60qIBKXtxC0YCcoHQkIZo/UfM8JoIOZRiUc7cXCaURdsxamJK5RE5nEfXlbj
+X+f25SXSuyJifGVcJfTAH3kHx+VRILcJS5ERJ634HFrztH9YRSvkYF28LLUny59
iSR7FdhOV9aIrfdEFhtSDlTrqaNrW7UC0m8zN890UsJcKo57U+lpMdI7kEZq8PUB
3/hIKT0puwq9+Ude85PA/G1XpeRDUtXgAIyrehmloaVUhEGFCsZQxgPdANV7eBtN
7fIipFiBfjw9wE1Y8P62Z+rwrDyJjwRRWcgo/YvHQKoRmUSoDuNQCdqeAShb8T5l
P3Ks5/+bxMlf2ZxRVcD4rmRfDoyfnvkR2XBeLVtHjfVT52FY0Ei7fCPHhOXztdiN
fu+b3VzVmYzBqh05s3CIV7+Bv1hTKKLAa+9YN05Vv1HEGI5gHcay3dph/xkZOKH6
vunxkzpW/Qtjya7e6ElSJNocYwY0Rj3yx9L+R02BV2697cftb5tqBK4CQlxwoaAU
m2oir+rHxwaV53rBggnhOfac/zomK8/QL0re5iukKo8XR69k3S+iTonUSf1BhNdI
1HM76g3w/TDGPCjT1FsCeCXVuj77sQIneBejP293gME40ZpyJzSd1ea2RO2c8MIH
dNXVH7Z8XNgdttdPU5XDloNFaEaRhoF0xMku6FmMU40T/kqnLlK0I6xen/yP/9ml
yrl09f8jceXnwrD9xRTCj3CcwxhUJ1Ja+W7gkWMuiT0iFHYFQ6pKUgEVu6ZnKWmg
ME5ySaJWy50lDwWyff6qAy8+w/EjHS7EBqCEDw3iAXzs141TYGpyEOzXf44/73vv
kuxT4oYTk+gOwh4rjqGKPEX10tcmTt1SxoOg3ufwsshlA3P2XeU/vLEAIMbCFq2b
ADCy/1y2a7iSuNJvTklXt7mx5UckeVgRAM8mUl/agKqOBinxMw/2uSCTO/OeDS42
NPrMEGn9SJfo2gb/NeMyLvEI0nW6MDf4AXzTy2cbcOHc7u+VbCJIIi9g4TMn5vrp
1Jfp2Dr+VKnB2/yZWyv/pOcTj4MhmDH+i66bXn9yBDtwlQy9wox7LQPHsWyYMlBX
SDVPl50IMt3+g8afn7ifGSMm4gfky5KqVMH2TF5UVceQXswYPFDkJc12yL71lJ/i
Xh0dRz+GdwfkertvYFzqNLiFZXTUQthBxLNvriAHfv4SHzMu0OEdKUQYXacuYkKM
wmbIsmxPwQWJH45dxfEXjKRskMbuF7OLl/ZlYpjRecO8IX1VtHE+cbSkRfH+QSun
QuuyCFv30HvKDx/vEG5Tpqj3Uk8X7lKIF8L407EZn08fW6sc07ecTVOw6/cgqzAs
22c3iVLMWT0cIKg1NrNNHnu482usoKqdtj/3J8Bh4wiFkBFUUb6V0DeBLIlmP2IY
hZ2UmPBHLkADqXRkqaZIJM6yvjJdi4PGBPoL+fVYnZTIV75YzoKs7wTcfQrf4e9t
Si5Z4V4lh+xO+cOvXoH9kFBr7DxXxpzarXEm6CIJUKR+2QkWW0haj9cMpTm5tpDH
CcY08FFTA1SdNzcc+3VWDiHnZs/unuDSTtirFFS47OWrFo78RUpXkdOlVKVHwv5W
FfCqKyCDlT8FNJPATdH1kkcmTvUJYPaHz+OsZcpvPd6VsUGPewcx5Q5aQGYDDSss
YYKJTj5LWXjEakaRt7InUZHSmCsIb8RIXVyZvHegfHe9RYvtWWw+tOCQnm2QOrC/
B/H/jrmvljEGY8bjBXUCvBfoCp/kjuj/yPKnsmkbnBFWHzxAQzA9OQy3VKpVYYLR
VtnDP2iFZh0a0cAmNMQd2gVCFEXh6ThaUz2L8HJTf/kBt3fszLLVt4E8R7JFT6Gj
V8ona8TrfHEWfuMqmBfbqGp0tmK+Fx8iqV3Es4Edn/0ZesmfU91CrOQnqjubJn+B
8n+YZwgIHQgdasXBS+vEfh/CowgZYw1P8U8c2bqJeT1RwlvX8clqTtxVnGMPPgeW
YOEgJh55tjPLeZ83r+PeYExHUTPp6ZOD9Atfy6OnMRrofbm8J2ONc9r8lv+0FGUG
62dhC3SWgQDpbGXivC6GGCZq4KHT+/qWBqu7LgMYyi4SVexj70XZHlTH3HBHGHoX
Bauzkibi7vQBxUkjJ8VNRVe2wGB++PKXZBDI6x2SkoxDifdHBbVKXXvchaM8Fj5W
Qxlhlwf2x41pKm2evFfUgEFj2uwM8gioVikpZMzWn8eVPPSsQj4wdsce0RwXmx6i
qKCggJloNquB5ApKM1VI1tgBq6wbpyjfCf89OgdMZ4TBpJCnsfratqikcPsvVqiD
mQN1sk5UOAQvDF2sM+EBpqVAGXuTs9gI6F1W4Kl1XrQhAHUp8f9qdjdRK/rYpTKO
EKY9yc34eudbFfYJCMtmpuNKugHR+hJUapjgtkDJ7CJnMt8Hw2jEpSK+fJIb1dUb
D78a1kPMHBuhXPAnnDjWe/V/EgeBEQ2CF1xZ73CxJY1RLadRkGSQJVA8JBkFv4OM
VBCeczRdca7iKr3quKniaGXqmOMkruQ2Hg9r5bBUrbep0Zwwy8jyZkhxHqRIy38f
+KtVVjCu93FPOReJUl6dmINZF2mrzruTfFBRFZb1TSxlJ+Wl5fvSbsOCHh2cJRPM
InXd79NUUCUmOu82OcSARufCOajf0oIR9VS0r6oVRvtWFV92+OPAr/69svzweOD6
8n0OnLR5ONyXWW9mTjbsQYHWBTfFoxx2bm+daQbAER9mCLokv5YtJ1zbyv6QS9JK
T2Q0ZlGPgF1Q6QA6Ptrg04OR05+TUo9zwBdjshB53AvRCxyap96+IyXEhdX0H6hx
9xgTWMB8ChB2vo5sfrE1oH6OrHg6poLNfs7Sf8bBpbyT1KNWKDqRZKfI+zaqAAz5
CRodhejTaNDVh1VgvYxodRAtOCIpZJkIyB4Anjt8wP+576OnnpgHDkaXEiSmaovM
7Y2TvwWG8u+8ALvFGDVlhVS0iUW2jaY4MEhcWda0nikj93k22oZ8iFUxrWwq1i1m
93jtxNrW4EXg/7R++LaR5m5cYofx6q5gXpYlWDo9+e3JeG6EmXalowu7Amqex5Vl
/+tttRkRiVyfJx4jGq+5sPIHTfWlkCU0Jvm78nFKwXCVWvHOMU6hC+GNQMP2gXs7
6Z3JIe3/OpiXdIfh2H37TLDtCtKXQ/CXVFY21fROHC47hwjp9eKyNaX7cwWvWa7K
QSP+ocwymaZMxlTFARZXNksMIEqJCMqKgmBGlHzpka6m+VdlIU3XvN28akvKH80f
1XrJzEG3r198xIKXCvu+iqJz5DyFLBeoK7Xw5y9JLjUeZoNisX2SC4ePB/UDQnzF
9csUkDWAPut4pamblphIphFyEpClSU6O/kgq0KwHoStRP8vduXmM3FNgGLU2nDDk
tQghpYFMKpDR1XaaF8jMyIQwyD8QVg0InooqY69CBmPy6VI3tjtxSk5bGd4OC+dr
Dtg6cFI425S3QJJqzLtNPivndntjDd53DJ+yosxRRvV3/a0qnD380/HOroe+Is1P
K4PCKfvFkeYRrJntp/kr+eNyFH8oh5Y16ojawZXg6iz2AJNXGLyy9b+kbNd4GX1w
3Mp8ePj05XvdTXHU3RXY2XXOtftejgOedm5A6Fk/vNWm3CVMITSsjamViWdaw3U3
QIDnZgqg66pIHfa+6K+ofbs+I9T3/wnVUjvpVux5G8Tk12WFwz8EiJIZkVuJH2se
r5mw/HU3BW4fXPJcgSfwzsGI5ZSEVCA31Cg1HdxDEtQsVcYne4h7Qeo9hmAaAx2F
WwVOm1VWs+Fag7f1TWVa/QSQ5mXzaKPot5pymmdaOEn47kG1RFuRcfoYLvfvqHk1
mvhSSWM/04gWj0+jX8um7Lrx3PuGRNmVUFw9iSOtP9FEUJslIIJ1309XZ5WWSQUb
Qr5iKlE4vU/NuXE4++aR5BMvuFmA3M/1uR/m+li+ew1NT23GHdnN0hdsWGMVR4nf
VmL4D8Qp7m8nZT2qdFwuNaQAuaOsGaA9s7MnBmLNMciT8/6igE4M2uIHHNWezStF
2ZxYiwxZlExCUFalj4JIqLpFjZYtQeiZl3OUJGVNEDtw+658fKtTji0pBC65n4uG
zxdGIOywrfXNg9TYrbtm4SWnyseQwjJoYUYY/qHXXeiHf6CiDql5ivP1pKCOKvOP
K2FqNpbYLpnav5ThhNbxqM8kIum3Z9yUbI1/+NZk+gjh93bO4nlvu7I+pkjQBCsv
TtA2VHhvXyGlxW71FYHnwqjlhpngB55wdThHlgfh6BtGITkI1i19VGnm4m+f6wRz
f+2dG4XfEYETWvrkHx0E0Gy2dLaLGHKZh9CCAgFFOB8kMlWs1ureqfMCxJnA9DS6
ICEcTWZiETrnY0kb2yHxcbYZjlWkT0DWBAJuxcMuIYJbtW38cEtYpqWVHZ1V91tK
Gk9jDmx/okvW/Yd9sXXqx7twhHFR2lWXqgJW2V/r5d0poHYT5hogrxK8uOxjBgtT
yHMyE6QRcZVLQ6eesr+nBXMiFQ2cpzJa6jsJshMegUzkXnswpAQ8ZVBYdyLIoqJP
3Q+mz6tCum+1zdlKq975850zTa15Uu2ArbsfBXobhz/RNMUM5Qkili+I+UX41B1K
ZqA4ybC7SoBNk2roiI2YJiHaaF74ZjDHT54rqHMgd0RuKj4IWybKpOf59g+Whr8x
Zo7yIRul9sIruY3DOp1fdyfur8+p0HKUeI+1D2VmoGqEwpJjEGiQim1VyNBvyvVs
M+LToii3P4skOTsq0TndwQHfuBhri8C6ijhbbL3Nd82MWLadnrPk4Ak1B7OlaIal
K/QIJFsVwB7g0/pRMamBrR86PeQI7619s24CJ4gveAtQ1jkgK/B0ckQk0GpW8hgw
KfwrJuAC1b1gbmsCzU+2PK8RzPkxnQd/Pg9B1DIwRZO60lVclkyHdtI2dX0LpA9z
aSqLLD+SsmwQS4R3msWAjxaHIXUMMs/tHWRFodQiHXb5i7P7UXBfR6dZz6J4yiXj
Yp909MlYML4z014E5EvSViCsZLBnc8Y2pCFfIz5Czwi0GEpURn80FJcj8JwgaQhC
81W5gtU66ZXtYC6WNzQ3bKH63ROgU6y7mocweQO2c1ur7LfNLQavRvUX951NG+i0
mj3NXbaS6NhBf8mb0pzowAYvQ/AOR79ppxeLXLX/hmHlLkljzGz/veJdbltUTlqO
Aw4urKe5RSdF2nJshv+WsJExOpl9bri/LTto9tBtvpspFHCyzh45YblGGEA6Vyve
NVJPM3DHllgUI4a/PBy3HoD0F35ybCs5JLPPH0n5dwmlq0pkf9RP6nvUmINvQxtZ
yrlxkIBzPFBWfR41uGHR0w0Nygr+dU1YdE/7R74SHnJ1D5IXCiCHAk8RdlgBx+iA
Fm1SEsLSt64QnhYK2KP4kIE4NMUpCdqrpSTVMkvEVHW0go/WDice2y4G7dqAkuCe
hcpIWVeN2Q8Z4GRpgv0l5exvG2vTRQQbLbzFxmrTOWbpxmgCL4p67Gx9bna68jWi
x7Yqh17iffiIBYh3CkE52+Z2i9ioT4rHSfLP5eBK673pBYfcLVv3M/rb9BK9OpN+
zfpVQtJSCRuQ3j8HrIaVdql0giRMkklmpHNuBmjd7txaEys0eTYzHA97pywqK6uC
F2Y8H+eZ2FAVjGrIE3L94ZttppC+Jwd5A9ShHbeUCRYJEy3qX+J3go95E6StMCRy
qkajgmu9BQLlRfENpd71eQ+KykxtY550/YAcAt1YBw0L+u9SO0lT2tU853uttnHj
D8Je22XOjmtY5jYliT1z5rY/tYeLl6KSG5HnSO57dkog0eDWRfs8JqnzZQ0EcS1M
Qov5d5cxpS6fF0q2ZLXWVqW9p3V27cLPgpZXBjoLs+tsQ+FoycR49IlqZdAathpr
w7YUS4bdY5FZ+cx8z8m+Rn1uZMwtsrgaktxlKbHIvto4BoZ3gynHwL+njppu6vHo
/E4E/5b9+YGMNkYZEoGS/7hSPijc1+tWFUrcfCaE2EkuJVkElnyaBFCmPUoKzLpv
dNMEpSFQx4ZgKBEzkVJuRzPhEiSMfUyuRs4KqlMovuJ7yqh3br6ElWUIpNeM52cl
0/WsYzLpVU3k3THsrCNKDUaBWe0yDFNgQqSD6/P6TH3VMa5G9imQH0Z2yTgj961G
evPXsoLmtJwKt2U0Jdeg7veNmTzb1lmZ0Bvl0d3WbShv1hCNB5qyhuMsjo+BYgNx
/PA2fYj/Hebsc5r/1QIJovkRh5mKflIN5IBU4p8lDJIce/9EYBrdXPao966BALNo
47PUAkzs7qcC+Q0jqIAgoy1e462ingSL8oEVhdHss/2iqD7Ohx51neSn/+6W4B3Y
ylVEDq5yZBi+wGQUnpVTS/GY4C9E4Pev6za1g/O79Lv0l7fgFVcCY0CvpzbEHHM0
bxVNEulEDCtJuPPVkICrijMLs7W1BvH3zgQQqMXXbQsyHyfK5t+v7horm/dvjIzx
cwa42WcPdN6BctMY1MhituRrlz1L82byDnkOEyHGBn/wYWsv5wyp3mHfh45dE7c5
ObMWo6V7J54PwgBuzvsawNbm1DKcqOjDWa5gY/r3PhSb7z0HT9hQo0g/OaH0w0Aq
dn6Xb6jiY3xqzleccA7IVENMs8YZvhdNt790bvMhwK3wCr5U+07UAmHFlsbu97Rr
tcY8gc/icyRMFedEDw+HLp0HTPYXj0e1xs0TLn7PMiF7bf/KgJ5XufR8yxj02u7K
/7PBzT3tEkgPGwKvsZJETe6GAvPnYQ1oyxnpEAI1W7E0j88cR7ygp8EgJKz2OZ/D
bdiN7D63KQZJg0uJQDYjs64gseYHymF7N+RiSZb3ZVf+n2pQHD3qjGaGUa0KkEvN
s82h0lhZEd8suO/hM7cSCAhX7JAZKgEa/BI+iscaS5bSjVjVsqg8qKCl6Q+Rwhzz
HmlgD8MpoC77jBg7CrEOaPjBQB0Q8fkaauCH3+vJCiF/KM4FiGCDk+egV5/tHfra
qM/nwLW9yzBqqUv/9+geKFkXkZ0L+W9FCfXd4NHrGqT2IxpDnTGgNRFq023lShVv
pYocw9GvyGrT3vQE444sYbc0NZLsQTFUquFu7D0jEbJYKzLG/rwvwCOSjKnw2WJc
HICHrdn8PYeHdjoSd6N72wwdZbpXsd8Rj1U1vXBjdGdyFo+hibkl7Ntk/98tgoBU
HCw7CBPDCpPSgLru4PerAWgcirctJPyTg7ofiC5ImtGEjIsvp+MNe26r2XE6GBOD
XyoAGD7tThXaF9rvV+5jPEj02d6f+ZjRxprbSo7UFXwDXoXmX2I/YKvu5QQDKZI7
pqtVBBPEEJpH4Wlc3t9hL4DbEQQ3k2jbABxjmLqj2Bh3CmHVvOw/OU83/5hoq2PI
CmiETzIkXUfjxiinioXocvUmSKeZUsj9RbOHTAnqkT5xtx/JB6Wep4DKAnJeiIco
G2QuRHuKZACcl0sFcl/LTz5kToZuaY4PfOuEb+emt9WKQDBWwqzdqsQEjTeurPKX
5ea6rZPQsH1cDd8dQc8uid088pJaVNF2ngXfbUJ1R4r49PiHi5AEwhqF7+0wYMt0
QZiLG5PQb2Z9u2qoXUKAn5O7vrPWtSJoF3s9Ahoeh+EvWzKkrZXg+XkahM9yu2KH
Ld8HuECo7IgmWkRPROQ/IUpJInKVqcxh0xwN5WpbJNjRJ4wyBe+oiTSAGqtsEs4i
+eFgUOEpRXsfauntGqazpAYRcH8GDTa2lBROpGHGucMDTqhfANAG/iVtrMncwWBt
hrcqL8gW54sqRCyU1Ttx9x4ElEh3uptSl+VDSgBfZhEYXXiyMx4JBT6yh/L/nDEB
Y7jh8NhC7fb5up9xrqq4LYTv3eYDuIxI5d+5UeWu8upruFQWig6ZDawok2KObZnS
eVFFLMer0mogPhqD+WOhalVXArjZOTmYhSY1OpjsENcv7bjQITF4tZaEJloCmMaM
U7GAFtZ+nV5HJYwhBcYSty7NRinQjmxvFMwaMl4oByOgXGDstddLMboZKbW0dLxl
L9xI5cZuidA8V7Cc6Q/U1xpJkvJ89g1HqKAtFNT3ynXOm0LQbpT7wCc4GxkmWiwN
GCbm871Mrma+N/f3MxxVLypnaNnBrXotkEg+k8qWAikCKTZnA6AiBkwmkSh7sltq
9IItkNJe6YxfceFh+gGWp8i+pvjJ65s4ciplIKcIDiSNowCfQwT/sq8C4f90956o
tXOHBztvPIp1D3AB7R0iG4LwYk5B+DfUtP1sjWvcAUvxS3yetZxCqFmkkiIKGc5c
ZrDEcX37FkgC5M6PVdvzebgYpQYFySUzR71q2Z0uDSCZZyTSL5DGSgG86rLcopRj
n2BCAkP5/C7v76DPuGO7q7k/q0pRxqrUIBrOht5aqJZI2QcZeaE55wBh7mWVaSKM
sywQE7NBSjIlStpqL1BeS96WzLVmQJbSfAE3JlAtKfCvbg2mNPpe1PBWmZmIaOtT
JYC0tE6n/9TswHehV5Zh6X4uwxOp/vWL8YF7nv6/s4VrvCM+4lErQjxkR+4ZVNJM
+umaE4Xyx+pUfn5WgH3b2au46gqIhrTegmzwplq10UR55fmsQ4JYzspN68E6P3Gv
eTRONlBNkL8hGrJPHjUUPbZ96TsFf3yzkOOFhKOjdontVK0A/HOhELR1/uNj3ZXq
QREaUX8ykI/sWfaUUHCRMKiPpxgLiwIVjjxJdZtR83bTXZgp0K4f9qZtn7gQZjT7
mqsReSatDHPND9tydLKjpHO4BW/oonL93kqaL5rdXJ3OcOllIKbBnn3SETZEjpHe
qHRSM6Flno6V5x+aqAM7ELPO9lj8PE9c4Ffmf6G35bfNkm/LHLzQXPGB1lgzFNKa
LYNHfIWttTir6GasgE7Q5/9KN+0kOHGOXfrNmod7A2bY2ixDcPEJyu6J/HG5/Mex
kGs9nBCMgeHFKqQJUxlWxuAq54DXsziZ6RFTaSXu3DseAdZnJaINOhTzolns5mOG
2pMlAERl6uA83TWWUSl2y4dv3s0EM70A0b6mxlSWNdb8qw0Mr7MweHzx9z2Y01SD
FcgCvIFXTm964xj2vBjVQDqjfXC9Pbsrii4OnqsbGy9RvVNy/mO8xeRIyf19rLM9
eWeFt6NAHF0vSw2draGtMh1i3hYFlj3hiD4extWBC0V+j7yhiZtNcigtPl6QDant
VIIpizML2LmODQOtNsqiR0OVYACW6alb23rchOlvzY0GWCOiGHU8irysfsSeiLAj
dw4N9fRLh6/PUmEbYMBYaHJxI3gTMcm4G6QJOXdpBL0450sYUu28/YHMfgwymOp6
7kEjv1xazWMmq1cqbGmrGLsUcFMn98ykVrvlBocIxjZ4e0kMVpYygKyvnwn0Ak3K
p/jB7TXglELmsWTj9+fegXDyJIEuC1C0bS0A6VGB/l5lyygZG+d4fqBBkmmGlA8V
5xa3wULqfXPi4U5mraBUi4Ui2t7zHgofLItWfgpkcHGonRWO4R6U/1TxyhmwYM7d
40aIspaRO0MVJuFsfD+EC55b1nyTsXYEZHAsjgqAF13CJ9IRALnHpgfg/Yl5lfIF
jQlTZNzYWAhAvKfC0k5hhlDl7x0v4QLSsS8FBb7R585stOYN7zOPG6ydken1Ve5H
qVL+1+dUrEL5pCO+s1b6vNafedDVmCl3Ou/CqCapV87gXctr0MLMJI+ZJaUvD8Y5
UKAGShdLQZADnJADsSzgus35pw5ylNiHiqOlEpdurBH1XRoXHA5w8Ix/5amgM3Ty
f9doGbYPSD3t2Tb/0v1196/lGLIMBZzzgcNKHw0tUAgaBsvJrYAjTT1xzQgg0JYh
mV1sFDaCqgRgzT6nqYjOjDox8gD4FfXvzzPTDjO7IGYNKgpBU8yJFRNbVV0OiOnU
9qGGCyCCRmxcoTgYCWifWi6HSiPhP3MlVlh8MIm5qPt6SdbYG2uMCpJCRXxRWOOu
4Cw6Wj+JkOol2gWTMXl3yAa4+Xiao7Bo5BFFc1SdJQ1g2DBABvia+9tnevIJSYlY
wlpmnybygA+1hnxJNJ8It3EMLt/pMV+dv5kD8cC1Nt58tkLsGjLDt7FcRE8qiHIY
y8cIXNfd9euF8xu7kXTGmRdz2lBu5S7dyWzCpjj7aL5Ht7Wcgp8a0dkSvYreXPNU
52lfvsXrDfYWQb/uD+tCijObtrW0UA7nkRhYrdGqtuom5323v2u0koOUTSSzmMJm
2QJSoyCN8yqhzedO1cQLFFaTzMNmtyQptTdgqk1IStZj+jX4gGjMOyIPmtBA5x46
SXH/pEN4uX86baoOebKyTZD8PnE/a2R5OE08Xgp+smB+uM3ErJH/na2pgGVYNNec
dbVHJnwLcs+Iw3pCbC879jhvR2fX99ubSc2AhuRYHi33ldGjZZ7IA6X2SG8yxNlY
Fma8rsycGex6Hp21aA4shyniCESbOVy4Qeb5vA8nsRiNL7z0uBqj6avfolAQwtqp
dTYXMWVqK0IrJTr4cDU0C+KhGqegL2RdSt53B5/XufL7ASDh+t7K74r/Jd29zhNv
tP+ZdOsNwI3AnzcUYTU8gEtXJUdrjvUJwDf5YN6vPfY/2n74sIq3iHsyGr3559QS
UXDspwyjo7re3eYvOlglbBiUga/BGs8Mr+7WXhfn5l5/XP5By2AI3VrfL+mbsbHq
YFOnYlS+r1XMyvVXm0OQEcU7d6pJ0o/b21Xxy6YJvMLM+HRl3T3vfe7Grz7IphzA
+wcpwG4+l64SME4PiD7sxr3hyOltk2anof0YSs4NLi3F6LJd9HJnfGWzGWZfMfFX
EkMBLocsg6Uq71A8ItUUtJmjCE083hfp0ZZtxcCqLoqRTyly4heZXF5zAhfc2qiQ
x3ns9Sc9LaQQ56HgPS8C1+Lxb7gUvKkcUc8+8GnBOL9KqkC7M0XQcJrvrpL5zT7e
/KH2MziNcJGRACH5uCbNcNEktZZ3Z4SxBiWCQW1qzxYrOl2/RNQbpnvElqFSVBuM
VNVqIrsijF7723bpXZ00o6F0DvGtSYozT/+4dWh5CcdcWBuTWmEidP0QdSdh6tkO
YqAdhaYqNOHp1OQfyLbGmMsn1Ifj4RBt62C4+Zhq7YQ8gMXkBNYIDzXwo/IgADRf
e8MA9jQ9evNoAZCzEnu0tKycFnFdLK1bfPfMC6db1VsCuID2ODaOu3LEruOe3wwx
CgD/IYSDx+X6sQicJGS17KMgSu2Se7U2fPOEI9l7SSOz8PpXPFlQuHoHOXeZ+OMT
gnPecGBei9CMtRRYCcOMVeiiLWP+dEdTCYJZ40El+/EGHdrcgqZSXaRijxy++746
jIsSCcCU+tVrbP/m4cRJk1Jq2b6sFYkPpN0T7Pf+hEb7wAT9FSWbl/PfrIiZkrE9
pJVhfenvhhIkFwEwqIcaD1RD3UMiq1mMos7MXWkSQBN5d1Ch1xd/X35A2rlelLUB
VrUbyAx3pWhCUXbgah5NvdIxFI+iA0rpnulf+qiwW5kvJwZaIveZdk6AQh9QNRsI
gF3HIyZaGcfAXcsX0JiHoDc28zjQF5E/uFYL/NJkbBsjBPQ3OS3TXVIAuYdCtlKZ
Kliwivwgmdh7H3TgkU+Ky5WXBDxeuKFzym4A4abEF2pVllwHw8q54DHyomr4O+zQ
lGHHjAf8kQUfat5YKSobugb4fP0GaC7OikBSQF4vjynNO0kQn0KL883qiiLiOZKN
OU7hQp0P3QAn4zq08W8TjB2V4bPx6WNAh4lf1IM8ziXMJHMJIq/och+GG3m0U10N
SwaNXn9YtseM/IlCJrhSDfZDcQe9Kchl3drBreLB5KARBbOrYPYLiU/c7VcSBlR5
NS/Js4AuzlN1GlRA2OM5jfjyKqYD4W8RBBmItiLwU0NnOx6Fp2QctlKb2XW135aS
3f70J7i5ys+HtSw/ne6fibfuRhEboK1r1ABlSjELKIN4Vg1XGILlaRT9mTjWauI/
55DmXK0u/hw00rvuxYBIaryBgX9H1MDR1BSz4rydL8JgWg9JsvirPzBuAeDugIRK
gFNSkvW6tsCU/r6NY9gIbEEKKR0c6bdS6oSvcO6tBGUzv6of3RWNYdhdQbuTvotv
CPWjJe7aCfwJ8fPpAs4Bs53h+G/Zlzpb+gNLvnY3HQNcKuqhMwwKWMd2Q8cAsLxt
SlegRo4t23Hljn3kAbrn7JYlqxOoVcDPU7S9LfzQmf5lxOaEJJznB4CpaFkUuibX
4UEhPD9NtgnxJuJDuw5ycjWqz3de79R9TFGRUTwVq+E1+xqLooYSVyXgOW19u4In
DCDrGK9rALe8hbwPBqjcGZ4GGEeRWa8TA05euCJDICSu/d5wt1RBpl50xPsmVEIl
FK84XWuMLFjGopHRXOtz1Mu4uztmnuNBHBsq8UNGS9JTeBbYY3WtMXxbmi6C5prD
uYsPTVoWJ46Vco15kFgt1/17MlKam5efjIkxmC+Kgw2N2NJnG2tvR/no0OLD4la+
dmuHCMBeizKZGtlI1D8H/6XGchAiFFSU/TZfFFU9qbGdNKBL2lUx3qYzWO9QuyrR
KrKX4IunNRpZP1kKdY9CMsERjPMdEZhGUPUSAQRquCjPuowpxgez6grqYTmZtNFe
v4Wh1YmgSTCvuo4GMZ5TPSbtoJRlfcPOGmP+QGfHHrt9gKSLv8Tbg4Em1X+DCq3e
ZlpEaBpb6bEA9GOndOLpRiOInm5n6c3A7uuqJrdBHCAwc0cyt/xXRIg5RugIBZQb
DahJSNh3rUVW60Onos2AOEicK94NBRo1X8CeIMRYxtBFbO1YhKJXui4crBWEfaTe
zoZURKJ0Vc37DlDp0V7VJr1l57/uTp2dG2M9AC/QfuNtTZC3RqlmcPyn9OcY8RfV
ELpOicQK5mFv3vXZKVhzNpOSDxXImrx5+xJeeWuKQ4xTCGZZl4gi6xAIXZnfzfSZ
rZtEqUDjvjV4RDEK9oUEvk4zdwLTdn/DmjDfQ+RkH+llMad7xCnyRdkUoIRbydMM
MOx7/QQ4QQc5CLLp+Z2LkCw5uEagDnpnrApImYDEFcmF9xZQDyO9DaaLy1CrXOUJ
DumkqjNEHPz7r3oKK2Om4Ljz3Uo29gbm0PR6/lR/mNfjwqqH2BpslkL+QLCJvHy2
lSI4FFNumEBqUvngeXcCsT6cT0mB6kZfWCqQ+ampHHBhDAzkBdygsoGdTmJkfGpI
F/I5/7Nu+dywSj64tJoC1DW8xqFs7qyK5mPNslH2pW/rGK7OF7fzKX5794M+uq2B
q2ZEQD4b0zIFllIbuhKOWu9+qz+laR46O5uYaBlaIoC02aEomziXOfJn9f2FPImk
heHymG9BbZDAadZzvWMjFUgnUg9ImIhKQsnu9dO+nxID5clKeMa+IgXv2ubh+Bq7
HZdfMSZFiUMWgD2cmjqTVy2+JVnosW7XUlfRCiIiAhI0mcjxM6F2B/iL3Slqw2UT
i5WldnDXC8zCkGJVhYn64SDk4mVWOgLUYyts1FCAl11ejTYA4JVDBR/iC68/oeeX
DExLwVIGxzn7oF93NGKk5iU2qdCqrBBm5rIPR1snKcf4eCk67lqMyBEU+3nF50Uz
hwwThuidOHukQ2/n5G4lp87E9JdYjlvplgXmt8b1j5rHU4bMvYatjxkuHYK+jPdd
tGDxgoEkfroeilq02NoYH9wIjoUIf+CEtbwS/pUzsf2mW1x3n10ZnR/WoNNO2SeJ
n0nZR7GI16RCmuMXpnuBHOtI/NpYXYrwDlM9Zf88QuTIAHB2GcBq2tJGg3WeowWo
RkVFBsS3UhereiEFNJIj429AlFBFzz2pDvvUmJul1nAoies+VFV+vEYlPiHo7Ov7
r3j5Tu6wLY4NVf3oPmqYjaZPVUgqiNjC4ywusJB7GrIVgdjeMld2YqQ1Mp8TsdrT
+xiJk1hXJ+Y9BFHo7mpI2f3QxqqjWBDDZfXGat53mX+IpCjaVEh/ig0nxGLPqg+R
3N6Em/f9LjdirN9dRMrUtpgyH9rj9uIUBd+uj3znJukKvR54bFnxv/eTn/qHJ35i
WvljPJwR5B9QxYUDvp+n22iFeAX5MpFjn07u+m54sfrSXdMZi2xCo/HrJtMEf1Ye
RrOcGTCv+Y7xMosCt0NWRN0Te9iLXm8ARZUBbhg/522Pg9hso1+ynkWjlrFLou8d
qy/8uBsbOxQDbkv0F1PBJ7H/1/NVQUubiV4TybjZ/f/y/tCTwe3p537b8eKN+FZp
Wfwfy3Xh8FqHIay5LsFYY4IM8zfJXTkZfmtj0yjy3QlAFahSyi69lpJMRBqWnHZG
6c+a6P4xBODusEivNZZEI1OyMp6xlR+pOO+hDRkKaFkhzNlZemouPSCrOvc1ppfr
Oto8FMH4deFYeqld8xTJRa77bW5OmHw925DeJme86T22c+/TvPF+zfxmcmuLGuhm
eAc2PlvAkc2c/dBUp2ydkOQprHCCsnhaYVgWdZt42Fde1uSGzKV4KMhJImGAoaYB
nlMmmzfwP+zrPswxfxkVYyJMNHRYzdIwf2CZZ/UROP22wJaR5vTq53jh1u6mQvUC
xV9hUyB5eOtXUbT2d+EgadfRrWbaR7r1xF392M0IUdbMZJ2FPEeZWDVw9bkymRgN
HlOIy1SqWZEDsliG0soBWGj0W0i3eKuh+aTQbHr19k/R+RPHruesI84beeW0j1aT
7ZSvjsR+x5vTCQcn273se4gdyG5c7ECalwECHpP5O51tlxxy2Ypc9SFk4DtRueHj
iJNYdxqjFIz7xMKBCnjrNg7wTHtN24+Q2xa3M98MyBFL6JdQ6FNVTxbxGB3fBLWF
XApFV8UlHmqolmQ5+DV5ZaUVtCJMiacyNcx4gZ5HJgCuYROjRdAKOxMaHTGii085
uM6Prb36/INF2g3fXeYBrJxn26fiQlPpZ1QM3R4vcG6/r/eFhZksEQByG7M2c8ah
Xv3AZcJvVXkhP3tNMIxllT/8GJ4WhmmA/UEIK0wiPQJvs5f6gA8ccfgkgDuDMFJw
dTOtwnb6PLg5zxsxwIifz1whzDlBfU3ZkpxfAFF4wj0/p3itRuXcqk/ymO+ccR2j
12k94tawXgFqRAWRVz6cjh4WLAk/HRJACwwrWKiIWwwy2UXiSjCUO/HHfEE0VCxM
/I1xGhQgwFpBxZYaVQuwjmtF4pRDNXPIARiRiSSgByT+Xi/wZDFMHwX9i04YJS4h
IVndzyFGWda9waPefi7HRKuIQDwXVXmNtSH8lh3MnH0AQaFtVgWFK0AjS5lWmMDD
W9v+HZLygd3x39MnEbChV+CeyRZybd7mpYIlD9m9Fy3y6/J6wZiyGyRJye+7E+jk
uSCF/VnaqOhnjRRcLUjPjThDvfyXU5PcICp1/TVha46wtSvK57Fnfwp/oFhfF6bF
iQqgbpajc5fqueSlweDljV6tO0XpWMrz+ivB30utDGUs5RGCCbRHb6PBRmAwfTSv
Se8DwB1NzG1nYLjHN6pRz4efTl94FeF06ocOVgdJB4UMXPGXsFCgwFTbvF9Zu1NV
rE390ySYJmcR5q4792QGdHGIbkIg+/bouxVQ4TM4M6wdBUWL7TWah6g0jJuW/gCm
uaQck5IVxdcRRZZGulauj5TqmqloCPuG8iJgJUqE1hLYzrZsHb21yf//f7D1Qr6x
duQrkSTypJzt0MqZZsql6ZehEmOo5w0gtXWDlbrW1a/APxgdfw9Fm/JNvOq/VXSl
WGnYvYl/qpjKd5uBnfiu+hDYPMpLVhKOq9Y1cVpG3t6tHABTJ7DG2Ys8CmFSp2Q9
uDcHEa9ecuVig4xJh2Tj9t7wUTHW/EwJ1mbjx+NCPLsZ4LehFrk6lywIUnW/WC+v
3GFMQZaBSe4fGpK2oonaeya/20pVryQ7NdwmXEiEI9X/iZSEuEwh5JImT6KALnIH
RQNxfhH8Hbm7IWjNm7S7J/I98YD1PV7Qq6Ry/PoYqVrfgMgDzS0uMy0UWIKSFLMU
zcUjLhIQzkzbUaYL71nYRrQmVdvzC3hSbn8sh6DsTiEhmP3+L2WLDL3VlPb2B35k
bTU8wWBgfVa+iZToVE9xCpu6PrmgFVCAGZOoXsEsycBUQsymO+HFImgM99ArEwwi
d/BWBYxXoifsPdvDfqXviG7Fwm1qIwvMPKORRMxe9H5m/g/ihjUG2/kKb/haAVM4
StqwdudORFiE+yiBoZCTMyE2t007cH6e6cQiHQMD1P7OvT/ziItGd+Ue4nK9SvAs
HfmwT7c59/ZlLatJg7hgKgcwKz5pdNuK1pQyD1rdEtrBORDcbJDCnOlyUQkC9xox
AvtND5ooEUSkh3NF7y41jTACqKSvrSq2NT9ovDnb1m+ZP2NigLp79KnCMeO9tFeU
BJQHik37PCZmlZZom4kA1rE2uZs/8ETnUIFk6K0UsdrTMXOj67OZCeZNT/mljDNv
9iKx50jsesm3Gg4hpcbfl2A48uYh5EPkbOnwRxU+apZ0jMVXTtVJlr6cx6cUy1Ge
so2NJPLK5lDSy4vWbX73NIZyiXz+lPiDikwX/0bVWQ+IEejvfM7hNxO92dCr+2z4
lDMBqmbu/JFc5Obhn68lZ3lI36VHjTlfpVgZUndwZefvNVz58y0VhmhHLEPergf/
HevrzdmqngHig13FAW6YKx7l/YOxF/2kaoj48I1YDGPYMte+21L9OHn8Ulc5fNhL
SrFPFanmxMvLXs0wbla818yeW5ZIrjWjkjlalqfxR/6E57gNPLQqCM0ojCNT5Nvj
EuBqX1wXYcpk/zWm9IddGSoo0ruVldfmIGC1Vvjs8zCWsX4lBhHBTpeCsKlSJi4h
7TQ3zLEW1xo9SNtbh0uqScqqmXtwPo1V6fw2Bc6Fqq848dXCXzq1KZ+3fJCXHHuw
eSGNsA/Jd9fjGGgg9Kd4QmDbAf+cyhQWghbzIkf60MSidC32QADTDDTrtpBXPEeg
Ulfshp8bK2LTyocw1fgiK4AlUQMIC6zxx6/XOFMS43wz7lubLe7Gu2UWkqCqHn8L
hqJImybfLQFKDPpFE5A86Zz1p2Y8H+Dw+zJKKQtHIRJ487VruYko1o5IOmTMC4I7
yAFngSFlRkKl5x2lJWJsGaZ5Yu9gxbKXAu6UfMrTsyAAspPMEip5sxEseTimRPjZ
GwSAz8LpehqHw94MkhDKWF7XehvrmhIk356MfoBNAjIc4obsx1jPxb12hRnHaEDD
g93qSzhrSWc/vvAZE0S34VN+46UPQVGUsDPc5SxjgpkAx4rqj2Te+FNwfA3lMJxg
Lt9gFMGRrM9EX1qBmfDd5sMrVSJymTOLwrBPf/HneL3bOpUSv52aTbRm/L+9TKJR
MCOplkNtzxUHn21ClNXw31nKBnfFjlEWWlu/T2f7UIBi8idVCTD/QuA0OswyI0H0
/FIiYRsiY3ztBk9m9yanVnrxrqfrQW2nt5vKF8w49ZykMZEM8189KnOZBr2IgBRA
ptxASgp+xxngD+8V0DgL9I7VmoC2wDeBpzDdfVJTzqd/qamqJQ2i9dGnjQ4I6ILq
tT6rkzvdTze7AdfwOG+aj9WM0B+rHRPQc/nVhUT2t5KC4W75yZeH5hG07vK8EH7C
r+qBkdHvYCNMLO210UC88VQP6IxnvS26Y4ytiiSsLZYnBizq9wYmC5F2RO4jK+Fu
ZmbybQ4Yb1K7pUtkvpZeuhV3MzJQNYjtPXIj5DTojQ2wkBEZi7zFD3ShrASjqcCz
tFXGygbW8eUeEOwrdKAOKaIvfiTmYnJTYME4/0D1u2IASRijrApH6kjkuU2l5hD2
LdjlDXG2Rooq5gkcXOXRKYUS3P76jpTng7UsG6eCVch4IX9pUdhKu3eHCp/74L2Z
CKpJggM6EdA0R/WXPkXVkIC/hyudwYcZjMlYH9ai2/IrdcQikL+fQrK9RjLn39vG
VhomA1jMt/HnbE2M+kVf72QviwTmf0mmq4pAv4u5DmfarL1aT/oXCLj1IjLJwArU
9KcLWTd1vfWIZFylCnNK59RMv+akhX8WjWyHdSyG4OHONqFGVVT5KEjGxH2iB0fP
byzR5sVrrR8EcIg8ZzXB2giJqGZ0+4vsavX8tJ1HDw19WDwsOM/4NDh/33Neez0C
TT+CrxteSl54+Fc88m9qjd1LLlnBT6TVQ1XkZzbJ9HsLiOmk99T0Y9JQnVdySLPR
iH5+bkTL2SGRwLZuUKZL47tsDz1fgboWSdadLyymQCQaHx2CXGG1IaI1rF8BQPel
fI8saHDmesxu+GgSLhOuxkzL6qrxkFP3cMM8zo6Q8vhTA1vg76YM6Tj7BnL/QcK/
/7YcDuhuXyQ0xdfSo0NQqwctWxHmGXMK9gC6qOwO1TOeL2TJevPL7xmM0HPxn+17
8IyaZLr9M9SswBOzNFAbylN2g8kRfRct2uPhhnRfh1eh9hEFDk83CMjVIflAWrkC
05uXLRv6/XJNpPqhY/LFpwKiVCSp00eXqy4CdZ03j1WcQXmEmkMIEnKtaHIvVJSX
kcSIAmCcL2Ng0NhwtDFV5lpFHwLWwle/yKhIBCdTz/AfE2Al5te+5QkKEpy8W+Pm
IxB8OEoVdhGZDFmO2u0ogPFZpJ1ZKerF8lA8vgdw0WlQ7Ni8m2NzdbsZPQ8nhB8d
LJvL+ndir9fNdkW+9Mu8Du5Ac6sJs3dYpK8Ql5dpjWjvKHt99dbJl138P3pXq2Y8
Nudaabup3io26SLjBDygMw5U526oYPrsDSTO0WukykNjR7d+WZWFjhAV2QkoEdLO
TjZjq0ddnQWyDnEC1DvFKkSWHl3fCfmMN/6KA6Wq4c57DBQRyO4Lz4nQGeZWGBt/
M7I4UP19Lqw0d+2UnLC4ixp5kwmztsMDIw/2wwFIGPMSxqCrAVu6wgao03xFUMqs
hLJ0+DT4MTm7Mqe8qhbiVAl1lG3K8Xn4vrxu6hdtwb4HIptTvhRPBmEuyoZ5ww3A
cj2nMmr/+jBBTKv6NNQmkKzaU3lNZ5TU/DQSHQghO+0Yhqj0yQgSmtgUnxghRbYj
mg+HzQI4z513ZMDEaHTA+2XpWDadSC9NJgBznECfTTBF8h+vJLnsyst1X+UMrOdo
UzOsjVO5Tl5sm5CDYb4+0Kxwplet83EoaUBUxRXtoaHBnAJ8j+A45HmrWPh3wZhr
wIclhM0Y/RgOuv+F1b63G8ruRy3MhKrTug1iPrNwN7CouObLpktdNTSXnP01DArC
gvVT2elHWrx5hL/AP25fpOKvdHpWFhb6rJGJmYB9qV6ud4wLwsz50D/0zSW32knQ
g18bdqIGuVJ9CymtRRWxe7fy9OiEO4F22RhxfhqnOLiUQe0OImZzlJhSBQr7nCnv
Uz2D+eOUZy7MklbOeiMx+sw7st5uAuZlGvgcTRyaSXt8o030YhIJmBF07DBSCKHy
+IoHmD25+3Bz3L/hahoppAzECECsuAY449OwcLJsPVG9TSNVuAIVXq3G6dOLasme
/2mLHYx69HKjpqP9JvwpJrClcy7pKX6vRQ5JEewx8Rm3w8cJv9mVRJpNl04tX8qe
EVap/+mYkRFTgy24CNdkkQvKS055brGl8mWb3prT74z0y2+x2ULhXvHXJB5DerAJ
1bJKzEwrHuPd1kd4nV2nrTrJqT+LunXGtkqdecEMN/11NgnI9liuhoujvsn2Cd6S
ldvoq+VwwI383+PdlxpmC/riAfqBpj5xdiIOWZQhpOewNKCIYXSo2SnlRFcGTTRU
QrvSyLIcqJTpDOX/n9Io7OnurzPC6CYzUaFcczeWjkkpsEVyGGDrd3dwTM3qJgj6
EVL8zY2/8XXF39kjIPSZmen2KUYVD5WNcqNH0+b+PO1uGXr5l74a1nowTtIU8ubH
ZG26L1Y+tgvJULK8hLRvj2c3t56+r695EA6/00NQFCa0I28oX6CkzljA9rJylOT7
ATTj0qaJSTk9jfVi7ik5/q8LdicmPyTBYjCGBzv3B6BmTUWhvtVgqGxZkr8aFdQR
JH3C2WNjYtfk2GeUS++iPgC1o28UmAxNfMGIfeEHe94ik9cesGxNweDZAwZ6cg1u
gOqB9jQh9Gs3mlTqqEyPpf/ldIou2DZBw6wX7OAWePuOhrxwBoGV4yFVre4Yypha
3qJbFiV1qDNLMZaf8H+N3/ZG3lMienwaU5UXBqFa//pg+6pkCe4ZT8oAs3U/pwV0
qqZRGnoXL8NTCinpL1Jmcwim7Qg2isyVA7OY3Ykjh2/1+1B2vXOYMismGxkcV3Yx
tqEDj/68aWHbjpde+xpWVZcqIhx2LM0yRw3I+tPOiPZwrSHUrRNNK8pBl+FV6BKs
a1z11KGcubRm/X75xTLifTvScot/HsOIuYp0snvkKW1temI0RgNaQESPTtazSJw3
PSLE0cvjZhjOh6vt2EUfo8JhDxWvRZkqVIWVXVmbOOoxY40K32RSAmLHJkW3WuBR
fyXP49d0dJ/8+jZeTrDwf0NG6kN7jm0vLvRyF3pc96g6/g3D6YzM49Tkxg27/vNY
wZcRYwMcSXwDDNWkLCCQ+lCuZVMzQaNW1TDuKcVhUCsIZIS2FhtC4qms/VGr5lYz
vxhtqt/LjLImin/4VY7m8cdsAS5yC6g5LANPVDAZ7hKr7P3kh0fknM2MlE1KtoEp
bXjGOdEn2+y4Ff+9VWxJ/vIBrgCYIlSd209kVn9lGrFEf5EkAoY+vuQBfCiOebep
9MyuzbovcXwC5ly+eaSPBpogZ5zCQVz9yyVtGI+yAGVgm8v96AeJcN+8lNcDfH6X
EvUBkVZ+IJNvIki6ECR80mJFHMm7dI4a5DlwIIOGAYcdRdC2PzRAmEVlgu117Cag
sBGaGsuPpEaE3x+Wh2fkAlbRCwEE59OmSB+vHDY9fBZF3e/hrSOU6qTbw8dpqPV3
V48IQb2KKnk4jmWfOvfcsSwNArxuabLHa1r3PQHXBweJMLDIPR2BVdqdSxlmXWAh
K8FRGbc3K6IqUtSckE/ChnhWY1n2fd5RDIurvFmU4MWzB2le0zagQqEsgE8wH9dM
Y7rg+/poxKhZvBi5MaUPAHrN2poEsOaGVzsxBrSlPZ58vR1qzBvL+MgAngJTbnLG
I4e3QXGXqm29iEpivwGeIUY+3hUnDxJV5Z3TsfF2JTV5T/0yHEekljPIMfn0gZAB
hYA/3Y36LO3m88hGZxhK2CJVUJ2JBgLkpo55HfyWx1rEJvWrcEjLwnyQl5pChkuy
3teyUs8KbkSqT5XArI65vafZ/DLnJKHuw1x0WlQ4JgE9E9pd+VLNxx6io1udmnyG
vhoo0SM0yOMjsia+iZGrI9n6yAQpJeLLBJ8DH9gUQcSgU0j11I7cQ17uVsfDzoxZ
HQ1BsFmZJcN/D6iOpOW2XHWm06Hrp0gRfMt25g/Gt+eeINGOfa4f2f9JKXzClizm
rkDQTMkYYP510zhzUCKLC2an0ZV+yLktYnGaSZglzldaAgisaviT2CvQyWl4saFi
PQ8O3/tEjjMU3Er1eNCFUqXIT61EvdooJLI28Mj6Or9VkrR7g6NfBH9Mmqm6BLc3
ahedivebedrg8PJBlOsKnbAT6RMowtobO5HZ8mb6PJG8FhMUArzH6e611f5TkYYz
eTbyYmXvHQOfuhpOVpsayj/DUMEMQgsQ04Y8yvKv0k1Q4dKSV4g7Rbciu9Hc3qAW
Ma/MKek7IRDTH2GorT8bLCk2t8LEro6NFcWbkTOvPACXbgWrt1YAPj0k6KDQubpq
D5sbdF+njK4lph9v2De+5gbP6C5I0+/ERQ8g/JfXtQcWh2CaxgjG8OT1VUpXNGYp
ExwXofafdCpvFsQDYOMjK+dWvOCWVD/aL3WkLc6QheZbGDNhGWf6D2m0sa68eCZM
YRkkrJUEI1Q2jwIu1FfgEFc+6DJRkIAypUu3llwnl7/P8iGfCDS61CtkfRkeqbu9
M18MQ7EvotA+3aqXocffakoQZj7ClXFfZkemYhWyn/YN3qbgQ8U7+FveuOgwQYqu
zh7ij1DBCm26aGaulROz+csCbK8+Qf3DQ8bEBAeO1p3AFD7dmMxAzinhUdmUtcEO
P9BC+NR4FpVSGPcKZSRIt91SHkxccWyjU4NYqMC7LNRh9NvqqpQzBhjRopbMgX3+
GTviBWKw+S2gXtrTbl+H4B+U/Bx6mhw4CL7A5Iy1WV8l8WRrjw+D23bZKVJkSpNw
O00J9qJZzswqeTkt3VoPmnXgJhEI27ioLxv88CCgUzANW/wFMU9o5knPXnwYT5rB
eUiY/eKiwWpbwQ7Joigu/IVfTCS7/EERqIKGVrcUpncfVbc6rA//XdK3u4cUWIbW
Dc/RADilLFq+baVTn8yxSf8OkZjHy0MdCATV5PyEKJKiNohP8TW3POyPCsOnpvMM
4Rs+iMHP3ksZ5Hs8XcT3oJDt8AVmvwFreh2xQsqs5jq8AcUQPPk9ma8sL7T/BpDt
6j1O+81HYfRUHkDR1uv/rOcl+7iwh1kF8yINRYtZCbs4GDS1zdpoBgLH8RfPvDxR
FMfrusRsHMOCrNcl527TwuWwUG/DwiupSOzjwI9wc7rWspWNvPU4h42XGy8Py2/U
G11rJAVAXIryFOsLi1nnMb2iNQUcWyktIko9sDLvvXlGMu8UvSZgKk7THXP8KeaQ
Lxhw/mg5n2nKHNHuvg9QbCP4NuKaFBPGwBDK8sqHQO+bXZipk6xcw3IgLppzp1F2
b7ncS0JUE2hynQobH+qA+BTkEHGReUxC4wzSl86aYb1mMh2D+EP/NtsbH06kKmGz
d5PXDtCVUQ+5H4V7Mgwo2/A3wsLxx8tq8er7Sr16OBKp1mTYMUMBlJYcwn1eymWA
KBHg2X8aejdKhbvrlw1RbtObWO5KI4nP6dMCVGtPuGSaxkLEwqtJN6VQh4+UplHf
BjJ545PDKvLz4r598p+6CMAyhOjn46tiVQ/qu3d8L8nXX9CJSK3+798PdcmcPvuO
P1jtU9OG34Vo1V3w5iFnA45YO/7SdTmnmgSmQHEx9820ofyksDNpXvdxr98/ryfM
5vSi1JuJbTNe6oQt7aYt+27G8YJu7XjMS8xkSE2PWF2Uo0mAnXuNvL5T7UBuxj8K
3W8NKiexgLJdjz8MJ0eIT/MoLc+32RMcPuG+fcG7tuAvZYEZmrd8c1rH61Cy8gIj
mwpne+AyQWCOOnAQ1DrLWZ+Tn826ErUq0DPF38yPpruJ/DkznI4ZStgkxLtSE8af
UwSpZyRxn8e3SLxGIF+dTA6qLQ2vemKcdABeyEhi5k773nZF5+HRDT+KYKMeQn7G
NKc1/mL5c2qIafPRXuvp/nG3LJSx4cDYux8ceZdOpW5VAc2zPj2daFmzQxAwswL8
yninq5SVGi45+ZaHJgsSj8GIpccuXrKgthiOO2gxFOPEAVHrVASf0B2CBjzdZ5Lz
+vHDMeQL8qaH8vkQj8TbMW84oLhN40qJcpp7f9CVl0hpBCMiyCLpJWNOnJM0kiWI
YhsXEfn/7UBfi85JcoOgt7UZCKGfzNv+8KV1pcTo5AFq356xbICaeGAb7afa9c61
8gSHsWN/qsFZRCcbTSKB1je8ORkT1vG2znhnYzwa2JiGpE0Z5BPpzJZqKo56NSXY
+/MRkZP0Slgbj5fzV+6DCBBzO9FMI2iK8wBrwbGzg97xpNocFIjIFQSnt1E5KsAc
35AFR7ixc5cDQiYVgEnt0dBCj/yseNwvTN2PLkJnddRAt/PO7b8c8OGAzB2SGpYM
mMeEVjlAddQwKuSRb1CEUb9S2lfzuvGHM14pCArEvIqa2aBDHvaSHTsiuyWM2JH/
UqvMkiDYbnfoNmqIAvxqCaUXlnCMFoBiyLgXNArJpnlGMo1l5uxj+n98PaER6UgB
BSqcwDJ+5zF/fQTCYaZkvyc77EZ1+RCuZgBTu85blUHLlF/Wci0BWDfHY9Vd8x8B
lPRMU5ljq5b7NJQLRwCxmGYrksN628/0WHqSTMyGfdjhObyVqTyGB0dQ7keE4Qq3
pn1ga/1F6vkucvGM9hgvAVjLIIICtdo/DjJ+Z6rA4fwRQSun4fSzmhq9MMyfXJgf
NGPnhvc8ust3AH1La+uSbJtoGc9i/NBuosikTukgfpcCgo+Ucf8RY/RLDQ0LtpT2
GypAs9GFHIqLMH406TbGz03Cpzwy0OugB39jNjiVP25IILYIWxqwrRvbJxptnLPd
lWnbsLNQoXovq+1wKCRy2nhNqslold0pqxUNfD5yEivKDZL4wgYdrs/HwElneV3P
hiRhItp/vsdnNqibw+agpKwlTOO6j44QzQUPlDGqsejYrC/4TSnzYYYg3o/P+ZQO
rwseIiNnicsfxZ0JCd/aBPE7WuIo0i5c/r/Cb1sPXht7LShVVzZuAYmsCTYiocLv
Iosx0QEbAsVAbJAyEgYDIt87Ewh1J3Hj7LylIHUFK1NSir5TMiJ9DJctW/eakEWO
tDr37nWCJY64bf9VuIhWKHEWO/WMxOk3bW8h3V6THcXGlBa/gg3fDOl4GVa4GLpH
Axhn8sd3G8US5hmodWMZLKoB5g17nJz2wafuC6BVT+ehfozZvps1FHpbkFvXTSk7
McEJ2ra+H6EQatYFqayw+LjwRoTGY8lHU9wro5N5jaBH3p3qMCqzoT67Eh9DRx65
uCQ9MLA416LL2QH+5DnlJmtFCy8StKoBXon9RzVbVLMg81lc2WMJlMRfYF1q9n+C
R60HN2Gd3qRlJyQzNPohT5szBRaduHclqdvaKk6Q/rgN1c6jZiM76EmSer98dEmB
Qrjw9ktJ+LY7NkA88pF8R1SjbIjmorhjkceCXCC7sW96Qzjd4vYaLnhQLBgtvzYc
t/GwtOTbt4OETEeehdwJBOMrIxZkmUtCK2NSuJcggj9jHFdnZfnIOiXRBfi5SqyV
0RIMIyG/FAZcNEOaiXLnNYfFTNj5+cjHc8qzYblZwBpYxTNn5V3e6Xf3qIfKUFti
cJpY9TOgDkfiJU9mmCRY+rDPzvHb/xjjjbXXZMJicWu0ArW72CfMawxTQ93yt8QV
7JGvUs6xG56Th9EmDF/zHCwZlFMMYMYWJTpoqh6gAT2v4h5+Rn8EkVn7pOtxmsqN
qDc/oMC2fXChAULqWDzDJiCiXLF6qIGpXAPoYLanZq4pI4B/VD32rmcfEePDogdI
4MbGjaZeQ4P1aowJa5xtfMAt2/boR+zD+YMyjBfq6hgjfB3KLGwKCMHuWLKXW6Cs
HyhCRalfmHTysd1ppHFU1SF3bdryrVOOrzAXSL15B144fwRMY6ogzrLFt22ZhO5C
exdJzKs2p3iu6FBFKT4cTV5a5j2i5JJ07WhHKErminE32mQL/ORgOaoFvf2edSCB
2k2SHpC4ta1331PFMCeNK2A70lxLtWhAffS47oTkNxGghZ5OoOTjUg7TouBFsgq7
hKhKnNoJR9TGtH7E/xeK78T01P6c1y+BJIAY7LcLXmmMfS/13NURuv2x+uDGRfL4
H6Snx0KJBHUfcsCuzs1i6ugd8H9VqtJRrFrq9JtkxXEPH99SUTXNt9dLZjnOUOH+
YRCvcSm9TAgWTJvamI56Nyg/1l4yhBnj2x+wHHptsV/euSpIRJgqGuZIrN8wJLMn
fP3IQXQtC4QGwUrS3LOwterqYmdZzvLGv0k9uJYpk3qVJ+evr1ObyJoGFDNhtW6J
jXFebfxFKjdEPa2xzvPj/Sme+sSX1+yeTi6+QVhSt2swyVOq1dkMlQ+JwfhZBKVV
ugwjxymvgxquQswUetziPQEBeeKJsgh0kc0o6T3bDkRT2dwyG5XgAMpelkJtZquu
ZSlLM68NoLQC02p79NjKODXa7ZrqdVb1QRrqWAOBGK+oLqyg4LxXxUBvlGnSVHax
a7+ZNqzzyv8rbb4iITRrePxko/VH0Ac2SmgcyY6rp56alGIhM229l6ShhpNrxUtZ
5jJf4mdTkuR5wsnCNWB59gYNKHdiszRD0CCR5N6KsjObggP3cbE/4x1kGH8OhyeI
oLP9k1R+VGRpuX+CaC8lfez4COGsHHYaTsAL4SeOmegjO4ddpCc4CjJHBiSeVl7M
d1OwQi/tyMp5jEQKOpuBmn3yL4CPSCHauaNfhvh8l8KD1kbdUZCKOeOl9sK+1CFO
HTyxyZV8S0oEuIUR8UIvD1JjW58dOK+pti+/TSqMFFIZpKXeiFnLSBFyz48s8Lwy
TCPkL6auqODDwxrStqPxEMXr4W6oSftRPZ5qx24UWCk68uXe2iA/SJLGqBMtvm7v
zakmCnaOOP4/CrwvYGBNHp+J9v6s7ZpE2w4aTHCrRAqsLPM26aOzWj676rACkJ1i
GfLYKrJhFtH6F7WuPl7j+3ME2dhRxHM+IxlXgJB/YCadZ306AhU1iDFLtV7Cvru9
aQfDMjIDJNbU6gHsbSMVib9SO5R4lgUWnOPVXW7pOtu+QAUCLt97Xp8FTF7nmJLK
38eCVFM1y+kfyLbRbXBgOIW42k933gRUtuGE10VMaiSf4EPuK8r3g/2s7zVHzrsq
BP6uCLn4b8aU95qvwTccqYFfZ3hc0e3usYlrxcah/rEwIJpWA5dwR6mUzu3QzaKA
Pxs1M03yCy2Qo1ySJddVHFJDt8e0H3WajT4COzbJYnUYj277JPgAp1MaNOq0Rz9/
0KzGJK8jk7oN6AOS794BzfDNXXNGZ/DodlVCeiZZsb/7Y7xHlFlwkBVT2nlf+ajS
ikynXwgI9sA+K4joq/Ur17gnQ69AHYvgxbHj6MhNthNI1jStiILbBzMnKdz9pigY
G4Rxnr0MRHlG4VxPQ1DFw/4wpfjARkTNOF9sy+vWeVOnaCL+0qO5AV4I6jKHZKE7
+nNjS2aOSoqaf7oKbCHBNE18mvZG6QYmioPUzIDZI+peAOnSxz+nzGgd5Fy1HNa+
kzVH93qdWIZsNcWEDTaCxpAEavZWwO5rVkQJ68UBsFvK0u9mjnO2A5ifyrOWZvPW
CFitPU1BnwXyLPEC+rlXr80rtorVSLJgpE5wBrWBt3mMTw2Z2Y3bTmmNxwnYS0zY
c3BHok5+Imsd5zCSh5q2s4qEa/KR2cdBOXDeASaxEQl4+/vdhyWsetj2okvHiu0q
LucTsLw8w/tNGZG0XubbBBf679nIcS9e4VaE34StdJIf3EWSbDDJ2Q2/1+Szvgu6
LzIFmzlV49sTXpWr8TP5JN879XB4o9R0TYfTB0xnyaJyeNuot3HWAO5nSQ0yAzzP
ZX+dBWRHCOGEG/AFDEQBcTwF5AbuJs1jK42HBXwPlp287d7b6PblSM7pfh4/te7o
5RHPChXNMi9j29bDGdbUukHRXJO+7g3DP/MEE81OayRXzSpmRNTv/ACBsyD5F6e+
HNxx+XQgqQdRgfWSqFK7pOSTrR/8r3+thMdqQSKiferFzbdaxX6AyljMvyVWoF+g
ZvxjnZQiwhLAeeH+zODeQ7JFtlTDNxvO3n09OhDZkYm6VpI0+xkHLyYVN7RhsD+6
lxoRatOSvHHgOy3W/5NQgJ792lXAR4C1XOLSrKWouJ2Z2tbWd5zyvNkCJoFz5dAq
g1OiSN3/C3Ghw2L+y8/+IDLCXTZT1c30ZqaLZ2JTl0SFUThjhx6vKJfpM56aTjFP
aqU0z1SZdXmpyvrNXyW3fHQ6NlEIpwBvXCcSMdXOjRYI6oGYTBQoakiz8MIXAOgF
SsSv6l/feOgFMmYXjHPpbQzIgGK7fOdBZOhUq3wuL2zyqbUpS75xCAI07as2NBtG
9gtYpS/poIC/faF+x7eebfsP9C85tTrk4t+Au2e2GbWw3BHBCO51/8O9A5P/G0Nd
2z3PzMnI9S6B94WK/4i+XiE06kRa8WGCgZevFwnpypt5G8FOWdx4a8ReEGvYtz8T
hpXkyCJZDOsxM+Kfu1TBP5raBEwoIKekY9f2+Kp5VFtRtH+/+uKj62gfTfBl87GP
cD3iAvHzNfM3ksWGVbl9szD38AXvexVL/+pXG66FHbvh3WOS85oStvfYceRxzU7K
VQ1qvk+JIrsKQfSsQaMwh8lxWlPtpCPAjrp3DVGSRVq/c2V7Wn+cbMrJG3JapclC
6pC2k7DOCAgVoJSNMPfbbps4bLZp6hFJ0gN2i92cIpI8ep+FfuvzsD+usHzlDvhQ
FwlvYJ75IBDBrdocvSwY5U5Oq8A7jr5GrGeoC1SGORbDVOG5Muv8vAs/Di7vmaXe
3V1DeReCH7nO7JbVcH2+9tyAJWeN8yvnD/6QmMOwqZ4jvW4x/Pz4lzUIug56KCgt
3yPt/VTBRNYfwUlgk+MdxU65f1NTtSrGhAlOuXV2I1oeInRASPhkUx+GH9AuHXIz
JDmDaK0iG6kD1BQ4B0MKirM3cajIWCQJprrGh5TJs4ALwJUVlz66mNLTulUI1ByU
O9Boi+rY3CcAWc7h4r1FsftPBg6eba41J83u1JOJ14xiIlWZj7bLqt9mQyc55A2O
7thAN1X/PVcu6a8ciGSsecoJq8hFFGFZTcFjMq94ZQ9sK8MzisR3e8tkadUWtebn
H1u65BPAfoi0fiSAN3Cga+/iCg5mrL/OmUL9rt+a3trDGBiRcuF1z85zFI9saDqg
yetLB6OwHdV9ypDS11fpE6XjF+ScRSY6vUXGeZNMc1aL8PfLZZt5er5G00w8ee+h
t06TsAuGtiIBzmaxUacrPoMfU++zyr3TQE+VXzh8dva/rXqicFjkpPg5WINQq/5n
jRbSOUsILPS9Zy/E4sOinw/EGGyG9tb486aAfzb27tyUOEXzqqPrvBARmvbJSEUZ
7K0iIXzPnSSyoHFYdwqnZsXj0AOoZMHVOHAHcLFfAC/WxUGu2sLQv5jit1Nqp2ba
lg8MP0kRyKTJ/ATbXCeWfobx74uWJ72wvohcUNVYga7bJO0pSIX9N+ZSAdXF86PC
teWAvQTIdPkIp1LJCgGv6Uf+hR2j/nQr1z8g9q1WLZa1HHsNaxK8fxNHkADLM9aY
/Bg72BKssrKig+m6oHWhbuZdJnP9BKr3fwIbqyDxfNi4/woksKYOGT7hFf2sYygg
HFWx/mnmsOc8FZfphPVXOB5mz1VpnF3JsWIvAPvoBhaI4N15UCTS3b94VauKlzgO
qG34O9yzIa5yWtJdz7l0efljSz/XqMvFRUnJgUzEpPwNQJJBqql/UADAZwfcggzj
6ypI7nCnb5dnzXbz+T4emiF1mNqpXAluz92hyQVbFGWT16H11kKLYXJC9FtkUtvT
tcM3DRw0XAMz0jBqlCzhSRVBE2FMz7a2E3yJOArbIusUyj5Vn/tzJlmeZ7+a4I7K
jIMVBRFQjuZZmWPgn1zcjTaqR1FAkwVSZIFjypaHnX8u1iUfJ8eJMKB9kV5duRMl
zBqAImwQiZ43+Uo1LlRzTG3IdL6dWZDDZ53A215HkWEEbe/QrumNW5h/+pRC/ifc
SPy1yeMJhM1h5ZCn+XG9I9n2f09UEULEZTa9fxSJxMiKKwbnCVQCOez+qSDP/4wy
WdIbG95fRjuJ0Mewuw5rccEhTeyWtGp4+vLL17dsG/L/w+xldJpcBFsN15vh8EqW
OdE/AWTVtvxbV9YdFruckBSrOnC2yOa48gmzPoNJXBWH1gCpaKP+IUzZGnN1kEyr
EABtJa1DqX+Hhqamy/SULMh2NvDr0aegWJK5QejCwg/wp/lsI+x+V9WxcqfE6AxU
hF6lZTCyG2N79jwLHl4sHzpAC8yrky5C1DVxzrVI8BuxA29yv5SCh7A3j/ODei5L
zbYX+9rp4IG0n4VYoTHEBXNXLLxUOmHBZo2flUKK6DMttC+gzOBYRwf/5pikroOa
bvQt7hDNMZCyvNJ2zhy/jy20p0ncexjVOM2XLPKgdg/XyqfR4RyxgnL+17jYGqkL
Ur0ZqBlyHu2P1klyzecHCirV0FLFJXORsrTaXuPsZdPr4zAJowJnbxeZrTgR1RuR
j1ZZ+PnXz/6e7LyzsMBwMRnxTXkLjHyr7sQsbSAcDvKlerdTx2dOwXqwno5YB+To
UZgDtd+EAQj7s4L18Q7Al7vAZkaQB6LtMI3sgEKdOUf1tsRsw2OAzKFkmKbBv3xH
VHYUmYwwufiy8+mMomTsfWkw0ShmidoDNn93kIkk7ksOi7z5SU5wWjoRdLzxiKpz
OJEdMompGJ+9VmzITaM91kEP/18Go/hGWsrEkQh4RbsWrN/jiQ/HD7HN1n8lSuUN
ZcQL3bgQQZpmz6zrz1+z5rA3r8Azn15bTAfzSA2MBE7fEWlvczC+bMJ7APuYoOnO
4yIPkCG8Ja36TRgWUK5v8ZoZ/msdd8Vkln7ChIt6Hu8MVkffvxkbV3R2kQkFemfk
iM4QOWw/VKcjmLXFpdo7Q47Pl8KMNFxkzlAM943vLcrh0123N7ZvjX9EV09s5pJR
jkWx6sN0nETlAb3moxZd2CCWXe/9jSGsLQi/I9AzFeuQ2mNB/rAcCTptl8uS7Z4d
6uUWgQIV0POmokjv0E73z0JazKvNoP591xfPUEoviRO+tFLJH1kNtkNiVTfMAhzZ
IYkjxtKoMRx/tV4AcM84OltxLQ74/4kKomwZYHjyqBerwsIMG6KIIZwHwaEMM2F3
hI+Hf3cQfHEYxoLOxCDx9T2uClD9kPFWs/yDZmvtlTbailj0vTdoRmE+2sliaEt3
+cykWiGZHqZQX18/0Li2efERKEDNCV0NopbHEkFIYXrhXSQJilIt1M+/1wh8XglQ
L2y35oVZX1Bpsrk4ssqHrhWJKwV8jxuMnfks2lm51src+gYl4eSPi4M1duQ2fZt9
l8cO38xwRaECW4KDdsuBO7NOcGhPjDQrJlbRfk+lM5RdqYg99xmNrvRJpfeSG5g2
t3kUtRXwqMRMpMJcPAfSlpF0ysrDYSKPIp4qMw3dq2Rqn2Sy0Z/xdMQgYX1JeLgX
gddY+VQYloNGy5wkAwkGD3iG+p0ZXotcL4r1m8Ow7jM9yhcDs8Cy938ElurOWQIp
AM+E3bgNB7vKvfgx5S3RXlOlNDEFezGfUQ9zrVkJA+DYdtylL3Opjjwba4A3MGxO
psBaIVQVyN1GszORu28xaZJMkOpmOLIuCr6ijkO0cpXNbrJ/TCtHOVYmU3wbVrwM
664Mi9uKfym4Q+Gj5aa/TScxdivkUUVktZUcql8BCiL/NfRMzKZAa57aCGhcLhTU
W2xSo3JLJ2/B22kxAawcIxRzjJZc7U4zwru/GAdRyQfQbGICLK3aqpvGTZfsnZK4
juRMO1Nz4dZ1T+zbBALgkLnhj65WFHDsCpSY73aOYfZLKboAqGd1GniyehiM+qcA
pJMFM1cwJUxfuzcSI7JgAcNdcWli5WU7uqSQNkOCJELTQg71cWI7K7O3MOP8+zW+
RxJTFLsDQ9Wjb5VPSq80afJqQcztapWtkAQtTAprOO89iAh6Y8WqLgzDBL+tXKUy
Fa/2gO64sLyO4X5qiNt6d1rtnyRvHa1JJmnWMlLOB8Rxg9W5R/7us0PPvG4kamMW
BqK8PS9B5aCQkyh3vpNjebUrLUTT87Pu0qg1xOXdySGzxGYGCr+8IQhy0kyKssfn
euXS1/IBCQeTiAG+RP53DwEDsDTWk5roc+8zyyjkzyJbbkR8tfVYvZX1yDzbgcEP
weNr1/64Gvf5ka6dw/Z3Ap7fW/LIFKdNeAjpN6aEZEkcvbq21n3+/HiUVit/R4We
UKS0zML0v23YbR8ftCir7P+U3kfzgGLby4qA6OUaqYf56CilF7KUjR79IeMVyASl
gqSrJiWMSbeUDhBJcGka/Y99SZzJj7cH46m4P3EwYWiHMQGsNGb4YVH7ESiqoeHo
HmmutDTAUtcKse+31o0JlcZsGBfjJ10PzRkUmxv88mrOeu5R6RVAEH9Gjz/ewXgz
iapd9iMIynY9Wqk2IxpRL5IPpA2jquT6IUiqViTXqkerPFf5qW/zH8oAQt+ZKW0j
JkKpK12ZR6kzG+ipZkxwEhdGIyCn5/zQyEtDvNioVD1MoZ0UCXSQ7iGeXcDTHSTA
YF83eY+sHUznWplNvjipcqImou5Zo4KkDyRCo6CpI/P93gE/P2FfwixTu5j2XVN8
oDzOlJG6+iUIGuEkq60EWyEX791yxJnr5YNu6xq+MX0lU9faOOipRemhhHbAFdyj
+2QKQtq9X4skgYWfA1+TPIvQOT2oUWK6WSb8C5iToKGbwmUIsyM+fCH77Ef3ybcS
6TyLz4gK9LobI3nd17KOjsykAVW/uXtaZU0dmuhiEevPU2HmOcAITi6u9o2kwI4Q
eFzpBN1wFXXcZOLR6VbvJc88/WxpDeKD6YCjbfjmLXnhIKSU8eFcTgfNSNHl0Ozb
CsMxiM5o/s+qd5tXS0bOePXmovW/gxEeEdBpxYKUjiEdAN5N/RvhQm8ziQ6GWa9s
bXpcSXvYvvuo9T7X72loMR3L0j62hRMlzMVF3Esa8kZRqlNMURoA0BqQyA9Dqn4C
Domi0/teFw4k+/gEWSFEAvxP7PzBnT07yz1Spwm5CELSqH+t8Cr/PjU3WSrmVMrS
jb30QJRqEwgejTq8c2WIrbRAASwEbyXe/pXQeiamPDFdq0QQBI3SrHqbZh+l7lZY
oYLY/OeicZMzAidA7YFoC28wopPDfVYD03MdMXt9yOHYVAG2yVDTWuhBVHI1LD3f
9ByIHf1ZbA5zO3G2QDKrxH3gULYgCA/LbOQ06C1AEy7YNKecA1HShkHQn1xB4lcZ
F1WAaaS9XpPtaNP/ErFdrmmyL1Yr9y39bzsOdXKGTFAd2NJQ95t6bvtsEVKFZ2vw
/lsSGHmrsJy6g2kSqLCbUgjqv8h9cnHAUX/3RQXGLSAnZpNaeOtkyUaWJpeOGUoN
wyLFkeb7kaW+YU0SMEth/0JUqf4aCAet1uXEYgCb+bLb9BYsz2/amLra+QzFMZsG
wsQ75aAM9kOtSThUVQf9SblujBcdE4idQXnRlla5s9wyZdWPEdoNTwbEHntdq4Rv
ey5IPRw83DdwwKyH26TjljrHeEFwKOXYHksNYsOv5Vz2i67j7JUHLHWC/F+/zOCu
jBlvOXnxlWID4ceTwxzT0bJ9X7VwU/fdAuer+BKKIKiE51khpdq0oYx+eZs17zqm
2Cfg7Jyt5bfpYCy0BG9+dLZZrILg+hYKqGOhcH3fCj98xv46Jt3C2aEYv22Up9Ht
GdGhIh7xjA2hkYivRUDkerik8MRGfUnEdQoPPBklXFgGDH+bMwvkwNI7BtzKyM6g
+54y8UzKj9MhrCpdpYvoL3H1sHsDpl1TUIjonjKSWWWL24IDYMHg1mf+glKC3xQl
JNorCedavl2MIddesTloCbSFimBdK5+r4+xADSn2+vzxqEYT729pp67ZktkuDSAW
6UXjLQMZibslbtLYDXt4ZxhWFN1gORIfb1rFkSx0gf6uPM+cduLsvc59IpDW7/Zo
3dbDxdDAi7Mgi2ghjQPdrhjXHh/97f9q1Y+rln7+tJcFzDd9inPnIWCIXSEkYqUZ
lwjV80wauXdHkxv6231fWYFC9NlzT2uwsZkbm3DVtDPl/JwSN/x7kbWvc9TD7Nii
vOjeDtS/8pTDENlPdi8wXxJw15KHPL+1Sx4sOK3hb7DW5UhxCdOvqKXPmlzl9B9+
sfKAQSeKqT6Xv1RC3/vHduz62Uk5DxwHpXYN7KMoAY3/MrTTiDsCuuX6MriLM9OL
WafkC/hSBI/Jod6/PsaUBtBqUeKHeHUTeDnzsLJHcdXJAaHnYvToZOsyi3h7EPqk
QvLMz7VUE7tAvd9BhvkOQgvgUbv14Bhb9ZjoHGqVBgQiu3K/9JeG0hI449dMMJ4x
tQ6CrxzIIAcjF+Lt5U6qTnHvbYTNmOSU8Ah0y1eplB7gD+OWJL0yLh++D4ZbEdH0
ZGiQUXuiU0oeXTLYgAlgDY6+wA40DhtKHnHVN0mlzx3ek79m2EnpGDOuTF+gXPpU
aNfu88YgErdMo5cURz8uJ6oJFcOAVHwXmeKThqZr74yEAT6Wb+MF6OcBBuC6WGhR
FRYFo1M2+/nC7zspxEjeTfXjUai1eKhl7mlCsX15VgdoPSy1EJ425LOhOiaj32rr
71orMp9NuVYAEjv/kIpNevcYamB5V4r7RnjpEZdlCV8uYEkYtIQwuHDXKQsoLIHg
PE5/BObHadFMS+I4Ghi0sqa6JKeT8KzahrpoLuOvPE3rZkhWs1rTRMbb4kve4zQ8
Xv42+rPdBqDtgWRmCwRvnMdFbwp228gCQrWi8FenPBID6R3Ah+bReT41pZq0K9+d
NttEUpnXjBiWi6O8B5lxt6eeMwo6PyPADPpaP4UBp+gakkdyCZwgI12NHaqi8y4q
rQEtJYE/HjWC3OyLOEXlZx7E3egRdWyfNAT2INDekC143hypveETQjW/MyDAtGKz
s4NFMSevvnw+LYHGemjHncqjK4bVUkTrkEhlcv67XYLJDGZ6XxoxcY90WvQeuYZ5
7qTG+XDO6bWz7UGf3/Aqv5tnHvVybONBnlQgDUsOFg040cc0PqLO5+Hstb0S9vEk
ybE+YI4xp7Jg1lFagt/2J053fTqUU0+O6lXkCl/7rbcaJqHussAGZ77JrsAU7TD/
RnsPLt0t5uWeIPjo5TNOJkIi3VKm/EUppF/+u1b8HNtm2f4lAT0dH0cSpakGwPDp
cKlwQXKIstEdJnededfbwu9iWvUr4Zh4uuf9TBMmDUwur/jRKE5eemVPFsfSKAK3
idTtQO+RBcrD9hLajMeQiLLjnQxAquKbpaPEVGFOALnrbZNxAjeTepcwtJqR7B8G
iPccLX+zm2pTo1RWce3ru8OU63qxkYLkjb4kjGHuybI93i7V0bXYdfBQp2UkwOMi
/oFbjbr62dblByPRv0c4zVa5UKEzFOYz7oCYicZu2AqMfAuVcpSTfW0AHQKNtLmN
XfIb5AIax3CbGsSBu/yAURnJhZIup0v9BFnX+qgkqVCf9vY6xRhTKa5ldvW3E5po
17onWfqRMKhzoydNwlLjfm40pvqOIf1EQt+vBQYDEI4SbylC7u8bOWdNC/C+F+6o
+xdInV0SMKrB/k4w1HfCnrIUsIqB6xP8iqhuzLX3b8nvXSaucTSfG5V8oI4eNcU5
q68478W8hZ/GBjkeoq6tEXbb6UkXnoJh4E55eHdC8GxPpxeM3SNZ5ZGJFLigSiTM
x+Jlm+aDqbfOBvJH8h/L+QaGdo4ZtFpFScuEwPmvNX6mWMVTsyW/K+90OcF8fY+d
vGynqnuJBiVgPWG7LOj5AOKB1mMQVbRPJFn+3mpQUppJHgEP9iwomX7mhajL+Jm2
T/Mi1DVkG+CRcD5ZPxs/2T2I6x7XWIlFXUDHS7Pw+JuL/gkqnujx7PLUmPOGyBJ4
Jnmz7jDr/girFP8f6qQ1Bfkza9aMIFqrQCmWQlYtihjW6zFrSbiarDMJRMBUP8xb
rbUyszKCz8C170Xgyt2mw73cSetB/fD8YHHQFDQ3id2e3D3IhfD0SgTrC9DzWbCB
Ot+byUFZeNHZZmoafDbvaz68kxDMYgbX9ZVbdJ0XU806KntPTeItQnCnbCxAjsIv
l693Hg9e1tp6NsssoY+8kNFOJPltZ4/aW8LI3Di8vb2o32uJLdAND3gRHzrtdzxy
H8+B43p9wFUn9CAG2Y8Kj1ldAnVC/Uis/rjUJDOXlGX1AUbsBlT88PgmwQAXTE48
I2lbVdvQrOGqbYQec4LtuE1Emab6NoEZtA3dNfdDzTBXbdKXVxR0OIW/CmsrgBMA
y6slntdms8BREXUnu39A8X28X0BpgXRiVL/HNMOeMMjDh2mFMD7uwWr7LnaQFTym
Ri9G6GHEvd6SkXK4C+adRsaJOHzHAhC6/oKfijuP9Ho/fR/RNiWPQWHQmWPnmy1f
AfrbaEI2cFJoRlf8rDcufnwc8ff9dA2raIqp7yMvGyDYYiGaZPZ/JS0xhWNEcvGR
BFcqJc+fAa7tMJJOSUx1L7WP5zfRE24y4i8OIthZFysgmEJH2OwtBQQYlG5uBVPb
WoHfvZ56rTyl9qbmFtFcK8yKwOFuslt3TiodVUvHPooThEy+WYfe9tlOFmL2hwkl
mQL3uvJ9fKo/FOy4BDIS3UA6LA7Sr2sk2BOEu4rz+YqvKGZz49m9njvZbs3WxWWi
+wz7oSmuHHw9IQSotxwkMMpRGC62MEuD6pfvO7HkYhKsXc1j9LGnZZ30eX9kIR2O
w3UwNlH42cocZzF4Oo7KgEDkojaEuhCR3LW2zLGF2HmtnZG8aKQPCx9k1mrDCbo2
kqyGUV6X+TwzcNfy+XHKdpbXAo9uWmlMxM7+m8Anng/JGNE5nyvluueCBUHAeCBr
KU48DFBt+fQggKw+RJR+F7g7xOt1d3sBm/Ic4cE5vBcyWRLKQNZmDXi8kojv6+2w
bY5wybr4IxQlRBN6mhHoPOy2xqP2i8ikqocvN+oXBuDuAWZIF9GVxCWZgHJ30rDG
hkfsEWKJrodoE3FES8SjQeW3PEZec/3OpUp95WX/a8WpmoFFevwpmlC26nlLoPvY
xbNLbTYkj/k8zaW3ERf1/89Nd8TokqzpnBlZD0PfJ5WBwzRsi4CGMLVSak1lMGdz
3ehzKAihWpe4sEvvr2xjxL2IVJCvA7rVIcCxH+y1b0FQy5NFP2rHvMUXPyiWrLt2
rZf7HAOX9VBmvv+WBaz0scLn3fRcf4Bu7IdMrsJYexy1MNuHzYjvLbwe1S7LgNIs
4E9mVcfCr7UXKu02PagCgg9wYk1rNgJORW8+2CAgPlBm5IQ7wPYz2n0JM+77FwuN
tXKjdP5ZMGNTXnw0pvag0mZ/U1meTV6rhsCh5HVqKjmp9AU7OKk11NxHpkkKWAkv
VQPs2JGJRZpr2Jp49tmu11J7TulzmCt8bDhY2gkdIQHv3AUJZTbxm4xwH5tIUUeh
aOpLb7/WXyqb/eXYaTDjPV/LAIG/YNa19JkV4yX6ProVvjhhAkTZpPv2F3yYei44
I7Y9knwAc+k4LckNNxBsjieR1Bdqkmx+A/Ub4CxbgmlDdm8OCzN/IIu06Kd7Uemz
dnwufZuRyBNfNbID1uVN5QOUMmFKt4D1bjVxnPUYBijiNBb10Fp1jKCJtJAgR7W0
8m3fO2TS5J0NQ7NxT918e6eJRr9tFF1G8E+J3a4fMl5rdxAwUuFl9wRkcv4JkhNG
ZByCwEOuVvBeI0NpwO/s3Q/w8sWVTzAkjyctzYzlCFqwtq4PmZD4xLpoRAfY4TTE
w0p8mjU/SFYNUuiHB5Cm6SMXWvE+YyxgPXoGwfquwaYG/UWGEQ8oPTHayJHCrcmk
UGbRmWyNWPEyCnDLvl/HmyCXGF3Wv1Go6rC+b6dRur/bX8QQfcy/PYjJDUlFyNOG
9TOjQnfwNmmj3o3fTXoao6npt0AwbZtLjLAfgufFBiDj89Lz+SvJSgSQfhHnRmDy
xbb4G6WV+AYi/DrqkJZNYNqfo7pzoWXANgEVu1BGDLA9FSw+rK1lds8J/ONh6M7t
c/PqlmP2yzD47UNoZ1RqUsD2EGQl8syJFC0QDHwqPYvljJOEoKi38hz1zghY4Pfk
ldAxrvGKwZOn6qoxeL15ShE/1HNYVZ00e1Kzrt1al7wfvXTtiZeaIeW1rL6oO0jF
BmXRuBxMQ2kkS0f6mxIZTsUCzJEVQBPb1gYrlDq10vOp79cK8shVZOTwKoV9Iew/
5acGMbkUvGGLf747RL3gzoy0+P5AUbSVUiDzbBe/Sgm2E9S3T7CvbGU6UMSVru7O
eiTsuStSGLhztSUgfgDgTphCaK8iv8r5zuG0VIcQsc4rmDwE9dYkLTjsrTle8q1w
0AeicjpJcFcV3B8U4grCyA5tu8f6ff+sr9v+sveukiesSdZ0mP/C8qM0AYqlhPTc
5+0SDhErzmYR7dYG/Gu6XHq3UkTqv52BJ4CHtCEh7ygXZGeEaIx0wMRIG2UrEe2G
tYyU7p0YfabkozllLMan7ryBx9uSEQEtS+tS+ovRwkoe0GBdbQUrXLUzvYxs9xlH
mWLNceKvogpULWzp6QPHgaUX1oxfeKEhABxuDpZZULnDyPrjl717vZFPn6rc6BAW
hQHP51lYnhVJNaFD/XWNKP57Aee3BaHM2rAg+jQBD/di4xxCqylLCUZo5JEaeVwI
r4Pacox9vuwSUERAH5oMy1OThQRnXdiZXcAuip9bL7bNGJS6hFEydkhBMFBty3t1
VlXESWFHWppU7Y2Xo0dW1msJMogXHXDREXAizIU+iqKYGzcFyOMtM7t5K3ZhfkLn
T6TghMXW/Of9wqEO3WEZzFY7tzHDinMHZ5VAUWI9pF7+gM6/fRpZ5ryfRSeHyR4r
ckhSmwngw0ll8YB2G8a/zirQMFO2c1Vgo025fC3gSaTsnQgg3Xa6D6M0aHXvn+Ct
KsW4jF9AywYqgzwuVcQCLvWfyTRWbfcCWO4fSW994a+U9i/dKVtUbkBZ/eQw/eAp
0gwlKiDvEJ045x8wMuLjOx8TPeNs8OP8JcJjjXKLXb5T7etfXry2NpZGjMHAKPCo
Q1urr0u0g+ktbj1tWHmFVqZCJMoWGTMtjAFEmCnCPp7TL4tPhuKbnlnHU2zr8m0h
VS1u8EY2LUt4CzgGMQQQ8JUXKkBLEiFfRN+OiYQsd6Iv6AcN5pTnhKyXXC2rBWAP
pO8R+0r/zJI2RQmwIYNs7UamLLOfqP/+fAmz/JgbuXTU2A0PWvDeYqsYalIcbuDh
pIzVQKXiIsOmnVPCIl3V56qm/oaUZRFcekgRmzNjQQ5eHigmh1ZdNaH64AqYEg2Z
irbgqlN93n5QAnacy5ckMOX0hJXwrtyQ0vVIompA1ew3bOt0on3HeuuAKs4EBnlF
fGG5YNB8viv3z5ltObyqixznfQLE4lFDI9+anWoDWHpnICNJUcJcM21vsaw8/NM+
LCUVd+ttaeUDH7ypNaqwMHDLyLXrn6ZoWhaCTi8iTciPaPpxP4bBzD0UDAIOj3ND
Ki1R5EdbtDr2Clrsaxg6S83WIPPUl8B5xdBYglkIruwNZDGrRgUdTxD0HY2SQ6w6
wrhhgdPjHY8aYMF+W4X1L8rkCSxd66lEUtTWHVTpWOKkizbbNviHu0yz7UpOLp1j
RK3i7X42Lp2U7CmUQNckpFf6uUh+DRRmvyfFESGOy6tLHKzYNi9mAkRl5QGaw6BP
b+msUl1PxzaaTxdHrmPuFIKoILkksZkASq6FEzRE8gNUo7hiiwYNxIHJkIRT25H0
wHA74n+TOdsfKMRqAdYlS/jaQ5gGP0l2DivXJLQIsNrnzSGm+xJ7f8vjx78YuqUh
7IeHsqQwqYNakncxsXF0e4uI4+4mrUFlrmg1/G/TSLGZ1rQr35sGtDvcXI1D4qwQ
1zsX70BnD2TePfGx05R0o30YXsjxqwUJ+O5egrXcdoy2l5kGw9NjScjjpGvo8THP
DuLL4/55sOln+URCeSGmBxhzwiLxndubQadBpjUJIMdzji+JnFs1S8dzq4hmVw7l
Oo45ZMiLVoj4NzUp7VoeqDnzJ1HxVgdTFOhP+gSXW+qvoGDwBy+Qv9Olk+QJOpM+
Tz7mm6Xl83nd6Ctj6GDULov2SUGChyiDBhCQUBwyDSd0mozlkihI6h7ELmVExKF0
HGlcwqNMXmiVsK5lFrqPlrV0MkpgPPhbx3ik7wY2KELrdpHmIlvHOUCVZ4taPA3v
Bt5R0YQTR3srMBXkBCZfKIUdMItDu13ih+xUH2N8stjVSIBaxF8EqSHueqWRoqxf
HZat8KYP/hr0br6mnQV0/Nj5vUCUpywLo8jyLBVQVCq2MbXF3U+kY+N1g/CQZglE
Ge/jiWh5UvyNsTwErPuxJBAx+dc03wKewYLUT/0536XLhI7t4nvKpj1xGEP1Epyy
9uXJ3VQakEoKWMZiBxgXqg57sm9ZvRcSs8Pui++DUcW7kOFlf4Zvto94zllbyWSJ
JIuYW1Vf02rdct5CRA6ytpSHG34t9/KTdd6A8RJEpy1xShUkIQklb1neOL85zuHU
W+w4T9hA7dQc5ya/Kc48xRK1qfM8Fgw0ztfpv2ebaxXq7VRujhj3zO1LnUNxbGOs
GRlVROmGszSr0o4Q0gmJRzFku4uzIBA4seKkka5T7JLwNma8oDLUCsNWRuH+uCsX
quKhgZzW0RBUGq3e+GOHAgPKG2OGHTXEy8gw+qM9MdCE797xP3uFYkHDqVJjZM7s
zXqBE66uEqRiemYx0WTDVSdeuRtbcyhOObL/ujIGHryAvP7DgqqOwUf/gPGw0Sdx
Oi+FjiPrjIDNsLf9BhNAdc/T5nMiv+XnFYfEvVakYhnNuMI05O+LOxgwxkjCQ3KO
N1iF3JkC7vuiMr6htmg3qlaQMZ3+gvopD83kCcdY+49S/ViTfzJTDi58yBtO9tex
U2u59DTq+6iXfJBbPlEGVNMLrHIlEUmbDu4QtGwYGgw2k/QG9mbeb36rhpaPecQY
8uB8vXGntc1cUJ6XeriOmoLopHRB7sB96886KYLCjSXPR6Qh+5sQyrn8/CwHZbBl
kG6eyAhKfaAucIA/UgGezxieOT/s84QuD/sh15BJLBrzYo5toMZy6m/vGm1aFJOB
saKXKFh4JC4v6Tq+uCaUC50gSfMG/H3h16y1hLd4LYbPWOaiwam1OMNVKDSwlwQB
Zza6OhV9VQYE1dFfwuvmI1aCBNjh4VuKrZw+ZwLbbDWrKIURmYCGAUO2Cnkz+7CH
Iv2V6dpFBaMx4iinCv0SbrLeT/DPcieygrfunFFaOPGo5HuD0znbuWo4DiYUn29P
Bt2Ql+em6j6UFj+eoo89Bvq+kwwCh5ovk2aYFqxE7i73ZNHX3MyT8QyWokrklcTV
KsyoUimCWUZJhfOPYYlokH0Jm7eOmtbxu6JEzC/pOzusaIuCB6HsN10sy4mObQTP
H63/7sKdYXqswvjijFagH+kStSBJzzvkX5Tpa9yjCezv6i6bAxrC29tiyfe61v21
OOpquq8Utd3bhiF22mIJza4iX9GfKv3h8tOYCP/0EKzx7Fx2PVAQ4WuI0E7zwItu
6MXsBguzmjLQGsav7fAd/b1+C0SPFusxcqTBOPJRhzPCsQr/kP/VsgKkdfHSfWo2
oIgUljm7D5AuHIOCzlMhn94g0B4Xj2FhIZczhNLPDn/nnMW1Fl0z5896nD6NzBsP
rjPIMrqypkh3dd9iTVyG3pmYLPvm59iF2Ffnx+N08oZPWpCXhaHHDibUtq3pVSh/
F1RXqnv71Cn1qXbfLM8zv+/N4jJUy09m1qaiuPnDmmdvldcD2j8JwpyoG0Th6PcB
hCmDoHqIIIP72A8g2PAP92sRknK6eZxYFcWAmCd/UswaID4CKCer5MZf+uzfCrua
QT1VgTn+9UzXQO/bG+N9Xo4IBYHDAzMYzCJ6huq2pXwsDcfwkUaoguLBFCgjGMbx
7wJTa594VgaQv/wV2RiCArFdSq5LwBS43cTP5n0TdAbud2pwz6Dn8bU8Hoblm+w+
e/RMFuCqa+HC/eudtpLEJlAGabM/cws+htYkT9rXwOtPnk9ucehQnNeyc/aybUrF
KXZZZksa3rWZUe4XY2awbBYOcEeEl/ufb/zRRf63nGqM3wkKWzPGuxR5nTDCHcUd
WXG94ymDPbB5ElCZsZAtb4L81QMP+Qr1x1Oaek1Y1WgNefrrpdwqBw8pkqN6Objb
lMEwRm2b/Wjnz+9vz8nSzQGit1UV4VQFUzeMrcEWZFsZ+0t7+1/90Hp1Gei24Xkp
QuCOHVeljLtiK8Zr3GFerrzgtC2QSg+BkaFeiwBNEsqviQ8551+yGzajjGcs9xYN
tT2ohTrvOP84UAD0JaOIjEjSSuyd+SBCv0odyI7jBMsHetRL3n8sn4ZsG3EUxWOD
dTXkDQwxfIuy5zjdvo2OeXMfogCGX5q+XvZzkuErWUvXIEq76/CxBO9QMA8RBoig
Vj361WILT1/ODKXQid8mVR4RInGUKpgLgGPuz/fTI/7Fc4lTkGbmvfR8nLh1vQy3
9swomrnAk2QjJtQ7FYCM9zIiijrh2vpLhAIwEowsfxplp2MbzKYZtlb6V32iuMjS
eoGXCiT2zte2wPN9Ru3dxYNUbapP59DW7eCbgqdiTyAiJU8F6kXwc+j+F2wFyJl9
+R2PsqHrWeFTZ8oe8oFciTagU9BPCjhK3KRH5HdHE+TE47p5VuhbaFivqlzcYFBn
vBGhw+nMuOx9hGHiQ17lFmHtqOSbYChdCgOfQ1fVIsgKbTjy2OL+8Kt5Fcetd5KA
0gSQXor0Z7u0nIZxlbVrk+k9CYa39/Y2hpFL9pNrZ43yEr0i/ghYjAURxXBpbEHV
PqhO56Mi1jTOtm2AVz1oNq2MYHlYQX2fmz7wLtVw+XFfxNfAwhNsnQZK/H+ZL5g0
1ooLolrvMoxnnZz8pgU87S/aWMTkqGCPWGDuLZBBVJnRR7yTV8nGPYFRI1zrz78+
1V1rwkAXXnVx5XKAfvH40x0ohpvvP6C/duR6mkWSmwwlNuJ+reFv7NfAF4IQm63g
jFWnyLhgn/rvmFTm0Pec8v5Tn9Ob76zNex6gaTY3zf47P/RID28hI/mjt+iibJGQ
nnSWhgm5lQgyISAQPT3Q5T7euq9PHs+H8yI+DyVU/lDaSwvE7ZVoV7PElXs/VtxT
RknF7VMDNKIUugK/18b5si7eF+uxDNi06ZQ8iPKYr8k9Ni0T9jbpHdyP/kQwIUw8
IGnEuHMQvjNj+mzd4usEcBbr5qiP2GWmfgpsExSZuqKZxfNORZpVCk/2vNALlP5S
T55lG0MCNGZlMyEyUnK7EuQckRqAn3j2viXUthejsmvZz4mz7qAh813q4LAFa6Ia
Ycg7xWvNKESdZZDZCSRSG6gviDLeXsNSQith83M+I9WS/zywnedIRBydHgfzkuxt
deCp9vMOoQQSwCxRNerja/ZX20uTtgHQOajWDg3FGY9NhlWwkbJs2dGuZaceE1qI
lE60wT+TxXt+DQWa0OUci2QpyqMkLXUEIWLOl3IzdwOq+1oEiTpy+wplb6hvLGrQ
GbyYd7QDohdXO2tH2/i2dJvt0gP7zT6i9dXeKsC0cQNJillM5uNnxAeu1n21B/Wq
A9d5hqD+btMUJHgeL9vkwVwGrXeJjzOANIY0M6iqpIeaEiGTNCE/GKeIB55KYQjB
bC0yyflcJyDTBRLCcqfLybHE0q9nezf5jAs5M02v3RvWAgCRJEU8GxCHDlDVjYgr
38yZpD/sX8of9FLEzPumcYdTXCWH/2RT3spzw6RTxDgwSYjP0zj+qJPZbUKv9iaw
M3pmNx/Q3HCUmB/Y1BQTr8nFsOVsZAG6kW0ckFXgwiZK+HCcWjQsMWr+fOQZPbNZ
gyxkkb+PdI2ul1i7wFV9jdVXtc5JQ94c+qmNEVvNhzOhfT2zsXP+QqMp9RXwvy5q
8mhkhTVNpGG4/DZ0CYmcqGRlowVUixrw1BTfjLvyz16Rm+V0PtJbh6cMMKMW96W7
hFMlmbuyJVWSwsFGHIEcRzVR2AyhoxQocGUJLJ5nuPKVr4Nu0jis2ScajouN1ipG
i4p2L5OMPxd/7vm1Y4eDOGOa4XWLVjPp3tSY2+Rci6B2nwMZTN0U/XeRiB9JyBsY
BHETz0BkUSyaqphaG6yOZ8E4JT2V2Dzm6yojr72Jk5lfpHP1g5ZKTo7sqsc21K+l
4vCTLMtVO4wMPZQbivtazj5sfBoBoA48FO/aN+vAhaBA8wIRJvxTCBzPvypeqXMM
QjswNkKpx2cOTVkv5i4lLIZXihMPn5ZWJ2aOamk3hDfqJCsPK4lMExaZq2o+LGst
vgcbKZ7bysQcrY+yih70gS4inTmb1WWC/jrHB/2Yrf+xaqUKWBmP18epatLeUDpP
3j7fhiafFyUkqAulJ0l/q584AHQEhWZpiyP9p15XYvjVQohRUUzcb1r5btbHthKk
7AENZk7m4tzl4F6kp4+jPSzLWFO/TifkU6mkBKkdsn9CR8AV2jMBGmA52Be04VJp
PhQpJ0mDeoq6gR/rhqHIoSzaGeS010jnjRBW87/4+Ongj7+nc5KuNbNOc4bmUuYa
Z+OJ+lEdAHHNN0EBeTXwK+n7kOj6QnPfJ+0Bv+42Y8vIiRhJygF9ZIe7mqiI0lpj
0WaNLHq2xSZOOZFOmoExJPNQHSODAHsHDAZL4shJYZL9yWhrnGxEtGlqPu6f/o0x
2HnbCNeiKKi6zfcSXiurm2xQn8Jz9mUq8aJTOkCXxb4P69zpx2vtyY74E1ayBRSz
1RralLZepcy7uxG6yiwekVFsY3/aNv2A7ggx/kQVF0Jn2rbtZTy+eFW/SRW3QuCm
TUabxcDQMsqhyExXhA7nu2z3cq2ji6JeXKkSFZ70/eNGvARe8KJE35Ma3Kis7RK2
gEE/L+c7Nm8Td8pouwdgwQ4OTYen1HUXf6BBkjv/+xxjnKS+nGxSzFFxE34sHJob
5YN0rbVUDjAectvNgY/KB9PawGvTywvb+Q3b2SOHMWaTWUdW7RjfYxXRWyEGql9N
qnLjptgB27AZsJUVJCGs3C4UitswV2LTbsLaATiPGtw8tEjq4lpUaxqE+h3dei5T
RKiDtBhHcUM3VlFqGELWQWK+OBrj1XLIYC07mOwjBN2GN13CxXKsyhcy8x+4icag
gBCa+C9YaCHODls8cO/UYzj2z3ncHyMRvacWF/ZUHxmujHvime+isrPeJBGuZshJ
0ADPtCyvGG890mJNebr64LkMHddGrn9DsbSatFltr1X/TdowiQlc8pk/VpMF3m6/
19DDYpL0RPvIDbGYa44+24eYr8qVhNp5oryA/CkeqYaJXXW2aXOmXtOCgiJtMRhZ
eox2xIPs4oikab7s7XP0ghA9yYqyvnLa1NkRywBJWfHkeyTR/jVppuN8ZUdfplGe
B1TU5bpqDScDurDf2+FUCvy6j11hXsOsEHhetafRvTXOkOlGUgn7dY5GzNyy0Z32
sgM8mQE04Xmeqc5m7xFicoDUha4Z3lzFJ8dlxI942dXhcWiNyJvxQSLarhbEichs
AuKvPlZgN3EwbQsnNpCuyiEkbR0ZvfXsbNiYvjFaCY1dJD5DgAZMy1feaCnUq+1y
OXwhTHNi4WDBSttBAV6RH3LztQBBlfxj/590uQQvcZ50oTQPG0uotZzT+JaC2xpb
/ql0+HtsKQJPXlsX7ZSRp466apDcnf1IYUhfQ6WlMcLNrJ8tivarBhE8Lg1w4n20
Gh13+YCLS9DQSvKEQY6t1Fd8c3T/7RkqZkrMoO1YXG6uD82peSOgRjULpfbvEWcw
pkMK5KNW0WVSkmAWBEKgZrG5tzwkB8QEp1yNv7b1eOVGZOM57dQi7N3Xqb7ObCOM
WV9kYbTFb0fWzNFVi9StyUEtZ/MiUBGzP8qCqhTXM7j4rEpKrGQ9XW22yB3fsEi6
DsfYLmuPOKeeVCmevk8CpFFnos011NjAepEwxWzHlQqIF8PpkkDdHXatu0+wnON0
tY4s2mh5kDLgtGS+CLGaeGjUOMfHJeZeR9/TySFmQEiJAZRa7NkLH0Wj4iFs4p8z
sXdyCnaMbT0RnFV+fD8tEoqks1ByusFoVAKNd09JAZHPRpfD17Yn4Z1w1ZMBRnQK
KmkpY7nC8ToJK1gTr+QGYUvUjYymtnyrH4PDTf0DkSZ5OfNJtFAp493ORG4Yv5Sk
hvS1WUuTGrPkLw1ONrH9D/XnbVilpeZtCb3LIIPoSJFvPBJ8aIOW2IjRWW4ZAWQr
SfsL+waiNPlDMg67/pbXjtgiD1j1lHdBpTKTmBwMMjTFrwuVLUDGMaNwCBB7cZXV
x+zPWHH8B0b+rUbnhPztby+DzrPSya6fFCIs5kJ3Koo/x1j/Zrpq1BS1jxSJeBou
lF1r0pZmFhRzUf6ymFMmH4S1dtD/33qYb91VV0A5+FMVp1bTpQwWKyAiwvzFCT9H
zfkMnolg9ChQM6hsTkeEPxahM4sgGp2/4axwew9HUu77D4tj3ambFHYKBpkMnE54
P7QCkdzWviayLByUODbBHQrgQDgmmcqj4wqWgjdoZLBuW8YB3aEp+Fq7l6ag9bdc
cMWwvIVDquLI4cFjWJpGcc5Xo1s3mMYpdI2oqW+SFU7Gbt4fHtuZuitk/nV6JfF9
0RaAskwFTed8RqtTJuufOmTOYIqIm6AuMdAuRGWpj2sGR6H+wIayfT2BqgE9gQRH
0QiRxpsZ4lmltC0RiU4sn3ldPuxY2103lFIEj7HuzFiW7y1tQym7ro8jH5wx04nd
VA20DvwyY67HAWPHisJmVoXDxIOUZBIsCFowwriwLZ/0MaltJYU/9+9IxKjyZ6Gb
AeQhDtZo4aqgdGB3P1rPxlSfhRrT2YVC4wmwk1oQYd5OjbRCOwFAAMbXR/xAVL1k
65/DOiuVxF2FH6dRH5XI/a5Z6SZhPzXGgoFJBCOS9CrBvEncvGjMZvkGWShqa4g1
7mvHCKlOY3Nu9ZWnnGWCR+Y2X5ukZcO8OvBvoBg4jEHdLf140znsXs3E7Kh6Stz6
2R/L4P54CsJSZ6kjp0BI2WHeeHixg2lvLC+cEyQJCWgUeCdcAsg0EjnTCTsq2f65
oAcvH35ev/NY+WM96ZJP0IBhcONgK6Z2Csi777dtMNloruPhlhzYWqM6QttZW7Bf
1q52i9jJ9HYUvYAx3QBfwKOIV9FqqXacfz8w6TKUupxgIn+ZKqORq3m+uanndbLF
hyPTP5TMaLe54yVRtU3B3zYTagUsV67rGyweI6Lfq68SP23HVgPOcnsqLYrPnzUm
wXt+jJlko0RtQmKuwLjFUj4yx4/acufkJPZkjYtuqAZ9t0B56Zo6gm0FexZa+AEP
3VzUcsDmwX9ZMxuhXHozTo8IDja7R5uQiC+6cfY9eMrKWG2/cwqmtsI5++AMjkgr
EPUzrTnPKcq4idmidHCx64cwU5KNlsOxBRzu7IMRSPXZXLh7z2xDBqi/P0evCEbc
PtiqiURpx/BvE6Y8DwKwNHvzxzGrkeG860oKD4tf6+noBf2wY0Ywlwu9w8yHOi46
7FigpIsXvAxtLzFCXE+AQKWCIp3ZY22WdTPzs5H7PvrjOmiVIVX3Yf/LR1q5sB9f
UviW7srwKPKTn2ofId7Y1tw39V5Wbs7P/exjQzFKZYIL242zcr9w046IFHN5KcS3
gHBkiokhjVWFGl16u///2ReaUFCverNZKwDB/qpkyKS1VcWEppEoLnwL2OXSkd1t
MowebEJmIMSNIVpFPiW7aLzhJ5t27jPWB//NQFotLSnFubKeiKslrT1FsxBSKSir
DrKYisS89BD5zY3XVua34zBBvYUKryqvTC3PllgDPrRvpeQ37NLI2aY4OBcM+N2K
L+RTn+RUS0WGN7N653oE0a0ecgTd0fAUL3YAFxnqgDbcARgM55h4g6AExgeyEE3o
08plHbA82dT97eak0MeNZ/A/EXwHuNRhgxqInPjU1+XXzBtSMj59Z8B/az4CRprD
wrGDvNjgvI1L2hRfYtQeUfwy5IQBgc8DHN9/1WgkjT5fyXAM4XEoJA5LoNEu0vHG
MihK6sXDWsNeLnKaYdubRspVbVnXKielis2aNHzE0RhsOalIe1cf6LNT2gbzAxAW
sHDKZYF9MIsd/trVioJO09etETkLUjjSM+fyWHLZpwWV8lYdBKcxf2qQKihmgNJb
Hn4UBqvRZFielSktbQu3/9He+eJPouTfy+TlLk9/tx1BvcGpwR9HMZl2cqHwSqLS
7UQAMX8U6Oxvl8SSApvF5M8pRPCy8cOMlpAC42JO7CcEEYYtVylU9IgLz6rAx2LV
wzPZM/zHTZEQxwB/xNBSRKXjFCkgjnsgkrGB6cri0zR1BsvWERRMeU3SjzXHUjtW
kFJUGuUGMspurEF6e4I0DplldGY+3aGyp5r+3kgD4nZTbrMM6pgT0/Kdm9fxZkr9
DML9u2ht7r9KjKLGIzqOn1tTrwSasV6oqREIQk9Hhm5pjcsxIuJWeS+ePdnAsr5P
DLasqWDNG4slDpkHf927m10GfpfQMmUNWU0drg3St2jrP1ivyGmHo7K9kOCYR7G+
0kmjnMWTEUlMWyuASdcCXtPcPLQBhJP6E7q0fmCN9xe+gTWRG5Kp8aAhVdC79yIf
EMhCgLX/2LGLOOjsAr8xTm9FAO7Gf30u8hyHZbJNwJsYkBWGOnulWTOK/bA0IcZU
vKGiWvJB8j850TpAtcpZmCY0xGA0c2lxtKZJC7UmKTiF3YRzDhwiqbcFhPci8r1q
WK2ZOLzciuI7pQ8JG6rWU3BF/ZcTVq9MNnYSsoVO5qdD3AG2gpeGRb4EuJS8huR/
PWLSxXORoNoc9zJKvXSdZRl/nyEydscy7TAcoQ2h8sa3TJfdmWr5RJJ8/nt1wYiM
IciRCDpkcaWr+igBreHrkr/ZX7rX99lfnk52tCmQu4nyru5gbucjh01fg23ZtYP3
SvJN/DBLStkxMiCT8utkNLxx1axtL7OP6wzLOyoaBemctFpFik9gFKKz/rZ6CMC7
5c/C8k7JoSC4GL1LnNTO8Q/e/YILxxjGSUxXjk+EKH9B8aeTLL59Wq3TgvLye61S
dgZdKTgu1ve7X2A726Zbt56lCKY3V0/H4jlZ3YhF5V4bYuQp0EwRnrmNUPVrJ1aw
QWXaXFdTnoXo3GLze4UlQJDdo4smbPlWgBYv/y+SXvhsadwo7uz9aYMA0AXPYsiu
g3naVhGYglxJxAFDf6Igu/nIxdAo0Ao9WaeHT9dcYPARMjjVW8GsfS9ZTYZJgtxB
Bfl6AW73LvF+lLy8b3VUT1jIc50cLlOVJKQTLm/E83rB56P8/SNP95Dbxfd8yIjK
1aUMAG4fU7DXXySi2vZjWT5rX1fl6NQpCK5bnhya3Ggk9y18DKD8Zeyd5PzRxLMx
N/6Dzgy28Ypc+MNTDNEFgzNoBtE0tJl69+7qDBoIpZDlgxbJir3GaLN6wvmWhPbk
Ucvz+zaxDHlAanEiJwvPEo/+62QohMTU4obkQlWnzxuWMk6tB7L4Ovt5N0oOBV8I
lJBHVI7hDi3ba8DsITZ8TZKN5ENm3O+eeBbVwWbPlURy9T4W+qWbX/cV9z0Jt78i
fJx3jEV0DAaToEqTxqic73crSix8F6WdkstLNPfay6tNzAmxT//Rth6lP1X6a/SD
j5vKf7fqUXbuB1JsN0ygRe/RHeF/NBTsx2PybAzmct1ydPJYr1RYc3MDequkJx4W
5oZJaZoEGNW0B7LUNzBR3hFenX+jq9uOnk42mV3qhTn8afOnQqWn56+z+7NdIq4r
HQLZjAVamZhQX1JwnU5Rt8goE5Q/z5oDYbY6CsmM7g0ukfsddEGL/nKDoSuVw+K5
kihndohD1N1jpGP8AZL/law1dPk7iAjzTQEPqL9Pfq4VD12hfIaiYh3pzujlQArK
tSv2dMFoBGgbJfArOGBJLoXzn3RgnTHtIj1HujWZUfRZF9mkFlhCrgaaphQrHYdj
hIIO70h6lVKJbHz25uX/5aC0WhFvEehhqIKH/uw/mJw3Nr75zpaFP6bFLDGwZNd6
RhuFTUY0kSyWOHkosSP3OSIZJBhw6FlvrVlaxDEeGLNiO4BKMUfMYdG42sh02ezb
LIgU0WJhzwa3mC+cVmHskLqLUinTlyowPwaIy7ozh0fn/NTdg61sw7stCTjcr0J9
iGsPjcW3diMqOizMucGNI/xnss68BgPHcsSzVjJG0+62woFueWQ319jMUw8iKYv1
JDQ1pTJd6cJQ/V+s9Mmcw7CJnK0lAS1zs2pyPUOFUHhvMhgmliSP1jZhke5YoK3/
iz+778ET812dM6wVAcEbeF22NafaIHatmD/lyLjUWayaByumpZiwdE4MvNKQgPv1
EtNxfRnIAuG8kxOxOiH1PRZAyXjAZr34wbKlncuTxIES39M86VuweSf8YXzyUmAM
H8haxLnoG3RsYdB/soVyb54SJ1T1ni9OuTFgwiNanf/Sbe3HFz+D7NliBoMfRYvt
FN7TD1ZmIXUYKE+3tlHOMQKZlzqF7dx0QgiAjFsm3OaRr9f3cns0B4GAVH+aevqJ
L+tCQHOEI5vvHHbqpC1+RhfZZPCy7+hqgyO37yzMAO7pNCuXboB4sp8GRPp2bDra
bMyFEDYepHGMIeibAIK37B6wyuFpFQH9Jg8Ht0WI9TqsyOdse8qqlCYIicUuce5b
ykZM7MmeRsofthcQX459flEd7/GBN3mDLg5VZpJxjp+VahJPkw0qIR1UPoXakb3y
lmGFltKFJnhV7M0m4Gf6iXPePX2fF3XgM940Js9PVqVoUUd2ASrtteq2N4T2jbwc
gpc2yEksfg/ROtZ41LdR3D1BNNJUb4E9ZF7o+qDOjDbqyFcHkZ0JhZFl9EPW/A/Q
R/VjsLn2bcpWs97T7A8ytGRoCbZ+YfSw3M+z2VibFBAxVYVKPN7uXd91yGcViEz9
waSUf/YVNf0k9mfIFhK8hGlqkCQtRnwHhugdGiPzfJrpRo+mKlsOyyTSPtOYkpzq
L2xbOTk8jAtHxJrETF7d/LPtxtZBSm3gx4HghNXHxv9iL6/nKgBeZzJ8P3+Nv6at
SvrwLztygCBJ3UY5Pv/OAN3GJyKCXN+HNlIk8URZKia3J/yZIi1GTISDL4+DR1lW
+vy+6TFJgC0K63XWXzpiRpKmL74V/q9da1L3z2OmT+e44/WzvyHUj75srYCrbaHl
a3/8OfjX7WNJBv4Y1wrC7lGUneqgj59HNDGqUgLyLs5tjCDB3pQOZ69zoDscBjTh
ikvyUQRACy3SKdZ7sQ3Ds0nv+uIsv65sTqlME/77TvyKyGCdwkC7PCc7KJfEtRSC
6zqJ4ad1qR9BC2+BlMkSXlMMKw1ny27G8Zcm4yT4hagrZnXPCg6gWsnjLHot4mE/
1vPCkmYAwUsGUV8FBYHDwTf+Hoe5aT0dWeaqoGAxk8LIYE1V/x7E/ddiaKcWkVcu
Y5OFWSJIjdwd+5Ja2t4koVLzt3Jn6zoo6nsG8t4QpNIHOqo2P85F7sZJMqYFwjP8
7nS9+pXV5rPbv/HRqRVbdRDq/Wd4X5iVxH10maGZPfmvApskFZJ1xVorsS9S/oQA
XASOv78ISe1ZVnRdIYP+tojmIohA+vdjW+PoNgVFBOClHt0AMv7QxwyPbsJGR3tH
JDW0azT8xsazXWF4j6jmWGc0QcAzy8kpG5YrEFD6lYQJ8UmqUkdifba0wd4IO055
/NlkY5lgTgxDknBTwCXmTRhodyErIOnEW0c0w1i3EJ2PghAk3yGyb4Xmh49V+XVv
CYlKiqCYvzCn28Y/yIWyU4PwVgMePczxAkd1tOFIC7Ixbj5KAzjRGN7u/A6vZeQ3
0nYMrqYrottiNnsiSj8TELUa9cYX3MYDzepoY9dBW/p1aO4uzY6cJGmq78xZWLiN
KnAJ2j+5rB5nTNVKo8C1ujcWGebZSywnQwm0GuAkOMqAMTv5e9WpNnsRC2vfJRxP
omk4THUrHvat9UJfVrET5HkKhC10Ie+2KoF0M7f1XA2/9VqzASBQZ5mcngXsue2N
nXLUPxLqY5pbMhGDjk4P9LjX0ejtu5jpHPsDRcmtARDYvMzm20kHWbEzcfKrbTEo
6gR7Q+iVopaqTvIlxBDvrteNVSoxzBToctV+0w7HIelG9s5P6CBrgAe9tsT0S8M/
l0TV2NOKPRpWjlRNPvHENIUxk9M0nYp6dkY9ziOoSxmYb6biJ1+LbmMGt0j9FP4l
ssrK4SzlBJGGFLQRS8oW8i/plQ4U442/hryP6GL3OmXSDfVKNzjcBwtYnK5h4OEE
Kgdx+EQxsU6Rpw0RwVxuw7R02a1V7xAKk9Xh1C6zgviftOApVz/bYmvVkrF13Nrt
vi00o+wYHjDczRmn0+EzOyakkqPfDYIqjUwa4gbIJmVi2/QAOlwhEG05Fh2wTB9v
roBcLI2g4d1//CZxUS6FJy8efuGWQD4QBX2uKqgNHV2EoTk/x04kEBFveGnHu637
aSX3SxV9XyrYXVFL2mfdfWp0jwozjdMuzS8dhyQQr65D9f273PatuqH/hJ6pPGiJ
eoOiVY0x+SYJo77f2BhS89N/ewlCpZiDfRHSw1QhrxN7fDOD9jztueg9UMnXrduP
yuyIH96+14HaQeZGCcuxjIrre87Maox+b66/38Bpw+j1xZePJW40G3aHxXxqDMjR
9lek+jM8cyUhZYsmm0B35evyfXRgdojxnEkhAK8Vu/2e2a9UD2YqsxHyC+qYK1N2
HLXAYccyNW/kqzbmI71Uvul8htYxinM7hShZUjztNKTVcoMGfiMKescXrAFvZAt9
mKQuTnxLrj4SdFPqebLAfWCQyfsImCrXpWroj3k0+kv6dqLCGzWb7aFFMtt/tPbr
xMdPjCd0JtuMU0ZhmIBWXCV8OsJFDYzxwrRSQLdrIIvSl3M/VlEUBD64OlIHsCR4
nVTJFcMWgCIzBsO6Fb9Z/0cundz6ORtpgbVMgJTQYmFz/mW3qmvFglw4QxpxpYOx
kfkPkgqEJE0YMF/0S2PfSp9lbcTZ+5olCBq4TS/wi00QBPeD69j90S2PjTl1peFh
vJYShEiJKvLxBd0zEHexT42ETjF827vPFvc0q5d/ZaIUaxgXXWsXIceosANSiFJg
reIxbPECZ2SiwT+Nx6c+2Rvq1TcMdbnspGwV1yFOqlZcYzKgAuW6TQyaayGlxvFm
cl7WOS8G4hbpA8CE3vh8ERrmFIBS5ug2GSGK3Q8+XV1/rLTUMnByFFZY+r1QlKMg
K/TkuHlwT9xGTXLCJAtlWhGvwUqZMdFmClQa+7X6WVINS2kTJHglcwRZkYWiwB9F
QWgOsiDDYPBmZ15jDWY45Kk0pAA9iWDu700qkz41uaNcRilnLFvJAcGp/Ai7QeVG
GwsGVueepNzpzuwMchZM5hEgoo5Tew+sMCbdR015sY0/6jaaYfTLYS1yQe4S9h2S
KKQL9921y49nTlZsGZEcD2bv3vGS5EkGmPVM8J1MLWP1Rfahj0m5ZN+A8pRjMlKh
4jnlsbwGLW90YOhCbOSw4YFu0EpNCWwDG443uB9aYOvn2VPiJntnoef+qdcfAznx
ZGVgVPNbARfSZ5MWXI/l+RVgob/oVcj0l+4jT9IhkLf5RTJuV7tKTr7L9EInk1Px
YKeKsVSImAs9qXllKUDjk7lHkClJhoIrlfBHyo2XtZNx4wu0ZiFsfIdGo9RD1Kar
IClvxQU7fkMxs5vnBc9mb6mjwCZzRTJqsUA/Ox/TvCLlUkGaHOY7/qz+78vZI4XQ
5hcslhzZqqt2KyHwr0yhoY2Ui+GxXSvI4Hr7S7oEG35nGqTQaTEDwN7nZ1yRUyvk
OaXteflmE7dqeP8fed8WaZSs8qZ0F5Bb+Bqmt3q6fL6BglPPFqiXcaq1yZmA51l5
G3amUqTAM+Wc4EBeWkW+X3ytxNwCoxg96D4kBbzlTkK7SAGZQr79klxqr7N1eRaW
0eewLsUSYNwWt+f2Ry5x0Mgj33U0qz9cLxb2o8oiT/v+n8o1XMmODvPF9qcSVH7W
LkR+ZOvO8ytcKEtccRF+2rQBWmfjE4Hxq96pui2epHgFiYFbaRZ3FhFr85Pb29NG
yffUcmoPtIy15CJawBjRTBQ6QWrPjZLMAw5ZlECb2vwMg6OMXsIsf7ce8LyStnoL
XkSBlqpnxQqNryGCJMKcaBXjtRxWnBd/birsinEko5loXsxNkbhmttsfybtOHXlZ
1vgOL8HS67+KrDodFbR9dCVTM4nY6Lg/uwV91KmxgJCdNncmXXSaeCOV/DPbbQDy
LgkzHyR3OtmjidtAAg+mcZmpKO/Nf76CRGakwVfH23Tka18mEJPW+GaknWasAhCH
mBLqyU2ZnpIAig8EVQZ1uDGBtnfBoPcF+DJqcv3qoKs5EwG/mk+8WvNCtYykAksa
wYMszXtpiWPVeSYvDq3qFTNNfyiY/B0XNpqk/EevVFVP2ceDqIUrRnGc/uCuTGoo
wlkQluais8wIIF+0zC1g3u6VCd4x93xM191ne2nfg69OLu7Ec7G8p6+NoF2p7RKe
SFrcDQX03FD2hP30RI319dZhe5O3tu84PLv40LPDc6e5bXl0k1r89Ms22AyeE3gj
2k8EtxpWWcvfCh5hv6UMKGT7JYOtt0/qGe2+FuCFgUPZEtOr/VstSrUkwRq6esEO
kF54b+LJu3Tkx4/xY0hG3zdwdACSiu9Vmns1LWsPQEqxKYxKBefiN0ybvzkHJ76W
XeIEf+Y/+bhivl8GTeeZuUGfgYWRYWyAihbgf8tfRKoUsRCBf+CHaG6HfqChN0WO
9QW2Jvx6jR0dztsuvuRhYEdYq3v0S+wqxqSdQHORfAtFB8+OuaUkUDs/oQ4uYlbW
SV+At70wWAPCh/fzVtoNA1acYv1Vrf7Q4VBS3rR5cU/hPhx5k0M6FHarlQiGvDJB
dYX4vH5Mm+NRaxtq9s1EAqwtpLc1b/5Bt9T8IOk66kcRTCZPLBq3gpqP1tkkTaUC
P/9sN/IgZdLd0dID9+g+ii3shHWL/3r80n1fkhGLI8ISN+KDZGQsX2QpNLCuL034
OjE++sB4HbDxVCNEfnWIZTNMuit163tcwnwsMqFCgFSwmqtyqPZngHpNtxHa/uWk
fdBJmix1EilPxlvurhb07qk+n1c4lXU0I0ljQoaSXAzodxkQq04i77ixD7qa8Un2
Xdf34cuuXjAtdiQ4bcUuzFmWK6ZuFghtB1BznloD/wNp9IMKdgVkdHJ19KSvtko/
5v5svwB20TDxs7LeuRxirl4QppTAY2qX16K8MRWHwJgR0RsXdM4y3MlHlbwxlaqH
QRN/CBwcBaaDUEzEA2jqbPuy71XWEwysj4DH92GL0JguxByHdjjH+ZyUdK5wzSYc
OdmwGu68tj2Rj9vwjtfxglXaJrqqXyZo8Its88cYWURl2yNT2M+U4uiInnruL5Ej
zTQWR4HlF8OJW2w7WbewWVnH7SasNcgQ2PtTzV9bAMNDCSA7j0rRioGcJB24ttz+
x2pHglvzVEYMPcLO7oIY50YTCuxhkn3IIbzoapHibnzYnsrA91GSv+rcDWnqCR2Z
zR213zFu9ux591tP8tCNecUPqxZYe3RM8blNWsY3E/7gfIFzFa0CG7XDNkoRd5jI
mPvWXDDukdsvDtaiakt1qx+Vl8EBNYePGajdOImZnBoJO3W4xvXWxK8lVUpoU9Ci
4sOcduiuhIBHiW4V6QkKwDc5ikGUhIZlXm2bbsYriDU66/jrxymNY9hpWo8ots4x
OmTToO6xjsBiJj5LveRt6LclerZ7gqT6ycizZAJVnMQ2d8BZ35BbfF/5Vwoy1fom
D7IXTj2QLVXAlPH6LVB8OrOziCMftxufLNgX46QivO5OQqWKDlgw5k+VS9S1bKzL
Om/MB3CPzoyivFmscQEhCuFGaEZL79ytwcGdL3o54+moUZ1kApDx571z4Tq5ZXgU
SSQQehxYzvb06ysPn7xGJY22OY3g15seV9h8zKr1mGcnsJemubTe1XQtv766tKIF
v3itX4KfKByjxuHNBk2dScgWW1KSsfPuz8eE6CcOEN93zzW5rtsmZ2kauz0afa//
9xrgnryeWxo/cCF1WDb//tOm4bPsM/RgMzF5yUr1UW8y0mFLctgl6n3GRqsLzSkZ
jU0RxVERyY3NjR9D08LnWjXW3QNekeT0Fw4/uph9ygKIn66oAllq7lM7IF8oUUz8
NH71dCScFW0A4U4ct5Ly/u8MDdDLLCbO2F6L9kY4r7VVMh4jX8M/nHGLkrxDPJqk
hlLehVRbeTL55O76oISPikR6zpedIe6XBNWhedMsozpHlsNYoaL9qXIyD3zXUOMz
/d4iq492QhIqOhg6w3Fz9TyB7g6HU+no9VOdoeDFLo2ph9Y8a21MWfMXsvqBNW16
bfuWev3vTJ1JwOmZeTW+uQdDIOhFYkjGM3W48J26Fsw/Hbe8vSJzdH97tPSeRAb6
DF1lo2o2OacKpuFDmT4jNB+M+cRKK7pUDdF4CNoJsP6w1jCwE+6usj0T58dfXCcG
aYq3fY9RzYOka0Ln4DfJGy4daWSzGWUEvZkMQFaHvkDdY7RP+oyxzae/dEZmV9wS
n3cumqX/hz9Wk54l+pWs/yGQKEQ4DDnY5/Mo2mVUiOf7ZBMv4zHsaa38jzwBkXAc
vsIimLA4D6rEJRKP+JKQbr6LVQu0Mc17NJLK5cxLvGs9lDgdXxwV/i/UjuPj5q4N
Pf73cef3vkYKHsaJJ3Sgylbl/3kBIZmRsNeMH2rCX0jV0XRYquAGpqzCMnGhuDdt
HAh99oF+FdF9x8HM9y8RTLhoq7bn4pY/lGwRsXOwyndBuGfYc77C6HL1c0zejb32
DsNuHUc9/TTzPE5UFhqOXG8gSax0dAMBaz4XdZGuO3WS91BOEw89AEq8JgSjScf9
VLsE0eZ5xHxyZlfVir1zZKKR+NpVXXPL0zQ2noT2myoVgLLn5RsK3k6+BaOhfiXm
e2s5yLkq4n3Y65DplXFpvknwsQz7BE3ZA49gAMkPZE6Uw2KlDcBAjQn/qzke0xsF
3SWmIiTJHTfb7KqGy8vCWktHbWGLnTGdy9q8jWopYUWLmXO8vzqzYlh1ulf/ETEt
ZfZG76b81H3bdhqhe9u6nbGLQOFLC74zuzXV3w0FynxV/pzC+fcrAAQc8fmtrhZI
QsCAZKV2DetLKAw+VVEInWI8v6fkmdKdMfGWzUPMnXRd5BP6VNV1Btn4lYeVGriI
sNVgsnPa18eLLXEPrErcVscUMXuj4oo95VvrRq/SXoEa9pWxxb/Ro6WWFA787PXK
x+/ziARLUAghtCvqyV2KLp8wy+QGBRNDZPIceQrzMXcGDu+g0zV38sdzrZgztsP0
3de4fPIeHDmDtI1MU/oTYGSPQyhlPvOcu8/PVz3EA6bhZADdihApt5LkvFfaKjrm
Ecc2TGRZ+atn9dhXu3kSwWfE/7phuwIiGzianYWMkGVdxFiagUxaOHdx+4XQ/bd3
5OT5TOCx0In7stafwrE3VT0LGdwBchCs4f4lDblqqqBjNJ9G4qc85rC8PCv5HlhI
TqIaaNPAuEL+kWqrIeFtanJNVg5Ww+idyKDMB+vf5M6gV1HFNj/vY6md+Xb3Wkn4
uYH2nayjmcZPb1FsOxpQBangYcwAzMcqlAb/3/FgrRIOyrKWSV163Iu7vWzwmqFw
lIoiPsH7sZxO7cEX4In7u7NJo9kKHidrr/ommzbHq6wVKiiQQN3pQB0SdXzY4OxL
DT+eQ9Iv3Z7fOXiR3jJb4fKNY5xwjDVAnhPsX62wVgltvATjLp9dZc0dyFMizn7y
W5zEqF3au1EAllRym0u/jboX13VbRlTNH7Cl5E3VfAzX+GjBkA9Vxe4aokbVpLDh
1K59x2p1xItcAs0FvTY2GPyFHTOhgScOUxdih88P/wfq5Jl53Wy4y6v18mlXd3La
cUwUELxBkDC6cTNItoCYi2z09WAQ2XY6mt945t29JxvcqcUlDxpEIAFkXwB0H6iY
dx5wI0tsqIi1FZd1kvZG5wI9sSXO8579vXdtreIoPlrJdxYSwz+Hkh3Dkow1UlnF
0ZtV5lu31NCjOIWmHMB2d85pemG1TeOqQaWQ+uoI4Er7Zi8gFveTmZorDvDX5HvU
22F95TSEgY9Y2/80iqjMl8Zd2Z0M0VZBjKgsmA3hKt8TrUjwdEXRCwh3pCmK21RT
9AerNzN8a5EmT8S/8Eq5CdMDFx+GkAnlg+2CXWBUlm+t9roLJB1u74XnRMbmMf4E
C9YSxaBIaOeG3j5vsprLsDv2lTyEu0or45S1+Y2ux1g5prDKnlwYlBeUZFd08oUR
s2F/V5Z6dXys5Nr4YGXXuCS3/Yk0NxsFcnqgkAq+FXh82DYTBKI0ZXVXPt6mjmbj
iP5Pl3BWbLv1LO9WQ3GvUpQncWaBlVobVHGq1VViUiFR2C4MdFj7sz5uhR9Hlv0n
uuPGqHklRaqM/zanfDDp6NLBAnPnJK6SCpYZY2Tr3ILOzlKqz8uroB+7e4abogxI
s8EPgcTOdVB2bpXSfJ5xqJ6W0UleKwE9xgx+anK3a0OHExd55vgSs/iUTlWANuly
eKwUstayznxLcYjT2Iq83mPgShah6meDP1Fm+G5/wKrBwSYLiHFMHKQMa1tp+rE9
LrrlP+TFQmz9hDWpVSQBuJLbArHHHD1b8BWok6gyXlhznPL1nehJIStYHonskH6W
wzJ4GmaKPynJqXNwj+QsTNbYCUvlhynDu1g7mY9IQ5X4hiWQpVDHtHJ2iGJG8Gao
1LCQVManC5myK9ncE+HLvLVm5WJ3CDlMlVHs2CHEEOe5jcyM9qS/BlVc1t+PhM0c
ZWka7lCEZRAe8q6krxtG/cj450mnXuwTilw/XfglN3Tg6kcxOzTmA7prn0Viwg0v
wKTPjBTp5Rlv6FduoMt9UWluY2vtp38PS55WkzQKJaiSWVhzvrysupZMpjIfM181
uUBdqTNpKXCXji47ipBBePHD408GMWTPF/3IKJbRy6T2IfR8P9aP/HQuYvij/x7Z
fAqHC5jhVnE+J4jQbrIogr4A2bNVfUpmEGbcLW2NZhmicfgzJepiqR9uklCtqvMT
NPXd76vXMWPPg91vH4sUZevC+FQ8lcmky24iEgej9HcwXhifEL8XYVm1dqnHt0B3
DSihtqS6ElSaGEkLsluf1f8sfP2aEXfjJF+s2amSH97wWx+uF6qqHu/qIH4zWG7l
DMCy5Rlr7LqkOmoFWmcKGmICRHAh+JTsbm0r+MoDDHmxDsvRyYlFXC9GTCUC0ybM
g6w+BF8g97wo7BFCf+QHmbyrJuHxrSo9BcVwm/WLHenxqA3j3P1RlzZogpcQI4lN
lQin2SlwI0G7QSwBurBeJbeCtKz6ULOxnp7ivR229mif2pfDxUnq+3XT7MG7rbRB
3giJIkBmsw9as0b1ab7wpuPFsWY9mrUejToPsdvy6YyswK8ydahqEign+LGf0s+5
M6C6ke9NFPwmCeKxb+bVj4wpStxdqvtNUQkI8vML8KzYd4Lz2vFg3guyIFfjf9hI
k2X0zkYVynrezkYAtv9rB4ih1QzYO9wA47fxFnUBWQNajIhO593HBMvqT3RwS/F/
CW+4I8xfPdZn4Mj7JE21k0AKqPvJlXagw9eZb89mXv+kDFNZrvF3ByAzvQPcBVkv
Os+h7OqujUJBbdaKsooHoecC2OzKWTnI2S8eFptaC3KcabGllf/9ndilgTS63LLU
bBmkZf1B6jn2iVkcBMkWaIyQQEGvBCO3pwlK91+ritOaNN+2Jp9g6F+OVfVaXhMb
/0wjsT+2TDD5c8j854vBga/aTk6SUwPbaMq+1h1Z/TrK2N/Q2LVx6AlSG67q0iaf
pdKVk8Y6PkyDwW72NubGn/wUJnLKmEHeAx3fPZoa8XVC1x94J+Z1eoz54iuKOdQe
2nI6HoO3QvbmEqJSXupYcb9upWNGnskAOE4ZZdqgR1cATwApeLhMHIwkpITloiGZ
CdGsHgMKFT1Lux7OlhDiE+7jI5EngDgybR1/18aTRN0q4CqCsiay2DdfWied/Ve8
Nr9KXAqSaiY0Xo9aGjmNjrPpdu5mYC33lGM9Mdi/FHcrVZKriLKxdsyr0UpAU3eU
Zmn0yI3o9DkrRqsaQXGvCoGAbVmna2o3UZi1vKmeSe2l+wIvmKgxo5DxymKOXSy7
3+/UNWiTxK21Y4rN2V+lvml19a1hs9Q4ygVp4/hzcB6k7aW2S146efCxMvQTlufQ
K8m8hzrhVtUPwGwamKrlWIosfJNTz6mLr/JjQsoiJrmJR92CT8mBHA1B9mThM9M5
/s0vUb1uYfvj0HhzVEd5ZFmT228LChK6X4NyBzgD3Zm/Rb8cFLYxivoAUbcuPmcA
4HIEvvSEC/40gjB70yxs/keMcHsw72lAu4lR5p6tENnu0Io6XB7CMTDfD08OOTyh
7IVPa/XhucUMnMfdEw+E9UrVrV5xTkXz/OryNOmpJ9OdJnvaA4MAli8sBPQI59PG
nE4QB6UqGAxuYG7/2YegBFmD2lVcxY3dJe2rWxBG8/WpZlUuvVIrfayifDuBV6/i
TqsjyYfZA2z2ch2aSjiawov0mcWxEbeSkeVCnxmJILccf3E2+YcAG6hTIOggvmYu
GFq1QXQoDzfGullmGX8ljYQC4EWnA+ujPnboJ3X4ZCUWs50cT0Lsc2UowjtZ/D/z
5Xibmu4GR9vm0fLew0XZd/I/jXB1Ao+dBi4DGisDXFzVhhzgrha53loM7SZRIYGs
qaNM4f41vtqRcl5L5P9l2uc9OtcexY1kfE5MZnu++VUTc132jIntrkBrgvz9VK3i
drZR8cVBT/ozXz/i5vF5AJL+j0BmZ0EVUqeRLDrUBeaLpFkjt6Yl3+QDdj4n6r1n
leI0Hhf/xJCawiE0bFT3sUx26W8Yad0ZK8OwQOM+CCyiFdicciUC90wKyNYG1BbE
r7EFwmUEyc2Ut1uJZd+1YWU0NIcLj9X8P4eUow1wCA9DdemDuWubbbl972yYduHd
QRl0V2DsZcXrrKhyfMZYU3Orev0Oifakpo1/eGSujb09qoWXj9jncfmxH0mw8OBz
L2XhPR7sVBlH/O7GVeOPj9wTb2ZPsZjv6j63p4Dxw4mtIR3K1fH18c8HhkRujqgD
leKAagDUBSfWhyUa7+aYaFa8LcW58zx+j76hvStInPSAoeQS6w1mvPFnmfHwDlW1
X5e9i3Wu0HJ03H4RW9OW6nbu9R3heRxLz2C1RQURlePHXDhG2FYmpgipC1tA0nkz
JdO10KFyWICIksBs+rrUg+OTAjmamAoKmvEOkDSPbVXjLXH2ubkLqptKVMNRM5g7
F44ac1DYsqYo8FUlE2oKICzk2w5F7POuiu8Zm8Q6NSi3FRBaBO5FXHwLIeXRKnhD
EU35NW82OgutWtlNH4lfeRg+WpDZ18JNRa00b/zlgVHghTcejkJvtIDd/4xyfbHl
APrODwL3KF1i9aYFIOaEktbdXYHmUZZwL1es/OaiSHcRjhqHBa1CjqfkwCwtC4B5
KJCu5Bj6mCbPj575TQUQzu8whbX4ZZVZANgzYasex9yGcdn+CWnvzGtyyvzkO+m/
yLzLQNT72jNnpUm3flFNGbqjKOXJ3kdpgvhp0AdL3NyYUOOox56EcyjchK80LThb
Ozt1TxNPMPT3xTy8JESx7DC1yg+QuNMRowUZpLUsT7PYB8IITr1ILvkqzsUDcv9B
8SOMRNQFdnFMUgl81NRmv/MhSdEHY9GDtcVUEDCZt2mnBeR385p2R3NJwdIFu2KB
Bv6kLc5eV25NlWAfSXuh5V9VUbmrfjD5gQI36MKY4E1dhx0Gv+5BUHOGjBQgqXWD
7Lh/vyf6fLa3HIX6LVgLltxXa9HOqWIlmtPyeU5j+gM5U9HXfjIcno25ImdjD7lF
uRP4mnuZoMGYmlW13m9l8CyzumB+cjSZdDg7zAP3Z/MI4sfZkeyHR0XjLApqvc2S
4QUI/mj0HgOJ6QzcHUT8XE1NR2XZJ62FSHyvLmbgqy/NEsIhiyNOjZ+kEWMXr6Ub
A/VDdJlwKXFfGaPL5FLAISCWXqij+JNs/wT7fII44abMywSpUHNGasR8yDovY9Qv
wPE/AEff0sbhmihAbNkvc0ga6N+r0d/cFsH0EbHv7odTQayduaRp2ngSo5g80FfF
L+myJ61R8zv8FGEU6yq3iwDYnAB27eZv/cRMRADKv8ceRaF5oxSC/AADOzINftUB
HqkHuWcwDAkpWpRnIw8/LQRCg4DxW2CP+6hYR4udQ749jWA0jL6ingJ5O73vrfHN
ZhI95NVA7J0u6Z1P5wwZmmBflNCH/7uY/b4ukS+e3RHC5nJ7lnoA4gi8erOwX8Co
RZQnBin8IiIa7D9UsOXJNRBpp7tCtCGWnZf8vrADZrQ9f0mHzCZXvqPAoLhqwTmX
uirN/A8c8JpKqtXZVbCSXLV1BnumCo5k1iIx2V0QmHlNsr86J5G4APsmRU52yyXV
lgeHwrRNRCbHD57FKMH8KOngp5knA9sG6d7CmqC2UwEijnfek6gwYLvCcq6zU+Wz
BEoQsxcZwCZFzGuVqHzwu2EvGuK3PlAC4iw+ruoBHah71NZb0jQLlE/Ayv78J+Zr
p1+sy3p9lTIHVPOB5301FNGOkTGl3PyQOikMo6pqn4iqxH5O0qDUQlYmP0b3nUyJ
cLazbv9bOgo/QvAofiDLVQkhDn20TKOoFynUXARRV0eZwRI71Ik5Z0ErAbCXeiFx
mjlcDrEQj5+rT/Yc6fUjtxCEqgF22YyLGKSvwEtcTuJqjvpjTqr/ywOEyIqJRhEC
jRRMF6QNTXLsZ6eR4PVUDvut+GndZDzk9K+0gzQOMQ+MRoJbvo0uchfmDXefGA1X
7sZykiLy/jk5xW2Tg+8NhZPi95YPUezdIlbChOuxxbLKZ/t3gC7xBLQwm6UgSUKl
fAMk/24RM8LjPHbGH/daFJ6Owg93pd42XY+hNxO/D2ECXxSqWDbkr1g40l/Ld8m8
RkwFbKe7MeIZiHiGVXnSSmgVNE9e2kCXjplNHugznbdF9/sgrcEMRTmPv/9bBv/l
5F7yZbMGaSS7A7WfXzYPdGi9ENZkwQx2emvfnIZWiXuT0u3zj5HtW9Bm2rF8yfYb
7wG72kEz2kdVY+1WZv2xN4dClfbdrDQ0zDOngXlvjZZGq8aPreIVxRb3yFZ5H7E3
EBlDvcj2is8dip9dvB83t8VIyf9XE2wISMmCNIq0pY+xEdVk7QQMD4PSOOh8Grfs
m9P0NmDckS/Gseh6YSp35JiBHHpXpJEzhbyPMlYfUa+Bdyx8zx0g+Oh/+QJL0faI
rC4XjoR1YtJXjITxkUoBw7BGwYbzO2hpKAVUDNcUjEZsIrYRF5lPnWPt0IF5Tow9
CaPqS57cIU1UFSbbzjZv6eMVnGG8ZC1YyaHdKqkJlNumRrxrZzTwvRh/IR9PnVkR
J3ald358BsNH8S4E3fh2hHV/EEcSJiqCo/JSDNrbaiCGxwCKN3lLtlwN0FWt6SVt
ZoBIzOEnuxmrqeFm3nRWz+rFtCdksBx4czhANFFJLMZd17NAQoNbQLfnDlZRnw6a
cIXxWPOs/7vEo69weiDlosgybuN9uOpexQ+c8AFCCNlImnEmqM0AtDlfGDLvOTkZ
VYgnGO09XfsmpqLQdxm79lhF5iBJxIUxj7N4p0K6yXUzp56WcDrx7p1AXL5Y8K53
jUTmaJY++dUxo+K7cm3lNcwIzBkfV5Z4xMySqOdY1wxwH3ThpXcWa9T3OcHlpD3R
5PuR46WbN3slQqzkSRZzdsmV7BK3XcnycJ/eH5R7ea9rMBnz8IyVaBew9G/upGet
I9eGXD/lgxlaNbZKurVMJSMCEfhI5LTyOEnZFeUqj3SZZDBA11Ftjt0zYGWJbeK7
OXzz0ukXTYUNv4G9cb6T00ocGdPN1L7OgviUQbtvHRJzRM5Ph+33SUspNLF7fNkS
TMfC3G7M+gaE66Qnuu8xtfx49sxkm9qXHz9trYyd7GaSlnO4YciwdJOKTC3PMs2d
Mtlf90hx6O/RqStJiFUwN9xKa9Sbw69ViDkB8QDTcnMpwbaYapW+WmeH6GdHEMd4
RydzzJMYzgJeruoPsHs31KVk620ZnFKtCuaeooG2L7lS8SYeMKgRqoVOr3grj8nQ
cY9BxhWM1CNjBSPna2oeVjTwenqtpfqwt0lfuxPKpOfG9KJkYs6cN4pOzEu5/q9K
Qycix7zGiscR8zJydoZwGTWyUwochY/4ZKPATqYtADaJ4ey1xs2npXNSbs0JeIGx
2n0ahkkHhsGi9Mfvx9nppcOxRk8/6jWMz5r8ttJf2BOPwQnb0svDYtVReOFzHcxF
Y+bJKKJ6rak684BwLKiWTU+HGiNY4lCuvhnzbQLSoMCc7NesPbPpHGCxCxF7JuRe
9GmEdMyk6Z2Z/hShpaL3r2jN9aIaZXbdE6jnR+sSlyZRomKtctgxpIDVEwxizLjT
JSSrZqn9ySLLkv1fyb0cHheKCgLah8xS9gYMsp0LOHEQbfhzibSZ1TR4rMIMgEn3
H94CCUxNYZmGHwzVvIz5dYDrm3sEqQEmslsSlsG8KiIioAN96RZxLOm6WKhyvHZB
3T3gZRBtKXbtrzY1ghja3mlKXNKLZ5aFftEMoI/qwd86f7MknRzHICSXPt0MPMV7
UXAIDPPJ7MFhm4eLtw0GubNCxEg8NIdNZSW8gij9W8VvK8BDI04NiK8XhKtdhGyC
fNKlR1rFksSqrSe8Mmkz+OYicTOD0DwlaSHm7a9TNOxFDBcu9cIos99QImpVALy8
LuDMdCpFFF8/xJNRCT5zC/qsOZVZV/ysxjjZUnau+Nc2PNNzZuzW3OElOrhPktxD
oWaY8QsOimqdME7WZOcpSiAmIJe8ltsQd4l29qwL4jCD4cHwAgYU5vl1V1v/yOSs
YlxJqQx+OAvjIL6ouSG+dJioVGWoxDeTPafolqI7ZK9OlnNRZMp7QvOIuuCGHG+2
RpW3x4f+OPh7zFHY55p42/Zil61VCeiLUEw9f9H8CmiZNpYNJxERWUDxLLFm/HvQ
04aS0T8nxPo4spFcpR2J3xWicsIkhxNgsgo0aJECjoLQSby+6ufyLU4JJ6NXIaCc
6tXjlp00WmceKbqtnuhnnmWzNwROlUhjv+Uh6MqtF7ip2RUViOb7CJHexNqcwe7a
R2FJE+UdUsZaV5iKxlMl/MzIZA75B4mDrs+/6ATWH/x7CwoOFpQ34fFER3u5KKSq
0CCdq9+aVMtL5tUkS19MfWvNU26skDTIrtCUVWcai8QNo7hmfxKnnJvciU2cTcw8
nnsaEJjIUUzhcpNJzV+pg6iLLGQ5Ho3C2Nl3rJIonTD7KoT3G/SUI0cqpoV0Y4/s
FrJUAjq+jFAdMpmVPPh6gk9a/I01+e7V3SHLW//kBgLdnO1Q2O5uBXorCn/g6o7E
8WC2vFYvn/GMeOjr2oWc7gjorSh+dIfiEb0xVd+vv3J+mGbVDJs/4do+G/eWvxlC
lWyh4nFzb/XPRMmmkiifSfd+RPTKXHLBmIYVZvS6uNfHEBfwr8ypdPc4g7zciY2w
ZEK4Tx8wpoA2JVhTnonCf2G5sMDU1R3CqQoLLPkXfsTI1lszcpbgXaM6PduXr++G
CgV7Ne52raM18leL16aEdAiG6n29VlY+f3vaIJGX78NhoTztzQVDxZHB+VCSUPfx
wNGuvxVQL6uP0BbghBnKHgL2rFauqKxY7YoKKCotKhl55r6sPZvAJ6dK5oLTl+TK
i7OO4cum4Ia2OlOLikMTWZZMUhSNjGDuoqUwGXbUtxSV5pYZTZsg0qWcPRucI7lD
ZT1DyONU/zmXTenBEncMLIKeQJ9hlf41v/3FxwDQ8OYGzY9RqMTJ4xt0grUAVItB
Aspqobj4lYCW2FmhH9JlLdhtXhCffXi8avLNgk1WDpWNomORMSYkBsIlp0YQyHbR
hUJi1BbEduQau2KEUK0/4oZdKTY8Ze/URJJq5ppJG98WG5/KxDC8G6gPOz5BV8ts
lmt2bmofXgEEDd8P2ZcJeO36g7RI81nqhbBVr3lsbGFObOmmTf2Exu16grOFA4Xb
p7RgztF0YPTLbsjnKAZIDzzdB1KrlF5pJSsFMAl+JlhPuEDCa2fGQ1+7jx1W2gGx
lqa1cuG/sAyIqovXCTDdxySWy6NigGhnoCBmDW7mdThxJqVV/qGdTURdhBvS+OPR
Er1x1TdOdeLRf5WyIfIbe5jI5b67LFZ0RRl4bN3BvIbC0Di/vTTAOQwjD6Y1up3P
23cXpNEA/du9wlcI/09qv2q3E8lX/0oKAqkt9sQcqwg4puxHtlUipEI0wbaTFe3+
pqY1Wn4QW1sDnSwshFIEQZpKxXyU6tW2Gj5aNQ0bHFafNliBTiw5JvBr1/su355e
A/6JLuNWFR54uVgcHBrPGbZubwYIZX/bbn9KA5rMDLfyhEjO1yxTjvuU7Y+lJPjJ
SCn0eh5JvZezk/IXhdc4URJd5KYrNMStKvXWMVNaLXGaKHhhQOID4YagFa8QvwSi
zJ5FYVHnwAEm/1m0xDA1ix76p+NBh7D8jrL+tpeEn1psTtLwF4vPmQwb0DrSYeQw
QFCDAK055jcNThWTah471KTDBTWr638maOfd1lrDHmf5sReZVor029bBRu1Ey68j
Whja0m0ZMdYXQJPU16m9Z1GhuX7jE+JcwBfuqc4A4SF1sBV4HF82Hk2gipjwUMIS
k+aVWKpe+x7xRHKm64BSLQSJXhCVosLNgfTux3pK1LsWHHXe16taTqh2mksopcD8
acvqYgZXJ+hPYYuNEopgo+wWVJBGJ6VN0QFPyirrJkN3agjE/HKuIWziEmFKtXQz
OhsJGnj/ymnyMKClLw1Q4LX8fCjHqDvdUI6pZ+TWus3XiLRGe1gHFByrq3G/2Rns
oIMy3gmocUf4ChyZSN4H0AgtqE7lvLcl2rLtVkKZ6/rcgDP+0I0igIUQKu76RYtE
6fcTVvgBQWjzorIMJTJpV7Utp/lPymJ8MONH4ocyJKR8E8Y32FA7v0Rf/HYWB9OV
vnriGMs8gkXyYU1ot+VkZdbtBYhXzsALhcCnUeSQZfjatjEXuE7LtmnKT7XlA0+6
26NuFBEmlfC0hnWKNkdjLLHNHvoj+CfWm75u6Qxg201tBO++Qdc/OWQiVOZ3z9mG
cfQclgllYugUiqiNZXs7mTT8bDO+jmvwkuKbeaz+tz1zuRjUH0VQzR5Yhrmj5hNL
c7NDfebN/PV4+FyeTEZpxRLhYVJf+hep/fhJO2qRNp3hf6w4qDh4FHzmY0C0Xqr/
eE8BTGmkweTgqGAHf5y4OComMjULS8fvQcJYvXHs9INzr9F2h5wAPnPTOzqNH5HB
DCmyfsS6UhTa4HC+oxqCWK1DT5qOf4M9TVoKvAHkE48bS/S2fwoEupqnvDexk/Fh
Dhm/ehra+ZuPf1c3Zztm3AJsaV9Zd+EPcqNLmkvHfCDTO/ZZPWkMdENWkre/nG8c
r/HrAkrKzB8ZEtBi0yoGq54FjmIes9P+em+JTQui0jkJv585aGM7dIdANBSKNw+I
lIFAjgdSAvXLES/XZWtzekqG8Qc4+I0ldseTugvsh0Zq8m4MRNLa8nly4BORIvrt
6jUWInW6V3T/D7C0rUYQSJyf3mHZj+FF4+cV58HJbSa/8JQPwqoXXIaJrYQqDguY
h5Rmw4tHhDiDzVwh/yTY3awU9WKHYa44R/6Maor3aAwU3K6gqFCs2br0FzOupzlu
xx569KMfPegl078KBNmU7+op+q8O8IUrPuxMdizn0+MZpJnA3z2xdJhbmVsp7Fbs
fRddHp+kQtyMIeoX4lB32qc8UGbJSGOvn9gUIGPZqSicO25/UnSdriAJkDCmBIi/
30//C9G4/r1c65M5/HoNgSgttnvu+kICDdVj2bB1HlGzqtIQNKRZbJwV1qtHnwqu
5T8Q3UTxShtV8NirWXLaodWdTV9fB+DF/SQVBF4tZS0kY0FEOWkXIL8VHYWnAApc
5CQswozeZDnLvG/7V56gt+bp0nmbmxqJlV9Jypenkx2rvYrkqKBKbkmThkzSKugV
AGoZT5VA1jZK5KHUrA4Y4D32JxFT0jJ39UPvR7oDrh+NluaHXB711L6rPSwyuB6L
wbYI4fWsDKlg9VOaP4Rnl/fRV5Y7eI0PENgcchVzU1krV+kFa1Ky81avJqj8wKwZ
CzVRb6qd5bHgkS6oVVjBlhJOPQQk9rfvI7GSk4H4uTJZLibapFLf020XCGVf6/o4
R6y7OpzBlJkflz9LFfHdL/sxs0ZBs7p6SZSpkmSvn56s9vJ1g4os5Yjj9H4XXJb/
syENaBgKsVe6F+l2Wk1Y5essLUUrXG/FRCF6SEQ5ExlH4STTCDzIc5oC9NtxLFK5
XvM0184+lb674YzqxgwpTxl723G4J//htDKUpWagpbS4A8OUeyuhTw8eQKMIqE1U
MEJ/C2623sPRRX5IY9wtg0ztO79GD6C1x7O24YtX22Zbo3CDh1WNxp+fKZQ6bwlT
+kpG7fh2yYUGfVlRI3IbXKVN6SFR2VDItuKYGeSvmzVJNHMHdz63tMEy2wo9LYd5
eiVS1K/vHETtF4lGZXXTuRZECZah5v4G1phjU4pToIrzkaNVLediLicXbp1IE+ep
ym7FVkiXLUMYNQiMAVObUJrQrCp7ii5jV500MQRPuux/HQnQLOUL0kJOea5XSsSL
6lVHdKqulMHYkgTQjLrNpWAkpU1BCuyNreEhGsUL9p2wXPXboUbps6L5DS5EBW4C
sTopEEzAsiWRCIpvOSuBtQ8TvmJ98DvgDf0sfWB9idkyJx0YB1bgpAoKOKS5AY6+
bh3J13EMZH6t2hIO1/LTA2TCvrqHL7g34sRof4IgFtBjITChAShwSyUccGEzFLZ0
jPHIAJLmKAr7otpXU2qdrrSISyIpv3yNiIQ2eki96tEv3hVpgeh4KVRVDBs1s3QH
jH1gvKELP44g/1wqVrjbRvYWZse1JZ6VKtKJQnyurLkDNas4mCMlTu9eX85Mv6UG
qCn7tt0NTPHjGnNL1TRX9MKom71qtvmCVgFLY8F88rpcGmH/ywwCdy9/1ugSiX9H
hqDXi8BQR6Wk46YGbub6L0b3tk8Dh4/SdmgP3CocPrhv3XyJ7UTI172e1YZJdBMl
Tn6A1KKlzVbLLwXZpDgiSVnFXzj7nTe8RSpvlbDMa0p/We4UrdFgzawOf0OQiTfz
0ATY5m+9MUFEsaXhOid5rMh3sArpvTKSNdv+vbTLkop/GnW2sQQ7DLQrSjKDPVCa
uZj+HcHowUkuE8eRG9A/GIp/RuAIsYOhNB6cuMAkcOaLzfguA9jknRMiIYetuLAr
k2DhAhsPkroY8KeEfwPjqRA4bnoDCiEpxuenTD74SNT1BJdFtlLSV+AUu1FCznp4
ztcG2C5gyedMNt4KG4jz17p4Iey3hO6sNBOr8Uk06550lT+QkNLHJ9LO8+ZlUyTL
pozbHAp+wimHkNjLAhXWSkZzyQfUuKKepSDejXzcEG6S4pGnUX+b/DAA+i9sv6yZ
3jt3iPCZAyKdeE6Svr7rA2aJp9M8h+O1cmb+jMhrNWdxJ3oLgvFJDnmaCSh25IP1
gC9tYg1LHjtrFy4qI9js908QoTfMReYYUMAJ3p/G6W5oCJ4XY9ft9eGosDORXpj+
z7qVyFUjojDYrRfnZyQ0IuuVUrpw12P+4ivqueYqJTl6Q1SqSyQile6IDC/7rD/4
GcKqh24VAIe5vOBN8bg2fd2Fb7EcclatUeiyXvtIKoMaxQ7tGEkHqxFdQiEI0Td6
S9E6rAOCspXhk9NsveoqncRyaDWjPqIZbqXbjiLDh7uoJoBaV3yJdtAWpRNplGpP
lycTnpk7RDWiA223HnE43x3iJ9skG28WQ7X3yN4BJuOGryq/22UPVj59STJjUrOO
QYvqOeB+otHqduzugtqNcjFOsLluL09sgLMSOYXD3bO1Im07EEOpfylbbFdWgQIX
6PXHVE1qyVtZ4Bwxh9Av9SAlSXZpGCuedHIIW/P8Kak60fr60FWBUVuTMOnFVrlt
GXJf9PLXLbfAFdy+B9pTVBSpYpDy5YEyCdmpJcXlRSoj4IcxGNd5xInomuhjljwV
E72dkHl6hkbRSxkOJWpPoKq25DAsNcOLq4cBvGBskUS7LICTeqO/yC/10Epc1hQJ
BfGbOI055ABM5tCxM4dphNtZ0zdjZDmMn/r4YWbaKj2KIf8KWwo/an5yBE2Lhp9m
CFILCCdOQMvQidVZsvoRQR901jcnwZsJRsISlB6TpZfLOKshSnfFsgmr2CvA4+i4
qQYckXqxdKinx42UdMu0hz3p2lxE89ViZ1GjXIKP5Fha6HimZ6gl47YhOLoE3FXP
eEtEJfPGeL231UrD596GkT5Kav47SXuQgMER0HeBdZW6KEFaMF8bleJLS6uX1loO
LoGxFvBO5O4hoyE2CEGbXf1+eF30t0zATIygUK44+GKTtPZtpt1myR02k6HcKEax
iaiFgKsKjt/AGjoATwN/8ZiJ0t7lglS7IN8oOUYHcWOtOVEk8Gu+Ydk6/L3J4mV1
xbNLhzMvPVt1XelvTh/xqHzz3C8CZ8DnupBO5TiuRaos98yppw0Ht0/PSypri0wV
8Xgh0ve0zlX6P5v6B1StB5U2hBwpxxsgkwo0cRU6uMgJn9SWPnEfHA1hpDb1HIM4
Dcbk+IqaYIJl0jhsS6slZ0hA6QjbF0sIDuVEbh/4FD4edlfwhjHgsXOAQW/hFCjB
FgjzrzFxYfzWKGZzu5uSbr4bjF2MFvBxQhum79aVIJtq1NxZrg8idCJ30OPUCrmE
zVVvGK5fAXBRw8ThSxmJVE/ju2JYY3OchMGHgx6rCqVgAaNioAxahhRl4QvEh0rW
3FGrDL74q2NowbM32q6HWhjBcQiwv8SugsZaYcVmyFVetf8PY2qXkZP2PSn2YCZe
ErqKGf8vTRHhMsJ6POhC7TAxRCE/zbnmUxckvHBkKZbx/7I4H5W0DCr5xPT8cZWX
PM8hrsn74YMN3Z8IRLQIVpjovN4evWBq9PboZAYLA6BBQrYhLNiFgZR91fcK3WFT
rWIsAsEf2qbWHQ2I2Ybd5FlCloHc4kC+r2K6xr++0ByydAXO5y+x4XHpKkAHT8a6
rBMY/TYzdKIHObvx8KoS+Fb+4zmo27YIo8l1vtCs/AEB3GNZToU2EpokxSVwBZmu
gDNE5G2BACEyfPrY7PpvUzLYNkNb8yMMhSd5n+QlN4fhf0GiOKSGL5A6DDFIZIZN
/UIpRog7nMcV2gaHqHQUL9mN+ymmRvIP8nUsQPl+3qlkop7L0v+rA115U6/sVLjr
EOdI6UyX53cpqsZsww0rrKb+wIpPLJNB3XT4TLGCa7FuUecLrbmj5iFe9U4LGwfj
YBvxW5M61y3oUvCgg13qmFuE6yo1ctq1fRy8OHVFlUJcwEO6U82X6OKCG9pxuATa
SxuSUlhjVh3eE2n+g759zhdTkvPFShK7k6YlUHG1RPJGSwIk/UfEb3HYeEBIgYzb
96olpD2qKsmEwtc5K0/V4bTdaD9inNfeiipY1M5fohxELZUYct4Y9EidbxLj8MgL
yLEk+/49lnrFAR84z8dtLr+naLig4vThs3lc6OQ6qabRFtyd+c1+DoCz1neUIT8Q
/8mJzef4EoC+Rpmyb8zCXaEE8Bpy7PzeRGcEphHI6qUd7NY8wE6t5/lVkTkKYG6x
4XBVQBMioAR1J8QSwyOSDX+4oIzRSjFoxtUUrbiPphQc4+3gXSaIdndjLkX6axFo
yUvD3+BL2x0U2KDa8Em8CZq3y9VjzNLtW+l7lrkHCP76uBQUNEJJeCpaJhdPbTS9
Zct1TdM0dwEJWstkulywZ4/BIhAfV3alEhfGQbh0fwOjR0JpJKWpnnTG129NVWpJ
0P6Nng9ZhrWdbi7yHaXnoul1zbMfWMLruhvlLeA5+j166w+I4YKgd3jJXU7c8t2I
wWvl2YDJ6KxgtebaKZ8gZ+YPBF2zL1QGqvAWCoveHQhxXiWfS9D62UEOVFkakSu7
C+VmrR0x6GnvoT070dTNQyOtCYi00Z4FGQcVeKMaAwOtFVV2dqaWv4Ec1UvZCY5B
T3tUoMMwc49Jj0i0Kuqy6cu/YuSNxUjfjktsJRHFRgpLQJ7HwLkCtYU1RATPvFht
Qtz83YEHJp8JMFEVoB6567I6SURXc26CQO05p02dbGuTe3tJQs16S/YREUZ6dh+Z
wXo+4bvuG0D9oSvqJRU352V/klEdfT64XrIc5BWz1Qih6Y0t+R9rDb8co5IBJ4ux
49Lv2osFYZgD7tnavTrh+yEQjjzwkgOhBFLFdron/GgEt/QT3q8m7bG43GzXVMEn
4/2BzNvF/3jXkIDLdhONsgh429g/9gFuirC5YJWCWDkmL7UAz+DK1ZQnz8KASsov
su8o25bttaJeW2ZE6IMe6+ypxwifDywsDTR/GxXKdMwWE/+MBEY4fAUj1k3BlvU4
mfsGCuQlXq4Bl6Sfu3gttgYTN6zW7Od9I3pxxZm289RG5tfsL73y2S6YfHOYx6Qx
IiaPwNVEeV4qZe/BucggXE8EJERz7LX9ARLpzcZLSIZTuNcG9PESYHAlOg1za+OY
pXx9FvlfDuEJDSFJedJoODvfOTYLSH5rYoj+YxN9kVu1ZTefiToHMKATyfYMFTNf
rgw8SJwCBVtkFZXG3H/DS+qpg62OoDbuF2Jk1kOFHyOuzlH55sYH/BWfCqXDTTqE
4pUviUyN6SIkRlssrlXEY4YcLgHm2EOX7zHeajA8L+cfSGGUxRR2hFL9qiaxBf7F
TyhcenMi1jGsTUNzbTqW4rokSi4jB7e8gtlinguQDrjb/piltSCDw6w5s+vwyHr+
/VzhiDyhUdYS38qCV7keptemDpqaqMGAf3GrRZhIvh/dC98DX6fpKQBgccMUEuSP
Fq950qPt8MZGisPBW9P5z4kTYLPMFr37TsYvoTJT6ALh1aTF0gvF3pi+5TtYOZSt
4vuxWyB1RQHMB1G0GHsH2YDidnY4sAe9XeMeTBHMAg1JNkb37WcxEJ4Pp7biOQZN
IiS6Esr6Ho2za4LQaj0rI1NSXZrlrduLhuK3mDIpA/TXz4PxyJqSb+Xr4CnBznBJ
6tTgTAABjsqDWPn2eBzSxQQT1Ob+TFxuQVDXmRasHAuEWi8UPAlShhoKIgbq8+nD
gz8Vb9h0FT2MB1YX3O2jgCs/LS49EO6+nAQRFL68xKBMd7r0f9WsPwgKKHDvHKR2
Z2qRhV+iNJOa4cq4N7htmAjK+QQEVtSxqtWjZoaaeMgvOVDX6nn1M+ZdpJfudshN
RjvNybbl6EVLfxNuyuBASzsHXGrmn9tHPe1uHiE5FleMiS3TshaC4iSp275K0jw0
qrBMtTx1bQ2BeqRU0Fh6c+m3g8R1JPxtf0XaR3gohihxtfJyZW7jL6/zHkbe80bZ
dTCqm/DYRBz0tKo8Z3RYmNnCOQMY+HxUjljzUxSKV8SwSXoiFQ4pW/ak0dTCwzDB
nncV2wue6Pq25PQe+tZdWxDLppguV7qkImZbqFpT8XEXYgwww1IjxboVB9LxevLA
PfogYLZSysn5lMPEPHRLKA+9iZsL0jZGuz/ed42HRBMNkSSigzomajwZkZCTVLzW
Cbtuy0C02mjlPltpAVFdv+Uh3B5geN/WcXyp3OgjcFdZovDl4gaNCfUhaqZx7iBh
edPAkXwnYjrjCLf+FpjQW0dVoyAviRmqii83sWtBJ+D0lQTw3yvNC1GiqXOInz4z
sJQGMuQErm331D5RD52aVzpzoLO32vgr0IF8LAM5Qs+t2mrPh8E74ipIZu3f3v4n
PDQ56wAIkbUSIJeSNSgA068MdUk2z7jZhbeZ7vJTgloTL4ggTMs47jLLDEnNpiKG
3pz54U7I/Mr+k1DGak7GlW0AyRShz+2uOxUUejxfgwcxxZFZDPbMNnG5n2yqDTeM
+4id9yBPGNDXxcxWzzetGYlD7EPNfbBPTrEiwWB4SM2bRuoFVza2UgJYJ/JiBwyZ
ZB1sIPbgGovyAM8FDTl8EEp/MsloEe589Q5dauCVW3oUgEqWjonlswaHbzva1Pg9
URohb9re0prwmm71aodn7vjooiTcYBnKf7VhpFzpYYowKwbrNbIzKfn33O75QNax
KCPG/oOdbaiQr6KyqkyfSXhoDd06msBr0309rzyml3UFIzykMdmdprmE3SASzrRS
naTggv0rdxZPCAMwcgl03jGipNjMQQblnr2JDvXzRj1c2Hky29kwHcPtRV7Z5fRY
LtVJrI4Y1wDBGN7R8BEvG/R34qXOx03Vee34OdxepN4w9sudq0V9+gVw7Js+lkDz
pJwdNve/c+a54L6M6Pqn5h/YytkO7zuvVFi8E7jgkvnIhh/oLTcsYLIPypAtbigY
L83Isi8qz9XN0vhJicTE8REOhpykpYxHRtzj4qe3XBFfmj2W7LVDc3QLMUzou0eY
msYCKL7XBo7H60NHwu/W9hzubZqyAniVchgUFDBCbOdiB76wQTlhJiC3QCQr4Xyg
of26F61uYTd4pIzCoDrapOzGLSU6x0SlW5CpK5L6ZpPzWZK9r+02EYh6yo/I7Au5
1i99I/ehJr0UdCgaqmkkuzaYQkYWqihRmRi4Egse7NzULTfJAg5+fYghVDTIfUAC
//YUGt4dpOFAA3yVek+820KgBwEHeWc+ZAqmMgdUUwJcu4cIoRuRSRNB20tyuXQc
SmuFxnWssW6qGeG3wEVCs3hzSEaF6H+LfjOEEnG2esymcfcaDoDyrHgBSnM7RDh2
ni3TlQBbt5KymXsD59pFESjhvbevDaSKi052W8aJywpEq9XbRwxPL8U0oM8aSyDC
8QohCz3DQdaBwVqntkdN8maGag6sS3uX6MF5fXhjGeQG5ERVxJPfZA1EMgcK4UF3
4IoTJon14GdHfLDxXF/tLFAkO52aB9e54lRnEWVet1qrb0U5P1rROV/nCMhd5G+s
Qc2mhqo+WOrzDGAzml+ACNeY2OrwnWqL7gq0jOpTjfNJaPa9+sri7+4EOmjKHtCL
mysuzzrvPHE/uUeS2aXTVeJRLnWtB0ZlyzXaZXozLMGjuEf+gMGTZTzdzaSPz1QO
cey4g/ROBZklRf63r0ftkxkHt5xFeQ8OqH5DGpZZY53IYiOHJ59XwGPMeajrIU58
kvsM9qZuLNXyHjZ+4+hhRll9i5oo5MH8ARL2UX+4JwxwpeJrU7bF/fvW8GtUua5g
P93F94dp2I5yvT3CTvEf4bxYnJWeUCN3TRI8D5gEh9KUVvUij9TUmv3r1UQU8/wm
2i+f4otJHhcMyinkcnmuWNk8TbihIk0ftd2QwzDmmXM1SbdHkBjV9DMcjoWgM3JR
0iYjn+z2evslxIpIrrvJSHMiVJaaSiqKM/ZtbGN+La0HyNGCll2NxpjogoWtnTKI
Ou4epm965ZbuHKOY70fTBevc1D0jgFo0w7vvmjHVPjbx8TtEuNA/R+WsZtusYBcb
ZbyMx7Qs2ZB3+W9LIhv24X5D8rBhu6Qq7FWZwMo23P4u2xPdg3aS0RaqGv8QeSBd
LOh/kr9IzP3/WQopOmu3wwB100hEcaHtcUmweQAx2jbjSsEPz2nlxIlqLxPMVnnf
rujVQIueXG5PZlDoLG0gBFDQd0DtFuAQ2n5wWRbCPfkZh165mZ7WwIg8+lqH/ULw
SOAgTb+nEgnE8NhQrOvAFAizLI6huJ9dOuZYhFmKiO7hEONNfcUNPd1YxPFNoPaX
1zysIiYveli2v68p/rI6cAsLal9HCp5CzBhKvSXkf9PYpvOncqYpVZy0+nGILZAt
xsOXims0D9F7Wkx3P2Xz5u1jEZRjPPG2EJm0DFEWkpYMdX8lJjFOqQiUnrfoAKVl
T/0NjCTkzu5PuMKocH3L+r5LMZwSE9KX3UU0xHQ2DiuKv3ktNLEyF1R6FN7XEg10
v9q+HPX/DgB6X3zJcJ3dnO6BTPlrKHFqWLDSxMHW3cSLuRgTlmFV2eJZMRte1bXV
SH650UMACnVUaS2yDMOBPA3Q7YB7GtueJLZEm1vohHuCDaJuryT3G5X4FV1uQSYN
hfylFFfOeGrISJi5AxkEm1aWqp+O4iLlQ2woRgIsUgJ/oYXpCv5urUPQBKngqOBb
lZAzMk1ytfpeKrSdU97ens+05H1F5KuhlaWLE0WSbpjGlAu6WaNlsHo0ylAB9t58
Ban/DZJuS8tNfGJlpVBZO8UgGgVZbjrrVrqP7KfrgWIAuAvvwjWDqBMcFMYQaPAp
mal+vqoeh3pt4sCYe7PXrOO9F5yW8iAC03nlnqGigXCwQGazeZ6pRwws0Gcn9lOP
uE5atmR6gb2mtlc9AtInGxv7J18bJbhjyOYtTrzfA8wvf5PEDjsuTAOCD65EX+/2
7i9Spu40QGw5Ba+kKV+aJQdDk+Bn+7dnUpZ8qsDESOjarlnnLIIBC5rSCFlp8Gfl
UAIrECP7S0cYszWhg3u7eFoIrRdELpzQscrv5giZwHpo3sSJbEZtTGgPzjr8bHwH
XrUNum2BFu38CF8NGhK+sz2wNDOlnxaR28JBVikUyqMvh46o0+3vQoKJlxx9mAy1
ZVKqO8t4UfuDFIgxbGRWGIn7cNxg+SQ/OIhv+W3g9/WGoIX/rkwmOnIAch27QSwR
pK6d3iINa6h3dilwLgKspu4YHUlG61vAkNbWPp8odVWvoepe4xeLmTqugeMI7MqL
MCEZSGhF5W64i+50qoSCAyVvy3PXTwlHOw9c71sVIHp/qXvR5/9LIBxUYAlKxIC2
gAc0zqW1d44YtWrXtnWPe21D/Bo5mzPNGCPd6MtCsV5oOha4QnOuBNMK3cMx/lXX
flEcbwoZ7MSq9MTMeR+6DtHMc8pnQFuFGu8jJd1qibyVVhlJOA4oXk7dwlWamMWr
2MIdml2+vV1Cj0q5tN9VupORUrCSsML3SrGm2vwyUu/vqbnFDNXrv5yc0VJnulWA
bKvGQ9xnmjMYwgktbaGQ9eNX2GeL9CKZ+XMeOXVLOnXM6ko5Qo9WqNxkdCel3OYq
D1j0uQv7XgsjmHkjCB8fnpXYwc/tNkviKAyATgNtkD6gGTnCDoAiTAST54m2JMZv
7/M2ZD24Cw1ISrRARG2kxoqREujakDRkhiQLmLhuodOSufp8V4ZVKpI4wzWDmC0U
kOAn2MoA8etdZvAI6ZmHkZZvERAYvBF0C/my8iyjRa8WGvt/q+CJGJJT6GXrt8fA
w5eqWLMrO8Cl+3o3iMw4f2udka+7q/huxCYFXCZA3pRxv15XtIhxvBHtRiDgo+EL
1rhCVkCYXKPSr2rAnTzNEjq/LdaAq/1EW4Yq6Aw7H6BdEJ4VgZ7EFaxiWPle3qX0
JG4VojfDN8z9JfFb0f3EAXtOsEyRgbTwlvEBOf12SnND9XHNDDNAlTTqmgAENqHn
sMehLHeVtvBDGNpkTno3C8PmFE6Pis8aJC1YbQ2et8SSwJgyjPRiPWio6Ma2bh7j
n7NjunkmiRLt8ti46qcKpMJRB0JbPGHS088XOPs/dkD9Xng7Hl9sE4Ny68ICCB5+
uCA/0LKkOJEZkBKcrckUPntdR2dq5hSD7HEqEvCv1ITyR0DImylwRohjLTscVWnn
WRKLniE0QVWVP0pM1KufR/kj//UVSspSo3Lw9+k3mWLbCn+KZXYB4XNim1jUCQen
iz7Rk1/IqvERkLMhUenGQkp+Wv6C2+F1KRJf8h9POeWcnPofJjQTotTHoaj4OLvS
NoBO0vcK7xj/2qj3TSK3LEoaHZlJ3/SBts+CqqdO23G+GFCUgaDDQCag8J7TTiRZ
m8o9HROWZ8auoX5OqKPSdlo97cFIRUwYRqRcW9KyxNcHU4W4e5mzjLK5YuOD7t4B
sstfeQITS06XjNqZftypHXg2pDZ5tBTbwFEsylWi/drofBjz8jFNob7Ys5nbb57t
OLWW0IFxTfHyLdwB24idqshk2CxRPLuFUISottMFTYBmoxQfGzch8F+VS1Fyrnc4
CPDlzpAB5IC+nn8v8TJpJYPArnmifZh1WQwle6ySil5va9EaD98OEfm0vgiRkfJK
9Gy7Q+H9JomkGgNrtw0YcHMZB/J/Y8Ml63H/uXL6vU7Ka0h1RQqA2KKdT1LNoFMl
EepiJA1+GKt6y7rSAXcE7TiYJcdt3w/zZ7rGVCOJbAiNCBnIcCDNW845Qft8lxSN
p84LNikxH56nenC2bSknWzP+hMrIumbljM6h/gNA7ecsE4OSwJrg+wKEsFYY7FuC
0Dlvfh2jHLWpSRqgBRBuSMyOM2Y923IVH6qWibeblyzg40+Ph9nda18NfMvMpX6i
G2TSpS+1vtGXxdJq9Yx3CqkhFhCXJ+cKSDF8VajGxnPj22lPlBDxXOO3y/etiLJJ
zu+MmT83VbLOkpGZYOmO4GvY8KSUi6O41FDiDlmoxCWZwMWeK2I2N4FGGcygJY4l
aeH0svrR1ysatdxNnvKxObl8Ux+wnoLH184/fP7GlT7YuSctsI70bzcclYSkFJPu
Q9osR8IBJdtTPupRMGuYVnyWuzFJ8UrIBzJxPdMxMzH7P3cgVDQIQlT9sQxmGSEA
gtqBMf0tRItVIsmH8y3lVlW5u0FtEkyEv8ee2/NDsUJwM2Oxh8EO2YQmtHk2DYfJ
nru4d6mMOgB2ueMhGv2v06sVreP6bzoqFHy/uYjaST85s5qgncO8IJsPRMtxqHIC
3JMU8zW82XN1t8VeC4+yrQ4kPqEsOjfDeXUrUhEmOP4gE03k6vd6dmsyi58wGIL+
vAczh/eD96fee1maCYXnBRnNrDIzSpcG+uKciGKVRzZp8+EgN6pG5NC2u+Ihceia
bbvqCMiLdY8SwCxym0/2gpQd5WKNfqjkqrGORo2pwJeOrCkjex2cK4Q5eBmcKPOm
8+CPkqwFdhTOfkVgC4Y1AesXIsO6e7cq9MsQ65fsV7us0VdBYo+XXnFPMwa+5l2h
cFjZ6fORwl/pntuCyyGHltgYkqfNyWthu4fkMHAR52gTyqyj/uoO8n2SjCSOjL19
KXuAAdz/eoPQnu8+MsqHqMxollj8CVTAB9RHzhxjSPLc5XIhfLIdURGMFC7agRwc
KDQelarEx5ig6GzXsII7WhsTYj+3dFAlWOlLiKElKc1eHiePjIuEHbWVuQ7xDXLK
LSv+z/8kdIcgVXQ3N73a1g4HKy2O0ZoS9/wVqYF8tYnJIhUIAFab4sjD7dcu6VHT
rkjNf5nhP27BFvDZDUKJY9vArD/0vUqs5V62nqVxAcCL1B0aWVu/zkZIqvlh9Jbr
wuS520fosisyh5mCP47/Zdy5CeEXiQlbdueDtW1BVJQCl/A/Zr4sYIL5wRHpUp5A
ILYvYs22wPhtyne9VUufXlx17jq+7EFG4qHfC7afey9v0OUgLEPLcDyZK2Xu5gnY
Iw/H0/8Lnu9w5gcmWUN9EskFGFHmOhF4U6c6ns/2hA9PUX7ZMQbALY/eSnksRYrd
6/n5PQV4FcKMPQtQmDdMLmrRMefmX5LEm23Strfk7bAO1W1YtdrSZt/QLtZZYiuR
7cqvbOCuQjzCzl8vjxMhuwrxerAuXMz5rbRiLDRkNV7qc7cETh66Et2DOD90FIqO
vFCQw0ZVuj29BxiUxkA4Znk9XMeHBchlEGvSIrU4P41mfj9qa4hOfUfj8a4Rth88
9RxioqMocXkrFsMssEm6XuV4Hmv5ldDGEqkGeEOI6obHCXOT7m9SzzVxGdLJClyw
WinkjP2Si71bc1XIiGBhqrzyPJqKFPwk7sDOsdR96hfM+AbrF1dDsaQyhwfUtqAy
y88taq5gxnTOvqQnNnDC3UwiuzfrgnifhVtwl77BelGNg+QlPh3VynwTXOQeRBTa
ZAp5bp8NXDt/2BhiPYD4KrkAbbKjS4BKJCbx+SJp26SYUEv99P9UrtXtB5iIA5MK
u9rl/gj+1uySAvmou7qnph68nWHejNsvBPWje2PiB6yeYX0ZC6Vp895t508LFuXV
6aHH4QtXTXN9Ajd8d8IGb21PIL1WI1PZSWuWuDVTNX9EDuv+vWkPuXlXbBwxv7eN
EJ0N7yBUmrLc3rpihN396axNIQmjrfvXhaMc1sqAj+AgyKeWHZf5L1fZBT0Zbvy/
6HtQsw9O4WDHLpBrL47lpCLyvUwfD00xca15zQMDiJQxTa3vQP38eE4llV1ZwItP
I/4lTFnrL2saa+Y0uER21vjhCdzK+cXcvXPsZSvWwk4LsP2Ab22teo96KJxrDFaY
2VQc7fO8cA6mA6BmrO+w6mOghekklJRlQdNPKu0glfbNctem+sUzz/M2+YVSmU2E
kikW0ReIAXSh9bcaoCafmjNFCC3orWqa8Kt83eQ2dhTohrY9t8Z3Vaws7E18V6bA
Zf7t0Y6yFcmdBhskPmePyG00SM+38TIpq8nquY/G9cKgBL6dFCTpV1OxWemPnQlw
TEikOHBpiDhMwIzbRCj+5BX99yq/9nDmMbCt9kcSF8qm41T25SCGqYOZ/IHtKlCO
9FikAzaWOVHlxBSqrXova64d/f/A1Hs7WreF54IHh3UMMVAIwWKTNjZZHhGMJO7Z
4TxnXc6pKC8bQclTHh9hSeucgfEXEFJcswVn7Lvdhq6gk3DMGp/yurWyT8rPkTDA
sTq8IL7i2hb92V4YF4k4xEwkrcPIQ2Uo8SLSpc8wkGPFLxpXaSF7sdD1WtrrpHCh
jkguawikY/z6/dnaWadcvWqatbkPVeG6CUYH2zErY6jI+RuMQCgNZ3KsUmckN/63
TpEOfSH+cIhKsbLjeavOu4n2LllAPaFmAjnTJPTlAl8ncD3pElHjncMQdXqoDoFE
FN56NJ7hHz3P9mLYv3muXUoYzA3r1G6YDiWpqfj4Utz9Tj0BXr/YlS1luIpdlnHA
Ylau67HEJNDolpPDRQvVT9xg7uED2dXjJru/NuZc7P0/YuZ4L15Zrv3gUnuqZ+D2
dby089oJH17pHzhvs+jMOrrsSYH3JRBl5JuD9/Tnxiz2Imu8qRTJWGdFkMGMl9yh
iA0V2VaAtzPsVHJPVyhcmauBmvdLnVAA5HEWBxybpu63r29qzhy3tsQ8Av3FOCJA
vM7epnOK6WyBSWMZnAQJ19CtReqiNOMh6jVsO2YVbxspWkjZUiopklm+vuneEteF
ki3JxxTSjr4tAtb/DwlJpaQiJW6ljndYsrSWz6qIEtCeKjo/76FGP9YGFmlJuqVb
AcreQXf1Iqqje8ZxhTJviT0IDXpdSyTtixWyajOgOnlCZnCaFTPIE74A6ZIN5fOV
w6bfGd4krkpkp+Id8sXGnAy1OyJDoLu/wrOUiimsoGK6c3MLVbN35EN29BoWRjUZ
Gtn7gyNkALnZ2ROrKa8TBjghzIpJeQuzUgvZTek/vyPbKc0KwOFDvXVbunxCumUG
zaR+k1CNwfoTxG5td/GF+K9YLFJ+p2fgAUQnJeP+XLvUANTas70mGCpAvQydisSD
hYSpr8vLbzYUbkzrKvF1vkouebjGVu5B3yKGL1PZcNXeHYilKAEDHPZz57a7rx+v
71ocjuDXv8pjCJHUGUKAydaT7hZB1f4M3sslO8R0wuRffq6qcQwEk0sb2KBA45f4
MyiuDMFTOQBArr+ZjQj9ZLUMqCfqpzAS/9T/3euwXeXc+ZPt3drXBXj6Rl/mTL1Z
Ow3KJjv5s5yCJZecEvmZ1dCaGCC9CJ9DZQI1BPrAM0+2GtGcyGD3KjyJVSMe39Gr
+dA6TJxutXMI6Urg+g4vKXYUzqnSZlvfyhNJgiQSELrTwJ30KL6hE7fQ5ySmo9Ih
IffKVZA/gP4N9Z5yXrWFlOxYFb5v2w+oOv2ZM50BKek/6drVUm49eyNW8FRvmTCs
pO5KO4Jniv1t6C6x/TtoZo4AbOewxY5ijx4nj7y74GzA4GxP8GQF2s5xAzurwiem
Jjl1uhQvdByEvIaT57hyk8vHjTQoDDVdPtW9k60TZFjvQK+bjbRVdI8BG5BVsHOX
0jMnbfcA50AS5HiewkuQh7+sLSDONPINuSrlt8FzVmPWToJar3RdXn/sAvL/Rsbd
ADFQlXVipxGMVoof1FM0ESk+wYhl32pHVkcHh/rszAdgIFpR/JVO6O7dGckH439k
rnGfn90qXptMLhMRcjqZ/FQQcyQjjn1QwdQ4sEmyeIw50/u3xRSUUArFou3gL6NK
6xms8O3L/yUsjI+pMUAD3aV5O1SLQAGj6gMouP+8jAblcOL3yeRGKDpMf4t9e8Xf
AGjs/tJPoTL8W/lalqaKfo7lmG/aO26znstVj41WSq5D6sRSZgUdK8aawWwO/s0X
UK50B9a6xzivtbmuNPhAugLLCS7mAZ8GcFC3Do9B6fKiFsVu2iJo2u7sOLhRQygu
vqODL+a2c68pcRIlvBkrmE1tHFUH/Q57q2Iy2FxaI8s6ndUbbRU87LvT4QFyGvFU
hZU0o0luKcVPjGpC6VoWkGT60EIf4W6kleQ7GhRYhiaIFLtahfkD7pGdW0HHFXw+
2og32OVrfzLLnxomi0qTAqiHyjwEHW2o0EsPLw474nffftcjDW0oeEBXAPAeBmW2
hTIn3RQ2lybC1Lx+xyS97UTCwyddzoyoiU3M4YU1e1KCJDGVMqPdiMQWt9LvqzlR
PkDVC4EmbHEshod4ohZyiYUWmuHWXxHWZLQi2GO3qw9g3MSFAeShQC7IL4AvrZBi
BcA7N4XAFduTmqouNUGclpNv6rRTXh/ETtfkP4dKD88hHsvd5ab7LNbVG4wsLy+Q
jft3gHUTr3B6ARhtXsoAvcmiGg9WEXqPJ6qFypFKE7fozMhtyy+tG5cVwmI0XtN4
nIphjXuTvBidvqQnZEojxJG0QgGbcIOm2snfEpjvmPGmttib+udES5AjTxCQPUzd
fHlzjG2LrkyPR4qzkGyD5ccHM1C9TBUmnnS623CrSQltNnDCbyxNpBM/B0ObuF7s
NOwPsdkvLi5W9QoiibpQgKodO7M7mBYICj7GHnneACz/mtnNNJQCwZmUGBS1DVFD
SV4f4kbygJ+CSvahkEPiC0XkkD4/xFY5qJ+n0T03xGVEPt0gZ2Xj3VS1BxZAOpbf
ds7eJACEToZB2LYmWAHUIJT3OasEMc/LFmZUQeI5aZoIj4u3r49d/s9uw6etU3eL
Xz5Q1jjGtJfzEg4VLYy4t2w9Dcdg5IiofJ1d/pNgHuZw403ZqyqooMymVxBr095M
0il3HLpb0wl5/YRh1DjORyVwHMkxkfsSsxYrk5mUPMz5/eKV1rH0q7Poyxk0yU+q
mB4pDOLvpVuwGOz3W/Yr8nXyvhml6dWn26iqYVV5tL1nAfLzAEWx9S7h69LsNL6/
f49wJlpHzxwnUPUdm814dpBi/Gb2KAtqafTjDiuXBkRsBX0CnCUFkEwPCkGAY4zo
lQWuVvbPT/CSFmi7SsYlWhjMLvcWxymL9mGrY4SSuIzOSKfXRY9txHLQA/F21MzE
cbFTp/RJrr/xYPWOsrRvTOY1CbnqFoerVjRu3l4Ub3GWCUVGw+1GusLZ0G1kdx6I
mO/x3KDh5WZEGMmmvUiFWCpBGSI6qtUET6Ygp6W2ijyyEWgyE5og29B7eyDKnYJc
GJKemgulWps3VVyE78+v4P6wef+44j+2zmK+uER5Vg2jglXKznrX/zOe7R7TnU32
ty1LT2hH7A7R76QlGmfYFcmEdxJ3HL16HBGONpsIMh7k3NGG8uwtFfQ7/YHe4Ups
kwUN6bcF7p1L8ut8XWr4v2GQ/GYtF4BCGUbPmJR14vetwpA+YPsDnXjcvilB1P8J
wdm/6WJ2078+dopgvSqGwH6nZ9Ghh+Ras46v/F9ACPA/R0q13q/bWfEoIrh9Z/lm
keoOXtE6GI7TZIJPDAkdnEVwQfN5eV8EwtMtm0UsskrUbg5LMeccEi2Nf05Xf5+S
MXdTrQT2zRxElWuBob6/pzErzBA5BMmxF7f43TuRM9vI6UYieLiYrAPtJNcOLxBB
Szqpq32bgHeBn48UYU6WFAoDiW23k40gRpA/7s09F6Xdb1jtXfGkj8vVX7w2QYQa
VhzZaMLErYxdN9PqYKGxgxVyX376Kk8DnagB2g07ErKPUi14LcXl2KIMGgWow+eY
yr1Dhp2Alab77y4Egb3Jd6vmTfUpsvvVkma2l8Ywq6qeKhCfmjNR/lsB0BndUJjQ
JVSNc/prbk0g87rCfZEI/ki9+VW/yh30k7QZ4a6Wpjo8c2seh353gNTFoYaYgmql
HH+ZQ3Br8D3PfbXkYNpmSgSgqeos0clHWOUVBUosP13k9Ck4lOiHYfxIb8xMM1Wa
ctiCZ35xSuIR7O6jlHA0/Hf+2RUHuYm0y759N2S7mUJDhexmivxrwiII5fOHFcIY
mJl0e4gUo4GhwJkb7juU7jMGo6R2HcdCnN1aJ4dlk0EUq/hb6X5ya5Y/KLX2t6uM
UZGy5LqIxBYEatB1iH8G3fOC0bcd0CmS41i6YykGfJ+q9kVv1PlwS+nmQe8jpJs8
vZYMU0jNA8KQGJvDN+yRkPTyDzZJPP9ha4C4ITwffYFLF+gk5BGbWvK10da2xHzs
Q6DD4p01+XmMuLkjw1qRr2846JVpb3GpEZM6/imnROZCUGnpBIoNrdrXnas/PTky
mHayJQfmjO32bTz9AkOvG0P/O8B8N9rbWjsr5GRS5+/Wz4HBHYhATIgiScd71Abp
kSIDZc89YeYdFUBhhbdyBgvbEJTkmEgG0pCdw8aCwGoHbUIaDX+iXlxrzdpWVLiH
hkTqISRtGwUsULFPu8EvcMVmRTn2RuOHpVxENHndvYqMuta69C1lV57Bc4B5LTTr
HVRmEEjD2om1kpR5kKC71e8lrXodqr5/4w1hS89YO0KH5Ht7834E9WvLdLJqdX2J
XYzYN1wjbeACQVBPh19+2s6zN7kV0OlTOEYOV8PB8AG16n51leLCDYf/6yTNDROM
jCgJInNwMXZBuTlPoRgsIWT5XlJF4IAuIw3/xWlHK1YA6XbM8FoUDYps+N1TDqvt
Y3qZ0g4gHJd/voRAjio8ZCMJM4KrB8z2o2TY285reTPabSq/Pc22KvcCO8ylQoyA
OEdndBy+dpHEduenXMcEOQoVpYO0v3nmV5HOnTXmcdo1Ghzc5iuavQ642JBXFR67
kFk74v7taoLrCbYZ/fyDxlS8PAO06yZx/pSM6acfiFKl1Cn/D+KLCf6j9anHvz1l
tdn3nJlhGKo4hjLiMyq3ZxVjhyYO6rGSoAzahS0nSo9dhq/cnxSGOINWb3s+/YmZ
clwDeobEN5eud7whSBHKAo0Wzs/iWtUjNtE6cI6iy+IfnnTzP0m6Eo/h2BYBkvfx
eUsf5sKrv5e/io88ZQvEw6uVvU7WSuTU1UelRGQCegil2AGzk475Ixbt+v6ypKS/
5Gvgx7W/k9Mkh3gCdiDj/bcBr4GXybYnQ7jSWqiKZ2qvAveXqbANSYu7f++k40OV
RM2zr+oLjj/HuM0I+pLIw96u/vHdS5pyCONAqiUrKTZSQ16pQv0x8Npl1iqz++3x
1iGuhApPl3W83Sg/wADdp/wBIw5gN9DfSg1zi6MbJ77rLcVSPNzH5CiYAAnahBxD
cOB2HuIgL+QKL9Xc4BiEAKoEH1NU+aJd2YXZuiEnmQVUoGGci2eqW/dr+OZmLwka
0dzpW0tWwqEqO0j+85+FCNUYwL+1enjSjMKbEZl/pB2h7a96XNnxzbcR5T1tqTPz
tCKCEUD+MNxGyfDtvG/ZD+sOXBOsC5EK9mQeUo7TqbrF7iLlBegD+69HDMnMUSGa
ozX7VLVy8Lsd4AfO0Ad9KiyNX3SnXYw+ohrsJR4sRDi1vBBd2GuyruEP3ww3IRM0
gpNs87P37vzJjMND1TGL+iF213gxlIYwtUy6iOODIbupaToBnEn+dgYXFGy7/lfr
z/eOQYt0g7X+HJ4iFl7ejsBvEc8RsqKvGHXa0vo08L6i0Knb/kEvitbMA+nJp+xS
rWdrtbnxlM5SyquOSXEKCYUnAbvGZiWStZSP6raZr2kYyy14msaqNiAoApTK9qDW
W1HM7jI1qL4X3dv3vCytioBfsDizbdTnXtxVEwgpq74eLLbTS4HB0z5G1yL+N1U/
22JATMTxYjC5js83ykDUts27pOEbnr1g2z1cJrhCKJ79bRAgKjiOnrQ3Z8PPaxs7
1u8+wuqeYpVi53VYhO2VQZEvVo55xc8zgzIeJvfOfiV9pi2fbhJ6jlyjcUSbTBgp
+HnSXuzKZkDKl0FhTx8fTRWraSe1uxONz71r+/HPdKJM3dNXSlXBLZ773mvoiJZR
I8p1mOcgkcJsnAJ7ml6bEwZ4lYkAfaz7ksHd/xOrBCxvNtq8XeThatETy2OcuEFk
xxzLjabHv0H6xXZxmedMzmRgvVZGWk9AIJ1kckod/o0OSrAGwlJCe9yebJVkHUJl
CFOiAKw30V65OiiJeRHWx78LOj7dIePP6tFCRMyRxqdlVwl2xlV6DbDr8Z7pasiM
kOqtgGQFQf4ETmkdp2b1v+QDE5DTVwFOoivhcFoUXSUiQbddZt4QY67KlA6hnXQj
D11VyJgR+IcLLXhDeoBHM4R3I/pZdQgd3CEUEYJK2kHKwFRJZsS29EHhWLrcXnCc
OQgg+w2SgxIpmX/CvgxOfYs3MVS+RE66HRDgJePYtb6Qkf/3EKcfCpjhaoOHFHsm
MhGRvZIclnqiltY9uDMWMWeRn6SPJlPQFuv/aos/9GH4gIJW7bTALgbV2hEcbet1
o/zjec6lIPHzA84gctOVZxrQ0TesX27KbTZUW5XkylYvzpkkgiabFTF8CWelrxQN
0zh0hdTfBby7j9YwvwUQ8ure1w+x4lJLPrTAgpkEa0RBPBZQkljvGWc4US0V3A4t
19ZXWlpC3qe3FwS+SSwX2RxVLmgCiB6skYKkHPlaq9XcuoCYuV1L9NB8nFAGJR/F
xCRvFwpp+Ubn/t5gSJhZN6CAHSdydQQAD14MBkZvAP90y9zVhG8FX8d9F6hlZGh9
XkYD6zD0xwrFTdIoXH1GB1+6fwsuN1FKkj+Mk1uS9gzQIb0okmVjMlQSmUGBjHXK
RnEmjriVBRkrcJAPlNFR+vBAFyz6JX5EBE7NS8auE0iEyrhO5uKloeQ87k8Q0elU
a3OuFPRfdo6w5GeS464mssXSdjSulR/lRl2DOXAH7fdg65zbg5uhZ8bryRHnaqGZ
/lZN54gOVq5VGR8D8DNE/QjxtXB5inuohQKue2aNd7YQYlpMBHd1+wFIQRqtkGll
aL4N9WZZjFnyvD747GNKBdFGa4e06iktfXAN7MJKIbw3ydV9aWY+mvfSUQ1N0mbb
VnMarw0qUtCkUcTIBZeIS0n3J8hMK82Lez1AWr/ZRyWWyXiIgXiaaWXJ5D/3qkdV
ajy64Ewh254f7/Uwo45+CdPDFACW0C6I7ZUV1Kpaj83RBtzXz1zKnHdiuAIgxOW1
X6ptl/yhtd/FZQzh6lLWfOjUnQlZx6AVYW4PfsuG4nqjeEbBDPm9eudosF+9qBFv
1g4klgMvOgm3SkChsu0ZQnVpb5/d/FBjgpuBod+srvrcGyfaUyobYTV8W9w5Kv4i
TshcCaue+U5YWzNTjkx6DvkA8gMc0TV4tlkW7T2UtE26FZDf9mzutvnz9mVGQx7e
2rOq+7fb3/Ns8wm/O5e7OgUZpRWV9Ml/4RUGDojxW6KqYZfFOwF7wR9htXt+8DqF
fooY8NKwImVmp9XcbU8jQ3OZZLfT0E5amEMeR8XP9Ni4JjCjMm5WYcGTm5pStOcp
IJQuHhHOCYh+CzpuKZCNDbaET0Qdt3A4A227Q0ktbbfFz+lmSSuWzH/t/j1iCPDD
dUjQ6ptzeUJllaXzfXlUeZs8+g7xskdk8MsJjINv3Kmkjh3BJpQliVL72Bjd562p
O7RmpzkM9toCu5YfqOefZ2XT5kG4WXgHwRDds3kODUsYvVXzF5YSskRf1uQ9GTaT
uQ7dSxhXWwdGNpE3iLpOfc61bEGNDD1SlJeSxAYnXYApZXGjXScZCDI+ncs4pUd6
S/kSBbOsH5h1Uqe29mPDmm/JnX9ZEU+LNuyIZaB0c6WhHqNmKujWaHmeztCitGNF
xjNcB6PL1WmEEo7c5m8jFo+HWL0vVkf8NUCs4dQKsXVl1b6nlt6Xa08jymZcN4a4
u65Lk6fqQZZoM1tcUOsddOQTBKQYZ/YVhlMLpVmZpFUO0M8VmyuPK6LtSggjjstS
9XbhT2kz3UhI1KByuaBwfHqf8+sA+DqNGwmy85HaDqexzU1u7v9deFK/U1NCuLEG
xYAgHo5nhZbl3RoIb5wVcCa5NTr1l3rtyK8oETCtZX81hOmODkONbDhjn13adB9j
TDlTkRbuFfYP94p1EKA52umJSx+3tau86WKhH9NDVe60Ydd2HUCwrJZPkedE0va7
FA81tv7Q4aSP+c9SjYYi3tnXGoQMVi8MjGl4zUrjAcd/l74QNkO7VnHrCZ5T4qoP
5rTntxrTwlygkZBKeZeyWVwvTH7FQi3tx4QR/Cg5BcH4iFXQjHB0kRY56S9GPNG5
FVIloYq5isj61wtS93hkURmKDgXpBrGXthxKLeRhdnHbRj0hlZNQ7dP/w5gytKkn
lb45tEatYcmWslOYuXBU+zg5cA8UFBoP3DDYfWFXqFYVzf2EDH9hlNqpAg92L3p0
aPR17tP13ZNpzYqscxRuRzw/y+NPsC2CoJmveVfUN5v4iCb5Y01KMTZyIJCNh9N8
ze8U9eHt2c6JpLCU4BxgJbFhhEBJ8xLchlqS3JnSg9SJQU2KOqL/SgxM+vs5Ufu9
z27VL2cAJF9piuk4pAZ5JjLPEPngJm9JS9VZmJUW70FpS1pS+EXLTmQcx3RDGTQl
TQLUCrKin/Aw4eW4k83A7SYwMEeZ1/a5HNBhvgcZeTdCsnHXaAkvC3YGwcQtw9Ko
QAtLkiflczEwDicuQA5fY0QdHBNXzGKGzFgG4bxovG3Xj6nzgOp76wqg6JujdjDC
DHUYPPWTABSSa8Y6NKm+1LcCpydoZALOs2YtrdggKMq15z4P2D+Wj9SKTYGe+bwk
EKx17gb1iXjzwGU0hy7idFjE6F81nyEGiDqRdhpJMScjzAW3luVuJb4clgyht6yJ
6cCUpPUpRDJBk6MjO05+r6Jb5fLJkQhmcVKguS5DCuAqMf9qFdMDuN0B5bPU7VCa
3X95lFEP5XTH4cUgtq2pdyGuymK7yHhhlZ8jepmX+Has3T9CnRkBgJqzx4leQX4a
x0pOFZ4dUlXSX3WTPmlOXt+sRQTCvnOMhj77SAo9ywuv4W1LR9rLuUO8BFWDbJvM
JY3yqpAp8fsns4IGsx+Ac6NEcDoCS2yJ5c4YWj+14VLEj+cnTo7snof7lZKbYaRK
qqBAAsDbfVjp656HnVZz7ibb704C5P3ZMxCGnRNTzxKW+TAVPvwew9Si5bw8Y1Mh
dJaNe2z84izouxlhcvQJjyLrVeTMQ0Jh7hRXTVWpcud8EU2egbQmHn6I/NeVuCeH
yZ5t0SSnhWeGK1MWKg7fOc9EIxUXlTXuRXTzaLE5JV7vjqwJMuWFHvE1GOJ4EgF7
Q9WPefnF7ESSDGpRFfDCxHeY6Y7jIG1RFrzcXs9hQpmDBbFHXE1Yuij37/tfUjho
TETksNUKbiZg62JCrWwaZhjmO3rQiyVZ2KoV84JcaV7vkxTl96X1bZRjsvWtpmFk
daz4zsMXcTRVInSSFatXr/MTo1owEvT0KmTLqpdXW6BjTziKIeyVGy+A0TcSKuvo
rsNC0L3QdGzmrZywmdkbJuRCF785VGmKPqJ2JUowxMhnH/fV4fLiTq1DKfV+T4DX
IB+1iuwbFBgSfC2Nlao5FT1PxLZt8Si+XfA0PDNq2YyF4wcfu627YV+5lNu64U+G
OddkJ03hiPL/GIX7PQw5/6ny/FoDeqIfprJnvYeuTQY0SFlQTKDZzs1wntY1fF3q
6KxObnGsjHm/vCdQeR1IYGlZr/MjMnyWVrRQvv3YBRuZMUqQD6YhQexLMNUM9Wu0
9JKv80GlFFDS2I1wyxrYUaw1XEbndmfYxNGsEl3KygCOimYdWhJSi81PoaC7kwcB
C2X6FWF+wG18Vlg7no/kG1i+6tYwnqoTKQQ1VtJUvMdNp69nH9Gl6fCUJ/gHt9Vf
qs1ceFsZdjYVo5yOHOCrxgLmsQ9uMWKn7vDh0OKOgzFK/FwPaEio0GuYCUrFJPR5
n3rC4PSOGkRS4yYbX943oIj7mN3ZkTN9738eMK6ZDW6q4pyKAKMtSFJr7MNVX/AI
QMGToHScanmniL9tM7OoapZiSCawFiC3C/5nbp48Ql9IciRjrqafrst2L76P98/U
FU07JEU88bpEiCS8fFcvJqw7wGDEGpJmkrV3oDVGIuKsRGPjlETGudAXAwzx9A6I
1ZVLLEZNDuJB94G2yAUUFpjgfYY9r8QoEoPiLakAvQqKt+H/B/c8KQVOd5ESl8vW
1n8Hi2V2NUyP/8g47toAY4kTqtpFNGjWPzL1iQyyNcTpyceq4YpvQkdpbyazo0jn
TnY4qiemSCOrpSFuCgThiCMH7CnhYB/hF5wFlz9o7+nS50GJ2g5gzBD6QliOeWGJ
EUbPGi1StIYkcpjLS8Zqp4E15o1anesVXwL9zVOACEg6MjCnEgktaHrz3Xa+eaHs
dRCgRU9hUyo26CoFH+YZI2oaTztHnucPa+ViQ1OxXyx5an0p6rF1L+aKnYZSgF9b
05tgq2lKrK2QDYqlUckBWG+5V8tlMLJXmfMwf4FjsBuWkw8zEUveT9FZU5fS3o8i
ThC67K4iXIqr5wHClkJOhhfMT4eHTbshxIJRnxN0SJeKvgY/2jWeTbjRlzQ2IXVw
5ho8DUA5e9b0xrYjMxjjwXmxpdMGwqKVEKhMNV11+WeLYBjPG7gqpH77JHadGnf9
Nw1wdM8fLU9REI7j0kOPrUhij8oX076iQraL18Etpn5wKtw4hW2/YvV7qA1kJuYO
qYtCjYjh3/x9NgiAlnawbEqj1ObYhO7jKcBqZVBFZJscGNIoCg35K+ByvPo19OjO
92KWNJGWpP7LrrEGRZY9anBQlGC87Vqlu9Z0U0jRPW+spBnwYB3vqsYtvlAJKGUV
/ObIZD0h1oQyO3iVD36xQdPiBU3PrME1s2aj6WQHBCwrfPRIiyvFHDxh15hLNKaf
tUoqlCoxVTLyTtzlLO3YESuWrA50vkPJa/UibzuLO2KDjF1aqkfz7nbKrkg/zm7b
vSDDfw0e9Zi9dKelMg45uVIozTORYq4ooM6usiydnPp+7bE8nIaslMUz8KuIKfhU
oO6rsyfUQq3rfpp+oCTW5KSbJMw6aO/pMhOQXerNoDitM4Fz8vkCKoOG+vqvxAzZ
cwjYBPCAmJp4UASGlpu6EnrIdvWI+HJCsxXWoIpFeRy8dAngY0OBT++CdKcWwfpN
ZfCKrF3WxF8deM5DgaXSOszBfR+Kp2MNwieEcNPaaFQJ565sRhZgfflxSm9XWP9K
hcoA9fBGtY13jLcPtLgvYkMc20UOT2BPCcAzu2R3csVX6xqigY+YESl044DYeoxZ
HfLJenIeFvP0y9f2/dPQkAQOfr0XpLubWCPkq3TVteNC0eDrOO53g0WkbWlEPb67
bo+ZtAyrP7w1RnAKlO81t2QaRbLajMf9ipD/sbdourpTZbIdHItmZ0rxYK+e33D4
lXL9Aq3MWUZDjBibxM98TEYNb6Jh51S3J0LIvT9fC4KTNevQSNIM/UHsO0A8IdPr
qD2LaJFui7Op0LGYQMvd9Yza/C/VPch1JZT4poJn8MxnusJ2am4S4/N9Alp2Av4r
ZzC4nkFEZExhMnaKuB5gi/KuAnkEoMhRRWabcmn/+T4CpdeW1e6Vh1EoElBK9ABM
RimGcvYcPamQzoaRslQ+TZz5n8qGHvEfkyQvbZtepdLgd/Wjq51FoEPG1dQt5STg
Sz/Z/PndIxLUvYlXTsnYxxTdRM+AyyfKNnYKx9xSIK8u1eEeNbdwGbSbli0QIguk
z1kn31uU1emCMzEwEIZx3sIsTHXq7H1Il05lZp2wGJHA/RnvEyxk6v88nPmwKCBx
kzjuV6Zq7tnbXDtQPH4A/2z4wYHyMVX9C4UqsgVNY5JG8jVbcjdQ45VkxC3aDwnO
H7NthOSMsqvS3xx8tDbSwD1eaoos8xXVBg2BYQR+vCqPJGvH3dKdEnkDO2XPv3mf
QwAeorjrLYw0BHXhsqkLLdVdN4S6JDQ+oTcUxifOCI3r14lNokgA5FkdLKUIo5RZ
BZAbLhAQn424Uy1W+1TuH8b62sWV7ESJLFXAGX+lhcecIwa7QrrFUmQYemtCHv4+
xrVeuw/jjp+u5UK/CD18kxoCS5BnovdMSfEP6Ug0TEc8Savqx4516pZx2Trmjto9
x7SR0zXpUhYCLtmYG41z8OWPTEP3g6Hk9tyiWHmpH1aB8cl6xmQf+Szy1GSKFLQK
DUzSihf2EyDEVgl3djkPxyPCpbpc6iL3KuN/gObUPkJ1FQLCI7vhSKWvoMcDXnbw
CA2NrclZippJp0H9X7m3jQLBpqzXpoqBrOkBQ4nzFQSGkq2HhSzWDyE1mw2Z5s5d
4fP7WRJM83MPjjAtNji3lbvkvl8NVB3tFK7yplV3ezxLdT+gKnt8RsvgyKBgz36V
CBFjTAFdABCScC1/Mqb4jNpE42fQONZAWcouKRWPPCzqHYGIBAFnD+qdGXL39jVg
9imB3GUVz96/NLw/M3NqJiatsqLxK2J3falOAZYmmfGvk9e77bHxVV/wYPs/lNNA
TNpIQW4d1ILz5u3ODPhiwy16sIl7U5W3BzvjLccnr2PeZEbfJ0GdlkzPLKXM/hoW
EKgDPVV5uKPlF60CknHK7Wf53pIbA0vdVGIpbYE/JTRyeeg9epazBemePfsYYSbp
yjJq+pcHe2FVP2QVH5C97C9SI4dwlyNA5+OZaQjE0P6jGPe9Cr242kQF94+TMUYs
WFrLMhePMoYgLSRD+CNO7Past2aceBtHdIPOAg+nevcBqKg5QNmcCvCNJLNZVOSG
7iYjLHlNrQ5Gi/sOGHMk2tTib++5d6U1HF/PFoFeVofgf7L0vN0tDYemJY3Ge21u
+aeagAxxeiWepRJbnP6/BQVjI7eIBhSb1KMPC3Fy5n9YrE+WFSZqOgOCxD7qTt5X
/JeTXXY3f5OMDklRlggEe12FsLdrOL/3d2QjV5ry95amK0tFBY2dGyeXbIj+y2hP
AM+PCnoe+90YsKmR95V05QXAJPNI7X5WWvtZFXJREpIjRKJmdomTbc1/WOoagmTj
XHl+b2XVViwGT3lFxAQozuHLilTeIsrESaxpJkoEuRbmTCFIA/oCjUyEee/Tmg+D
zobhHGNsayQ5mNGpv9KgBWqAmmt5r6uI+lKxZBZVYk7B5YjukQK4+PFZHlbfWVGI
cgyZkjbf6Ja4BWlRt8TAc6EBXNagoWWWZux11/lKlhc0bv/soAaxSoon8EwQrcN/
2+tDXxS6zXm2fuMNGnQkbKrPzmnq0P3chNxkMw/wjf+NHKx1Sw6LTn6IpjusAsl1
8LdgEg6pcwgE7CGoY7ToRJhMxc4KIB1wP/jTFkMKzsV2b/U0bK3dz6a4YBxwDDX4
XvOGdHcfQu4Bpt7oIbn5HpPm5obSfZIrbiRNj9HU71MbbowMdHQVkaNK+y8LksGb
rGaq/73hOe9LX44QL+tXpyVCn14LLGiq2UZcLFlBvTHSpEG08NxBdsYHlKKcQMbL
I8QwcgHyh5RiQoUF7UGoKD5RpPneM+uH3pxr9o4x15xfrXUwZw1rujrFddUi6Bzb
bqdb7LbCt8gfE/3sDg4bVpCtugH6ZYues5zqE4uW9CPs+LH6lkDZTitxEHRIbNpk
n5svXC6eGfaP8FArkiuq7tPgO76wDmr8fvJOoap4WSbaL4NYllu7fG6kubWr5fOT
uLObOwz7iy0OOaXFr4grh0afOWblsPZxg2DzKvjbVtcX+6hRSl5SrxqwyKKUfjNE
LOJi2E8evJ3AKcVq2pWxzcUUUs86TFUYVHKjMzrMcsDyF3JQFQb8CG8EYFiNBz+l
6ppOjiv1kOE9mYa5ukGQuwv60irn/iLpnUZkDtmidYwrj0jUkyq3y/8yxJ8Pb8Zw
Ll4vvhQFtPFWqEXQVSfOZ/H2yuwor77xKnQMnC+7pLWIUF0nYuFZk3EFnbl9k6Y1
hT0c/Q+xO2kgxJgrE1zjSEBiPA59wSi1dHiP2Cnul5FWTCnfRJZGGTTI/owZvyl6
eoIhx/SgYX8urhPow7xpzDGJMAe4kwZb2fFfCs+11VSUohjksaZA1P5Q+zR3kMQs
vpuYIgXELS0VfwvbKPOAVcdNAIbzZYRXfcVHqmHA343klt77SACROsfyMIFq0qpw
gETNkGDoD7ycC0AnP0nyMh38V83b48WOZUO7p7WAbTUbt8oHohewyKst6yWLN+Cy
gccdT0cV7ob6xn7UxEJm4H8v9ZcGhnZYbT8ead9oGKVfW5BnjpXJHB99xOi64uVh
oVDdjOuTjiumybl40I0n5QvQB7syh75cfek6JC5Kx9kbIJrpVKP66R+ty/zfHPXw
R3lOe87sS76KoAiALkoatF8Hx7KNA8EBV5OHnlv4VOyt5UfEqav859US+PM2uQei
c0XXMOMmNcpKTeWSJqUxlXEgvBOUxW9wzpqHQtygoOqRUabJLTmMV+S0KddC80OQ
3kuTbYLCdH7aGsAvmtkWSu4iaSIN+HNAbWwmk6NKN796ggw9FxbpnuFwrWmBb0m9
jCiHvXL8+YD47IYW6borr4U/OxaDFwv4mkqc2KHBdAD5G11SvHj3GUQ+3U3UpVeW
bHXgaNYkrhl1GTgnHL29ToyMoqR4p0RKD3y+1UejK5t3CoXDyklZLmG1NQlAenu4
bp2X6dcHChitVxfGxZW8Ws1RR4LwahKQrfaeXKzI95PeZthf6y4rc0X2/RxDcSuF
ankVZ5SBz7IRPYyl5rHIfiG0udM3WKfOS1QTU/lntT8zVSFhEdeFOlpdF+MFTNbo
Fb+PxmEgh2D0nzMloM8wEWiiK3bZGM7ixXh07+ALsZ3dr8qr9UcJ58zxsgen28YY
N8+vyr/+pzel+2J6L5il4pXYRF1tBVikVlj6DqVfbkf+z36qsAxFWPy0bWmC4AMp
rTihu/Vm2XJcdp+Lipaxwh0IsYWyTX3681hyU54ZkhvBT4i6DWYrg80GzdgyN5W2
qgZnSamUmuQuO2OfqrZZLJe2Lj67/GSPFx5mVXc+2dCdhR/NGIPTUGAqO6D4ip68
iyFpWXUA8tfGdGcQoaxDLy7fffVHrFZdXCK4BMEIzWazu65/alXratCLxLUZQZiI
9431RJ5LGEudH7DkQFhicYvQoESEmkhjODj6md4MyuOWNbyE+i6U7Z3gCAgCXlfU
IeVkMtbW2fHyEjtA4frLnsSW+HwKatzn83jtQkFbJcy+LAT/7eTUj7d6kHPeV2WU
JddDCaDCvNjXq5+ApPsDwssS4EVwO7nepTB9MDORoiarGTZDhdSHhSlBRGZGKGJ5
oGaBPg4H/G8yXE050d/euy3+SxRbNtb9rbmSgXAlEMx3MfwsgP+URIF4BXaQrT/4
5lWeosHa+K+wOd+MA3eFCrOVL4tDOLnNzTXUcxDmV6qMwCQbdYua4By8mwH6/KQp
AQEdfxuaxCcZFaDCCXwO3eDA9ZVaZxEW8Glzg+l6nzTfB+vB3T7Y7hUJ44VYjV7x
pYYAVAoAR7ay2oor98siUsSnSZwO5ZrRI9R2HJps5Y+WJk0jaNlvDG6i4clGc8ud
4xQ6ayd5yAHUacS7/cy3yj8gxw2Ik1/EjPJ0QpJVZqpbtVlvy4dsQdBueiwDS0N2
ddeo4mRKBsqEyg14SrsUTLMihVccYtuuyjODKGqsmEao63RD/CLvizUNzDfmvtGu
CqNk8o2cnLOAphjoz+9ftdxtwrzCZQUJFYLMM/GKNz/Xl+vKNZmq61Pf9Lm+AxLU
di1g/MxP5bkbTiDB4WHLi31beDTfDaxUpV/vbRuUSIKinDxhsboaQvnUg7TjR41F
cHRP2daiNSkgO0EN5g9h39hirstHaEH/aqRt5NCGowo7bXXoxRU1tp0xflfXtRZA
gBWCJ//v/oUWni9JnyPI04PDmDqTi1C3qbwLUCkKfwsQhHbYvzpZGlR3c6rU+UAX
QFnMVyZJF4y7FTan521l+0tytm5qMa1/ohHlLeSz7SyCayn7B5yCCv0wGUcYcWno
+8mI0puF4JgZovRxdx9UdjAYf3Kne1gM2LjA4n6ETX3NE6exqOHddfuAllPbrYy9
VxlDJabOI1HNuArBUa1hMzhayQG30WYWaLm2xVfOr47qqXr0cvwRMipsDw1nqydf
VciR+NxBCJgibuimGVvpRaU065QeyCXsVyBtrnGX1LLTH0H9ehI6p13Hz9u/gOpf
IZH/rboV6E8dAyBCiGFB9G+jXUlJvoeooCoM02dgY+8ixCTFStGkZBMvrtYrG6S0
01ndzwvhQHEBC1RxFRg4h48tLfNAgo10w2Kla+RiL2dbQ7JBIrxJiuOot1n4KIyZ
ynE731DGuHeAanElt2NrRbbtiSoN6rfW0eLSbs6Q8414iRolZDUoGXJlSJyPT5A2
CH8DIFBYLmMmPawhbcbCHdpFHVYj4PECDwjLQ0r4iuOGQF8fXhz5RnetinOwgqDO
V/6cZ8nlMvHvHcVTKcl4ROPKIjE5CgAA2uiRQptFr4I227chXPQS7oZ8UbXS9BCi
kU8tZW/rkM+sKkDSkfxQ8Rh21fcRKpqEdIzOsHm9wIojPU/X6qXljYcBHkcXwngM
UjWB5AnWWlWQWwvYEuo3LcPAAVOK5Yw/Dy2z+oaf0i+70ZAHPy4FODctt8G57y0B
22CuQn4Go4zS7KtRgkXM+/zXX8/gsk8kxA4cIqH2pgZDRIR6zmOhorznchEmr3nj
Btxtzvg4oYsOfgLBqJHv8vY03oEylYjQDePH9dBHftNgUeP57NnC62Q9069k/vJ2
uETyLOftMl9NjjMthBposPZs1YtJTpBYUyH3vPRGCaxATQskxnTS/rVmUXTSZx7E
GoUFEwmJCwoorLoxdH7BYyuBs6kO1wXGX91WHZzIe+3+4cg9UFa3AaSr66N9IVwK
pBlX9PeC/mMO0WcK7VwMYS22T3CFt5b9YiCsVkRXSZ1mKLlQAoEHKh90OP/6YtIe
Sq13yQc3c6wyP2LFquBCdrxGAKuKeiDUF9HrRZQlGrKzCsy7ATMlwTMjumK17g+G
W8Rufk5aQW5R5PATcP9mhmO0kFHS+ESUluPEe1nYpsAwmp/YU94jExnzvLows0ye
dhitgujACD5T6k23z0EsxgreAPKyCn8mfgLZ2FaNJClhTYmRLEVgHgLeqfzai3z6
/ft+MNL1LaA+ThHA6MEehJYzHddJxyZFqs2BI9PZuIqKMryqxmLPYftQQXSLgBxd
OMNz0zxB9YtN9NXBWIXCwL7w5vFreuJl7uIRz4wNGHMEvabts0w7/q5rwuX0Hn+H
U+T4D+ClBSC/4whl2GgceQXj1tVLNEf3ShwtRP8Lco0PC9ioIOhMI496yDIw0aLA
GvS0Moqj/9yF/K5Fy4BVM6yLnzc82F4eLjibTOJQhiOik3Bvnh0bNq9Cw0kaFuEh
2KcHOldU03DdCDwcIVAYFK4nqYqagU5PfnIYRnY2smxgEshlacjAqFfWoz3dg2n8
YuI+JroJVFTlkI8tkKtkusInJNKii7SKDwPZDW0A0olVHEqbCCbIgzty51INzOhK
AQAHoo8NPHMBg7FL3FdWKVg86PiM2p9sjZMqv1+jT2YaLrcpUl+fZMhQ16+IN2cZ
l2ya02RUojs+1M7++jYp26Z0APRa3gocigDUzkgvssU1h/83cNCCJ6ERMx30MuCE
sR15LCYAYHsgQRfhUGIVRuS3LIJoH2gq4Cwhn3FG92TydcjkEiMRppyX7+Lk4Bxp
SrB9heU3VH2BPovNKTmISw4PA7Np2GABBPToie8MT+XKsWsjoeec2V1MK5QQ56ah
BgFA3xde0dWkm4G0zghO0wygxOWHUEn0QFQAA/lcoH3/2s13epBAIm2FCjqgKVST
voiqSlvSlqKIXp4z8JHypEMl99IMtyGbToukYzFJIfHNO5A8fKZ3TeeNZpl/1pOf
PH1x1dAQRoz2jDi2maR5650UAv5x1gU8stx1FC+1S9W6f1N5tpyscbYm7FSI8iR0
7S7UxnCgV5puJynfTeGKJ9zxOOjAFMYI2QPBz1dJqVxOuAv+s8LzkYc5a7rUKw4J
6oz6sqbVTr6dE8yHypwocxcCB9h68pxTAw5ZuxMr46TeAzHB+69anGdpWbG6K8s4
K/uuyply0bUpilMjv8pO4W5ogEXhwuKREw5AyYNZTHSw5nL3/md7R8cfqNeGCZd1
Edje/vBZSuPZ1jXDcdDwuPqfnhJzVMqzTSWpzp/D30KYMXdA+iyPYqLOx/hEXnI+
UQ3TbaGSkGLuAgCUnQgVgrfMH69F1UJjH33679Kbr4lFu0mfjXW5VRomwmQlliGl
RH8KumXvDQUC+ABVQ7kRbTx4QzMt64KAumHMyID9QfwN4YqQ0/xE6P3iTIQF2gD5
TSKmR5u5etLAm8tMGiLT6k71V1g+b5aVfDDXqzkMwS+0BVRkkqXBUJbF/oYXCA9c
Xx2ZedGGkbH1s9vvOW7LXPOYKZGRr8MtgFcSuXMnnsBKSpk9CnHLsaq+4tepYk2O
RyfyNEAU/brJkmaY8enK7hrMKFb8BcJ/V1DCOQWTGL5UcnZfh/UptpUxHW+GNnuB
VWU+is6wYkX5mTCp3hZnwv1VUA8gFK/RyYGo8dY1nR8cec37Kk8kcX4EbIDlTKmz
vNAgyA8ens8N2twLww6qMpk3gY6/ozkbKUO3T5zWPnrOCyv37t3cAqxapoeu2Ez2
8/Dptq24rIrSAOFZOAoj7DqQKEkekLuMMitkykII4GLXBP0eMVr40iK1+iCgN0gp
znQLlxjiLLVvitjNImdC1v+5AWYVphrqCVOHUT7+T9NbYY3FHHxl62a6HThyRExg
NRdu3qz/eDHzF/0VsEEGkwOw+NFKwPtghjdvw2F3a4M80BkrCvVBIPV2RtaVuVlY
M6cdZNaay2j7YiVHIUdbeHDbGaS7C6Ri/Vh4eJqhxZWX1/6k8fQIzMAN32vBZ2w6
YFST8L4ig/8La6ziYw9Tv8s8lWta7SGCzMeqvVznJa196YrgrItqRQowRmgK55M5
glsitecwEo6R3wgh7+cdNrBoq7B6BLr97J8OqHPqkwXzNfcNjMDNDM6AyviYz69F
uNJrYBzvSkBy8Z1TRdLog2RlKoCpKiQ9LozBmp8U7FNHsU76rHDhmrfepHf1g3Gy
qErlrBAMf9KjUnbNJuVSQdIMizIi742i7Mhl6MRYWsv2CYpomQMkhoungQ5BK2Aj
vn/1aKe8i0NP7BQA6ycIaVqAQJobjE+LOBYvpIP+YeoeeDYl+rkVdO6jhCsRza0L
cU+Oj+gI7zsgpv5lPzBh9xnVeEVBfTatKHb9qBfe1fe0jhQakEkuoYMCKy3O04om
V0eq1AtGh556nYfW3uClFDa0owNi1P3cJZHKi3XcybkVAbYkmv8O/SlFZuoQsWvX
XEguFKO5TaiGZiHIe5y1tSUOPKSvz5RS1n1iQQSIeiljskFl9eAqQQgiMs0p4Tnv
q6jPEtzxMykOc972AHFBv1regk2BLb9L+lasd9ac4i82gtjJfANw8/aYfh4tLCdi
gc3B69pSd4wey/s+XCJj94NShHkz55MqbCjOFCD6D2KIOSBps8sGo9PGuT1yUk/B
jbdEejR4uhCoiknrI8n5AgCr4q4hPiiTPUftl52T6fme+3hiN6MA17u6o069Uh8O
e0zAhfBq9P++hzSKyLEXfeSuYsnzeyXzh5fN2GYB6AaQOWjgu2bd185YRx4n7Ajd
VIyjISXxae2JzBCxGVXr/RAxicA0MoRNiIRRhmM+vzAGmbaSvm83C2B99tPGLiG6
u4C/hDunUU/heKxmW64n/N7BnNoyoZNht8NjS0Y4ryH8Ab71lcDyDo4OqFXg7O0W
ORZbpD2hrodKBA1Pwc4BB2otct421NtdFxrShQvHUBwQRuHjreNiksrYKCN+xmXJ
O7nPeVP5gE18Inz4FurQjVLQO93G2Rqn3G0sJq5HrryVaF0y7qAPJ0Xb/lYTX70M
tYFB0VpZf9tOG2H31cQcGN41vuFQDt/tohAcPlOhf6HJ4vWpheWhswVOYXpau6cc
c9t6UOe+n1szdcINw2ORgBMF7N6X64cHWZPcy5R4IF4BTybt//sT2HNOL2betTOm
RyPcwrGttXAOHRx6QjOyQV3LqxKG+2WJYWbtR5sB58zOO5gFjYGu3RRMCyXFz3W4
RAbgjpOc1m7VMiKiyvzma1tS5oTJjkqec017snmZTXu3rDBHVuLXncEt/xYKLvA8
6NZsA93bH1ryOHFuoJrCWD6y0MizrDWCMsaQFshOPlpU5xsCFIGAhPZq6py9FFgp
4Bs9RnecnGgBcuD0ulR3MdbVnGAXdT6/8piuTpXplW04TccTS1yKYZg6sqiX+mLP
NVGpQN1SrRxa2mnOb+sy6oypTifV7H1u2PVUkyc0Q60mqB/Fmce+p0PSWpEPSzza
9ocWCrvDO5kaTO9pddM1fjRq9C/DEKmyFLt4kt5KLO2jp6VoOfWHEAfD5JXk5/9w
W09MiyW+UbjjCDpoEUakyrucvVz37BHMBEx1GO3G2hDU4kzfmzp/N+EfM+V4J6is
CC8t+DrKNSK4U7NSb7VswUubFna+Zm6eyOmKefxYDtg9klqMyv1vI80ARM/rIPm9
sqqpMqgvoF92TCauyAwKYL+JFnMOh4HiTVspfemV3OIx2Z2zhDLdEGyVRUhmyvSv
38luyzrIGLwoohuRimvbcx2ITE8h0tH4M/Haz2tiKTfPE35fodn2FZ4gEwRrVnqX
cQdg+wZCvlQXqcHW39hfJjcmKNLPGdcmCcSKwaEErEn636vKS/ITywOOJ7hNAA2N
3MmL5Xukl0Ea9OwbuckoHdIlFNMfy+aWnRQs65hQcDpDKpdgkuGkVjzP3pB735+i
iOrO+M37eBH9cCPCTwEy6goCa6IByHlx0sc9ljuW5rM+oBapOHo2Jmfw1jujx0RW
3OHRT7BF/VlmPoiXVAdsaBEnzVF1Djfl7KEBO0pAh1rxhD4YXbr4dV98WF0OyZia
e1ZeZ0FS8LhJrlyuJ1TdMAtPFITiCHjR3/PX9XYqi6SN2oLW70GA9ZhdB4UdzB3M
52LbwhM0FkE7s1Gz2bcCub/IhTUt6tVuRug+d528HDsKvKdYWV0g8fObs6keMpgK
RvYDD8Q0wnP8zqUP47QQIAzdhp2b4jit5xWzgduK5BAxkmMcSMlsslFP5W2TlMG3
8t77dG1a073Q/EwwcIFAIJdITj5EqAEYTxezwdbYhcSmE/ahaULGRTPumSsqLHHd
v7QxKIXZju3qyxICV2veAjTH4PYHiQTPdavI80asNE9J4z2FSSydos1/ebeniyx4
3UtpzmdJZgksEfdgdo+eANJyBwZxuw8pGImM587ghNpH/VBIxTGjdSqOH6q7xNZS
jX6Na+jDkABUaEa4gg4N9R2WFWPoT9PFAu8WlXCn+d7xWA6aHcd6XDO1qOGaFekB
+9VvG3T0I0xHN9PK/w4bBqn117wWIHlvSgNGjSRaCi1/vTPgdvEYtkyXV3J2vdM5
tTyznFwY1t8HoA3OZKR8jYe95bF/qJ9CIQa6slebChga8PUGfafOoYjmOyl053Xt
TOinviCVs/tpdH/EjkQOfydXITJa+mot8vGmFqcET/duDGzH0bEkrnuRkj4niIpY
OA/1Sw2IVuhbd/rOgVBWch2LMKqw5sNCOIZHB0TYP1pt9+xqNoZE67aC4TFQD8eE
KYdi+uKqkOSFK89/5wrUnWiGvREIauovry6Kximm6CteNN5umO7dkGw9045xdXPP
iU/7gTKc/t8tknGP6ExyIdkzDTv26G8PtcDbQx6Sf1YTPVjbS/DxPuz7bhMtdKG3
X8g5tjydOFbs1L6yD4YJ8K4YWQcIesOg039WRQLRExs9NxGJHfTLcESkCPFGszHl
RAQOxXNfk6FI4V2gz9QLGWKX76tFK7NbNE2AEXpEDkEI70uanaArmrYh7L1/b3Y8
6H9dYl6cMzRWf+TIapVsuC1djiY8wuDTCjaSXVj0yb5sAmWvOvTFiE0+WaX8vSkK
IO+76oboicd7+04FClgmW/WzOc3V4odRiaHAIjB/ExdtQH1DZZ5E0sHO2FzdYsP3
XUJGgW6jw12uK5fUzrsrABx3RLaEkyUuWikeRhVrhoeiBZzwPXxDlEZaaH89lYwY
wqTUaOJWCCqt/RR+FZBa9ERGXOdC7YZN0wjomyfQAFXtksbK+XeNjrihZhmFHEqd
p5qMiciUs0xxU/mE3Q+2r0A6+h70RSX9jTkuNTnXcmM4rlsKeHZlRT8FVWZS3shl
wS/1IxsVaXpgiu/+hR+7WXZPMvAjFkyOSTEmS3Ahvl0YRRru7I06VNtiJJyx1CrC
9ELW3GQw8pYD+ZPNLctvJtGcFd/1/wALWaE9CgEs+3HmSVJo2Q89mdzi8XulnqSW
hV1eZ4K4MBVXPdzEChZGZG+tQd2n7TIr030aBjHtz9pjsjEHyVryn3OXskFQQE9b
FVtWniz8XO72XpAS15GfJZ02iyLd86kz7Wsk3Clk2JNfeRJoBiar2prtSFff6AsG
7KHS1zmw1xygsVodzncELiAmQGD3CxtqFWcfp0hOeb9rl2dOCJqvp7iij7uFGr0s
p7xeqOhRCpV5BUK+kUVDrBv3T0lcSYYMVC3s8eBF2nd9p84DpQjVAiGgmB23bGIW
a0n73EihY+V8v0X6rM+FtHvUsVyRDj2ahI2m/cN6oMOHKacXmjTfXRU1pnd7/8RR
0eNO5VGaCE+bahpBwJBVIDgncCpljZ8gSe8x9zMQbyIWGXQHTvFTlrvkVaDFHCgg
ruDSuJuR+quoFdaoW3AQOHpw/fl3pzHty8WQ7qzTyffRnEINzUK7oI14g0NL1Jgk
s0KNo49pB5W/CbbTev8MzF6uS1cGoWZn/uo2Z5uNBZZXeuZ5YzuHYRJojR7qWwT4
8LOLS0cfHdCHebZ1ZljBrgIHPo1M3LSqri6SQv+kOQvNPWtHKQHdOcekbXNvQugT
GdYOdtVDgNFPyuJf5jRWymPZJsopqUFakQQP4fNcr7HGP1vssG6jFhg8mD2LXdGP
l7K63NXJ5RAGQNr3iMvenM3YcDrLjL+stn0/8XG8EIxtdn24WotlyCQYLYjRAkLK
Ek20y4UVp2KT7n5j2rtrQe9M6DtJLmIEjHDR89T+JRgHZvsdFpT3NiiynyNGEzGt
lQqO8P9qwmGB2bhSql5uYuqZKVDGUeXOwuDmpSwJrbj54LzYpQJbkgRWSF7uao+E
XDsqvsVzi4NbQOdgvP8LOUL9EAkzA3gE2tvTsgrCa0DqYGwyl4tmFra6d6qpumG4
/Mz1aeJCbKyRCEe7Eszv/SlwCpvKQZso7yorxXBx20HArquc4VUzwQsOGg8z1qxC
hNN26vU6pSvYcaa7nR1XuzKrbo8ItgFhhxP1lcrkXjOOz3ihNtmZaauhiP2Kv7Bs
TTR7xt1fHHdqj31/wsEUSHIM+2ZDwSZDEeY+mPwwTFaOpKsxIMnNILsdV1ISslC8
nc5Mr1jv4haGpbQXZ7Ly/vjxeU31OCIKgFW/EV7PfLhune0iodK6KZ7nbKDwyS7q
3q/Q22d57iGQglL36I4KgOs5f5kngx2YBm8H/4qMOQ3bqbcFUXinsTKSpQCKlfp0
EYthi9K1BvnIVeNw2+CMVeLOHW4LtwTcm+oWDHgtVo+ZimriiISINQ8lSzuF60od
HNKhiTyARvj1o0L09bR1gCccPQ3VfE0SJ811ycESFhcwB7RCXO5B102aatkrYz7I
KJJy+A6wJ6mpgqm5jaeCGRq0sCjs2egE1AE17BRsmNknFYGHvpE32oNE5r5AwCpC
VkFVnkYhtkrKZ07Qm0LJ8EOEFrvnusVthEu1MDAo/bAEF081psgafmQpbXJp+7tj
FAIXu/UO5XYxP519hY1oZ7H9wogldQqhVmSdVtV84Ckm4vrI/mH8ITQWeTPS5Atn
Yr/oa03hdbHlLVTDKXqdkUbuB721PJUHqNvDs7b+os56BKFXOuzVkQ5Z+tVSL90r
/A0jOjk7LhIU3t1pL8JHshGU9Fxz+U76tp9lo5LoaA68bVoElBRpUop4EmN59Pw7
ZgOqhUoiLDeo/0StpyvAIv/FeKtK4rjxBfE4R2X0wemhgwQiFkrAuAAPhWfnEECb
5I89qhjW7ThJIPj7qFnbmkWTEWdz5UqkQGCITq8gyRklLfahl5FPHTL/W/fAyMZt
2i+buOQrYsqP+jgf5GP6vwPCGx/Rx1ZJo+02BRoMQf58ivZD9x/FsCG1h+gRlwH8
Xm7D3x0zZtEIU1Sl0ejPBf0eAhuriZb7YuXNnUq5APXkdmrIhhTI5gu95I7qc+qc
cJrGmFAg/cGS0pZLCJX8ek7JWgyqvswNd1lcIp1teZj9g/JTAziHWde1pcE8e306
FiQLLbQjeXvsMx7tEBIlOkEAZ/MfqMrIxFQ8ckiKqbGM1hfPL7og1y8iEOvFE8JT
FhuCG5nPXT2hB0KWltnx7CI7nYANV2lWdxVqaJKwkTQ5b3ntn4IhB5iJwqlEQdq2
urVN9w6f4Cu4SSrk0rw+Wfoy3SdQCefF34vnGmDbAxGciS186nUJs2K+aL+WhC3m
L23z8x/OEfQjeBP4Iz/tT7V+o1c6OvCzCDnfW3somguA+Jujt3j5305p8bOv/yXg
N0oShs96ySEaC+yXhj5LMDFWYH9AI0qZch/5GBriyofqXv7OwOoCBLc+BfVaPl5q
4vbgBUUny+bQFL/7iTpgHKn2dee+I2xhSQRyEy+9mPwDhSgKSKUQNk3mV7ijQDLu
1DTU7gHH1FPlwkFMPXOZkCEcaVnvo9Ek7zHG4IX6mAf+syJA5962A+uolpAP8I+x
MFzoPzVjBgb5dxOA3h/HXev3Uc40i8xvQ/OdLRmGc5N9mu+fkm0WpiREmDRLMqlH
JCNWUFQwgxt7zcFwEblesKMLJnR07LF8cao++mWmH7i8V5WtkQApg9NLMS5h4zK6
HrcLfzfQu/qhr04YKmkkusKBZ7+JByaDfjvMGQ+YJit/URoTSBOU8nT39tOS+bwG
mOaoNLV0fBNJBJLVO+QtwI1JPCY9VNveHJtFvt+h9VgL5zZPUsPYa5PJE8D4DDx3
7VHaTizm8RY5IGoCRfm4pND5r4VfANYBY+WNs7plQfiBIq0wsQ5baCR8gFbqDlE5
m6DbEXMKyPgQJHo5zpocq/1Y2pj8zn1RdLFf67MQPs/dsD3Ii9imIR0UZHSdD4zj
vvGQJlN7CWgc1f+2JT33dPUB2oB3NAwYUSZq+p4tLPXlTfNdxnJ5+1nV1hZrqCFy
Zl7e5r7VyNaxBEuPYXyM8rAC9cT4saROv+FN2fkikMVbq2vsfiixgg1FE/G9653y
0eq6xrzsVXwXTJ4/BXZRRlO9Uu3BhZ5CQhMgHTug/oDqjXtSPxCFiX5adBf5wDt0
4BDbpppDCYI8k8y1Ya9MZUqfLvg/PYgJnPDUYHTydDz1FYvn99tThV+s8LI3MH4H
IJHizGUcvg5Lj0H7p6BjJBfZFzobde+T6bW3wS/UcF8nzYitj+5w3axqm7bvxG80
XD8Hq0jlA81aJCBlHfOtX3OrptxIZG4o59fkcUdcXqWrjVN8qDe8QUrzzVXRJYnM
M+6Txt0xwdV54UEiJCQl8j3I1wWOnXFvLJ9wir3phmIPi756IfjXf1E+T8rSsH9l
x/1uKM6CuRGjdfS8/7u5VM+YKqSJ1d5CCNKFoT/i7yZRi6xyAU/Cg1T9uFfkn0Y3
lRjY70/gh3qRt76ewOhz26L31LqcdB3AtcSv4QxHTW2VDp0vd0jYxr03uLaHVI6g
3IIJp5ihj2F5JS8a8OMwYUuFeoL0NiT6Uy+Wgc2Tr5DVgyoFoWR45wbUsw4C5dCn
7cnNyFqUPtiTF5pGZeFWS638/WJFZAxF8Zz8ejj3LIj7oIyp/AeFVYVeR6d8nsTo
ZqPmI6MBC3QrusoxjXttRZSYlOxsPwvrjjv2apamoRc0itQuz1aUCeM+Di1x72A9
QoVpXT9F/k7XDbpgL45vYtAGD74jYsaloAE2/j25U0p7a+CGh0CtdgbyZYmQ28K9
vpQlClQ2nNmg5Mj1pgHFAbglgPnK5dB+uiYWuBM++gF6HFmfoze7esmjaaXmQta9
UibuhtEOAj8g8N7lvvEtVyxnnVIoqhBTx4bFnpjU9GZH9J7RmpuEqakSzn38Upa2
8JNVSr0BoWt4wbQSLkQfCNFD+W46lXRgE9IrZka/uEa9sDe97i6NCF9v3HPx6zLl
2snzfhhh8jr1SLt1Ac3EmijB1GwZ7DFSoSSBKV/sQ19XnRSq0y33UMku2z42JBOD
7UHwhDyRcOh9P7zCPRn/ZLSxYFw2D0tJadheA3e9EG1suoUyBOrDaY6joTfjF20o
sNR6NiRJTWaPcQrXhOoCRrlNHtpNu5UfCxoNdP62cYt9m/kFcgr6e0xwcmeBhOs6
ZnFZGG4ImTFKGqvEB7CsoQgd8YXgeOUzfQUNfyMNO2EX31CAdYTPzkp3Ek4VvAgm
JdikcmFulxE/J42H4/xEUJHYnW68zS0eT1Om/zT9Xbas1Py/7sdOohJi7dGm5Dv3
u/ubUW1ExLWKj7E5cgxCRorIYkKYWgt9gS2FU1Rr513Q75dCa62y7vuR3aacloiG
SCmhS9yIgF76SlLnLPPpyt5O5eLzJdl7ASVkgGzf/NYBmV+F0EBdUsZ5utu1hAnP
hU7Ks2aBxltQ4W1HHYxVcP/ooeem0zwXSXM2iQJo/Dr5meNA1HidHtHIMzdMfOwo
va1y0Dvwb3EA+VNCsAiBnnxxnFq4ApZZje1YkbxtGXdfuL5q7lmhE9jq95ORyLzG
x7VzElrkm5YeAUHyy36iAcp9z0MpYmSsGAZmFpgB+zRLc4Fe+WJ5PnCDVW7PJ9Q8
K7JaaToJSQ7uVKqGMbg1aZBJUeYymrdWJpVxsL0VlkXUR/9nYu5lb4j5G2luemUw
yPDGBKCrYYGsG1xXsAPHwrfoDOj2AppocaRdAVeY0kdkVxz+Ps1msgBHosTvEyUr
JpuMrH83rBcdtKOWfl+FFcgXdKvPS+yvYG74jovVWGmp8w6YCIcp9IgCo2dbzI0J
RGC9tn5GrOBfdg08euL4FY/oR/zGDsNVnjhyA+NSMc76tZFi11ORlBXr+B2ewp51
Io//wt9WeIVTgG+hegePCq06tj53Qy70tnSwA5ZxpP4aNUOXIZwMxp/VoCf3nIIo
ZjMmjkTlmN7cVvmXtY2Myu9s2Hko5m5xpHcMA0PaxgOGcEJlRn3t8t+N+gMRjeWE
sqUp22V09jCmRwHB8/XUzl6sUwlQ3PlH7+G9K0TW+/vGFxuMadKn8FrHB+m/Ntt6
l7/KcP4E49ePUqgN2wZx9rxwPAIuUteY6FsWOGeeKWiFoVN8w0Ysxe3I4sLaQaiC
6Wm8FabYakHnwUThfD9Uu4PsAH2JTL2RyhSBST3fv4/SRezzS24cVPt3cnsJLKJ7
Q27WPyo3qpxW+R1xvlByeTxBvkE3YaHowZ+ZZm6hLLxyVpy26+Fd7nLK7nLJ3WPv
LjyDQFcZHQOvXmESC+2uT8xlk3EU1O8V8sHVwpuaL2imU6b82OwplIO1SjZxBZAQ
5VWd+SMQ9FWDyBvUaUEY4IDUVm2iU9nmMBvP560k8ywzXtS1K97kfK8lWZ4cGZq0
xBvt3/JMumzpHUwOfpJhTTo7JUduRDoFZvEiMxxO9OuHihHLTLSL44pUxoLei+4o
Rxgd5nJtBDlX4wciqZfTshe/irJD3KWLs10ZQBnPhl0zm8thsHdPpe6SAZYDAj8z
TojUavQ6Xa0rLJRaWC786fl4WX1zeKk+PKD+9Bqb4TYqxI3Oj5h7tVVnoIpiEWVz
GVc9dipJiz5kF5xgirJwcSxd5wzjrtn5HVG7xqt6nI1COdeFg7VcbhDZU8dnOErh
czmHw8Kz+IZvsOuPLMkMQmGSEr/HuL8aCQmyH2jpG2KdrK/+N+yzjUCoVK9BT4g5
O348iHrPzohpEubgC+3FmLH9tXXiAVltBBumBS4ahtSt9gBp4F3sUoLeEs2CiHQA
n4CKeahkVO6F4TRStBH3ZuHrQiEsfe7ZPmZilZ0dW50LD6Bh11KYIgqxHChVBHXI
Rth/ntUcL0n7HIbRH8L6NUrznpRGsDhsUQbilhJhKMWQHuEKH6llbENMNydSdh6I
cUX3yRXEjx6263+7FqfnbjV11uH/p/+nm2ayCf42CH5yJTPCgCv0Shy1+OTPY/Qz
oQI78DzFXklJcCqFbaU4UccY9Rks1aDjSFJ+PRHokQ7dMKinC5N5o+smCJvTYmtZ
6rufZZj7YnKZ6A7PqgIHSZZIIUpbfPYyY1rSZMlJzzQhYKUmUMUcu58kEWTtVKBJ
M22LTEYtky6HADf/CJLo0r0SKQMsDo/cLdesQOv6cKBD7uJ3w/CyHDdL2HioRI3b
TOlWZ3/hSUnjrBtiJP83Sz58HrChW494pihbSjdgDTiIQCv8MkSTWmOkSJXLy05k
+prcGSt96QSvmjNlb26Wz4TfHBLWvRR1DBzPVvpjWK1JYWx2ERPOueooYsWO3Yna
Psqsb++F5UxJDa5JVG9sUDTPMAbS11IGO17YSOlv29oFnd8b0ccOzrXh1pENYgjV
DNwu8nJk6hY8qn9AZ9lHwMwLtKABR/i872Pt/gUwVx8Pz0jqp0bgYhUSfOB2ADLE
6H0zqnx1Dl1gL1/HW9R2HCmKV4Km7vcwlpTCke7UEZ22p0/fw0oih+Ni8YWg+snT
EKs6C3KK6l0qWdOS67fZ5SJVzAAbxyE65b4Ipm2ZoPcG/v48DaS58XcnmX4c8HYX
4vpQQE5xDRqGcUddQclo0XQC0RRkfJRZqUfdq6SN26DttNDQe7TO7mZ0Sle4xMhY
6hy8aO8P+/KZGUaUNpl5RKECLWb9SL4p5bBoGWsROFMgv+uKFZ7HTAS6HQeJLhSd
yLkMFpK9ZbQ73qV72FvpXqhconHnw3OlA3hpv9tMTV5p3kim/n3y6vN+kNejAsUZ
X3vWwPaSBSwjE8bCJmM5xMKalunzXFx2NxaDugrewNJjN7Ul6rZAC/EyybNhHch9
Ys4sSSB04+PsEDDxniXNr2SCmHoMSJaofKIurbv6gtOw9X7/LU44C1a143cg5wak
pD77Ns6eHCE31+63pyyI7IXgrMEBGKy6ub5iXRjyI2VC73jh0fTvOlNJ6v+nnazt
uFBvdPvQeDSNQ6pEq6XnDOoN8KHp3sMtiLdfbWIBqNSPr3sFCyFo0q1CS9mVcqmZ
+v7qeDXSz0sE9A79jSy2hPIWI/nD3SZq/l1tiSF3suuMTZHYD4nAg6KeuSEc0jG9
69WbGWT1tZpRv/df8T3CQT4U93HDLN9TbIK2x0pFhV5N5v+Mio3eX2NNKA9k5CLL
n3/Fl3HDvf+PrUlWtPjw9Qvws5e7KTyHY8tbNAbx9LyqmZ050fc3aaLue7Vzj6GO
/52M/pnDloHMSo3eFhXgsnREPPNYqNmJIQSsOxuW/LGZm5ncAeMCGrYv3Li0eZNh
+a1YDLVdNk+NeH16IS7jSfQQwZN04aqbdWg/wb8UtJms3WlobS5pqn7UZyd8swSB
6tinuKhuP2tn8A3PZSfENW6nOSih3pMz1CkkrgDLLO+qub6lwsjoM6aMa1OU6gMQ
QE6lPVaRSrLjuHPIxKIGNden1wqhjBPQen2sdyZspL+R9wJr3w8tBczXjsLDUw7E
KdTsreSqZOrgxxWDpFkEc0/UwmvDDj1m89VglXjS1fbs2/H6g6d3PRxFYdsd3C82
SrDT52WVMrBdIqV3cV8NUrvEK4myMn6cwNQiwzTY5WqP4MZkt62lysnh9rcXVodS
EfyPNXb1bUaRCE9K3SGnVV2p6YHjsXuT9B1+BIurkLx1ig3pzFUTZoxhAx0JC3aq
2VfVfPawT19StKL9mT4eWL7j+J4+tU/ATD4E5TbTUtXVtISTsub+A+zp5p7vJR5S
D94EuIf0DJbXVAgLPResgz1bpnYMqtAo4r27Ja8qF9+lczEjMcKnBnAMUCXMHA1D
HWnHAF/R0z55uVEVq24aK4BLB5aWAxkx9ZgdF+5B8eS7PtGHxtx64cMEgepaJehd
POm+ER2WV2w92jCdt4qeivh26vkubouY3BtJ/OqBJPWurCFyA6efutIFkHd3bDLX
qPnyKVrl++BeQ9BlFbBlc8S2+ajy3bKOCa/VWMEkIiFp2AawOpYPQs9wRFPRKWnJ
68+GyH0ZKU90muhFebki5wFCqakr4F9iBgReFRpWfIhNHNr1VHmo8JA4MOB/65aH
pbo+f1tEMzokNlnXw5TLBV+iyu2PG9JXbBfmOhtXVxIRFqj32dNP0zmashTe7Sm3
fPogbrdAy4XTSN2ENMSdjRP8UF0caceVwIWMy/hBgdwRrfbxIhLplvf8Pykido9C
Vx3Nb2n4YZgSMq4vrOzCctGa4DT+hn2IIC1zRqYE1JjqQ7xgMMH8FGzfZKtEoLrT
VhNgmoUjEAlMFEaVNrbUdQFXgi2BGofivNagrLO7RJix9qmWVFzEdXv501XxprPX
xhRB+hF7fBIdviQbeB5kgmyL5fimy/s4B4vt1y/CffqWJoGIns7OteZ3Atek/L2v
yrd/C+YVueOnaYSuZ5y3wz1jG8SgZJGq7PN4v1U8bQQ3OKlXq0waOm46ML7CWNel
IHUxiZHTyq2FXGQqCyPgm0rX7Tg/8fZL3IMW2g1wtwYEd+iOZCChK7kz8sZIgJU8
Z/GnkT85U5HlnsK94UL95wGwXjPnstFjp5JnHKo0hO15krfsxu7+Hv46SJbF0csS
z3L4HjEOBRepyFZW3H2/nrdRAWzdBADh+e48gzL8uZBL4PZ+2FNjNLuA11QdCzat
GhyaN7hx9/YfFW0Y4g1m+0iYIGC7ggH3t1IoLG8pyrl1AvJz7/uRpAgZw6X/rHWg
zZHzd3oAJiY1tkrodTpK+jTUlgDhWASfqgWgSLO3z8c/psmpOoTx8pV4Rz83GG8a
MOuDwuxL13TZyh89AZKQwImVFJ72tuOhVDM0RiUY04YMLpl/6r/Swl2q59JfcMRT
XhIufcryoa3o9hgTLQZsdKZ3nLklEz6Q+iq2ym1GRKq0L6fpa7vjZ4b52ov0Qewe
LVUaZjbp44Z8xgyZ1MRLgeT8ygwHSGJJE18o2L97FP/JtLhh2onSSlet/qnekiq6
LPgrg/qAIG9eOdy/+3R33MZe/XjW89y2z5W4pd2OVmHRa4dsDPMik9kXF6y10JB7
06Jm7V3PNqf1SrpIZXs6RfLtVK8/GBi0yJU4K7nAXpIv+ADA5Kcd7HMsjxsrTUvd
GoSTp29cYfvA3tapaggkhQkGcJqdIYcThdxaAsaC5qsn5u62r5qA4+PtwGynvNJ2
aPcONbJEdDYtun5mwEcVKzabfqhS7PyJjT87rtmcug+6cRTd22suTgfgaXQQ8PyI
xG7CILCpTKrF1qmap7Pa4mqtmw+SVlkUKz2EySOyyqttfxcOfGKkZCoXlyFOsos5
xXFOPWaSOut8E8wGzLeKejisrcyvoyD4+2tgF7bIs9867zElmRMDz2krceYxC5Aw
0LU55T9f+zj3J4Y0u0rdoTXQU3DYGRYKNM/I0PpBUVU=
`pragma protect end_protected
