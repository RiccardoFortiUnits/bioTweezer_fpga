`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
maIe+J1laJ0NA0rYkuA33lzZdsD/s92JPSkK/3658EAHDlBJ0hTCU1x9OC6KdcF3
BuRL8v2VcR7kID6SHNMzx5A8oNOCIIm//z24PA2BUfrOOf7viTV37e9zYy6jD4eb
92kNiwRb0c0iPS6rYFQHJVsW8LRL9bFS8apj/2Hx1Pw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3280)
F8Cj+lg5hnhS87uz9l2sBgVmKEHg3+jDDo735RmbCUCxeFx57Ra85ZdMPgZzgufV
5kq5+g/xTdR6R1mjoGZoKt2AFHNexfY/91gRK4HeRhzW+UNpAeOHhX7OvVg7hc4U
5A1lOmM9GCWnSmMHD9FTYv0g8gghDeUnlK5U5h17M1SRLycvwj+YEXRUZNlTWtTG
IO1D8CO1CHY+XwrpysEG8a+hROeQTlxYfGa6K1Sb+HZ4xiD7wD90LYUKfoskhdsd
S3hSSPTxiLlaOWsRU9CRlU5tUn0nN7xqIB5tEIqMoLie/OqFVhZZH7oaJedw8TcR
7B50Da6jl4qWY2bClxwwuKLAy5RorxJbV84lNrB7waswezOmQPVmRMBXIctIVAvZ
ISQj4+eg42O6+emeyrEZbkWwizAYuXuUBfU5tsqy0nbs4p21pXTuNRRgDRla7RT8
YFe2MGTeamxwRrd+AL4GGmXlicocJ+fZzxOTGCuBFeE2NcG8fVYAr05N7SrX/YWc
mWxPW8uT6znEjGtlLK23J01Ge89XT9d9Hb6tz6b0RjHEmi4s/zYDFRjpIJhAXvWl
VG8YhZoY+Qh1f6BdqUKpKcSQqktyfzWmSDGkL7lt/YqcsU80j4hIOnvxGLlJzKwG
/bWPO7WSGcreX/5rsnYe7rp1HM7/g2OEBMItyJ551XwrG6gfro2csZNC3zENQCtK
BtVOkcMfVlyOPzAC42he05+FNOnTJCJ2USjXGvIPE/xjRsIJZhOQv0Fmbq4+jNw5
+aB2pteWl2r1YfaPhTMkyyEnGv56riA1arNp5amff+avgtkpw0tgzuL4eiVx4lWD
vPgK1AZBNPTEei0hnIUVAUWdQyaHDsYNGwrvtPs5ndVQWjrM7ZqfLNlB5X+Cb96V
0H5ciHuaqUtM//sZkVakOcSJIArb95Y1+u9mmVLqEqmjf1NhkYoB1I0zdRyblPTB
iNF2dNMM2JfHkM6dSRxgjAF8puzJ7sGoV+MlVKmJgkIESj9c0wEEs3iwYnhIyNYY
GFMviK0JIhGDWsskLnxICo8FktPtwMarDRJkly3igRdh52cMcob1X0EADgcvnPsp
Mly056FjvZT/Fxody2XYhuRCGMNE9zOs3b/P1iljkJHJ5PgNsiAnC4Jbdv6DqKLt
sUzO+dNePPpHXObCiiEG/n8s4dwnQJP15VXeYpLxUDiZj5k3s0PkE8Z17FTT2BDN
vaH4LY5Zv+eBjFDgG2zN3S2SuDAGFPBVNGrrxUBwNy+21nTUP+kyTddGVbGNqsL4
k9ZeIG4PPF9lGxVLTUdr/QCoGxHFGiGsSpAXQrg/OgjTrID7kI3WViGosFPG+jPG
iRgmYjJQaJdwprO51qamuYh+MvATUeHkckjRmbUL5AvngAYot2nk1skPAzQBH5KG
TOX4RwMOYGbRIhop1C4bqWxqlIlKYclncZRh5cieP2xjvpddrodRWMK7penI11QV
q0NeGB6BmXPrw33MVGFVpcNXR+HXBJcWtQ37DsGNDI2CimXt5Rad9PzxmDpulFX5
kFF/wPMfeZrSErXfsh6rQ7SKRaUJWttb7hJmtwt4hMYrVL3XZ3QLycd0VrecP17G
wluMJwWJ4HoBFcN3b4jstl60av1UM/gWJW7T9fzCcuiv/Z6MsZf7J7r/iE7VUqx6
Y06PHiibcHszkIu+KD5DsTu6wgneMgV16wR5LTtqXAZ0yprMrT0rKjHH2KPWm3v5
ZDOa/oGHxI66eJ0GFWZvJ181K/yooR02kJa15J1lMhoeX11M6DZddzOh5+qOix6r
kW44c8i4WQDgMS8o+iqOXEPnNK8Oh4EE79AjtTBHzyB8JiNXLUDeAixsJtl63/NV
7UG+ZSBIoW8CX0vgoRiMQtjFdudLLAV+6S1Yc2aO3ciBa6NiIHRmbB9/Z8qWbfkg
NeuL98YQazh0jFn2htQ+fmzfE2sds2wBSu9lls6Zkb/pa7zarFP8ssRruzlT9Nmw
oCHs4+1F+Vslb1MCTleQLRKbuq4EnBro8h4SSV7LzYbYAe1lr9FsOcZZfBuermkI
JybIH5H+oWXQdby6Tz6rRChukZKSUOu4TW0k+iMVA9annaemb2KFdrDsq+t6Xk/9
3HB7tnbI+MbwekhYEAfKv4aQwTDyBZC56C3uEHoXy8UZz0QkHnprrlZFf25yc5HW
zjcgXdaTAxfrjqycO7H2eF+MOrjIIJYiIlE3KP7N8dPHK3hD9emf+48XGatRx07h
CUg/sWul2JQqLh8IlHfmTCcQvmPkgQaoWkJUIJ2u2yqNSn4UQgBdw9ciJDWvxaXd
l3n6Hj2k6a/n1tZBy+U1IVon47N+JgXfDggnZWuX0002gj8W8dzE6LYNCd4RkEzl
ruf4Yg1flNgB1GQY3eeZQ2VHAA4pZbaRcsAEM2hQx+SKtCI8ESWO8NgzArhDQLAS
YEuHh1yOMwUgQTTqKfxW22urKvElbmxU78HkuiFXUzm1MY/FrEWjGOtQlW51Hcyk
bx71KMdduGhOiIZoxetwGJsHNUkB4P7T4sMFERMmClW0qEhmvVofDehmPIh0T/bS
N9ODZj9pDfMgnJhUiA3Yc8UqkuGiPedEpv04DtT2kfEfaHCIO+sccgpLrkRuhAGI
GKQBEzmpSbjSBrtDBduZPmTDe8IwhOH2jqNw/zQS6ykVP8aD0RXGrWMoNkQODHAb
TSlGPY4wA/8w/8xwoi5rNkXzciAMWEHKJBlNq8+lj9/gL90mCFHHd1DwkAlE2Q2C
llLT4g034s+Eq7Ze/DC8R7w3DanVVoZF7vK4pF34/r44z2m88RMfBlhYG/v+rcSf
9Sy+WCYAhQMFUMgYpwRCmAknpqHPdHTDNJesTo+QWolGBlqmCXUQp/LIlOzvdPrk
EECBzsbf1FglxfXjAhiX1UXEMIHJZ+nNK3IaKYJjOz4FEuSofJGCvEK7WWNDLR0q
N6uyAr9MpHXNn2ppJz6hq0lSaB0Ots6uKs2BAYj/uVDBVjEiwRTyW0vljHZaKBFQ
28zEweMufBK5K1jbDIFQXtxhUQK3xfQurVAiyZwP96YoD+XbdOepW+UgymYFtFWO
oMu72+Syr8BAMPUa1ozOeHf88c4HoX74he3ICGJlM3X9T4gEq3XFCRpbRF/WUSM1
ocreN3ezs0GdFgnsaQLX3+uqz+2J6WVIvHP1ulexQmv//Ue9Lt5EgnEwIybgB7H7
ns1dlpheuCV7nIol1e24O4hWwOkJ6gkhDZcrDeKlAs9RoB37I/O6r3w2xklBddu0
dM7uHgHzpmYGPIXLJcqZRAF38wSRT3MpoCdr3pcEJ5pBLLzmz5j8JNGOBJveKhiS
Q7TMDZVxkKhDzRRsdxCQhTGRCkXV86UQc3Z5I6yl/dn1bGyR+1yRavquJ5NY7f9j
hYep8/aHTVbJVka6HHllbopgKhposLBdlewbT1H2sI8NzmvHltphtx0RA/ufJRyp
RXhksGjkdK7e+QQhjmDkjBPUCc8YFvRaxdgrxrIzbGCSJP/eKKJZ3zMkx4xlHkSr
QyHoLwi7a0iUMm9HdxF78Fc08SvXGH9kiy+1i9HR/h/UVjtju9Kg2xujLJPiH6Z7
HiivixPPfZ91keKvf9KKyB8Oy22lxZEF1jbPNTwuAWrXVTYZyGVdKdzgXinDeyJp
bZdSKhUsmhvNWKE/aPp0rZyFL25euXXYmkkRxmv9IBLWYTyCqsa/CZVKwkad51ES
yITdWGwPodfq641KYfaxDmCSrX43bBnN6DUh+VrcjRA4yA31j3W2Kk7JDYNHFRM3
rjScGiKWiIZRUZrmmVQmhcXdckCY6uYbp8OoViSdwH630bOf+83hcOyX1elbkx2S
bZiiQSm8LYCaS0JCbcR4iYp90d/eeFAtDimCX4f65HGg6++6CQZqz5w9kBokNT90
NgpPkLNeRWeIvavY/TvD81tbsZdJ6B4SWdPd2KTjceqYbIyDfCsN1vPIxUM06KVa
LTwa5AfWOeoqthMKd7wacKtsOfzh98wfEkepvOJhCcqZD9A9yr6VvCmdXV/VBwPY
g6vrks2GcsuVlAVkCAZNwwIFXTodH9UK5lbNJli+hiIFMrx4haQP3bqqRh1O7DMt
f9hBPRHkKLwgjzy3mFd0jnBSN06sxL+/rojHFQ0Fb4m71WJt548KIc0Vqp/zoKLL
7aigg0/EDM+6wz+E2KVz5WIj3sPVw9HmSyy6JZBzHL1JCLYl/8WyPKD39djVwW03
zvp0pYhnVK3uB4HLSC8acAbqOmM2ARgjbCnjZzs2StngsY0uW1/1NJcLwLIXaS1N
G/HhL2ErzXv18qZcOFRMf+viHordFEFSgKQs+lfmcwX0aZlLXbWIHH7Dr89p3UQb
Av8f5ByOd0lX0oPtqu+gig==
`pragma protect end_protected
