`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WGRLYb0Gjnitisk+YS7Lq2Yu+zC8xdz0Tk5PbVWY7dVKU6vCkfIWGDMCNodohrvC
boU1z2hznLLuxPilX4BPJJZ93pJpkWx4UgAMZDnifAVoOQjwcAGxuvw3dj4bGMPj
dwfBqyLPJWVUOe7DuDah86LTXYvWULhS4QHPv0d7F50=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32784)
WWg64720XgfGzEfOgKH8oeYJxa5FhmkyA3saVo3s1Kn44gqfZh7ilgqU3jBZvMw5
u3OW3A/dPC4yLFRYzP/jO7JlA2DMDPqNvggFMjWJgE87NuZ7VDZy2VLuXwCzAamF
xI2VcgkAlqOz4VAeci6ytFYiZJo6/92+TK3xxh1JVMMHakRvDN6txxQe3txtCZ73
GMes7eYxkgw7WFV216gwbUOtmf2/GvdxPTL4KdSR/Li518A1ofOeL+5IVLL3KYgo
TwYvKeqDulAkotBTnpFPZ9so/rx7f+y8qIe5cHVfZGN5CeZHdfqvUvEmSVafPUbF
oqNcR9BObPH1lyvPz5zlAlLqTNF3xmhAncSLfdz4+otn6/tStmpZyh2YSFqDft11
BMRksvNbAmQm0ncno9IJh/rpw9NZG7r/jZFPVt9koHRIJ7GY/Btyj0Ba2wvTSJdF
XOYCOy1Yc1hQG/cIG37Hdp9r0lcMPZ30jloIj9yeeVH7ZCfRr/awl5xJNxtMQJtB
lajXzJ1v73DhZXdwkuA30HfvvyQPSmpOWC1B2C0jv3pM/Xoht6SyKwSghJ7s0SUz
ppFlgfBj5Xigul3Ej+qVJ1HmFlmlVMR68x3m/v2Op+54v6kEmjilXtWyef7pYM4R
WTcw1va3pt9cNXVmJlpwIbdtXtAVHr+VW60V4jknULDCKWhFB4JJJzIH0nfKPlw0
RKB0w9ka0X0grQMbEcleGT5wmlGYsyisvQZEyR55m8Z58F4RIOl0hD9LPZO3qCzN
8o8110bp9i84JDp5ZM0h+D+jOv13YKkdw+XrqpIMKJyonOokchJy2GzhV0uo+YTn
y70g+0EhsmbPGI5GDDPdFxMvwHuPuQ35UU9hMKJjnu98DUPSI023UnHfouQLTAI/
NJrnjf9jcLp0wq7v9SFch7mWce4fkdy8N4HgyXyH+TieOaGGxiMjlWaUZPCzSQaI
3E38GfiyQ5MZy11NNZuzA28rpWerMQTz0IWxhR1fIQkXrk30qeBqTlxVGwrTbZzw
iMlFalJIc6ljS9fS+/xyAT1iWGAkXYJFpwnsNSh4Ixof3efbx+d301o1ip2JGRvv
YlHfIBbjcQQ2dHhvTEjRAFDVX2GhQZmWLxAZtRlW23KvN/iShbB+5XKlYFTLuYLn
lUBmQwbr0cvdoK+18VXfMeb3WEoGeDAyUQUYob0udRk089REc6ejKdB1QWLZ5NLh
XT65faO29FxM/TSxSJsfhV/ZlwTJ1tSReidTb9Hrvg3r3BmnOO/Soa5Q8b/SsAPs
xBLlL+ZOFVj/gCzCWLalxQ/jKjbIyVFyNs2eCPB1TJSomQ0nwk0xF9484PqqiS3N
lRw1Ib8264gV8vYV30+Sk0uVE50o394arBCXK9WZ4E0W0CO83w/fy9D4Q+pQ6HYP
poFAR83uGHEBvZnq/alzBInRFvz89ZxwRE9HFTPJ0wHoyNf9mjXpxh1RRCYucmhJ
Z8HJxfaJHt/tqP0rCnfCfJiV/eo+AfS0aTZeL7Hig+q7thU+oqFnNVK6A5L8U4Zn
xvpX1P4LqkCJQ5NVrzcHXF01Pq6GGu0zU3EfpkIUhP4Ti/Njh09nYz5/3gdHsyCG
3bRjfF+F63Gb+41qx/P0jkhbh1ENZPOOGJxwQPyEysAbIoXh0wzHYZ1b/LSzkIGX
mR8AH8vpyAipR/q4xCd65a0B61F40Dy9afTmmpPEmt5R3jG8m6GWShloJXHOYGV+
FGGvxj9SM6rppuuEOFAvTAtq7Q0oq5mR2EaOGYCsBgOrvGHWcI5ppcUqP7gnMCCj
RYYPsqaX1ZoqUZWfp8/gdc9KLIjet3sr3qgFN7l/9oY0A9WbFvcU4ARfb3wh4wGc
IInaP+PtCFaFxIkiJp3w5urSYOooXOx4sJ4x9crrspaRziHGkqVHHCXDE+TB+Bu1
LHZVig9MvJx64AotbYzm5B3ow0pnGqueEiT0AKUEqOrwkTFFvXu2WtPeSBm0pxHX
Cx3kb4Gtjc5Zlc/Z0NsI/o3Ya54/syd+u71Hng0X6oyrv7btNnKo3AmtpapjFIHG
LPQ2i77HMz4krdXjoGf08iFwFfpcx/BfiWOaBMAudacVDM1fcOsVXsOWNoJyAIfE
ce79b/qiWx77i8HtkZhgEiZcgOV1J5KobcFsArGElK3RMPy/OKGfq8jw4dAvKrrX
RMY7Dl9WunDxy1Q7DehiUM577YXe3mspqJFVbyoQg21lynBXhNznG5RMhBrA4qA8
b/tJGv/sGoYMWmtVhn4Utf428ug8sWPUpLXiZjIW6srzvWmxyqtWE3aLahz5n6/C
Z8Qp9H47EqztNvSFrXFxxzzsyVe4jDmPwFI1TY9teYtyKxQfjncM/7rnlK8Ql5QF
3x9kSiSE2//owNyvydGhLs3XSdILhBhylSKr8PX30/Wt+FQW2wltyI+PZU3b81/q
ZTjpO/N2eX3uJJHgL1BglLCbirJyoN6jB0p4v8k0QB9Cdlz+FSeCbI7wZ5TzEb5u
rS0u9+zdwruOvayqk78MM00Qxiwk6Pz3jeO2Z8h4RyjVI2m0J64dWw7UHCjuT3Uk
H7SizgnUBWHu1tvmNQyplB9rfAYMyH2NguOfZswYOQzq/SXoxTrizu9eQietxGRb
zzk3RcfD+3jAWUqDkwn4KJkWksZlCKhWvVWjnlaLVBg6a5fxQomCdAacavOChq/z
N3GpZYnv5sEibFgev1SX2eq0Z5APZaZQiYH99eBgVF2NN0X7uZGGgJRZ7t5wxOTp
jKwrgoXGvdA/A5quovfVgIhTzg8QS3BtihL2eOxVAyvmjmyKReT9TeQd6jJgJ141
aFheqzxl9gRhl73gszWuucHPX9fr7V+FYkK7234jQKHdYJLt2ZbL5zEEMT7GU80q
kUNX1ZJd1G6jO4E3jwdoueMt002HQP0tFp0tG/2OJgE8F4TAaEkaCA/26A8Fn6cu
6CuRzndwkk5ehVMPVS/DNgy7Dd2OyIUfi7fmkvQWjmpyIeBBaPyptur1c4y6wSga
ycvle8reM7vKVQO5bnnrrqQL4QCSYQop91mdSQdPoFTsEE7z7Hps0UwxrJtYTAFC
aVMS2vYC5txKE4pQwZsduYn1RTSolUPpi/8EZzRYIkVVDn3FO95vQv/WEdH53Hlt
W5WJ8B07S1vBFK3gFwzSieMbKYSV/km9fPzlob7uQ1O+BCfAm1rj5AfYd1IW8TxP
PM1EVayKhbKUPcf5fkSavKCnAcwxEjQutDRselxiIpMQBpiqqlPPZjAn7uI8WGoz
lwBztt0SuMCtDrq1w+awbW3Y83M3K6vz1Mtw49QTUKV8a0ZgqeeN4cT9quwzps4F
5Y9xYMg/R3GaAak0kLyqYZCffYag6vmJz+u06/kkqV4NZbLJBO/gbaUVmCtyNPOq
P0waLZi6vRZhTiZXloAUPJrSLpZFXho1YHWLUzEm/Q9Ev6R5rbnW4kKfaOl0L0jB
kvvbxhY8PqohIjp71IxwWPhsaPe4Sd5GG3sc3XR/zdXNGKCK/QKPPKnfi4ao5eQB
cOHUrY/oZ9m30I8tFrbqQoHZEZP41RDN0zr3qXEMzdYu46tmny1WILkOSutFkKsB
1jVNUQ+Qn4RdZXaonN2/eaeSpC4tJ5NbdKl3+OJoU+I3IMwf1iCc2kxDzF12eSIO
h3vCddYMxoCzNxMRRLod7yR4vZsSYCfA7yrDfshJkqBVFLTnZxyhAvEIvWUIhk7L
ezDSbPLYuSF4Wht6WWyXwASTG8K9H275JxGstNx9IF0kn5F9S309KxySOzhHJKXP
c8VXRVX/GxubYFD9PNWtR++N7HnRTN6HpY3FPLDv/ky/UEoio1n+KwI/+o7B1bJt
utVRj8I66Jl4GV+ni+IsTk4IDd1yP/n/tXoSN2CHHs9CfHjoVszymCgRgehiAUuz
nfV+GuaeVyqLhAe4W4Fdc8VlOHLeHm76UIgN1opExThSVtvBTV/y0K5OburuW9I8
6u0eOwdjUCzhxJfT3VX3bEBlguPkoKHXEf9V0VKz82WRff3Cs5ILpu5A05f5iYHg
QZ21WqRC9BmtgTOaFEXsFYA6OwyC6CKg9SNT/IzCN3h2jULzwKx60Tplu1zFuBEn
Cdw8p0w+iTDndN9wYIUL3gHu0ainqbpj3EwXtH4cVQoahBYEV5RkRhufiNQG1jwh
Zc1IiN6NZe5mfl2De6drk8YRuSMFmaDWkZv7GcGQOZ9z2llTBWvZbYtqiOIfoEzc
5weQCeCdUAfosna/DZEu2quL7gC26DmksWlRjw9fDl3klKbIH70Cn6ulPvJHIwCk
QtPm7v95Ha9wNiA7HpJMeiUGi57WAx/+yfpHcCpu81saXHduEaddTX2LfIX90OyP
b9AdOOKF4nPiY4631c0P6slKAt24sbp3hGGX15UZtLljXy0IxApDQNO+2NOqQN+T
Zr9z0DL5nPdDdiRpVoMqyWnHsB7VBR0+qdW/ocFq4hLHtG8ZOCX4c8dFayQUaU5A
TgRbKngWD1bE5NacNW+/Lf/5FpLbcY5N0rIgJ0P83EG5LHtiZ+Z9Ti5RZ4VV9Ktv
W8w7swXxQXzeJtU7vABlhVbFox//f1ZxNA69XwYyIUnxpJAKCqWb9a9T9GfG14Ei
JMdv/3MwXHJe9SvsH8R3qWIys4sIH40nPly5V+HTCvA9MfQCyTMr4FlAsJzqDOsA
jJSIYVqRkYSVHYDfXRGuCthRe5XE65/q2eAUsME/JBQk//UAMbEvEbSKzH1BYZTY
kX/73g8664GhEWbLEXPw0EAFU9KyXGqhQd/SFVnOBV9abIPx3S+lpEWBrpRCrAzU
IHu5pFhCoJyjDpJaiOwbmVkBrfRFKdiKsaSvmX5zjDY0fHEq4qJQ0MH5xWrPAjl8
4px4yw9LZmVQMnlg4pV/YjZicjhLhHCsqftjJWYPgoaioBapWEevO54u9xhbBh7d
N7Bg+AF6cS4GEMceC7QsYZP89d3xUxjSHo9XOkyjxIoCQcIjN6oMYXJTVkLSYq3y
5WHGmix3RAIysl9lYYXV/+50GSktPRaQ+6kldxtcNx/qYHYSnglHE9dAoZhMFM+8
EVlZK/QyNX6GfwHc4enm/BhQyyEC+LcN6MpfBUrBb2Y3D+cmGgnfvimparTez/Tc
XiYsf/50IYrc06+VNOvxsGtTwsc1vVpIFpMoTq1tbX87YteWFvvmgasutJByKyIP
UpU2Yp43N2mUDb2wqH6Fnxzs1VfknzGPpapPqWzFF3rMwdKNq+o0tIYMyK5krWc4
lwM8ioum87IZIvb7cAODwxfEajoPpx4E0Gulky42sUgSdF5ujemy6Vb+hutpyFZz
Ul2WmFzB1z1eBzxsJGibNGkw1fONDoI5I3WxKVEIQlHoJHgJ0jexiLD7ge8wQUb8
rKVzMSlanuDj6n/4OyAELiiIsD6IZd74qvY18IiNj6mVDb+DR0gDPoLFvIcPXdYi
WASQl5txPK+AESJP/IEnuUXuxr9JpEOIEPnuXmD0aD1gNZZ72EGodMaFWmK6NNJ2
nEdCzA+sjwVh30zt7WliLYGvXfqPdQE5nsTB1SSXiy7xiEFronnLeC5c9ob7V9Ou
oURyN9ZJZDb4h6sceMvT3e6Y9CiaiVG2cKEVd7epsfMdJE+hO5cDtXOPAs3lIRXr
mjGFo2TsaEa4gYQ7ezov/cVqx/HD23oo14bpvVCPknyxtp0BNEZ36MA1sFoOjKAr
EgqMKIHTU/k0VfU30A8rT9qVJNdHtGnQFtwh0/adgFg2KzmA6pVdYG2LHZ0jFCoZ
gb/nuSN7OcUCmvtx0ZbSy9q3DUvoQkSpqGSawx6za+M2jr3QGJBXOoQSDOFVB8Cn
yjfiOrqOgHadrxV3DFLAiAy2pf8Yl5h3Qh6D68Z27HFxsB6UolMqHE4PB3kABSPQ
M3dN4h/qb8Vpe1WQWzXyNVu3EDKzMkjEYyxJGEm4F3sY86LsDnr2ieJLVzO6W1TA
poIgMfhES8HdW+aLfswkV8n5nADlyqfbOcXF+KMT4Venjy9/LSG8GCj5m0dveEL6
Rgn1lFSaqDTVIfutiktpOhkDH/8bDDzcjVmiljlJt3wW3i/NtrHHl5zXCuX9gco8
uuPIgKe1cU28zE/apzUEpSNoTvgOI2ZL1fEOQTXdKGNp40jrFgtMMA+h718t9722
KKU/8M+o95zbzVzrv8p25dc8jEfqLChQfBIvjD2/aRmq2WgKRocKLPmLyO+zg/oC
fimJTLdH1rSwFMqI9NjP8fyh5sSNA7JN0R5+vYGEwvidW1dNfpNwCtg9aqAvIslK
7iuFqiKF5w7005V8zB40dgmgm8lRwa0USZ0l1Bgxjas0AxL4fryraU/hvo/mb7sJ
nlHKmVGllJ+oVd6RcCZKPidFgPt83ioIziM5AcWl1mEbgtmhoWYpkoW2SVoS95rn
x9EhpzjOB7fFr9i49/iDA+dJBLZo+g5DK/RXS3lj2knY2K7Wu3uA2u1MQQ+NOd84
Q42tJUthOQNF4rqSqKeLayi9vNBjtEulQF/gVUwQWTxkydR2vLADdynnKMZZP8Bc
pIsfetWWu32+4bMAD4qRrIwfur574/+RmU/El2+8i+JZ7mb2d2IbVfEJ/aqosB2E
NPDkEuU+Wh9OkIICOnkMdPPsOVn9bTOBSLiune33GXxryHDS1arClq8Y3ARr50jy
hf75YZ9jsxKpE64gR3IV03RUmZTroCFBjR+OrOTgirsQTbZh2PP0pGes5WBP+sPb
+FIdqyQqilCJeFLMCDr2fr3c3M6yWKzoib2yXSqENZWbSyPC1+FXWeaCnYWuhR44
kbLE6vFTS8Zx32lNH86kEOIvihHs36Pae4qAi6p3DDBCzaz59BztJXSFZJU1sgqL
MAU0+yw1IHooYomMG9hJgATAvugYLhEXbX2PYL6UnIWYcG44a083cZL/DCTI4vDf
u78noKED+HdPIbD3li4HMvgmS1Sy3Jlpn3jsicpwlYw8teYlaX17dZjPmITRKQZK
4vOr4RqA8zy/VrmD2m+F1SDjF97nZNLcmVfbIIy9FLB1PP5qHnluz8degTVwlEbS
ZAD1ZgjaoFTY8LasrhYmTffDUB86WpwXQZSoc2YbTX0GQ3cwZxUaSnuebUg1l3KS
vvh6Yg2gXtNLpJiGS39DEXcjfeEb3Tll2A60EtjoBxnejm9eVEY/78Xq3O91rOtF
IqQATH6+gehnaH1kGfofyjxWt0ra/3ZluodEFq4BDO2uvqozhwLHYdYSVCTZC09Y
vAosCca/My046eNkO5yy4dpCmopF4Dv4aCv601IEwDtSeDFo5/aU2rtflxxPcuKj
gbdLFk3+hZVIDw05/Tx9Q9pjAZl6O8VWlvzrR22GxWOR46sQs8FjdwX4YSKHW4Fl
8ptCogm/UdUrVdE/0XK8/KL8uA0Wr+sXlq48JvBjqIslXhFMfJMnyLbzulVyls7L
/0ZwfvrQ1qeHVII43rq+SFy3+SOtPqk65P9ywzSTSvSvxrzSqpAajBECnqQqqHwN
USn6B4GsBCnAxLYREYrbjve8k3W2NoWZowPZf51KzM59PUUoOFCzgdq/9r0TNc1K
HQCyocs8v88tNauzOaF6NPBVcYO/9zSPO6S4qvWJJB8X9qrEbjEhe8eyxCL0PqNl
xduTHh4MUmnv5fXndORa5WBZyeWaTxR9UtgF3UNOfQuxR4SwrKVO39h0Mn0u2waP
kb9A1d1Q4H81YGMyic92XFlGwsYNdBRHs9ujAI61lN6YG7YOf2Jn2z/yNK7/xJ8Y
U1HERM9T/gnA5PtWsymLJ9lB8ter2WbfbDqPkfzBAsaMOhNWQjCVc41Gq8vZ3DQE
kvTApHUVoPkVgfkWMJmGPrj1rqy2fEsRKsJUHTPeKHQgfOaXFJL4oyyctvTKwuPG
VB1Jc2aHchM8k8Krm2idCDYhFQ41sD/6Kkw84/CTgIxYYIsQH631SBVhSOuq2dLn
+yAIlgLzMoD2ZFjAIQ9Rmg9r6XqAgHfky4eKf+nXmf0Svi/SsOaxJnIxdtH2lraG
kkbaRkbiFl6KFLzQSJ4N6j13MTbEHgj5yLWgHYdmOXxXWaQbdCj2gajH8UDtFije
Cm8EyfmwMyBBr/g2wEVaH7h0XAD0Mc6f/uPj6ZxAhI9n3ug0OTIpQquDkQpWtSFp
4A08OjXvhMnYEFO0thVRC6V6pIXcWVXU06hEGrnCKpb6Xq6PVuf7Z6d6DgiJSG/w
RatZoJx63yn1dxmWMfRTSOPuQX+lOLEnU0tMOqqE+QWUnqsaArA8NaU6weYfSb/s
bpdPCUSzlbxh0mkLfC3WBQJwyVc8VPt4qvkelOrUj/RedpO64rMihk3N65wYblb7
DrVYDln5El8j7szXQp6ibXuE2N3z6dr8Vvb4+v7e8NX26K/2GrnpJR8v0qvJcu7L
pJwnRaFYrgkDwwqDycAM05DPjiB5FN5UDneIdakoLqB696lbk3uK/95EBmAYpmdB
fEcaOuBIcp+TqlUNOROgWCHpXAhUOQ6RmHFFMiijQo9R4xrWTW5I700bxV+5PhJx
joKG0ihiIbUtpIHjI61iH7YJL3Y4RjZIP/zaUFoO2JOS4XhFcMzHMwF5Coco7DuI
WvzDBTuf8JaIGne0D8YKXHPXzIxMnkum/Sd3JWOkNNPDtYtXFf482NgnHMQkJPYf
bvpwrz4ABp5KhDc3LhCTT3XoOm3hr4CEAc5CQRJMyR3A97cPLzuUVQdLizSuedjx
oRZpR+/UU3pPiq7fz27AToYm0Kq2VxefwkQfbX2sdxxYW7BsSHtwaGF38Ec22dQd
va7dfEJb3D6TFtXVPTkwP3S0p7/t7XcDRBPxP8fLRGWuppiI2CS4xHsmrc5ZzXkB
BO3utWxothWLOscjVcP7TIJA8wJRSYsIuM/5FaaknV0Qt5UtE4EfucqTPseK5osQ
SwCZ8PQQDa8GadrleJEsFiP+SN3JbPk17ejoc3Ux+pbBB/uRGP/uzqXpGLcaQU6/
iD7tXu1SSxFNcQQw0KiP1ZF+DH5TPFqNsPxePDJyMH5DHZ+vTza+lJQ4DkxFD7cx
bFf8B5Q6RySL354u4zfjV29IsZcbVdnyQtlQFBksi8Tqa9HiZeIihl5CMPTIPT4y
nnb7hwmiWsutpvWIyjElH7D9Sgc8iCPiX3hZJUrvTN6R8E0cIOphcXB+aBCLu52Q
tMFQMNyrqRDm1Li1k2HzkOA3lxUCeyug9Oguc5YOQPc48q7cCtd7+4x+/KD1CntD
oBfWoKVur1rYggkrYAbGe0jcNpZIQmdTAmctwPnMmke+9tPdGd+pXXpybAkoeE61
1ndH0Lc3QRsuuvL9HSpp50Edp5SSaA0wbzHO8MmyjW3JFpIGXl/sTvnBxiwZJQm7
5fvAY1tUYTpcRwPI6SXqyHqLDaYNKzw2+kye6HLPzQOSxVN+yjiAk/I4CxydDcbr
aj0MWBe1R7Zw7AkVfzNvEDIpIZhvl8K5kKm4iWm41RqGrl6/p+33RMGs99C/DwXs
uwACFf8h335cnGy8j2i/54qpGPJGnmvRVmRuG9DO9+7iTPzgPrYM77zqpZj2VJv+
P0a/lYlPjlUWIhLfNSx7FEXUVsMsowSyZMGdQ8q8HyHoL5Psw1LQsNNW07ekfXhS
NhrsL8N4nHaU4IoSFpgXGVUZiehlCzfg9+9ZziT61nxOLPjM2NmwPsFYpDFaNdDm
NzbtZANtUS+aC61uR/8xCq/SRY0nGrCOisBKkd8YK8gb16GFdNbvvXfzRrL17xXE
x5l/Cougt3lPwU+cNMmOhBuywkAmsPjAE0/xgn3HYnCXw0wMaOK/6RFhTqIyDFE/
VYfPHuVGx8FqQFhBD0w5KXos5/IuzY7KlXtOSjATmMSjKrkYRkXozHmJOsvbbjh7
5mU6GQXkVlirGt7Hq2xeVChfc5fthTvRAsKn1o9o9q2aM/yeiw9Zal81mFaSyGjL
MsDUewVovf5wxfgOUNiSfS1eXCIQEsEhMTdn0QtvkuJyytLQ2SqUIv/Au9bwS+tr
aSbiM1Wp9A9RRSDC8ZSAstFDq1SFQmYg0yFN6BiyCSraAa05K/2RNHa1q3lyMv+u
x3l07EheM+1jNPHfqprFSABu2fhZK0jbU4/xejDWWNZSNBzGLJ+8r9SSTLvzGilQ
QornSMNMhTMukmWRSa37W2ZUl2Tz3SfL+Oai+NXizproZWGyFUXrZasBkgxzX8WO
sZAHuz2MVZt/yqm7uVtHJlTVpasJuX+DbUn6VxVPpw7mbT2N+amYu/EBSTVmXUEA
87cNYlpesX5SiCStdyahavHtFXR/3JwTcnpFQnKqyXGchwfhIoLonnsNmZ31F5H+
H/8yMPivKDWlM7oJAMUICdrVZUvGIhvxtBkF5DNvmUHL3ApgXXNU7Qz7Flf7i1nr
R3RoxZfh+7Lj2rgQ7eFTvcgvfjEWoik5B4QLtxSw19vUS8EjdFW0dEKU7aV6A7Bi
CZjcU8sUfs3V0lvwjpb86oOQJ/xEvrilFYakgLcR8F7T6ZLB9qTyoM5UZeOf/4Lk
JRr+BtE9GYheN+Rcg/acMX5H1wiPqFRzch7P+dQtSbEeqnF83yLCdkxC9jKNCr6f
UyQQqlmdQ65JF0O2/a1skSvJhlRFlvooMDfF2OpRmkhZgBcDxK2LpXt5iSnMXjyF
ejJm07+uVN21zZzmueWs3CI/Q7+gMhDmiEDN6FkYiCeMFxFmsJ2iQTkrtU/IcSsg
XX+TqR0/qZUZGVCs25UPISzgZKoHKCJG9fK/Exf37AyHZC02ans3z/y3NaPIS7Vh
8LyrTt11oI7v4lTLC9i7e3CrUdRkmNVmI+whQYebhWe+yj7eqjBdZACcPPW4jWyK
NgUdfdFi1cwGqwYtIHOX+oBqtu65CHYLjpVvW0CPX2Uv0FnHmuUFlcXGhbJPZ4zL
Y+8TygrY+2MUmHajxxzzOfTnTU03Gm3s2E5OIH8JtGAZSq+QLcZG9/JYvE9Crs2+
8waqULC0ByKFtoZr/LL76LDEydQVuziiVaSnN2wWwn1zKMfS5Kjc/URCcvykfl8Y
z7FOfiDwpXUtDPW4r0R5A7pvicMHFHEsTH8pZdAaDEF8dYzUKDhqvAX3uurrqwsa
ysP2glraVSED1AT7mpTmV65izVS0jGOLM9ZQrf4DBFBj2fWZmqkgofXqsBmox61P
GOWTuoBze3F1fjyM08nhdm3g/siDmJqAUB29xIDbwlOyuVMJ+eDqLWHycBhm7EUC
wqTOrjD2F3i77j4cymjGIgzq5vmU8UKTLX9purGUM3cNmJPCXgKGJ4FsZ+mwah+k
J4VXFwGDI6tLpnpVqIKiAGJWYTssbO7V6vmjMaaxORCVoAgdMscPPAUrifATOKD1
EU88LA6Ez4S6P/zPmV5wWlOO2YXAdexfVr50/4PnLtmWzN0mwmVUiwaxirvqfTZr
QZ5Ara6zm0kbB9DePQ5G3jZjj+Mga6YDkJ5tPZpO3qzPzIcAhDWhgR+6VFf62Hr6
VWYQXF9l0Wwt0UXbIkgXRzAU496EOYTTLjxkvcjnpxFyQD99Yt1dKzCft7PbCrCV
OWoLpTw5lDwWQ8bhyGshD2HrlDNwF53ISDtL2lQrECoHnVknNs54Ii1yJHjmJAz+
Bty5EGLU+A5hPPJdXedx4Zm1oYvHFGtEXCpd3Flwka7Pdvt26HLocKciv+SzHroS
WBHjY88qRUQ4PtKo72Jjsi9ZUDIi1F4FOxGtmUeD08Wnmn7Y2s3FC24I7PkLy8fQ
ysCdVr0bj6ROtolmXMu9xSa8fas+EAqcgbY2u7xO/OKpXXwg2o6WD+n9U15NT1tk
9nRbNJMs2QkgErUWyljU7g4E5JdeGJThh8xRHv/YCHfJIZfziNoEtRls7iVwK3Gh
/KwqP2j9d/ALjgm57JZtesXXvZJ4ot3E4mIXfJWpjyJnyUgfjys551aGHbO8ENfk
p2+B2loqSWK+a7+bdKtXirhRjRMAobPrfuMNIDfrpblsL5dpvAFINws9XNLvWsGN
ta63QIqJtYF65SkD2/TVzXv8161KRra5BAMqGSqLbjNNPTIgGkCdJBmt1U1kRY9B
ELqoLgGdIY1B2U07WKILuUenjiLCBZYopdX3Og7Gc3w9Q718iVSxDfukHT3vAx49
934bU+Jl9QzwmjUlBPMk53kGpTaZKZ5qTsHuK1uelJh1HGEL1HhpS52MQsrfEOZY
a9MYfpJCFvQpIg516l3yD2X50rpDi0Auj1haHvahTFU9Ljgx4+6d1FX/lrqUb1/I
3O6qYz7EIDBoW76erzVSl9MfDX09ViHJzK19RqN7ICu6HMrSsV9LgMSWweQmffwa
Ju/42DiCzBTre7s46u29aGUqkc7SdSBOzVZvf4y1DMCAlsDhg092RO4HukfYPiZ7
FRgD6ak28JttfgDUyHqwr7M6oEqyQls3rW95EIzGD1A9uQ3M7KvVFvoWQWVXLCco
VRi6vNa1g2llVsh7Qrj9dM2oOH9g/X6gkEfDjbTKMTOKPprj9LKtwkDZRP3R8n5T
waij6oSy0gYovLeByMMyoFsx1amL/HVEiJ7WQnpFRIYMHdmvnm7Ypgffx9VZTv8f
sqZb9OONAHeIIaaXQYgHwOogWH5PjgULx7iw5/csQ4NNT08g1w7AOr73yNDtepQF
OcaU5xvfyF+mQURtXUmj/mCcZDhsgVoB49NWj0EPhfVbq1ZW0yWvi6wuIJ2PX5SZ
BUMsBchflg5+APZFw8kiy1q1VccQiVPU1P3PpjqL/VCO7pq35ixY2OTNBfMvt7zf
lPRoKXY0/z36BhN/El3JGdt5g3nIEuqcDu+3faCdcEgW5qBE6TwDhVSt0hH8+EdB
zQ4zSQhMB+SAfK0Cb5R2rqFMWr6tQNjzjZXwKHoh8sPH68dPu4wc0y+nH0mgc6Oi
/8Fi4cM5HjznPO6ZSqOVn6lTa9Znwr0d2rgwt6mK4BeLo7Y7QEl6u5jM5crLsRPK
p+T8IS3Drd+yo0U8uq53HBtZNEzmqbLRnZ6Npl/+/J/KF943rErM1Uh2I/u9xHgi
ouS24Zt+QTXduDMwVJbVm49hN2EydjmkkDmaoYOyr0zjBfVAGKeqREG81zkDbP4r
6rJgYcNg1ln0l+G/JiJkdW2wYdKewRby56pkGenYRzfVdjDETNDd/Tfa6zNeDmp9
0syilotG90x1W8DZK+5AloIv4VaJUG7Xpd1ye7SuDKJermmMfiUI57YKdaO0CSqu
oGVffwS7og10sxatlXFLsznbcE76F9uLyLPH1hA0kFU45W3jLvvkt5jWCBv9w+9O
WMivXlQ40vKw5XY49yvnuOu+WBp1YbRNqLOhOifDpfhIxAHsT82IHfb3tBwI41qr
P1tf/5WpHXqqwdWSd/uAJ3lttWmgiLja6Jai/Pldvzz9209RHrDAYUcBDc9KY6xq
zqIAT7bXTWkXX/vF+Wey024ZdkRiKk5G8cmAtInO3AWFUFvqa2PtwJkMMU3Kvy6v
zdgQOgIdIm3xOjn4HserFmQf32Cu1nlbl8LqTKbgyrriL2VHsAj7WrG9jjFFH3zd
qjWLS2JgpD8rHbqMYZ61tWeGoQQCdgWWaF2KS7/xXJdD5Fwn+7ex1ITqM1gxlcE9
j6Xogyz+ZgynQO+7vXOFVDZmhD7jp4MwuMjnDpzytk+OUAiarGdy+0QWA3bksVF0
SQIZ/frafBZTBAUxZA2+IPidUEt936ARWEMTvnWNill1Eqktuc8TTKUD9ID7FtTH
ESZL0VdAcu9NJoVD8adS/S6sAbmYjjekIf3eqW6n+m2mTrXza1VxRzl3hEnNOh7x
iGN6wD9EoPH0zX+wMoUZ4sr+hCYjoSD5PEgR1sQGKSn+WYepLasrBnmEid8KmRxW
fOGTaBME4Q9/maJeIAhxQvg7vzc5RJjDeJFJu5bnZ+PM0k9Rjg7GfC8Q96mSTgVl
yAsiGAYHzxCOk9dtZQf71flsEl3bFQvYbRa7dvwyGdmy0wARPJSXWekvQUxcguWC
Jiz/5C/dMVoPmMcySj9mivsrlJnLB8coiMz2NU9SARy7ha6Lc4uSayLRbALqJkba
AyGbwMUas6Fb1uZ3vFTJ6JLNLpdpKqmTikUVSX0qo0CVRQc7YmzSE2J2ICG/dNJm
s267+Qvk8tZPLfxcD9MXbrub5Mbs1x82hj/EBOLdb7A313NIClKVqQeq2M4cdyxV
PpxMwuE+rmOAnPoWbQAVfIaL+KfhZ7YmBNtRuJWvFxJlIUq/MumS+lkTyE60erav
sklytTk+9hha8xeYKc/UrS7gKanKq3lUkxpS+ICpEvGuQcJTgYDY3tDwk+ndtNAI
oab3b1mni92vbELKpTmkbzH/+DfmdIuGBycchs8o9E3syvFwNFzcz2GEXL4dmMbb
qLBvjlltnV1WKFG1MTFyV2NVmSNKU/vhnqW6AghmfnddhXFwzvcg8pWyrtXnqvcu
fYVgZSkq4LVnz4lkLPQMq7qo+AoLTMRuF9A6Yifkt7BHqodegD3O9ptyBp9ChFKL
Rb6ZefxJjLQUmWw/DICuwTebj0lqU+0H+aVQ2zyDPDrfBxzHuV+rq3tRKWbNgQg6
GnkF3NYx7aEq4juOoEX40eDDmbB9IJIWMyeKI8N90TGO4uD/lotCiTvDe4GeQf9y
UtOKLFhO61dhj5DKElD9h5gtXNr+6lYaNknNACDlaaOzHMPYnOSRITuuugpWRzI9
wesFLwe4hioZ7NAYc4lcsya9EYeX1PTTnbCvAj3EO6GIwVJuZgr8Ko+t+mVkgl7j
o0bSfXDaYlZJBp6Qai61stHG1z2KOw2PFtWYQkvy769g32MeJ7slh97XMdFuNs1M
N0jxwfdfaReNxkl2bbQiR4NyTEeg3F1AvvuWsA4oxfraOQgGdgGe3aa6J2NCMKdO
G8rUUEHTBnIi7xCo+Y1TdLcdLUSHSDWfQd3f2MdCbIN9pUIc7CiLDB5AJciDWHvI
7SVp7CmpKnduE3egt9oAjshPWXYLVHeXsAfdbPALpo8JrCZGjQl8iojGWt11KxwQ
kjopuOZvGBZSOCu28QYoU+6wIGVui1Tc3D/qjCwEml17mMO17I75K6povSkXONrm
4wj9QBjuGbU9TK6HTVUZp9ZMBJiKAxwAxgpYNZRg7yCvbXsCGYS9fz8tjkVxoPp3
0Mkx/+xRQuoEM+ZYsUg2j2yTJACpwQM6I5HNqJGAOUvUfJ3CXjQO+0N/6gIC1QQo
bCWf8n1UF44GH3dXEbgG8W6ZNlv/GbYcHwtzNL7SN/NGHS4fJp7oayUdqhP8T8RO
oLVzgxZBkqke8PNhze4L7IDR0wfIrdohg5Eo4gSUyUCffx0PHhBBHSWMHkb2kE3U
UckLZgY5Fkngt7hs1hhXC+lqqyGq/8i0BSKonr56DFqigZfJSKqVZWH03xJ5Z5ns
l+lDfguVX3gyuqtE5eqfinxeS40IWwdWK/NwNPHK3ACEjlMarwEbzPdLHNhfy+lP
swSmY1yF8nsMKftdXkt3+tifMn0gYZQqIMBtosJXt5FvNA1OoxbI1TX2i5+Yyca0
B8mXf9yU6wr9BmyJG45eWZSAT11uAcg8sJMF+jFsQ9rorccBRyGv6RlY09JNsAJc
mCnfx/fdyk2h7M0BKcN/uk04a03JO2SYiXSkbvgCYdW1X0nlFo8izCs+6tx6ASYY
zHBqe40yZwy/yBQ/BljYMS5DOzNQEwK5nQgbyJuF4NXjPKK4OtgWZiXsAGEOzEbr
c+f39gjjQeWiA2PmFFZ4t49QXJMq357M+oBn8szmAhxqNM/n8Kj+NJRHkLGKOYzE
Yui/NohYJrQPiS8iKhYZtDRMuttVf+PYZjCoAwIK3KGOp6B2ks4M6hYh0SI36QRv
LvuF/n2mkKEN6dOYsjl047208Au2Vj8m7MmQPLCeAw21+yxDH4AQXkD9J1VnWtD5
7R76EQToNfKZIc85OfWbwXpL6bI4RWrtl+8+ilIBBSP8kZ6qb/sdR6CPvANMjmR8
lfwQQqmhO5/vWqYgjdhezrpBG7nnaJS6hJl/PeljLf49aV9lQFZQUS411QOAiBri
WF7CLy9AUJhL0z0JaKKIQiw33phl9SAGo0zKu9zFmgE42l198SYKseNHCbJQvAjW
Zw48Yoi6hjM4IzPynxkVQoT6KCCHIeUAmeZxqDkAnihlQQ33C19dDtpLBJdiH+h6
aR7oG7a8QxoDilETij0MwcnMMaNlfAzcd/R3YTP2o7McVLBbJYJxRoz653l9rljb
iW9SwWg0IwZkBcoJJ933vEjwJR4XKrY5AAVjbzzRefbDR0fKrolnrsCb18rSdhpU
rpa3ixvbDL3UQ/RyuWN8hFr/1/vewP45nzLomNq2MKED2aXG7DMyatoZqWhWswlu
4bB17BDR5yVA3zJUMv59sjIiJ5ikEisOz7vb8TvhlpCSOnCIGfv7j52ppF8DR1DN
D4j6veWSA7ksYjMRHPC6WmVdGkVZpToIwVVMvDMC/SvysjTdVugBe+pTF0a2PmhR
6Tedvz7tmfiBbTkZZ4AdDEtmb8Jzah5T/68Zt06Em2FSfpB8HEh42aBHH5AlZ0pC
aOIO841Kt8ro7Lr/43NSq0kcevPOCr9FzbuTN03IDTE82jwQHaQsXJsMowYuAnZ6
pNQVgRKQa7BXnBg5s6GUAxAhNfx2UXjWwsID4DFcL9eIIDwscBrmnW87yaFi/yQD
KrmBWhGw0si1PzGUFxJe603wr+SSEWUkYZ/EwITHPJLQJjOiRj7Ka2ThbH1cTxni
KCbSkcD1TtSPEcaQZHMvauYaUx2Lc7gj9OE6rgebZXtrcREPu+GsCdI8x8ptbh7e
cbJFg3SN8HURHwKaq1Q+mVRDdCpDghx3sbTf6tzNfIphx4bbvxSeDhSmyz4rb+G7
WL5MFUazHz6LxReFHK0XRCjD7z2gV+sGRFEnhIe7HTmuNARcc6e2JhmNgcgTO+4a
dUzkGlXk6vQbfA9nyimhaFcHi91UMHhF8ggeIKHw7OSyPd4xqVdKpg88i/5hCAJp
K3Ovp6YvssYFDoEBTfyeXhQ7BIhxo8wEOPr2tz75bbXH0h3NBV8u/L89bN1a9q3q
/1vJ0a3oimv4lDyv4KdBB4YsWh2GLN+aNVu0VJbg+nwvZ5/YDyRCZPktIPFIidpo
kE5vBP+XnqeXNRGmNUWXQ208EkI540YhKPOT6BrL/fiQZUrgRdA6qw/FnMZ1vw5U
LCUp9VLDsi0pvdM4F5L+O1EV8/Ir/9lCsfQDq81g2oEAxHT8PHFZ0D8Sbv+GIJJP
tAp2azrya5khUiOyF6cKiA/AoomRtiezJe6BjQ7xqpaujSsXqhAAoe1fyuXpBYJa
W58lLGLMmAjIy4aJ15ivLJBXeRWbNea9K15Qu0KiLo1+jG0IYD+MhvPAXdrGmBxP
yFivLmaJFKAgrF8i5VJX3fldDU6ZmTqScqE0qw8B3uYuNHjd2XZO8MFVBvVOC0Vs
UCCQlenzuq+rK6DP/n9XoTg/53jKlqK7ESvq0RYjV00odU4MpW0yzGYDK52VgrIv
pfH0GQ2l8fA1jNs2omMFrnlsGeSZ5w+tDpw1FaEKxLsrl9ODCoc4BFdeqEJJzC2k
/2zU9j9hKQD3uUrWr9VOPaHmTU2jdxj4PfOWsTL5HNM+m+jERrrn4hdiFHpNgpAb
k/bZGbVmg++mpa+J9D6BSAAKkbxlOGz4yhtYfyqZ4B3XlnWT07HJqebSYymrH1VY
Bw1c9a5dkCsUBTBZHuCeAs/oXHnQ1sorY9dXGfj3xeQPIn7Hxo3cTky5lE3SKyaW
3NPpoME4hTUo/XQxgiwUN+IyYY/4icgV1oGEBtiN5grLyRw6cYSQToOKMD0EFmoZ
VVdSQoFvwy8/qsEiPFyubrEYIeZ3naXpdOfOtFDbtjfSjTwMYIOBumWLg+uQPw3M
llLaUxzjYEfKqR7YtrfW6R+QgT4zk3YhgVm+pdg1RJmXiUxReKKwz0lCxlso9/Qc
6g8vdrR10ChSNlJbNXDBPXHtkNHwlvkmdISWAekC4473wD1y/QvsefSKHMosdtrj
3qjypJ/fxLCyPA50se1fKWPtpuSQVey8kMCj0wJLGfVaw3aKyNkZZ6Cdg/BzVRL+
lXXj7VlGbEaKhMmSDKPWzQ+s5wkK2GEWbWtREA9CL3eoKqVj2XV0o5VBPMjlaupg
Oicc8tl/XQ/1gpM82bHuR5d3EdfgfTQUh1xKdkQrQVJEjzEaZgCICIln+imdol7B
+7aQlIxYCBhAdFJ4H9g5pMVR1iUErLiYY3YDRHQMkIGke3Cfkq1ltliKzyAs0D09
IH7aEnOm82qKFk1fMvnid6oB0hq5u/HmuqPyn2SK47dgVzFI6iQnIv5yOdkhLxY+
JVFiGUKieQK79FtW8flO6URAGCA2uHuy/SgtMpmnzYAxMsE0bfT6YoFRx7hCIB+u
2o9SxGdToi2hLpJm//yadqj7c1SSSf/qLSFlilm19QPvpwBcyrUL/N7/e4sr4HAV
IsViBJ8G1wrxEk3Q5FdtLHnceRYvWt5gdMcQM05FBrQX2beVHXOack2g+hPLUUhp
dbWWI87gSXLg8rYXP1xEcfVF5sn/n1XyDJBkC5HZQYt6fO0Cbx7WHzfuqMIjMYFo
pWzB5yoMOZoKfa60qX1YwwtOGLzR0eCofsMpYbEEznxFgijft4C+vBviJfJ5bPjB
tVDK8HqrcaxnA5KDkaX4n0nD2tNj1X+uMtw6GnGjSyWWacFcNK6BvyAqXYcN3NTS
cwyfnvhlcAJkXLbrscH2aVt0k327tmPzrfC8RTXHudkK8ZttG+Gxw8yrOK50hehQ
3tqEITQL/FfRkt+sgwUDXQOetVqXdezURXVU4sm/DC/Li/LBZLDWEuCMH8EU6k48
iVv3jUtePe5uH8pnO7kMnyJduoNXMA4JeuGoNhbQShbKtWcs8iBPDYlvd+J9slbO
ECxz2reEfqEigJ+Jzu1hArD8fQ25TpLn1GnBbzBgFoUkNOFFsxPkDI027KDuKwGT
6kCLskSzePNVEL/62GPxLrA75JSN+Ro0smJEl+AjQ+uGsTyzhhl4jnOT7yxXQkMW
RtIdoG47VCIW350BZVSZIqqgBG5gscH8GJwc5BgSOFz9jiIOK0XnmgCZ+r0DdVa0
9j0/9H2d/mIv8ARtFDeoVn1375D1VcmcvjB3ZkRuY/PqwDeDUYEvREg9nzPBA2FY
8cgTyl5WuNMT0M/wSWnYONdWOn3yJ8askRRpMHgVsO9xTCWDlGjbaJcOSnGpVD74
wG/U+Cp3TkRGdn7qdD7nrGrV6vgaL0q0yCYKwarM7oD3T55JW8tFwwbZx1Kz7TJz
TOAyryqgQ92Or3oiSr1sHrd8iVex/+nEPCiqZryHCfHhQWRdjCEI8STepmkqefyV
P/7PP1Q8wVClLz7BYY8ik9RcRx+JpWq9UaeqHXP4dAjTFqS4EJt/+nqOFeDhM8rw
ObSK28L1/ic3bk35Sk1AuAfFIdLsXSuesvo8Fb1js1iiYyPAtMPKgDlWdzIdRfCx
9/8UOuSea8ZMwzS9q1kQa7jLoz4aCHMfRGq5NgjGbggBeEusQRDD50gkCwP3AT5V
41rlZp7lL5ZC2DBaslGuNXgrbBXQQWUYKQulivTNzlEczyE5eVmO238EqSG5fRhq
cmumz7YYaJtKDaBTrAbbxxe8IzmM/1cq6e6O7rSw5FmnhdhG+HyElFGS2iju4iup
yThZy7Vjj3/Wz/7xJndjG2h9Dq45MMica4ICPbDu00C4NmBst68exlrqgCbZDZlJ
YLqx9LJzd3HZWh1uRgMnXhnDbE/2rQiT++WeSgBIy39QiZafUxUqYN0AaVkBwJCJ
VKdxqIHb2Sy43lJF8oHvKfdD6KaPENWzGvRhifhFKVK2HJVnvY2vb7nBLg+hvSjE
oFydOlyqS0eLU4sfATTjyKQUDk+4Zo8+D+k0lMSEftlD3FYgqF8AfBs8VEoE/G7l
zFSGxkJAzG6iSRClt9WQzmKE2mZnAh+RTKETkndHhZHBQMQ/OSFCCl+2OpoiGIO6
kfyA0/CmnE5xlR0x0AgdOWzYXTwm8Uxukis4UFEHemM92o4kQ15ZW3LpRdBGyrV0
cnxcRAxD7R+1ui7kyQ5xSFei1b/Fzrb9xz2lNpg3AFCwizMKRlWlm05Db7UFOefi
Bvmmcep3+0dWEkwHWYB8BYcclzbp+9MkbkzgDds5DI5SZ9lM+llKi8+umBLGC4Nh
jhotUSY9Hg+1qPRJijICb+YTvTzbshcRJs8160rYkps29BHdaYlt7NfRDgGAvTyJ
382Sq8omUwdKiE2lRLDCXQGPWGJ1eQjvtYhFVVWoPBEJdvw+EWy7KozDW++nlzNZ
ZRGddo7FWJezLXappfiKhPgZmNSe80TqsoijbLEGmmmFZTh1lEoXSX/oBSF91p4J
KR4qSze5sgCAVbXjI6MUj1GIUVHut0zPqAUMmKkci0Bs5LR8olIFXkn1fAtel4/+
uvBkVUWdJT3ozD+fzVCn+pkTr6qRADCqI95wYfdnp4P2TeCUSea+DxhQpxF3FbLB
xehVJfLSdpi5MjTZgy+q+jb7gHRPVS2yJauxuWsxZoSMUja8mZTr7KMu5RRZORGL
D19R3Rh+6G1o8y0E3dTkpqcpdXKYaDp9K+qKMFF650PeoINvwg0ks2NoEoa7TZYk
m3wmBdZey3XEqEsH2rJl4rHk8FW4xR+0Q9BjwUoYoVeXwBmdlBpCvrkjNhaxZVcr
6MkeHDsMqAyHdgicRDw1OLD1e2Mr7l/a1pVPVdlCtwmAUuiY/OUfCCoYzzI2s/Ok
xXw8uxWzGqKKYEIM+loSh9GZj29r0Q5auVxqgZfPlCgmeONsDu+MAi+59bP+hxvT
Q1Zbtuu+tEZVMiVr9GJgk8e6g6ftkpVXqB+Cy2hZZrPa7KPnS9wrRzSDYnR1EpAv
pHcqV3ipqPOsh0oXEm9BWgPYFO9muPJNE/BiOj/R3Ax4j/UOrEtzvgs0TbJz5hZC
S6sqluXBmkYqlH29B4K1jxfyS9Gve6xPSbID61ru8uSoJGc4FEdVOrhTRyaN2aEP
0/rqRkmFf93aKbhgY1UQkf1mvngQysIi1Q3uN6ndSZPUp0Ut86XsyInxoE0a8RjQ
xaQIRHg1axpDXl6BgqixjZQrL40plEUFBVuVBRy9jO7dTZb7ZeSEPMKtUg+4Uzl+
EqvnO2/Wc2zpCiZuATx4GqntQipDpJ6ivxDaF6TFEGXCL4jn9aaAFdT7KLI1WfrD
GQhGfrOp/iy0NGIAwWot1cPOVxfsv474dlEvLIGd+R6LIDzodMMdcO3sv6/+SL7J
C9C1a1ZhxR2uO+J57X1uGno2SoJMdxtvMO0tfIc7ScCIXjtV+Phvy0G9Xq1trJsO
PUqZP12/w31J+X7fTfXpd/MDsNVmE/0m74GClOJgnE04ooIwLQH0FS/9+fB/gpSS
5PHukWl+0QaqrZAlb0OWy1fHKzHxrlX7Nkd4J7Hr8xTbsMNF51bjxCtZIFXdDCtC
ZZa6Fk12V07HvAsV5lF7+aIGZvCMLt7xdtZneRP1nSLH3KfjY9Vf2hXV27faip5W
D9I/t6W7EZPHof5a45F6DEzaUKZYIK+i5htwO73q/heHyHRG4tTxozP49SLX3duP
TczSqu6NU89oBxUCUCvcSeoTs8eDlRt3kfUU0ql+J+SutKLRO4vpFIvzk5MApn0E
kDCcmnxJkrkncYS57C9a/0OxT0mXTYE5nqbsqBfXuyoyLwQBdu5wPBfKMinYJ1ur
1X3o6gjF2772j3uNIKy0bou0QxfzyXd3Wd9nZw3nAGAIZcRZ0a3ccsipKUcysGxc
Lgd8ru0NIdIRBzVMXRVuzy1lp/gKiHI+m54ieQjWEZqira+jSY/PUs5NuOWmgIaM
fVli2A3lKzf63fgbnRNRr4+kM3D0MVw301BlIx6f1tPP2EhuSSZGRUjnw+Cqh39R
LTZE2Qeye24yIX2D9waPtgrWSx+Fz4M1A2SXK1MvTgrG7ePrlVy2atbrQ25zISX0
R4OK7GrHFMrqXJDbtoErn/cX00iXEF3NNQMfReExRz4SKKaZ9Es/L/Qax++PnLG9
u4PUR8V5TZL9b+1rdsetmhs4ImxHswexTQAHmRlo+LeSi3OhPADUdN5XUXnG5pkI
oDNkxHbSBYcsQN5dyhJl06jPIgdCoXfNOPc6MYEUyVF70euui2clYuW+tDY1fdj3
J8q3UxNrRK0LDBgvzh4cpXJuyGsFMWO/vz2efqH3Nd4V7nmsKffAwc42QetFnzts
LY8EObzY+eCpvVeIKJTKcrUbCBENOVmw0tMaLUWN0b5zKLJLcRkFzYFg9pP0GIPO
7BlTqb9c/IgA2wx7rx1VUxI81NZQw+3Yt0nsr6FQ0tm+jlJWaP9kQ9txyOO8X4ak
i4YSG2yxoMUHnlr+9S9ZYBjZbkSdU4sC+5AsYKNugP0L8ve3USO11UGkeVD588M4
/tERhZ2vn+5p1NhHCx008DJ0kVmE2X69wE8+B2IN5gojgp8oL01a9rIvCtdcJEQh
hyZNqNS3szJRu6A9tlN4enGMjlpv3GCd/aNwgoRK5qou5fz5VrFMcwbDycGGN4S1
8kknbFarPOT/kHhL84YgBN9UOvM7+0/pqEZ7hcvZ4UOObMUbgLSbeJwF+DYp3dy0
9b2DXwcq+tQktbvMVdLZGRZm23VeYaLuXoKAGcL4Vo8JGcZJhlvb5BYUklaQEpwk
viSOnYmLKowXWtqqh1+k20rlRjAnbaXYXMLjz+oemV6Q3ur57pqfzhbWSq5zt5x8
U5+L/nUsW6oegaU0ZpdE3TiKHHC0lHasPjQYZpeHL4SaXGA76yxKBtnLD5mhoYXX
/0S1405ee7aYL1wPidA75hnyB15UdZi3u5hIPQ/Yr/iXeaCEEhokou3v5AsePjDx
t9bGTwF15rcwWFEEmGydDdEhV3+R6ZXlhQdw0NOyJjaabuu9Zh2F29F5NrLDq+yE
vcNUa1i5/HpxSpdtscXJ6E7vd3+KhuXyOKyGqS1KN0gPWqMgHIHJ340qCp8QiBGK
YTvhmmHe6NnG7tiPkVHRPQwzEUpPBRWCIkUaeIh6bwytSZIi5l61Zc6UBo0b9PqC
guFYspQwhoahikri/XLDjM9+sEC3Ayn2XatVd0XqU4PCXBur/jws78/Ndmvhh1Jb
SS6wQqOSO4Y606hpq3m0eRBx4TUIuGKRiGV33I0Qb8WTFA27NU10keozYrQlcEKr
ZFj+l1wM6rDjN0GxbwwvclZqx0f/aZoQrMs7KqaW6okAWPOwlpqXOJGQwk/UcnYU
AB7zFBdJD3Ehg1OO+tIcowje853Vp0shQTxFsVPZfVzkFOQopnqzg+jGtbI23hHj
yp1hG/nClyzlduWObp1iqe5bAi4oaFsco0iZG/R6Sm6IFMtIjDknHnGsTBmo2vdh
ahVn1VOwvQoEm2ns0mjtPGLhVN9rcD5h1Hkh3sCgIo2wEchoN/k2tSdJlth96ZAS
sz6DXFCp0aPoJo+gTJ5iF2jB/xYX//sCd5CjsgEEZJpH7uXqC4ixLB74XzhgNCNF
Ijdj3SA7ftRGtBw6Y/IqeDK3YTO4i+14On1O5/dbD1JHvNSg43LAMjK6nNsAaxFp
koZrmRzCKXtnOB1IAIXOPujqJ5L0yyqKRMMjyFIv5D7ndqHYFr0woyAndQ06J5f+
hU1AD6up/DP44d1jQ9ErLZcopTwLb/4jf3psQmHRzV6x7VGzc59iD31kDdF56aMK
MNkpw6iy2VD0Nunlot47JdtHgJKSQ/92pZ6IzSvYqj029mIkbXCJsiJjHDow2evd
QEE3nhOl2cLbgeQkjHHEs+lcf5PHZz2T0fwghSAr55acBlDIsSilIohU1X2i42Um
iKTIOZ67IvwZXJ/QqxNU6mUHZNEnAHRDa/bGYQw0lvLWkA/OvCdKlK9/xejF+BpG
NgIbrcSpFIrJ+BC0+hNLgcxe9WjyAQxBmAw/UxfUmH6QJ5orL5y6NTlGBRUqxcJA
Ifz0pES9P2zMHmXIBWKAKxZok27Cnki2U9uCBmqKX/qE9CGy7mRsfellyzbolDJG
nzRKwW7rY0sdI2GApcYUDL9YlqlVlLBvBV1Mv1wfdYQPQ5nLtpTMPxaui76VsrL4
0gZbyRYL60LS73SPbGLXgMHK19NwDTdACfS7KqH5UV9IcvqQxbVwBdq+Uvsm/Ilo
6aWbDZckMzuiZAWAPPIOKek5oi8hkNkIWCxHI7nCyljjr/Xl+cVJfc1YaE//rq1g
e4Izv+nw6no1ziIhtI7u6HVxrmV8q8fk7fdzcAU/2p8JkFt5321edecUmDyVG3u+
1xsBnSLK/+MTKUvxE9fthwHSH9KI2L4sAzEhwrXp7k0nqS78xxftQUbUyOTFLmXm
asqr9XSOZW99V4V8MuSb/Rvw11t/zlaya01ZPn3FbOCbF/SveyD1gvj84WsERlZ9
NYLmTTI4EpsZ71QTOEdjDa83IbANYL0Nsf16BcRhkRMiM2vPOwSCqijUFXe5pd/0
oJGCH6uNhYQMQeJ8WWJRPHqSVLo/zpj+UvbleJzWWxNufVon9aHnWDzf+MiQLijY
x/Wm1iJ1qTVvFOsflXqzgl04huQKbvCNjY9w3LV6PdKHx8eXSctrdYshsfUIutwy
6aH1m0k8HruXnNNuaUwsopwhLYX6UJpY0szLq7gpikq+HXF64/OPt8uwrDfST+zb
XjhUx8ufcJMAHSmEfUH6XLyaitegKu1QJ8vfiAP4OcxMKFuSaYFEZDqx010YcUm6
QMs+KrAFj9zl1cIMGW0mCc9o8cu/e4RltqHdt0RvJEERtMnGdQLma3PlbVE5tVw4
E/8h1SuwwzzRU3gQZ4qgHQHq+dEBiwLDqnkwcfXJkjatFCPn8KOMD5Uwg9hdVOGL
HRTQNyR/G2/VmL6L2pDwRnirphKjt6SVqbAvOdwmrEW1BYbRSYcXpBfmS4XqVocX
17DlTEokxuTbiqAE0jqRQvwKy9jTfZgwl4It5dV/7WMWGs3dBN2q0evUCdiASs01
xDDpYBzusZ0gR6gEAaDsdCNYxxGlvCJmHqj/t7JcP3PRuC/CD1jKFhxOh6B57AeU
cBMQXHpq/y2NdYzmF/JKznJOMsYfzEXwpFpKh3Mc4JfnSDFBwMIbvXlqCkA+JsR4
cQucMbTiO++pAtFvReyU0rZooBy4aTs5/P6yNk/lW/boKLBhnuba5vPic3ZHII5u
F3KszJZBsMk19QuAYQAp7IyLx++8h15h68lf0AmZMsuvpE/b0nXPlUDFD1Y65kc7
Jjq0gsfJMs/g+ELNtZDc0OD92YVyWSiUhAwbmf1lXy6oYmBCUzEcM+Bw0Im2OOqE
oAFkmPWp+AWGpYzoy+xY8E54K1jNMEWlIhVtMDWA2zkzxsoIv+nWh8ihHh/fX5bS
FHGNCs/9kDhVosVb75NWDdBl65eJP29824T9C/nUr8XA4rSnd5+/CBXuIQfdipKF
suUempFfksuG5kn85dbMrmQOPaPjVQKezzpTPskniQoyVumMQWvUlcjVs9YMqYw/
kWzdl+xKQahVUub2r3wjAcWpr1MSOBEOk6PdgR8CJZRgTWILM2OnA7EEL1WcbC7g
OJ1FGJrh5BU+HbpXwt1Hsc5O5yvsQPX74Ntxxp2nySA5s0NdiMpSCu10/GC2TwdO
8nILTEVTZlblyv/JVu796tNM6JvPbyR94N3HC81hg5I/aMz2K/x89oNKlcQAqdk4
iNAf4lSavNadcdJ8++KGYZ7nCkKl9ZzQLUcq1iNVakt8708yHDXOG+OdiwTFYc0e
TsX74aNaCqQAZ3yhBFnpJpFnDqSCKKOjv+PQD+WgxzR8cfSKCE0BrtjmruNH/K2A
E0lKMUFxbAJMTeeEpPywM9ERQmKK0073cmfIUoQa2ZJWVhNKOAPWCiUcbTlx6wIm
Ru0H/3zeIogyLGlsdDZ/gJiq5N99cKbLnYvOeOIMrdimd8l3W3l/8WuKqnyrMjOI
9c4wNJximWBwbR9mLBXgPddVzs5uEyqVco/7mGeyXK0zyjVfYMW5oR1hfTScvhjr
0684OsIl24RbNdtqzptqommukUPvS3/HmkWn4mpoMPk2OBMnP+0hQcNODIgxl+tR
CqCTcmUJbH9B92jqegVfQ+VDG/PKdFeHEI18VkvCVj2mt9ahz9osweo0c07aAF6L
SChNlzFJgaIbK+IO1b0A2TabUoGW3d6YibpqUNQ0qZe91mYVbIhp/JYCystTnt5z
OLfYf37N9WpyKY7ecn2DacKc9nqfP9Bk+sYl+lY6Uv6m6OzUcKFHT7uk45XdhBrv
DM7eGyXAq7Fj7SH235nNllxS3WPx6noiUFTZw5N9HHQi5auypjYbftJbvgLaYEaZ
sVYocDwhjqeZQEHTJhQdnKNhtZYKf0BwfxrIx+EL3Dv0hmkHyhX0immD7lReAja4
9FJxXKoyUfrbz2KlbmLiO9G9/5+y1XI7ul2NbLpvNN8vwT+GCcB1CN7t7hH+140F
7MUYD9X99567X6MbAChuCUfDJVXTm6/0Ry+DDsw/CgtpmR5LlqdFZC6uJxj3KOOa
+NjYXssQG+R3ogaUzKE6HSN7Tc1Mj6KyA2d6qLHarz4YYUTAcXNOq5tLK2hNqC8+
DcncNvkawUAhnKk05fcQRrwo8ZZCyo6nfdl+ajQ/BEpUhoyWMjeNtI2aPamOmw4z
3gdPZPMOc+PXmAjou6bJt053UP+S8U49oM4tNJ3AFEN9X2FPBgBupBkTy34udXzS
YqPZ15SZNGjw1qc9uqmz7SBWqUFaqU6NUEUpNIMhRuDdDkvGwu+a/jvSmr44WeIF
WXfVCKR5u1GoVVCoirT8SITk2h/REhWI3M+wVHa0JW+nEjblq7J/dS2N6JR/Qo+E
fKdSdsk4cJYBQ6nisP8YER5aaDyvDSaeRLwyT83xrzYKEnCY+QA/S0/ZxFXpWG4V
HCJspOVyMFigarJF1agUbWAZTrqY1j0Ujb0YzZAsVcAUxi1R9jw2kmdNwyV/GwT2
fpGU/2OgX++xmzcdeH1LgSNzfdJuvAuCXtHiUIpuL9fdjolm28xvI1+OtCCYQII/
qwiT3A2pNNaAOtyeSipJFjuHlvn+u8xACSX+OKy97qzNj1VS4LrACOl+XRGXOePB
aveGwZWS2D0M5AvimVlm1mMGyKoDOXLkP0Xhd3qFrf61vd1UbE4Z2YNHGSEkaLBa
2FQTJc8xlii/nw1Gwr9a1qqtZGHvJKffEJUTk3QMtEv3Bqcz04PF33joUh+o2lAm
qblf82M5AS7qYLs7uTGuqKtkWpVySAt5ahFXupVf5Vic6QK94CinkR2kG7MQJZ+4
2v4FV6SqBNxMCSxfvy1WbyXLDqo398zGoOOO1SHHJ9bwiSqAn/vtjcTZ5C6KIgfg
h0fqdu2oLoF1LtoUmXaE7Kba4zG29ApuCXX9Xtg8Q/I7IWjQBu3ewtqiRbcop10e
FuLYxBA7qQ1R8qgG2XysFVRXW33Om03nXOQmz3K4vOtdpgxDOR+4QDjH25IM6FRI
8ME9U1yjCEeaBdQrYoj5BWYI68Zgg5Gc8iYeA+cktlSPWfrUSD4dYEnEnY5JDyD1
m0eybn+32yltspjoeDlQ1WsKq8jUOZSdiUOQRqdOLDbpOcOgUZqxbXb0wqEzVPT7
de9LY+I30Q57Jroy+/ork9pAssuo17AbTaTXKB68qdavP02eQEM4UxQG3E2ofSWN
6FU4k8JfmFC+Sn+lUAuAIJIB1KNbONnP5nSCZ9Ok5dsYMCSkIuZekzPYgwNPcrXd
Q24snJWhGJQgPfQJHix91CVnLSmVZlHDcFqPHVJloDpfq2p0i/8VD4p09xMcePjB
FzHrb9feZh1S2UfelI6Za5r4uvswAu0vpC2vg2V1LmMbTEJT0sL+Obkj2+Iqo+Mk
O9Od+gDDbmSUrqnxpqMFMiguL1Eo2DeImqcv9dkLftjz/utGw2vT7doifkwYNPTD
9f1nhkgEUQKJUh7YmeAcxW7eW4cuUX+vvfCqk2m3c3bL+L5iLN0oubXzemqPrHyw
1+gPaScjbapoSTSHcemv8f2n0uJ48HkEAYUEFe+Xs0VcrIdIorMXJd7RFSamAxNU
7d24cmE52CkPvNsUh2E8JAFVTf2yHjvhBt9emw24MDRgerFtFmWPIPgWwt9XMZ1u
+6jd6Vms30wuftTYMH8kvmuSVGTpEEuaG9/PaX3+tet3iOuzCnsfsbOM2wKjCaAa
+1utlHJqYfTuIuACTSAHEYPmWNmENyEPN+dIHTLuRySbwryJ3Kxgcan9q39+cOi7
aX5Oi7LJ6E7Ph8fP2/NIAf5y8mPrRXOKGJmV+ngafySwH7j1DRHkE++PM9cPMjyb
jJnf8pC7sAEnBkHWrdA4/72mo8XSTU0rTscwCNZMprDsNImRY5oXQEoMkliBmxmK
GVBXZx9sTECD2Eh4Qxik3jnjO8ZSR56ZqxUhiM1UVqMlZ3cZM4rdU+6Qe5cHHxQ6
tTyuWHCuO6/X8QD1aRAB3o/BcB4TtBOH3O4wKnqCQEL0Xij6qakVsJQWY9D5Z9Om
QzzMiwhfIipK7pemvp7L5FLmIQ0ZzaWU4QKbeLsGqaQszvGEwd2NfG5sqdLE/czS
zJAeq3EnuVI/S3WXrP0tEgehox4UUpABaEkgqmkWW7nbPjnNxO1Rm4DTYmCv7xlv
CbTndrguNw90nrlhQR4agR6xkunjJa4m1OyaoFKWm9fcS4OKF2cscvGwvMhSiabF
3j6VBt1suw4cK2xEq8weUWECy+XlanaWCjS8JTYSJdqoz0S0VCcxVJb/m+hFZlBq
1RhC+kLfOCTlVWNCd4i7Zh7XaEz5wqmM5atRGJc40Oe6orp/sPVphaNDDsY9JC6R
Bl8LEIzi6+x6sYP0hRvp1FaGypV61zu5FDAuDcTWBuRI7WYdoHNCX9CwL96LlwTw
sn98D5SIU0+oejO0pkL7YGuhr7dAICXwuYUkuYrXRJgTvJTzvd1HpuJVo69EiyLw
rnAFwRPI4nbm4ZizrRx+JjuLN2buMBa+JM0HkE7RyqFjQzItvIqnV+lRmGr0MPPC
vbrSMaPyseXvNMO1bq9QQpqTkjA9lgMreSWrJhyk3Vee3RqnYBpy3L3hj27uxhx4
XXc/RidC9DzPxIUSPJFWFtEFicWAg8KR0mVoFF/I7661Heu1wDiS0QGTjZ3h8jVb
yfYkuk150BoxO1RR9/tm8ksBA+JTphyx9G8nqtx40fi40FRwq4/A6++X6h413Z/z
2tXIHkKqVcpdw6JNmd5U0lkuc/3u6kyA4EBPWqPe+fORaKVNqazb6N0ubPoEFOzk
eK2Qwuwe2HlWnqaEK3dq6O9WN0Afp3oR3l9uO7uBZcQ65R0IqinkX/jlNbOlPw+y
rCTWAEvXPcJicidwHPrwB+fLQP5T50Aj1P42i4U8Y34g/DV8C4YjNuQARFCN5r4f
vIfloaJnq8nKAzSTFNlKcbWZHDXy+Cu0m08ilGKQ+D+79PeEn4R6QAQJE5S86uwd
zwlbho7RS0G4ve9Uc8kP2GYJ5hPsQLSw5WLLCeLOjkhMAB7jZf84K68/L5iNRorT
1AK5pIS9quBKeYDDd4iiw8YsvDwTp6sDzGiqjLQ5kiVPFMjqvRxKHHpO/R3FbjCj
XXWpcsvUEJV7/YNmQ2kKTjvLpCeSCdYSROTjcOXt71JldymqwTiuibqxV4leAshm
glsUcKC2q8RbpZkK4rtB7F7jRETXa5pgJZXi0CXdo4css3C7Mxl//i0Dg0rqUWq1
U6PLlZo5/VToCRIBFV1ugBRcs/i+pZ9uPtGzYY1WqqRgNDwthdAylopyNfE0HHWa
PNFwQNYyWz3vOgelPfLPdWcwyFFkSenrpHWzkKPvb6Dzh834m1DF7LVD8yPpuQkF
+3QEgj0+hydh6Dm/yLMtLmHDLRbukifi4XPL5yVBsjo881ph5DM0hjeuzL1r2Sy1
QWp+FERRRIOrhQEeRPFwP5SmQXcaqwJqwgCXq3dDi2J4jT7kZYRsJuxv3OldWFLl
C1Pa8UJnjaTt8Nx2RPxmdY46Y7ul9sm7mXmGms7Pm+rXRFCfn6ePCQVnc1hCf6ey
xFv9YNS2SBEzyw2kg2AAMFcte+RHjRZlrLL5nc4AOA/AagLwPul2qs8CbTNPU+Gl
IDtyaOJYM01DBuohLqYDEei7rarIYpr51bt3scTGTlJZf9SD0FUt28hYTs29/Prt
y7gM0hYROUAlOfkuEnpOCV9nlHbdfbIxEY+WH+JuJBsy7QUPRiAYS2SdKJBVlDTC
faWbdaX0fY/Cy2J69DQ6mIK0qmYvgagLQRmNDT9CpYVCYCP8PyuI8gdBk5ThBx7B
pYYTGyrBQz82b3Z5wMv+0TPnzKolYSEvFlhGVfzeeEP1KNzjpvfYg65cxeIhQGCJ
ILmHfv04Ki9J3s5gmtL0cTO6Ou/oDMrFWe8CvDUFsww1NgZdbq84E7oLM561bzzB
ccv8pV7jD588D4iBnZUi3phRYz+5D0tguSayGXdkwnzC1+MIP9PC8C7TNcmQVvgc
gBIxmpW8zCOeMfiqFVYTAWGyoGa/NvcGXK4lx5YrHcIh/4B0FWRbF2w+gL6zUYw1
dk0uUeZWEL8hI8PmjNehucyDrIvW42WnszUVDU6khK63lTjGgi+8oA/Gy3e1ifIj
Rf1O/TSs3aFIGUzfvvuSzTi+at2BkQWJKgA+8RvKb8cCMLm4HiQA/f1GegekG7b+
Uqvc1dupBOCqAVAEr78MKUQMnoCAvHJ34SMaUrSBweO9Rn341NacD7KAvws0bfK4
WN5XxxzbzXRv3+1Hay38ogsKSQEstGPTVpWXW+RZFUf3tEAlUHR32lYAxHH1Yeuz
HrAU52IO5W9NDLErFmHtKxlW74vSL2Rwp74dYeHuBhDftGYH0rzsk48KHfWfmFGi
YvBZL8CsFZxPLe8rSOJrLu6TH5whhY8a0a5sE809Mn9jqHJ+cI1zeOgZ3JAXaLYX
9XYfwN8ufEOjaO8KntlGzBSuHkbWPzug9CcwmkuAkP0t+GfLOENU7wtnBZgsF9pN
8SjJivvg5TuX6+Zxn6mbDCOicdwpLS3QKwniBMF54BeV80rTjHFjz93M3zYYPqEH
YHt7rUWBMgrdxQQJs/T+B5gJ0C4Sf8bUXWZTdCICuUmgt7GVeIUBJPz7SvobkEZX
VYgJtNYVbs91gYJNZ4Rc1ksfD0+kcqWKeBmiLvhJoobeN/wt/KvRE6Y8e8XhoI6E
6eibdSFenEdJpG81a5wdwreRMwAoZA9XJ7g8+hsRijukWTXySWjUuld5Qg8eykEB
ly9pPP39MWTSuH1QbmBhnd1FXq06NXSCAJwYXGjxdOx/i/idUydhW7VI9DxTVESy
IIV3UICrm5WrNjUXt+IEYnw07xulKpRleQZnu2NyMd2xIOva+DZ28VqdTwq+r1ZO
q26TQknk+ixnol2x+zds0aFgMR2CF+6REFkRV4VKINNSbiXqHtMzwk7uhObCzxsA
VCAwvCLzBeIM+cjF+cUks64jBlNHHauQwIo2stMAdfRV8upCB7vG+CdoTg64/aYZ
o7G664rymVwjAN6EMIJcN5r83HYKNsiut01xc21VInBJt6tIyD93tkUdENZEtu8R
wXE9NqEo9c7ALmjXfxSj+UkQS2JZGsGfFfrW2x29Ju8lGZ22VuxCIR16vYKpoE8W
r4jwvm40YOnr6BK9N3BwHaw3VASAB9C1IoOruJ8uY9QyZkwFIQY35Vc1SzZShTAW
jtA99gPlb2YeRZh41F0zrkcp/gXTiWHzJERIZAzILmbD7m5qTBnoVobN0fOn0idQ
CFbPHaS3eIe7HSKVRMJMQsMkx7oRc84bQMAs2a3zy+I38LAPnMkcsSvTdmR3rUJO
ELWzAS/fDwySEtkZBQLr8LQeUnPXWtYj45d/ta4p29tcF1JMLw7fUdFYvW1W+k+7
k2BfL12GNw+AQRZnk9ge/wys5YCaIKUU0y1vAd9t/kJG6PFiRwYqHjZxtMUvSJEh
u2nmgMo2aEn3x63NUYRkoaSBDvxvWW1YEIY/QRjwUdDsXW1hXSBkkkV898wvTmQj
R1EvbfQ4kgtm9QDh8YeNktLyKDi94Vx/TQlRCC4BzZI3aM2o00/6ZVc8/w+urRQ+
Y3lr+hq7TKS6/KhbfaZsxvbe5gDNAZPAW6ofNguuhN+98Mr1678ySMizKm7R7dxG
kUcbA3EJ+AkRxACV+H3pB3owpZW4VWb6t4j2yJj8tBNzxL4glkNk7vbXBTjhJSnF
QOGlfylicApdFW2zM25brtBxNSKkcvjsJ3nylCFZIVYcoFgtU6Fe5HupB4DI4Kv+
m65FH5gxiwt+KflLxBGrl86uWR+5cuCANy1F6snfcJBwJjwPTZRYXJAagYjitpBb
s9IWaDM9kzeWb14qZhp+tUtXgNZRDXjWE+LdqscAhl68BpZdF/N4Ii/N5W4IyEo4
AmETamUc2ACGmu0sCQs8x4UenthBy9+8ARfRxAWuU7dzmLElRP1T32NrezsDIyFl
Lga6q0+IBcKWq3rq90bqbjRFdDJvq4RI/dseYLY1hkAmBcebLpen4Y/MfNM+W69s
RDH0rV8DIL8HKW/pwG31HvwWlfx45mUhn5ZO84lL85j5WerNyPpBEtNUw3qQpI0f
xcIdIfcxUQ6Kkdsq0n3R282CnzUWfWp/9CCPUl1FyGFUvlWuX6BRP7bfV7q+CEd4
e3NzmLb70/R1UTre3DtKbMG/ezYv4AMox0f0072YGtIehnwp3OQxs7blFeEGoyVy
TBw/jBVaTjX6YUEfbzElEv8hYtCFc3K2HWEhSKpohp3SskDalnmHim3XshKbcre7
m9JTM8F/prYRvbN/QiQyzpZuUCLcOs5dGc255KUa2p5zLVWNVAGpTqBYVUKK/nBe
CEgTbjYF2uLEUCeJiuLuJsE81ERnkzBMvrBHngK/waLcJi/8aXr5iIpCSHw3Z5Dq
mp9d5PafdpAY6sZTw4fIBET/UkM3OQZyK8NzSkcrCc2ufl1eYbcd0jImqVxLiuad
4x9BUzd9PKDWJ8XYwWiNjZ0mZExEf1wSDVO/A3c0MFltHjBC5x+nl1P+qjWFk0SV
9WVAtp8xMOTR6LkCd+/wAvjsH06iBRCaFNiaoCIJYVkNOlfSf9y934NTcu3uz5IF
9UVJE+ka0sN3cuwgfQmIVT9NMHuIeSHEqat0tu+xZfMe48xrMpTeTNQITR64rm8b
5+YQr+I1PBFfpq57SHYB13XyeTsuxUoCOYhzyRkXckcsgOVD9W7mSUSl6PU3g1oz
1nl92tCB/oRDJaBiNOrXJURQYYo65na18w6TRBJLkxuN3MY00uiPydBr/GgtYn7u
00Yy7VmJ1gOadazkrM73O+9nMjwmTdHS757LoPdHIUt6kO37Ug2l9WIjX507pSws
8Lh/GGAVubVYBSOXA7R4RBRlwsuV3AxbZeu011nu1SnPQSC6vhvM4t8CbNvt24wb
J2j7ynEtdE24bq6xXfqMVLiU3akv1sQhZlX6mekaqlcNI7kNbEs9Qw7FrvsEIvsi
jpDQV4EVLjxOSEmJhcnXBDe1EZxHncI0QQ+la5/0cK+YYKc+u9Fj1z9HRVjuhqNb
jFujpqLQPj+agZGLRscLZbebaMqUq2IT0T/h3XiIDf1Io485CzyMlUwq4gtEnwC9
US96XgOCo1OehXUa/22KkmQjr8quv0EICaKllLR8GwX8JXPTJjYcUWbFhJ47VZ62
RXOlL4aKU9TKfu11gV5UiRXqfbbyUcR2oKeiXaANKepptzE9RG+BJ1XnI1we5243
0XNz07AoZsTo8AKjBAOSZVdIXqHDnJrZlM0GNhOeElxW6WJ0DtaI9IgVLxaNZ7Zy
rfjDzrjZ9+T3U1r6vvDz6SP0Dsdi3C1e2tm4m1hgqu2yllfLSaVzHOF7zTeXK/as
lXEs7dmAVOZzDgwoS8TX5Od3BDlw298k4TQ4Y3efz0uYeDKpxxiQLJwyAL+QDz3w
h7zJYtzd9sKV+fdedwrVbHWPtUq52oczl5a8ZdtkoIqShpqhKA0HXEe5Sh4yiZbp
9CTvPc3YrNPLFejMQVjddBjfHi06QEVzWI7HRjdcrJ7YbgBVxndbvN6fFHIjfq3P
y95nWU1eKzvZSdrWMe/6SxeHida+/+A1Sc3QDgQN2leaqA+y3RMi0IlOs8/s+ji7
aTn8fHVHrOzs7/L6RYDX+fz1za3g80h6k1quMm/GZMaVJx3pUGUmeRQbYIi0oVeG
kpdIww9qIeIhlipHfl1bY+ccZeyq5OTUFIjjoivUD+f2Is57kkCfwpOW7TYqrvgH
VmWkvuklTxOw3dwtwg4FaipgPCuMugZQium8/xEa9sXFTHhdYjjRjWhPcW/64g0S
pg1Avo3fm4Wqn63Wf2r9RPZgpJxCbth1+qrjjtuFhdrArSaVCvXlWL3ahWY6EEDs
scomlfvAemnpMzCKsWX1jr5pui0/DGOiRE47SplyK/dUIHf68nmzgLGpiKDqZSl8
NOz4Xk+aq2UZlQx8P8I68LcuoWevueyHxQmfEuUBHkVHZ3qE5ZK+NBa1sZGS4AJe
Lqb6tdE/1TE3BfoM7ygm+cLuwf1u1XW2bC8ihu0IC0ZrIR3Cve8x3eRJP0sA4au2
XOV0rgimRRffKnmv3yNShmjPO4h6H6ijWar43NY+kwmm+B3GYTL81lkFlIE6FxMd
lOnlUh7UkzMTZF3wEnVeM1S7SqbMCdU3WBbw+3bBYoo1ih62FBjGNF0JUhp794yz
RnJw7e9yUSiFhtgF/2u5bc/agrVtwu77pyTOjPSJWLPUFFc0itIQShcwcXZ88rNc
LsrvOppLFLRaRfgNV1cmXkQ7RtsldtG7xcbQ6wZDAfpgnVZK9JFzvE1slbIw29Tf
zGkUrukNNJ9S6/mIeRZUjjTWR8uSScytpo51xLln9vad6Li+hDOHjvRWXbKdZauU
JahlHYYMLoVIL7b4Gbm3P/z77y0WSagfzdWUXXbT8Cs/NN8BOTpwo6YZkzCy62jG
oYXnInBW90nlpTKl4WXycJxEWJnSDhkY5teBCZUvjIkiPlN0dkdIlcKIz9yDMtUJ
LwPa/0hQYgL0C3aevawRuZ4GJXvOsH0pjsWyIVt2UgfJPJSoe5rxTb4FBihtJV3v
WXrREvJjmtREB9a2ZQkq4mAtyhATN31gzh50ghJtsMSV8LqX8/MH8Fv9GbEcq0QA
cWsyEohQycQQCktLzJlW+BNdfLUcT6PgkE+SiAb6fpe7443/wEAn28mqu7206rra
6Gp7xnF+3jxqWbc0N7oH52phep495haXlpo5f9mWWxIX7kCEcjZWNahsmiYDDHNd
8X0e2G/KXjpFVIuOHIEi74e3jsQaPpklpsVN42dk289d0zO+qzpLGxu+ffcX6xBS
XyG+2sdH3Zlldp7e3gNn3Jp0/yc6E/ga2HSU/+iMPOdJmR5RHkyylERPHZP/LHPf
pJ0YPa2yftRBeBEFkQ7ivsqmA2CejaofG3G3kudi7S0s1tX15GjpQXTMI9pnKmDU
3LdMt1dl1WtEm4k9hU0RXMas7v6HyjybkMMACOnyZ/ZOtBKe/IPyZ/189zSKfNqL
FmZ8pMM51Vg72YcjaszcaTQbDwzDzH2EvfKdOBOsjyMnqpdCxtfOVNZTu2FkfN8A
HBdsrmga8Msczqs276bXQqU9ggn83UEYqtC9xtxpP2LlE/hllIW5pc3jsApiOW0e
5lkfJaVpEBX0U26CyJxwLxvTOEwAJ0ncRNPK52sbNBJuVJPsZC/a8sQAOFNuHNpX
FP6qd5rIe2vdO4zPiyCSik74yySNQ9m9SbR9UU7rXN+jjcaxRk8B0JZE32Cmwnr5
NnVa9HYtfEy3gqdbrz328xwVfvdVCWy9GUn0rl+mIQ7bo5imReQ5JNqsGuQd+2yS
ZAVlpNWe62DTZkl/sdbilUGiQbZdt9JsaW8PmfLBff96z97Ga30fMySS8qFDgWVG
2RzQ5Q/AebUiF1Uv3c2/TUXaJFYoioAtvR+NUZ3O9jVIX7wfAFNf64vsCpd4dBHr
c+CZnW45hiQ/uo/UhcYFnuU2L0GFryjozDhTDFgN07X999l++5QKdDKmgs6Qv9ih
Bstpff1n/VSjP3ffYcsNEkwQkYzOrl69WNywFUm2eXt7P73jIZy9iHkaXFS2ls7Z
iguVxIP6tfCLTRCG+qgM8UpG2IdvUiyZwVOuPwPnSA35wZ0oEKAWYpmKtBIP9Xqp
EL7U/HKwmE+YvQt/gxSZZ+XH8l+249CtZp97MK2gHG1P2U8t24XgFo2dxInx78eX
vxdQNbpaI3MG5M9diD5U9GGn1coZhtCBYBREVLn9jot/BeBOVt2jCYeDmfRP8r9q
yJXc522DodoCcsYzZzrNfQvgf+29dZk6YBJJOmn1iiNVkKLU9rJUk+YO1GJBpH8J
xEdrOjgSEviI9VPUPsDAcm8jSLidakj+TVyX8qX4vdGAG9wBSLpHMdXYiO2JdID6
Oboh9xVBQFny/5bksBrLZfjfyKeTKseRMBM0kM9TgDK5XsiKmdZuyECGcV5ste0z
nedlsvgKCNb5LMFuAqjiXbmGj9j2EME3k6TNzq5VB+SnJI+4GY60vbCCkFGUOIBo
5DI909AMBHoNp6+bVgGgDtC/gJ8DjZcSxzSk6bg55UEP8VkBDI5aeGgP6Zokh5lQ
yA60lwTKecebN55Yk5apdkRMsx/rXh0liE2M+oBoGQ0DA7yteS1NW8Pb9deKNBKO
8UlY0K4a/f5Kq//TAiV7nZ57M9qUYk1eCOtbhzUxlXS2gwMr8u0lwcOs4sdyhUDZ
s7Kw+F3FtChAeq8dDE2MvREUjtUX62bY6uuGvgRTiGPj1MdS61tzqPrE+M3mSeUH
IOn1gd4Fzexly3/dRYfFvyWIoVmgSCptBW7H8Ec/KN/CuVGBFSuX1Jg2lBbbdfqR
LT/l8QARX2mAt3v0nzkAhRxC2UOSC6sguCsvMsO/ntXRyF1+E8m4l0WC39aQhIV1
3Mt0HLwcK8rj2UXzeoF0OooYfcFtceZJpMmerQfg1/JOGxScuy/rIytiLDoiO0Se
2Qn0KjBYWiPEH9Wnkphbpsif3G4+gKbqevgv5OrlSYsDX5Epw1VXPNBlNnb8MgjX
47f0q7hC9DO1UaJ8duMGj7jK5hF/ETEa0Pxl8vjjKdZGGZoV2+qlLt7hedrSUeOi
Wxeo/4UoedrdFbjxw71/CrTfk9WUhlpFl5YQjBNh9kAafb3CYWP5Vb0s2Bxia0nX
UVqnratGNZCGwle/0BJYPd/USLYq/yrOcCmcLtZdawOluiDIZyBF2jqYLchAphIf
U6EGVr99Jqo37rV037gmRyX192pcAjV/GMgssdTnFj6t6jO+Et4XDEc4xCntVbdA
a7rip72dCxlxwF8d3ch68lQbbnoljJoPr4v5w5WjG64GEAnoI5PdeWeyhNZzAPXk
2bJLmg3fNGfveYZ0EVBKRJeAazXwpwavoc78zCFWvcZnl/fl8BH+BtsirniLJhkG
4dDYy4ffPWyNw5G6N8jg1Ic/0Ia9K7MYu6IWlo91xaCrX+RNP0QDi4jCsicbwbBX
5bz2L1aUxihF+CEKSwNyxclDHM1Qbg/xSzc/MjKNopwsyYwq+kPfF7VkOKbwuOpK
9j1Xj/p8VsqVJhdoXK/1AHDKjVMJzPdKJHOybmL78eBuTppa2kEQP1ZVZb92AVOG
RgaQkaXRAGwHLazeYFTpeEYCANBNBkUrbiNVr1v57mgGGDtkpcNfyFZ9DLRojJiV
ruiH6NTcDiLjfO6APtfCWQlv1WjNL/FyFQmrmrcTAqkXeMVRZNwU9UPcD2vtf/Yg
l9ztZuS737S8Uo4qJ8fJ52h4TWNCQ0P8A7aFGuI72pTsEN/VBZUCvuLtF1BihMT+
csmPFuABTLyEtiI4Zp+ziL7sIo+/zjrQZ1RZOlwWhRKE7DyQy1hFEbWqYbJOmMvY
8t9eeDC4O4wztnV+rgH+IgfZvQ9JYMWQEe1vnytN/PGSu3TWaCmlWCZzbp8POwK1
6M91Cudg9g78XJZ1PLOI6kqsOKGBfE0WljD11mdfTpkKm2DxAclMj6gAUD27sH9M
E6UlsO0CHelpuheJjcsxuMvNTuToS/i8nYy3S192yKZIXykuXNBzadvQvXlAwpgr
yz//IKSEYG2o5PZrWhIusHCwgcGbPJBRMJU93ROkR5WFQ6shBj3hLIwfbKB3fkmi
QefEC6LcMY8HhnNwFRHNJU4cXCS3gQeAYv7wsP0wWE6tbwUHHXL8Z1FstVKdJ5tj
uWcp2Uz3cRjBEg30EjJh7CHuLYV50m447nYkLy/J0YxV6Q4E98O3IP9e5qJ/1bsx
Yev2i1EQ6JT6adzpMp3/N9KyUH2VkeBfw6LwrO7aV8Sc0nLFZ/gdXUoEKX8LW+nq
dRVSzeot9c8mjLf50oQpawY/ZMa+1l5mpYexr5B+ZzbW3h6s2DcXcqd5/I4jmudZ
I6UZwuvub/oETrtwzzMpbLib07zB+NZVIfLZgH+8hDHo1fgk8UJGhFPe2b4jGK1C
SMx8NcCsMG+v55Ac5xljxFsCQsBC/NBrhmIVzDfihzTjDFBvLBOgfXN3wNh/fUiT
5ncIjcBOqnH5TJudhLIvHNYbC5frHYvdFDHTqBDIvDhhVWybFmuo11KciSDw8EfR
gQWcLB71K328badrVPhkYxpFeyglB8803JnNh34F5fGQeNN5U9mMIuBlwmemgGbE
YmlmbPz5L8CFmu1Aij+TDMYyrt+8DiEXxP8htYz7KZdtGf19Cdzf9MPET49zoypG
n8zrzffaCc9zkFJl5s2HTbvgWmJxMi06FrQwpaAtJuBqR7g8aus/py4GWOqP7873
rMHTzGK9JSkMms8jZiobrem/S0C2hicln2K1cZpLUQvnQFE01psLOA+jst/8kA+8
5MwCCkq94JO5FuNPY3sw2eYki4YWLF/zlKQhL3J1uUKJowY4IFQI2wTxUBPdiaVJ
J9qq6g4RvvI5yuzGj1hpESYD7VTKastIVrwb65LEse8IUR8alQaXyKno0nE96vpB
Sv1B6BvXEkLj6mmII4WVriQjkB6AIdO1zwjZe/+AZT+cZLsK0J5BClq897nX3295
dA8PajAYcvTI4QRN2nIo3+ZEC+Yep/z3vZTQmuIjsTTUiQ92K8vVVRI54RXu2E8y
656eG2EnLqNvRCiCrQw9e3v4ZLvAvurH4z+AHDZh/qY9g/cawFnnArBOXhrSKDMj
jgMg8K1lYm7c/OIGWXhG7W8JcPWAWW/8kWbp2NKsPko7X/6qS+/dcSSadOeg8G3O
p0cfpBTL+oKMxYLWKH2CJAmQd4Z3Rm5n8h9X/0TOyOEUXMQ+ETt3TCYsu9l5izmk
fXvIGNOxCO8TswpaKtIycqOnq9AB+xNk0O7STXo+V7NEsXOxrN1wKzVr6FV+TwiI
YHA98yuycVankFx7FeHVIXga7AwcSNVHcfOaJr4WdjwVAyt0yoGHEZpeRsQpnsgB
7jsqdXUB7pVU2AVcpYHKuYKsH9LWFSo+4cdARaDKmeGrTD7wJqSLX4F77+hYmBAx
Eb28dF3koVrSLM4GL/7i8CLvrs+BRM6bsgOP28f01/5yFVVH2e2Xgdd/+1X0dPER
E/CR3a6UY/24IV4WCdgsqHEbKAGUMQ5Dkw9VrgM9L9ChSLffeH8VjQxiTU9MKTml
37NOONQtof2bFHJdEkTnpNp5WjjHcxk+MoiZ4phrlExD9PzTItWOold8ON1I8dnT
EAQfktAlmSTL5lmgxUI0FJCgX5x+HEaZ5dR+uwy//1u5mi19r7Le8v7Y7e+VyVOn
Dq9+2zdkJJRNr0yxjb5zHXmlIpe5IG/OpwajJfeA1CjuDJNiTuJqYsSoNdwZ2eE9
ECymwfqf9BpG04HnnUoak3a+tLn6PCnPRz2pk/rCUmn2hM3pyzplRvomVZUypdaA
bKvpV2CRWqUk70FCAzon6jfm2KVQu34VuxQ46Y5KlIhgkhUprIWk78biFAY6hO5z
nCTDbjg5wvAgBBVidU9d3GcXJRvHIyU9j5pFwIu3Zb+gBR5ZT6atuJuIeQIpbOY3
7dHunis3YMtgtmFdd8YN6fRZPxW4tuBZu1uH57D0p/RavIqZTCkeNg1K6ZHpYBxC
cJMjTAx7KPWk7VS4df1fF0CVOyohFVn+z91LUeo4v8UYc/etaKd/BeYPpTwwMdnA
v3Z0ycla31lypLNpVsoZotwEqm5VmHY/4NpjlI3J0VP0mLd4LoeTWMvY4HWK4Gr7
ClP0qipv5HoYCWeyqevXK6rUMFI7WwIX9Vh6geOokhvYuugn2Iupre9Vq//p2R3A
TvDOpTN8BUTdFR+WcAkxAgkBCyyxp4KaoPjuU0UQnmUDPBvdAtdzzjXHkASC44Fh
YW6F/UkxMkALoESmmjg+HAqL7ygnmz9V4hUZC7E9CnLhDHlWWTmS5I/b/mrXo5QN
FdKVNPvk6JvCSHTD+xvlJbY2E3uAOy5fCWJqD6NODWHPNGIczSaof5yOjvdvBptf
9o750viF3un6G0JNmNlIzSCbj5AzLnbL8kjP6htmFqFEF+x0dzPYSWhrFEeX0oTK
sXQA/4wahbi3u3FDvIRKvMGCTZFr/JWbtQAZMbv53ImTpH3g1+5WR6LxhZUkWwue
ZS7ov1d1Zt6PkoEOsoSt234Ml1i9IdOl9X4NRjRAfkILII5PSTNHjo9yngWsb9Xx
WU0CdMwdW3ItPm7G9IIwNcZDiNeNR/L0tiXgblZMKZMspgKzQ7iI3+ZQXOrcbNr6
m5AfD8eXwpIO2UczUju6hD5vubF5AoHMZon9TGvvQhENEQICr6wyfyJete4/H7Ga
u0i0s3+9mog2gU7aoaNm7JURA1fHIbY3Pam6W6Iz2ugJeAFS2NPNJEzZsGMg6++T
ZBkPpBYu73sAI18Iu2MT3HlMJoyfim1SUplRGh/NBxQhc47Nfkudq3Un8KV1K/Ae
EwxolqLZy/CYTzevTjwWOkwu34OJn3zCllGhaYh+5ZiJ5pfjw/6SzwdKiJ+GZeSX
WqPWlcHPLMpOoEz3P6+ZO0QongaU1TKBfT/6UG2L/DanG1BL5EfOyHt616y9nsNY
nHNYHXkoiZGVrhnSlnVx5d9uVemOfWHlznp+bmZ68RsrQqZ7b1vyuOA9lXGLL+3s
RtXGo/XaUsGMRy6QPWwLm5/Lu5rfI4XWWJt5SuSxc8ZLBmEQ+sa3qR/vUI+D1Zm0
qYg1diHmVHt5ifjABgkstx4h7aiHlrQEqgSEHzhmJHysZhHG5dsIBG3j1ZkZTlP4
ePexW/vlwsvz5xSN/giJLKrbpRVcFKQP5ww/XGiV9WAfK9GmzSBq9OrDMOZ4CENB
McEKp5hvTivxxhLLq6LM+dLNF/0QNbF73M2z5lUzKUDZUSZLHjd/7/hg4nzEyR+e
mieSidOdBinEXpUFmPJBbmwrB+isjRba2ZMD1HG9yG4JMc44vJ6FsuUZUWqvkuB4
/i8XYABbJTR1GwFnpaYzHBmIEWxi1G4R9MQwLuGu68DxRf4SFNubTNUUSn18c81O
XWf0H/ZYRQFHkKRwcifAk+397PBBQheX9kuU+U3tBGyjfy2xgveFGLV1msVFYWvE
yFj+ewM2/9e4NBVYCg1BInGWyjUKVECa2KDzAO6Qolph3TPjl5fH+rq1qo7owtul
0yJm8qPpbKiZmB1i9c7oYYRe0KcNVAF4q/wOaWP50yQaxxjP+M3yd6n88uuKPXSO
ooo9AuD4yT40Gx9CV8NVHhNK0z4ZsTD6/5pKdsurXnZhA7MqYgaY4zpJhYVIbWMn
4KNTjeQal50s6Cda4CURoYJfHhTUfDqwTFfWc85bdgv5ATB6LRe+ZYiXNzgpZ2vh
9MWZimJEsLTsIGjHjKnUJfW8CcWPZpk49Z+ES5QDeyCOVOZ3RQKkLkpBVFtzrucc
yMG40qcKtZxQqcot7KgmK4j4IFHXkiMv5M+XPkEC9W/q/k1kvrWABwET/+PnX1fM
EkR4ha1ncnMiJGtiK7JFSO34skQ2gHzVP7ZV4nOkscVyeK7kiPia92+gg/Ffb0ob
LX66OHdTfRkM2TtajdGFfG/VA0WfB+2Ja9Rkkd1yRgbt1Us7fofVVp0SHvKaWjzg
f7kzJxJ+2DigL0XZx81XQydabdtxcIOG9oW0fO+DlHXFvzdJBIpnubWk1gIjyopx
xYS4xWfMonkw35iRhH9P/vMf7NA/pKopYPBbgp9KWtypUduLMs0E7tNdUgW0qVvQ
m20ecI3cfkY1qYsjsrywmDnYt3vS3WTxQQa32X1WBaKPQqcLDt8a7KHdAKMAOdbm
GlNcAaSiCCh+Xx+r3xWJJ6Pd5FssozC06CV1plhrtFTKEWUbfxQ3PziAAo6H9UvK
8kPsolej63cbbdK+i/ntmqXpXZEK5X3nQTumMBGzdY/zoT5SXTetxkVUqgcj+I6r
ow3+O2v+zWdoeZLlUGNUNlIdFi3inhFwOGMkE/0fZXt/GHShOQCPj8/idcAKgi5p
5MEMxSSd7IL2uUCANfDmwT+eC7yAAzR1t+4Ol1IJIibZzke/EhAM1HdxCQV0NgmH
U+6t5khiFBrMXHu4i9fpwZel8ZRMdKsA9yhpYCLSqCS3d0ar59XSvkUmZenx7I5z
vrSHjz90JjIyLhMr1odTfKHFpj66SU+qdwdbgWT3rRhe8UMbPYfDVHjmjIiti8iZ
rDv5KCT1/qTBn6O9IgoOR7gwn6Budqs8mvtXGx+enKUm3y3wiMl7c1uPLQHdF1Ii
CMDKX37YS2wMRRy+g/kpyiR6SsP6AlSBZkETc81pbjcE0a0PnqL6ZgluZjnPt4vu
nChdLy47vo4LQZcWeoQZqfvLu1Ypp5i8E+OqsAMY3OUrH2p6x8kilnaPIia6Qk74
HEh4cPJPhUEy5wv8X/OdUnraRo4bxoCAJuTYjYJiPHvBTTiJwdLmpwFPs8UNQvTI
Jbkb/nIvij82nI2h+P+M7FwoA7sVRJDk0d9yzPTpd3wRqNsws7bhCZig0EeKZ8IG
rjTgCOZ/rBCRJY2AeJ6aIRobpHFw8GgaTQ6d4zlKIO6XovYwUNrjKh4SyaU46WXt
f1EFpH8lw+N7wb3EMcwrIQttbDuoeoPatiOmfzRadkoJuGArWy8F7FGDarAVnRmi
Ridh+o1cPddfggSB8yQjVHXSVc4c91hnhLo/RLlf+fQH+2CsNN4F+Y9IxewtXEb6
D1eQ3XVqVDjolc0iCCm5VvK9uJhpG7NtNbdgG6DAyXtryJdeF8J41HebO8j7nIap
1mm+KLO0j6XhDeuB1ZNeyqFnEBqcKPaJvNSaXWbcydMWGfStrIKEhiAqG5X9wJ9d
Nwh5r7a3a+0jMVy+VwsGC0O5RifHo03seJbxUnbmoulTGlCVJ3mzoUJC92OA7y3G
jYvaI4Osxvmygs1hIqyku7AmXvleLn6ulK4qyTdEChf+o7UXB/9evdIT5HuGVVdA
2zK+WA1FSOgED0SBGVgVEmwsgyUAO8246hXsaZ3SgsYT7iuwuA/sk4y08oCqOW1l
UG99s0IUmrktx6NVPh4RvbJzKimPZi/8z1RjS7nqJ1ZaOP6WofQS13/Mskj/BrFW
NDr22jyxAYAElSWnl9/slUqxbG8UArz87fGQv7kul/hoXnFBGWUDlTXg6ksoyIWS
v0qzpR9iuNBdw+PXKq3DE4hG/cmjIygLZzmbt8s12jGqWIz09WyX06uIv1/jq3Bm
3VE/CBdOPN9EGlVTXwsqL7gc2H4aHz7PqFWVpbo/35MgZ3m+g2/N3QzVbkSjCSLh
`pragma protect end_protected
