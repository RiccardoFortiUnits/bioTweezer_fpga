`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jfHUIQcnwLqWyuY5QKw3V8T+e2OnMawr3BuoXbvPMh+LkU5g/6OWUBBXy8FAbmRO
xxCwrOgrAvJGy2kO/ak7DeK6DrfgxuYFgh2j1I3hmEXpHg+U4zL6tQSZyLEsfTAI
Uqc/U87Ll3RWPKYIEnO4b3e9Yp0GwNArqZYt1LkklBI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
xgHdj8YTDzcra0ql8nVuiUH/w+pJhMJFSAxBHKL2o3u1068Y3eLeSqPTn6NN23Cz
2IDs0DzAyDtWLNmjQCmv+3B5JAeENWtZs+s7HM305CPZiLg+jNdRtycx+IS+AQTH
3a1tfntUsuyY6C2CVcJjMVXUvQzekMwUAAph5ygdaeyi1D1mD2md1e9oD/X/Kbob
AMf347CQ7gY94Lg3RnzyBeqSQBJwWzT6ZTdNi0DIhl6q4dRqLWdqEWLzPoQf/UGV
3TxM96As0ZX8D1EB1lCaFFwzJX0P0m+D+QFMqwU7cPo73pUHG1OZpbV5oWNIdrFC
VJcbkD4D6TVnLDnXXqCqi80MQEzvNEHrMAQJ70BHpZtJOphxEBAOTB8zvZ4b+HG2
U/vfN1uytofdpRWKZwMNsoNBQuHoaCeNTvCxAS6kddQgLHMWNZ6IG6URt9rbgo0Z
3OVmB7dK0kBXx2LIcOwMqayb7057LxU7FxyLhYhDMRCPoVSjmTuNqtu8yUsHGEb8
ykEP/JTWmKTVsxr3XS8IL9jiiw3X54JKeFi7ThpkiaNNuJ1Dd3FP4GTWmZexoCjr
v6JZZxLNPpoYm2Vpu8PxIshs0kcV1306niozLbJKjrA1Xh65rZcgx0QGVLKN0W7x
ReZmHLk0smMX8c8bCwSX8XBBTUPQSO0YrTlwtxV7pzN9Zh8geO/Llw4CbYgLWI1p
8LX2IPCCd/6dxQEFz8aYGdJGy0jm8rcEvMg8YDYEBeTFNXniWNas2ASHBIMcc7gt
2vgsDzP4KclrXddeSRAFBka14OoXG+AgAIT+inDbW9vwiije03OIAWOXFU5WCUdv
r+i6jI23R99sgx22npwzY3b3cpb0QlA/ypIcXRUGaT5LEo9jOcjT28LKquiEXu8I
qWHeacKw9yTHP4NxuFvYaqAZRnnXd4aY5mLpeGVg4wT+FXv/PfeKYe7CCIHH+Q92
SrN+l1OuhELHciaX1eei6Yn8z3jOoCCa+tTgCTqhKel6OBHyXF7idvlBPXYYS/Hj
DpUgMgkq2FJCI96ca1kwlGmT5QOepdZ2uCkccIyUHhiDNCDJgg1FSomoQslwXo6u
ZfhtQCcLRJmXHw/7GA9zrw10ZsTBNH05qOAkYgNDT6kZWg/aze7QQM+0jzMKyi4n
0ZLDT/bjFkWOqQ8WNlzCSP+VQ+UNZfMkxL/RhHEQuRKf8VyBpaxuq5ZQTYDiCJbW
7JZkgzzp8PGgnXftfUVgoF1U37PRo2EPHwI6nAW7zI4gQzpqaHWQv3MteVP6gkM1
PHydKGP7rA6vI0vANOKlarHo1l8nRyWiPYiCtcYjkwEovkOmTyR2A9oFDMpmwOnu
xd0sbpmIL80shl3gHM8US+ftxM2xrgsI1b/hg1ckz7NZCfISgvmGcwDiwhDE+4X8
ySIf4Z7vqhVV1p8knsP3LE5AV9Lzkp00WsZn+2ZCr+MkZj6MBceJ0GOfNDLUfnIM
PMJQvEjFZlPzXiErp6xVwBa/Lyc4BqFG3YCOqRsElBkBKKPWgijx11jcplXnfDGX
o+mqx9UPsYWOg6jk62fgOkoqt2tjNFE2L0kPAzPSDdT8eMBLTQjPHuZf4krepu7Y
NiwrRckZhMSn3ZNFHDBQ7DCE8DmKZfxmMS+it0wfx0VuMsiGpRwVQVzo2ewUOjPM
/KIZd3DCPsW6BMyI0raAKHh58OE7Zo46vHqYEvMTwJguhI1aCLhUhg57Fi2XQXgC
OE7M1AwciMYwa1Umk3VAfwHk7EV5JYi2XnIA0lr7tTtl2Cyx7aAqcJN01W3d0hYS
AGOVS6T+eve27ERQQbd15ykjfI/WDg57aitOeAv85UWpqbPu1MiP+/j6amQbZr2b
KKTkqfZmuO8KqS0+7qPdAshZO6sVSvqX3yhXjrPhDnDcjZDjZhrSthof8T3R/pce
2LA0QBBdPmSA1ingjYWXJcOE52Ee6ywP+CvwlsJjD39ky5qTxIuFoDuVtl0ThwYM
WAlLAoR/0Zwm8sjec00wvtoeO+xyU8V9SfioOiWQuxHEH4qH1VqLo9gjityoeGGK
twzr+ixt9akw2v7TysdG4j2oXmhAADXyETiiCWZKAPyuaFmAH8wEo5GnaOlS7PKE
M/SbKIVRfaL1HQdk8udQLvYgWQ+YBg0e0OYciGNOWg/Pp1UJkDKkMj8jNCco7uOy
9FMPdfDfrCrRYLe2ymwPTtdl4JK+Pfh6LcP6jvnPxXaNUPJlJZEV8jEQ0+XCT0MP
MhjjqBPB2zF34Ve47DWivqv2ZxOW9lyTkbv7beDDut9LEkjbb2dJl/J6lrFGgk0p
pdXWO+NPZvFDzFWqBfdeUKtnJTd07q4JCzgb4OPyMnckpsuO7mfOy0862t7YjM0+
ShMCCMNV9MI1IlqrU3jFqxU1uUpvnqCdz4aHyVVk3HJn+yy6S5+aM30mMbiZQw9T
xpjEMTDqEs77BS8uwlKmcQ5PoxMaGjVYMmX/2DA8xnmdAGe6kwfN1dOTWwaoxN41
8w/uX8XKs4fY3/sc41kj3LjlxerSVss0OE/6HRRuxpQahSHjO66LIVbkJVndOB4n
wunHDKW+vVm/zOiqd32S5RdxMzNyuRbXgJJ1gJRSM1wt5gXF9z0bEdWTD8S0syG9
lBowTz8NYWH6VuLErNOxHFZxawM8/eduTrORAH2n6gtGNkQHsu2KDo9irZPq6Ge0
Wq8VMdzUoUSWxdblNSl3FJUOzACfTSD47KxZeZ4TUrgqwejkPReJqJk3hPqzFVXq
bbJd1BNW0Z9tescMjAqZYb2nHUk2CFSg6wp02ZhUYYkPW81ayOKLm6RjTPJQSH0/
Dg8z/pcXxBigIFwv+pJAh7c8upf6C80N/spQnJeCZb5/pZUYGDIlJHbY0ER8J2JH
svNIDiV4d0cYOVdPfmTB4WU3JQ2Yn83KOxK/xy4dsaYTz8KzQfvWoKZol+XBCMYu
BYvRt5Ff0Bl/T2RHtSWJ2Uprrijb+B72aNWrfzhy6t6dJRNixEdPyH6+gthxh9AH
5ePyzD6e+cZ0uWwbLNvURC/+CUS8Wc3/iirESkan1llTF1amVWyfMccyVMBLWKn2
vDf4AR94DshnHq4ZslrNrMKHBaWGsuYqplfwtiKpVqx6td/4j58wjEjNgVkhQZLs
lLGkHYKGA35ngW6GBZf85JfezbYN1cmQyVKEaJrWdyOON1hTPD10H9jJuWtbGFXr
oZWZj4Em2BeuTmEZzCZPt8wmdtNdM5dDmq1QakfLkGs3kRuzWCngXmzgFuYzDo1n
sgol+y+HRDjw5PWd/8SL/2pgrP+sTgDYZ7WA5gfDc/t3goB4BojOQDY+xLl5pEgX
YDTMiL61+UWGb1VoRGde7l9pzIR/rCpKO9iJ2d7qyqqz3hpJqptOu1Y8WpJA8Dcz
uvpMIsxtXeAkEfojGM7YPMjWWVTK3ZBVV6IIANrhmrpEbCALYhfpO5lxwS0n/Fkp
FyVsZwnU2RHpWehBBC86N8J94RBRfIulNb4iIA69leGvVoGvkVpyE3SiNfgtoqY3
rXMRuOH9VZoumOSDO13KoRgywFYb+jk/rNcfL0kCzZvnSwJp4QGBVKoSY2eKSgzB
n1YUbzMm44DvqNWPZH0xrFQM//qomFmKZPMUiSIa8JXfSXA2fKTaZPSUuhAj9qdh
mY4dC1MniYelwN2bwzksKpBD1LHcLU5aIrn+qImEC9a1gx6gpLAJstRel05XmIYD
vxy1gH54IXwe8QC183QzdF0DafbBWXqZ2YY8iu+DXO1Kq3kvj/jDIzCut4AmODtA
hiASVt0QiGY8ilVQnInaAnL1g3KF3od0qwdpJ1b+jd538hIUGZxUgVe71TJV+9bm
KFhZ+shuTgShGU7PAESRSAF7x21dy0BFhTaaHskG6kVUZzhAFLm5cF/rAan89+HP
CyGnyZc1XGlVY8KmmicMyeUchuLL4JTyYn8Tb6GcA2/xR0RRafcRcTGE/mLkdYiI
r9kqTadW/tacDlgPQzwE59E0l4ksY9aAJ/ojMtelCVmxfHRUcpUQqZVzaHl0zkQb
PtgHpPnDvNVB2WwnZTJaVS+wo4sQPGJ6WIMe9qF5dbeFVmo/OT67LHGDc/hy6SLH
/hHQTKJuTKpHx3gifipjaSazgMbR0kTwQ+Pdnvcq6a3Lj8LRwhabKjRXGfNgAUnq
EHZr1mUAnfOEBYfWMKbw/n/as7ZsUF2DuMpfA2++tqa8HqnO5ECjDlVEhVcpWoUV
pGilJB/D3DE3r84ty54HBHuCBCgxOO9joWurDLjrZGOl9vUaYHC+G66YW0dsR72p
MTJL2/P5y4ntcZp50NnYcspLU+adIjA0RalrEEP4Z5yYODvcA2dz0XiWlyIKHiY1
AU3aZkkMFp43N+SNQ5iZGMKywXABudIirj0SaDdD1lT1D4Fl13UEdm0s93m+j7ND
oGLyWKNpRNXAZz7wluGRPF53Q80qCMVb8H0iQKpn8E2n48vOjufvKIy4+l5CBNzF
tSZsRLDaOOH+4lGeTG+rnQybFHawnIrdPvKPHOshUOtGekiAHraLn5TnUZ4OjF8Q
61CGr+QB9GXhiPeO5DwDseFPQpQGpCo6iQpE3q0OO8rOTT8e1LlNwOocjgFQ0yFt
7jGZVdmFGibMErE65g8sc/qvinWQy2hufj7Zrf4TmpbD7TPJgq2yynFLKq6ffU8K
AsdYkukfMNpvIn93PjP1mZ8DIuJv5B9QBo9uht3pLLxB/duxKTMyErDDZkawkhyt
aZ6D07VyHU8xPCFHHYm8dRsdv0NlUZhGpxMRCf9d8G+0T0Gt7G5ZQS9qQQvEe+NL
a+WlT9D3Hp27nBC/rU3C+Q7iYvSze9i1Tiy1AKQxovTj3ST1nRQ1N/UgD/wOO+DT
O9pMkQCF75vr2wR9BWUGpCzpnFS39qksSiF+BShw6bX8ZosZhKikOhnYRf0k1H4r
z6FxNaZ5I2LjJ8WOkBT8iDau1AcFqk1TM9w9zkB46WtoWQ8qkcZ1keSGRgL9M/vG
nw4YKk4BUZ2G2Sp71M4aRmC7kxl6UYN/b/ZNKt8900Pr1RbxYOA6b+itA9BUu9H+
0xmLT4OSXIyhvfLo3x6DnWWM4bKPApXNQICaSWUgf9DDMI5P8/SynthmauXgmNnT
vxA3fWXmSLTPm8/RYrK56x9mIW9r0NWuxrMojAaQiuSeIz7VnQo0SQjtEePwQYfl
9AhSUnSIwzjmDFFuTGkF68ZiHOIzBMPp/Ig103o3EK1HkZundnn+mxEVa+FBCsAW
ppAoXNauYUzpny+BQzzSSq6X4VMwvU3+d0lZW4goEH7ugvgb0A8NUboWsBPaoMT4
JhKqBgMJkfnRNDe8SAh1pHc5TUAK42v6kHwPToZOmgFzX4yMNUmBH/ZKxji28fmB
UxqVFOSWxTnlp4pjnU/oYdMi5+mhCmqF/rItAlp7bkEMWKKNZmgw3/AOV+0rWY0b
23UniRTQR0CVZWTLixXZzauoMsieEtEMomSZEq1SlrRPiV78a6tLlVKdf/YMCjct
9dVpY4EzBEY7OFArzhr0A6N9wq70Gpxt/7UuQXfbddhpKUv2TLUONqyWd9B7RJQj
q+fpbEQtpUJbBp9/C9+uvJhG2Vquavogyk7ktuEAx7QjfMEBOyE8Ogf5mSiLECHq
EghG2OHQIP54f9ITa2L7GoiAF1y/GTyEJQhKNxAW6tCtf7dSichCkwxdq+LE5rKA
v6LSz9avJ+rmIZG3ObOlFx1Ia3qj6OLfuNtvgsl4T95CjKD15Wd08H//9GG2QSg9
csdQh6P8NBTPaqbZU42qbqa9oGionCIdGRgn5/6uIsjZlpH7gJQdYuhWXigDuoMR
KI4APDpuFWzdMyqPJ8mfmcmVmemzJNdszIXxOO8gn2Sb8xho5h9jcrBE4gTAwA9U
CUsJzLKRj13izHPnMzZCXPMwwV3nucK7FfnjBVCSV+JmyC6SoeYPwVkKlMvaAcpI
4Q8/uzKdfQf1XT7i/59Ns2q8dHn+KSl24b5VlWN0DmujdGWL1dnQzAQ0YBhMbkx+
nkeWJKsM29Lb/1NYcgsbFsBZmdO2KCHJtluNQI1z5Rsb8XP80F6g5Hymduq2+E5w
1o0rTe5CPBCfE6lmFSY2r7d4TC3mxSQLKsSjtKY06m85/HzEI2xvn4O1jQ7WJnJA
Z0Lm3YdqhMMjNWP2iamg62zjKsRzMdVvWjCqOIjke54TaFV5KolO6bV/l/MGC/vP
cjA7A5L4f2+j/KcYQAttqDyhKx+retU78P4uH7mOYHv0bkm1UUj5NtV3qYQiO8CU
G3O1o1C2eMsRebOi4q65Jnk2REXMmUw4uUCsm/dwJnSYJG78yxP35oVgek298YCs
jDE1NCqovHU1LOtcwuDruK8JFVTV/ryflDja6lA7H4eqZF7v/ubnUukJO8PzINKe
s11/XwK6BnokTlNoUyaW7NIwSymAo51ZBF/rA4l1eD3B/25Z3Fp+6xEFR5kPoozb
ELGgG+OuDYowt7rWSDEaPLgLQfcWhD/IeJX2/C8fQ0m9o9GTrH8PY6Hu2znkr8uW
eBkPBBjDumX9+v14ZxHopgh/SHHhCk2lUZrwZc0B0x/hasZzoOYHsnhrcUPkWHDb
EU/KoNPM0lI/veJa7xdnGh35roz7krOIeH3Vs3bBctSzJHqKin80QUCw7FxlLB+Q
YBcFa2rQ65cdskMu/4sJCm6GOxaTw9S8oSmR78L3Q2kvpVCXIzFqjB+7pDPZYDO0
Xwe5asShfB2EYpDcqS3bV+gFUazR7dBRmrF00pOdSx9o7VDlfH3hbtnEj9UBKPzb
0GQS7coeqsD+EdqyVC2DDCLNAcnltryOFT5463t+S5yrUfxF0//sbfJLZj6kg1Wv
33W/WRXP9r7TwtMRk86WBdMHdY/x/y2HqkVeKNPCXtbHhUJGI4l0y2BhWpVud7vO
5Go9ZKBWecG+p1g2yjWzbO3SpZ0AwsX7RnTzRFlxKCiZwEl61hnVrJPM37DQKDZ0
UcrqigCrFYAQPhozR7t0fnr/5KhSPuSRWlAdPTlvkrrxiU3QTrij3VWnTJXTeYNU
D4Z2xkbqloenclxQ1qmmJheY+lRp82J62D20ssVjDKcibFMP4p7Wge15eZmXAn+B
5kJnJYps8ojzhxjNthAAkZNgy0clVm8SJ4XVlCssMD/ms8pzKWl/ulq9qZN1BkQD
OeS9dXChYpyq2GEjN4q8yiaLMscga67iLhD8CcCtAvzB8C90RvthKHQtb7sVHv7s
ox0sBDf5fLTVmvllEnZQM6DPvp7gZiGgAma6dxapF0SZQxkrmyDEI4kA0VCnqgK8
ks8md7gtwTdQZOBuDGv3k23ZVt/JeygUviGHCcEH/OdfsVQtnDDzzYf2d+JroBOA
WpTEy3jdFzFCktfeh6NkjnDcqci3CPrqPRFoFZDS6nlOaNPQg8pGniXUxDnOLob1
x2denM4BD0BAYS19J60XG0bErQt+SdR+HpSZSQDUFSoO6HNfsI3jKUm/d00Fs9MO
72l2C5ZXjw0/ftiZg6/M4tj4JB0JCMUm8KivlmvKaxdwfIyuHbkZJyOZk5ZHPJIS
e6eyfMxDIYSmI9McMOU5xo1spe7bOhJ0M3qSJCzFDjSUNBAUUpBeRt2fXkxep29b
wHsV4Kj+0p1uqD85lvhRTf8ea/JcxShkKwUvED4J0z1zNRUB/bNqtaYV68p0yhTF
DkiMLZHkOxmnbcjaRhqSjbaFsYpMNUrMosVwcOAAWuU=
`pragma protect end_protected
