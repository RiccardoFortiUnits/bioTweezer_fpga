`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hMWL5AgJvhMqqMUTFxbYOLXj0MmrJn99eEq+RuD3m5W0BZOrb7meGS5tUbw0C+tk
MViF1mlXbYQVpVajguHzitniwM4j3OBFY50Tnolcq0srUKubbyIzgDALWGvfhbbj
HoJ9ucBXX9BLJ6LmLvEvncbFHwJd5sjQdaggzfupgIA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176768)
G3T+c8JXmFV9RJHgJ/bTnIQFqHpPM8M4NQXZ6vbfxbVUAeEhXDSfVxvn5RRsUzq0
wMxQZSvquuqpwDbY4brqXfpIVUnI08xAzYbji+SfQbxu+tz/9P95//RUCrQkZD7X
msjWMRPFQRxOQV65TAHpueEsTcH00+9Md++ukJDHRpxewj/SR/gmHiJs6NCNuFrv
buHEwP2MHzgPi5A6ZDC5c1Hve96uiFRDOuaZ38KbWR1GQbjEWwYajDRYCwRBwGPS
byjGo4BSP2yqBImg2Wt1RGwk+aaziFIVD/9JwWYqE6pWr61fcVX3cRow9btjEVEE
oUZt5ro1+drjhzBOsjM1zN5ALgmZdTQIDpJARcP/4/gj0RK8TWW1O3MdzJIG3IDP
6VV4t21PK080aj/Gjie4Cmm/FKNkLzfJevfRrDA/Wn/IJ2a9SXn3LTStZlVmyrzP
Ud6Gc1azblWRrmisbEIoSH50Q8iDktN/QQOVMY5JyGdy+ahGLPvm9xasP7jaZcLX
uijp6BGYvozImPNWozV2AHrdlIpwkw/WYG0UvruUXB3WX1pixX1oBlfVnvVjsyh8
i00xIg4E3CFcqtKkmxCR6yeKFcQyBPy7UuYymoRk7OGKWPeC27pt2k2opZsr7Jk/
TKhJm8J1A1bs6Giyh2J1HowMgR2T1lvp7+qs/HBieDGViN0oFMcRQDrTvTMMQJS2
+Qu7UnqU7grfthuikJlDra8w5n/dBtkXMZgoaLSeOHPnuleO5TLbUgLZwRWv9NdO
oWShCbdfWNXfKqW/KNsFqkbS/QIVslQSUf4BVQ1d/uteF6+2ZeylVhFRAROKq+yk
LH6abPUBn2G1RSjzIOuFB90pqlpUJMyWaE0XZgCXOCDZPbYkQ2jagOuQV7xcAb77
YiJtcCjeK5kOVGdJyV51Wlk3YOlv1VU34gPfHRFHcE6ulRVMy1G13hBJh6xcKSW3
evhaCczTljanPO6WoWBREYYOi4YxlsOJdaHP5jLV1kvcyWjLn+WG7IOUXrakrww5
dxCnllIw5jfEke/u90mTMUuDSHmrsxnVQ98CHAZWCrmnjVPWjzEFfHu7nbPsLhp4
xlhAeKVJ5bXwVS255sxNxl60YpZ4DP411/z2B3rniHKrzGRUryDr22Pzr7UHw1Yx
ULuVmAzpTHeG3RmFZBuJh0hvjiVYHgInwbLaNpuyl2d8WZmowjesiacnec/nSCCq
5tIaTO9e0s/FzQZviPKQuNRB284Vl4L5dvGdNoADDDvLKAoBh47IoVf/vx0U7JJT
soLUKGEkv+hxXPBDPZ4FTzi6oFtFyX12U+GlBlzuSrFY6qOGY2bIuFfSGfwyiI/z
N58vxygbfHmPB94EgBjF1kDPCbBisG0dMQ+G8C51fdPAkwQclHUduOD+PhDqsFuU
TW/v+Nb070kBo3XpotxH5/QefHQ+UrKtm9ka8JZRkdfpLYrVHWjQtDsQCtAxV6Q6
hllZR8mRYCsjhRywdij2skXNxTP8TbCxks6QCWDiBTqvBzHieb+7E0LkGC3GrruE
6q65yaLvFtGeVyL3OdKcSk5ZsIkPtN4IG7dqERH8j0VQ7I+QguF8TzeNZShsb+zi
zkCdyc3z8Brr4M3GsTmJOc3iCmSMahdw9yzCSi4sCvPB+dH+51GIeFT01FdjOicE
y3ezYrCRYguoFPujOIe2Zu0OUOHh1wYrC78QSqkX/H0lKGEpJSyFf0avKWZLiTGR
tFPT6fa2H4o3lSPKvDjvpSnVNmDAuJaiy7zxi9/PBCxvq9erk2af7sS8gLwBotSF
QMVYbIQUZ62J3xx1iyKN2Cu67DA7oKUbBNfJb1HWmhOCGhqUaJEoB2FpDU0NfQTy
+zBIZR/h94M0+/Iqi8w/btPkKJx15s9qG9ysTFGQHSK2vm+2foDq8M0VhZVxM83v
gMlelArzevsfYUBYByn0l15tuc9vyis//0pwyENDUA9eirmNIU0GnUPt/+DAZrvx
A2360pAw1kmqFcblY6SRVCdhy078Ci341HrKkp5XwN75FPGfLWsmap940LiF62xG
k/jg+Lpz5668jfa7vc19i7kJrgLEOMJr5Ty7By69cfCBoZzWrN7zomz4y8ysC8UF
vjAzfYDnzbNKbbB6FD92q/ehJln/b0u7B/NUtcwVlCSvY5OYoyMcOJFacvqs1Pkg
lVU6783xcll+xchyQWSpt7IMfnOMXvX7qzdUJqPQb8GAR6MpcOV632ASHurFgyct
kpOD7c3FxNgLHg52d9Ri6ycbBR6IgLcio0wGBLrnokcmMVehh2xvDSt5YHVAHWAZ
qfEfrcezDjOB2Q1XGncI9BEbhIO9P92UePMdUN2lf2HfgDr9CsZdysFdYwaYXqKz
qvtHoy9Ri6a0f0FG4Ns1Nu27bhqutphlFJBrFrwUxhhbDN/F8MC5y+yFIVNGjT1O
wFaDfQ1uw7wy9Z1+vkOSyeK9tvIEWOHylerxD3S+fKeI15voJCtAiRmrduYt1Ksj
BbvrBeAqnaprdII0uoGup12nc5TycBwvdcE42BWzPpw+GugMFD7AlTEUHXDb8+vW
G+WD1gdMUZiWsfc/xSPy2wrdkO/OpX04N4G1PnNgMx6bpj11O0AcJTtxxkxYwYQJ
B0ofu78+SrJzB//lr/fvaZoOWsa2O/pp9uH2aFCKl28zO6K8EhDuvT4OH9wQybfV
Li7gZouLsmzHN838205CUwtUgcbJGljuu1kas9OcCTVVr4GmGmBz0p070cQblNXA
XB8xWnMY6WD+cFMxPp57LC6HEGdrFfeYIo9aIEu37v8YIdpvLefP5jifIEIPzwPS
De7HKw85XIE3Rd6bdzlEnNkXUEIJ3Sw0Lu8/ulUfC+JoOC+DzsRIVeyXcLQ+dbfs
U48D5FcDptVYB1z526Wv0DnHjEbzCsEuh2lu+pFSlzvQGsBQ9GTI2QCNEHawK1pq
dpSu/omsHH/eJUPPsexddzslKWjwZfVh1HMg3Z4FkCkgKeXAV7KWMwj/5zBWSL0M
5YLaFik+zouaDH8sMwksKlCzAmpohBVopdvEK7mSnuhlFvl4kwHxXapqGon6UaAw
et920cNTGG2fI3Sptv+DB0Y58FxjZPmerCeN0IFM2gWjqGo7QHzCytNLq6iluJTV
cZFRzNEhh2LUXL58RQlak7KVebPxubIL+TNmptQPsNQ/3yob2ac9lCr1km3/4CVG
iLaTUxunkfwBY25XYXcVR8nuZO0O9eRctNdktdr/0Sced7ZxCII01UucXYwUu9cW
NRJexOWThm+Fu2GYe43ziWKfhePs65gAVE2b8PmniW8XyJfvHyiUFD2IMzlR24vx
bc3i4KsTte9Y9V5QE7zUmdw01IbJp9jNh5AtM9viV1N7Y/ejYelyQ+BHKwS3Nk76
rSHoagNkFdhuBDXD4VvTXxRvosdavzoVGURuV3jW9j/ivH3NWpQ0bKj5+gk4JLwO
fT/ZeziCcCa4imOFNWD5xjZWkcXmMAlIA8Tgd4V9tIdPUZtGDPszU+gMFcgCHXPZ
3lqyka1itOHLfyCuLCsQIwWs3AIsNcZ0sUjFVXyVcJSYfCyAvYGcFmNsFSmgBgUV
oTf3EJWyZ4mrlCocj1lGCWNq2NyTQowiGRBzW17P+94mEsFtSu8RrC4rpHswGtij
InX+xn8YeSUgHNk1tL/xX4YP4ER0cae7deWeu4BhgAKcVC4yWPI1zu9/n10Kiu/m
mjcR92KYmhzP7FAnqWy48nSo3Fct5gmVAP5YbI68znt/fLJiIe125gmL82CAZv3K
xhflfiYum920FICEYuVPCedIsM3Smu3/lPLA8Gi7/dBcKbnRjXew6T1ic0V9lduo
zn6aNYe0u36oYuuO+P1ZMuwfwbRkPBA3Zl9r+OPEG/sauBInK9AeoyzKpkMBuuWr
4cyUCuRgs6hLE9BtAzed45JxS6Q1HaMru6x6pJwxwahFwDGbvK3UJgozXSZdb050
GrhD5i5/eQPHa1OZ6uMWiqvtqct4I1IBDUqEGo17rRKHH+THBemhprINFeKRwd/5
26/KroyHdMOP+RftPyQgUsc+1o7/e7cPV7QaZEnNd5RisL6tZxelrOF9dvDR2oYY
GpqTSIM4qn1GJHmHIJVKnRoeLYkDsTZ3wO2iNeLDtu9fgAkbzGpPykZflAOa1uMu
pCobgi6L1+xFuk7qr68kaXwRB0IMaUaLuMeYZCP12hvxOa3AUHOvMLwLSm8vAqzJ
WlgwiiR2XrsmWyRKdo6zMDLdWk8DR5SI8LehEZerMbkPzTtCGWibPlUp7QFAjagi
X6KMbH4CnIFf0ZnPUxaoRvviwpl4E0pcwnzC2Y/dNLtEw0DL6xh+pVfqI3GR0Ec+
9PSYbipKWPHCvgeCvS4OdzxU/0dTooytOS9YHJH+wKFIyTX/oRUOXaBi6glaedVB
JdF2elcY0KbmBsiq3+M5yX9qvs3OgcI185FQ33+8BX4onGErZCtK6m1S9/vGkJSY
+EyOJx0V75+DwO5EDXzdzew3RJlezxjEa62AX3wgqtYbLVIg4u1pc7sxoMo6ZhoX
5/Hpo+G9hDGb7IYVGwzftizT2m9a2zB+Agq9IALZeQD0vprVHBbQ/rwmaUQIcU0j
vtywIrFmdZMtKDYNX5Xbw1ftvyWOv7o5O7wZx45ulwPtXoRnN7H6GVZlaO5j/fnp
JRB7IlulVwxcU5X9o+Bie9yATvDP/Ffk1/4uHqDrxK47bFjH4AXTorbJUmMPCbJw
WuUVboOOBywfh0SpS6yUr9NRsPRxzYOYVTkboAeahY0ImJtSJL1dFsTgEUbPWw63
ZjaOsdJzK6kjo5TFCNfPXnbUxKSKG3vFA55hI0zTaCXu7TbhSjir977b1LHkzVpE
OkRuR5838B1p1mo2y8BNVVYsbNIbIGU3K87fU0gEVWO9pqoY7+yefmqgiyVTUQuZ
gy6bP12bjixge4TmnfmWlmPr8LjVjgn8/uoecW+XHLES/VLag8qqRyMVU5+l+aGw
Wp9WPRC8q5LMR0wW3FcEt49B2JFsZ8TG1BzTjSCjS7gc+zdFUyajeDSwtH0Yh5yL
+9RMdsACEFWDViXtK3X7HIUEiLnyj+hKzCU4aPcBO2GCwvoczLiQYevYe85+TaoZ
iQwF2JgYZvnhdIVZknjH8x0kyQKzpbd03PmkvX3E1mN8pbbW3wNjJLvooOHm5OUd
wm27WgVQ2s/L8aKcE/FHhh6CytyHJ22UJiSqfY2FxlKWY2cmVnkEEJ9WSu+wCLrq
oO+9dBoq8oBOfLkB1t2UWU2LBo5ZyoIMg8Ok9u20zbrt5TIMWqRoW8zmFAluA0DA
z4aDS6voNDwIuLUPGvVh8hNctj6BtWstrRYGpLF/FrI3BwZQcsx6JEMxxQ43zuzR
gmJmdEflpYT/r1gka6T3+ZfEeRmQKaboAOi45dLjF//QGw1I36XH+9Mg+HjEE+/A
ASKniSw5AXLi6+wPWbgEXcyMTXU16CFfklJb2WoAbwnbNVy8CX7t41A/3MNKKYSm
IlVYn2Cl7ZoVmGG6iZfmhVnZNzverecZ3ZykMb3hNWM1XI2iSu7FmzsT0nvvRUcD
T+l7m8Sj1M6ghccQ4Ke2jTHPFvztpujkXUoUBwiVc3mx1HFw4J4O93Aq4ICl69lT
3I9sRjFNAM9UV2pMx3XhdMNxZE7CpzMW44xH11MXA0SCWkTe4Q/6rdbwoM74f1T0
FJwjwaG8dTaJwkOpOOUGUxWkZTzSCFiG6ALziwvDnd0FQmPVkoSY+ZscZkE4nx+Y
cO/JpMtSOXmAoPaAHQZZm191k5BcJ0ENn2MuH6WyBkpfNzzmv4njDdXKVMs5EGAZ
d9bPi427AU9vemhT+0SmEysZuyiNVUou4o0PDmp0up2boXqu072PjzL6Fl18ikui
dUjccF0eHzoTDNQcvGVUMqqzHGN0ewX/nWiG/YQS495S3R3T5HygOUHR8pM/PmH3
MGrjTwnrXF1T85g69dRGZitQ5M67eq46QcK+joBXftihCVXphoMCvwY2eUTH/8vV
WixXUJadWdgZel6Cg4pbmio7S+U5ebsyUD7fMAsEP2Ntz2Y1xhwRGZuUfouuZoeb
2C33q/1oEs0SSwEYajFE3xPWETMgtK8s/q97JzJpwR+njOxVj6Aj7poxRKjAVH8I
zWrtdV8rMA0M2BIgz6ThTNT5PYw/uRWJITjiNQzMGVd0ltAHzEGgPVV0uGeH+H22
e39z58oA0L4+TPOC1cZEEVpWZZelu1sJbYhX95/ydyYIKbIRKZk5/NC+1TlxAg/g
u+LgjjaN/BqQzu/gB/urkZvtrsQ9WllrF2I9cJFV3/TD7mTFFIoFTWBWtQvcuOhC
aC1MAxwEnQK1diS64B8l/tbm5VbJhQV9gewspqpMS8uvcsoEJ4sRC9J4dEEeCgRB
BAyK2WZSrE3HONYcpZi1v7jkgWVM0zT2pY/IL9rtkOmnqb7ejJ4UmYpJoxhjI//8
xuIQ/zeU/TxaTI4A6ifVno6r2h9f/MFEsq+elIIjvUYCogHaRzrLV4RBnglGAYdU
7/upK/DC8aq6k2XzacuRO/alpMuo7GAkhOduXIWmdqaJQ/9FvSaotR5W8pxiUZHt
scZibJck3GEXwUmwXnrQbq+y/rx8h7QmyVRgHG/YWLwpBLmONzkoRAOOENk39ca3
3ggm6Rx+dZoMt9GGBcub1/0YntZkNeIsAk4lj2yNWKpgs28MMP+QqLFJ2LE2cQsq
BNDcuFJBDW2AuuPDvlqI3dhecjEci3vhFFgjW2P2TJby3x5uwKsjetNsihxqlWXa
3xiCiELxE5CA0+2SomLs+UgsEScVp1fZiAnZUdzcSNJo6OFqw7TpsbfRPDL2B1/+
45b069PWa1AZStCrTXxWDixOQCkVvIrgHlLNs6RP68c4sX3nCCKDEXwQg4a6+sbS
2WQw0CEL+HNTsTABol58Gush41kx7uaLXUOMNa8ZQgG1qAUaLXOGTxc1W+R6/LIe
QpBU4UWsqXXkOeULaFiV/oX4l04pufc80FNadpfGhsqcWfeqHTTzLRj1LHWHVXGz
Hszb1GUKjEQq0IkKUHMS31NUs1dq2Qj+o6fL6PvFNunxSptvYqFhDBSdPXqz0GaQ
6IMQJFy3llZH7o80h/Xr653HoamlpRnAntMoI18vhiJjcv0p8vEjechP7teH0ehB
tBwXegRk34QIwKHVgDYkq4gGaJk3Fx9IMgMq56J9fhl/+p6tNeFBsaCjTCChMnQl
HtJjVnAZ3Cz+Crzd1vJM2ngukwsdMZj9FlLz6XuA26AwhaBJwUnCcKq6wbLjFPyJ
ymIfh9uEYZJgSfRSrCmR+VkmmIV8bpGe4dau2Uj/DImnBoj5pdCESETZ1PxL4PpZ
5laBfF2eEwDKgP6dB38P6vvbw/SbjtTzgsPeW15+kIBO7um2rleMQd5u8oLmcnj+
gCrgZSAu/rQWLBO9zJBF4znQROGrwLrAnYYydB4m91axpqlcq8KcFxbE+zQZHz1C
hMSPxWgCDV8XoSrIVwE7j54dxxiY8Tp9CgM/b24KomH/iHeuArJS3iODwFHYa3UA
KUdzq8q24CsR2wewl/0RVtRcHTsgOLrkMxL6alDEVkRRdsrFFw9dwXfPOj5XZlEj
Hbn8MgFgQWJS3zt7ci9UFgFF/vOBbZl5LFdNM0QZ7eR6nIPgSjk6RfzSKiuKXGSX
bg1ZyLxoHf5FBP8RZengz4EDIi9az+KvnkxK7hllk0M1HzhyCM1C5lE6qgoSvj1E
qnok3jmR2a3L+CCoRro1DhHYggAD8N9gPZhyLS1zqsJtCdM9xMYjwWAxe16OKlUe
tM+aBHRMDw7mHY/oMncfN8Y3y0UwyCM0Mmki/YoblyJI1h3CR2gL4zuVDhk/RVsJ
+7N4DX0e8lfGE040QlJMs3oU8sHPZGmEA1tlWgcHXaGvOcae8xsSya9Ajeo1zw5z
/LxniyOyiY9/iZBMfZORtXje7+VIAvAX/ZxApfxwiCkKyfgAr+AYKGK4gASMOKmf
JgnONLoLu18EwqqhXZZXBH9RdQq0F/qDadQ9m98beDHFtWPWaaBK5+01Q+gBT4GX
OdT0etf+aaZstqErmtSbrlqZe5s6tY8zDBbbLnXjayHZ2M6rcQgAbzkVPkWnWFnl
LGQaZyHcrJJ9Xl1cBAM5gtsmEj3PnKQEZHcZYnKwC1+r13mvacgNSBtMGt8E2gn4
HlIKT6W/v/lrh0w3kPF6LN/WaG5GXccdTgxVGONrhexjfe5rAzZtpFH/Mw7OsIwP
8ZqcrCWEfEmF4wsPsbw64KRaF+IlKhOFkCTN/57aD2DN/GLfSZhK/bexN508+WOU
6XoJAB2GO7uFikDACLZ99XdsCJkZkkacsAKbvj+f9vWEl/Nd7u+4AQd0KIgUHqMj
wnkq/M388IfhIzJ1var2PGAk4N/+bt/ldVGJurR4YLCzj9HpbbMxfXrG2MsRvskq
13HIt6heD34KT1Ea2EzuVQ3SUTuO5M/EgDyGoLNBeN9KQi2/9rmVAmnHvcXL/g7I
nk5fI7NdG1eaXdUd7XQZJp7Lpf844s6S9BScXVnn9Guo1LBo8PfjTbR5YXNDBmLb
SwcKlmnUS82btkM6k1X0iA+LD5rp9Ch1seKTV1n1v4Aj5s+rBDwnqKFjcHlh9qp1
Jh6dGNr8IOsjXWw9r9s21Tqj2xxQCkjJngGZR4B5OFZm288AHeEA3ccmGmDGWmFO
W5xn1Hn6gnLTwun2UQWtao662iRRhZlTraknwr2qxQdhBmS8lS+CPLfgeZGkPYHy
TlvR1heSTCdGqX4vxI7yQXRt135GfBUAQjaBnIKuOgcZFjD5Kbtd54vmZJ7lq1nE
2uz4BHkrykPqQ+/wrYB4bTnS7/0H23whzNy/zENwNZm4ZTEM7q3Y7UxE4nW60xal
ZNErxqM2roXuZBvLIcyejevFCAKVCCePjd0h2KkeBeLUq76p4DSJv4sglkTG8UJL
s2BiHj/NKWdw1PhmECZUt0vtdmkl9NfTHMvW87pdSsayNb1LJSGclpZ8EHWXOjK/
Zo928yCpxTq4goMJNyuNyzMcj6dpvLR4cg2at6iCBMAw6MJSf3lieCk72vbyHqTj
+WWrwVdbvEbsdvZfdUR+r3PBdwChyR7/Hu4/jLyq9Gs/xngFjeeeg5Fo7yyuW2pw
5SOqVUR9msS/IF2kRDX7tMUT9pk6O8hC/QEZ4mVAWq1SEYGrD53Tqce7oXigUE1F
drAzloGNqdZ/i+kQiLIstlK09EFEzqQD7TTqAyPry6nrM7A0bRei0WKeUTIig13v
Y23qlmQnnjxtchHxuerOsLiSsQLxk2+TLnnC0KQe+lt1E/x+fkpCqqCjQ3w0PlPa
yyc3CVQsPWPiGa11gNiOtQhOr9B56rWgDL/YNui7beL5gLyq/wLIgrEbL8t3LGLf
OkNL3m/btX+/X6aWpZm+RYa+E6WndsYLDI4ylGHjUIeHdEH2zmgGvuTDOyT/16PW
3D3Jh4v0t+s+g/IZygw3lKCCordLim8pztYhD4MbryEDP2u/LigbcTpzt3a87JUA
inIcWbAxxWhFf9apEF578WoMlz2fl3wOfGOclqkMCj2bUK57/E/xbTMTyWPVCg5M
zfLJppJQLeA8BBWtRbS9rPvPzuN9VjhXlj+MVirURQAK+k2IZdx9GFjvS2Gfn7Ne
GfqD2K+iE2ESDDjb8pDQjf2P9LVQ4EgGCSOFmhLk34/NuknqslGn41yge4Gq+EOv
Rov6pTiTgC8dikWcDvqzaoJ7YaiwMlGTNwqmlMNBZLaZZIrlOh4JeG6vEJDu8jsS
4tC4Y+iHq3nRA6BURUcOZMik+cFBUiJylIEZi86IxpmNJIYLiuMPk4Zrqk9tatNw
yF6C4m1Nu/tzCVjNqySJhIi4uiE7sxQo8pqTqxoPZIGkTZ8l1OxF+cvVDtcScJCS
peK2ZtEj2OkxputcKsx4oBpeo6vsBL9GYDlO6eP5jCjVpyPw+O8BT4Dakch65HH+
ll+p7rSSjhOVXw4j9UemdUE3BVQdbPKDoGrItNbaNu99BblfSpkNFV2wFkY4aB5q
A+qnWo6grwKoat4XKpIe2W9c86y5CW8pcj2BVOp+4+E69BMQQBLa7/IfaEqgKGyL
ZuSWRZO8fbMTqJoZBtgMKs6mcZvDNxSpLj+ZeSh7LkIUn2Od1O0RaAT8XN/t4Jb+
VpDEOCx44t9IMnFht2aiaNAAhXnHPfSPM2z/F1N1pqTfmZ5LDfmdw28s4AeDPwZY
Tiu2ZETv/mgJfQ2bIj0ptONCnAPSSMVuuDE78Jlt7ivseZMlY/Wheq14Khtaq12n
mee5E1puqni2oUjxKap5BpLAdBK+Jwx9UuYSAmefj7sjo4D/hZUz8UGSQ7oiiy6j
nnFB8HkZ5mRI80F37IEcLO57T5SooIpIzwTR1UQERiJWkAlPDzZQdmev6nvaxjXt
GZMr9cPFBOZInw29K07mdT/jmMbBMRstnHmkff0wjA1IhtJfTm2KICHcYzIqgPSM
8eZwYWHjlYsV4mgLHRBI+UB7SU2Lq0UuuNnXBUgzbs/qytYH1+yBTS4yiWEOmcmR
/cVZdMLtnUH9gO9LL0hqXWDrF572GT5xtpiH4CWPjeZz85PInSgTwCFIUTdJL8Sp
G0cYSAOUq/BP2WrUH8Wn+t9E2nButdzUp9K1ovHbQjPXjyDjXFP5EeCyIe8ZZl5e
TCU01aZUg1u9e0Q57qZHpSN+V+o3bu5pUsCDXzGzRC3nveGXNAtKx3ISduYfKy85
qkb700DUWfu6nhn+pDodduenNjaItgN9pjsliNDhIekKa0GQQ2U7OWpXhRvJ7LFM
wtbvG6Y/sT8YhB/TaGL79ymPeoLmw79oL09FdRuQgON/niEd4M9izxucwEclhbvT
7tMPNcCdTdfzskFJFNe3c5eBTHKOOv06vjM5JW9aOURVeSq6FKlv2zBc7QepnR8R
2Bmk1Tlq5nsP8dviExOOabRQ5Q4HiMHH0MpYk8wwI+CqGem05sOh7fOMUFWDAKk0
kUJCcpWT4sqDfZfvll7FfcjqNteRPlnHR/OJx6FmvJGbDB9fbKeJ6WDSduyZCoIZ
YuNM1OVBDjKcfBq52n2YzFE9IzxC7DLkd0imI2V9AMT75ywHOveDjSuCj2msgj6j
ZGIo1ApB7GBaIe4JJEvQpgMLgJrjT4Xt4Ww04AMzldLRdMG/UQmTuVgXNJqK94LP
yp9Xp9Rx7tZ9V9mImBJy23pImf9LI0C6A6ZCX13JZWK2e2dzYkfKaMXJU71fxIPp
0rqTzPCUQ+8dwZuUs/TzJtvl7UmISbbi4pRcbPwzp+pdbmHQ7wn/gxI1Rk9gq7ga
2yX5dtFWTAeDkY2b7yBwNYTPRf5gCYyJ19A7IuN7cNtmmLTMDK4zEv9ufI8eUL7Z
/uwDjgWReI59agWr/WhNA74RJPLr98hse5JVmenhIM114xlvLYt8lWrm50lPKg1X
dLMfS3JFUwwvHU+c83JO13tEoFjvtNNbkbw6JuQETsBiLTXASrQFL351v8Fqe0K6
AvlNQJL8Gl7FUgvqCHrB/yhv/48snv4H/CMZFRla12ZRyYhsEp/o0AanrwhUDC7h
xO6aRrcLSRkw+53/00AjKdpq2/ZqO6E6zL+EEoZU07EVcx+h5iioZ4kefEIsSycY
K4afBlPhmj0bUb+GhOXxxfwBJQM6x+unuwkOsAAnRmCfhZfqyH068mArzMEa0JtW
LiDmUrf3jVT5WXVyJ0pEZK9J7qfksKYwkMIgg4dQi1/Iz4LlURoI2XH0KzM/77bL
Ftwm1Rydu40pIweGnWy0J3awgXtx3vJlvGVntTp7Gm7LuseOk2dHiBmHOx9QVMAy
VYQkXeGQjT+KLGFnx0NdSkCochYMYBYeAVB3BfX8mXeGqLSODUrw8PcuSusq1bM9
N0dyvHJ84xWs2lSa8FgJq1MdDQugCO8WbkeJ0904nYVaTPr9+sNqFXxNekOVs7wx
Cy6jFXIESnSeYyYMAJvJinEWbTxQLtpCsvdsZB9N+LfaWOHdMoItcQfJuqqfeDU6
I2Kr6BlcubHwIo83XhOvSKEqKqzBfVWGPgZL4T3BQfQEteftByhlnBzYOHpwECIg
gzdP2nPK9pFq5+M4YYsSytjDG8Na6aRMNhVSjSehUN3nO+q7xKAbhAzBJ/8MNq5c
toBSKmiPOMcqx3n1DuzM7fhU49fHMzfdxDWMOhECHE/VHLaD+s8KH3oo+RCtdB6Z
/ger3ZXiMLCrYuL98VZF1xnxT6mmxITL33EqVww5RgT43iKbK4Bid5AU5Xvc4lX/
nWT/qMVoaaZVOH9dDAdKkN13hmgksHAO1Q1ufjNOEsa05FCmihhPMCnSZzxAbSdM
p+xneQGX+UZ4OOCS7PVcFRfBuqo9EdTMJG2n8oL2dcvJ2jr8C6JZ2JMBnjfuD6uh
aZ8C26cOb0VyKRh7d7I8NqjeDhwSljF3CZP0jmVqVUTq+rmKs5pfalos93qpGxhe
Xr09i4pjk+GsF27sIt7J78VsQnpq5c7DDUD529hEo/vG2L0IBL4oa+CVzfnV444Q
hLV/JV+DtNcAXmLo4/Ud6raTQs6pe3BF7ecILR9XDWQYy3ep43l356uzBe8jmUcG
U19QiWUHAGqLgeHOUvbFgfuOr0hPlj7R0pg00yzytuMV0cTCOka/O95xDNOMsWXU
jn1SJDGaSHDJwAYhU8RfXKMjimXcPFVmQHTFLTNadnrJadBIEBkcrQvpItFYWqDd
2iTJjMT/BW7XBl1mU+daO2W3dIITYCPKvodGmC/X4ZXEIlH7h1LvYyFX3Zrc0Jhi
uFEcfJqT2QMupFdFOit74la0nCSbdURxvLXMrWAnVr/uvrulxv2C7VdcFW2QOcbc
oj+cKEP978e4zb2qTvMA7/bz9tqxfLJGPw0/7AJL/iiS8AV6f5oV/okB2pQaS1hX
phA+fmPgdJ/a1VJM4rrsYJXPLYDuMgdZ2c3lzaJxtmJ9XmJn28zGklWW7NG+uNro
nMIjla2DWOcWCzUYZycmoCkKqf0WCmnbjSxev+qUq2POoukImMXNPOOO4a1Ei7gO
hslJncLHMsXSUsHG8hlY4FY5n6DTLaPK37H3ZTDkFEDV9AiAoexZK2iE7Qaq/Ftt
+FK4aDVbml5CEAJSFdXYRagX1lFYA1mfO/ddpkuJaJcyozdkzmbEsknGPMERQuiq
qXAqcGdXGdOHzWPQeYY5sf6UjFBASijXv9Mr//Zim9t3DfzO7Cgs5PjGK5BATjcp
BXy3czo9N7gC+8l16IOdMRiSo8yY/GcfXYsggPm9+rZzMPJ5QAysQDngoYcJnv3e
4jpdPEhX6b9/raZT+5+6FZ5Ef7Wu9mDMo0wPnWrtt73LWLq1RCEAcL2QFeBP74Ut
F0CWaAWwAm7q+kwhbbVCkd95vCLviN+sxTj++AQmXzHBpNGDgRS9HQUItuUscCII
0dk/7lURyZHUQAqzdYmgcLJ4x7Un3RM+j6+40mV+owPqMkqYbj9bOxmwljDO7dt1
tNkkvlj5eOYaRwrpEFLmj0YhKBL8TFqdZk6amJI9KJjcJ6LCG6gPb8LlPCPJfaxU
AAXURjNxetN3EPSTAQZAvVgVGpCFU3EJR9hX/NnUDqjQwWF8Bs5gDHkZctLzmHGU
e5sYN2fxvK+B52IizvQkVfpzv/E6G2KpO8hCMh0GhAKK6/8QV4cqYy44S/iZDtxI
wTLVKrBLIp8fczCKaGDTA71Z6UUA7ReFl4DwRY19ArK1MxTP022/yiWhcJ4VpBvt
UxvxFH1sUegIiT+2FRScsbocSE+IjOZaqw5b+WrL4cvJ2EkvqDhACD/qTOolR8yi
7US+uoM/mxLNJ7Ie8DWHXvVRmxhd71jxiuB6ZAaKFFDXrn/xnzcYaXilxg2+Ky5i
R0EL5y8m/POhLBduamy6MJ3MJr5e/ugkQA7Smz+wCVY8sF3G67zqOfG8FMeIlYzA
uqnlYIloGSWq38pDlMQjNbCdIJxi0B65hGbX3KlXex8GGa3YIR78eNQCcofBCMCW
Fw02iGZvaEtm/w/xtD+tjOXDdg2Me+t1x1i6L75sLR4N5zDnaK2ZwT8hkp5Y1F6z
8rYNLBUrAd7dJ2gTcfxWq8L4xniZ/TUSvI3pgTSy+MwX7Yc4MGGGGncI6/P8DIKB
DcHNIzWw9EO4whgtMtPinMZfksVV5innTZK/B3pB/yuZmbkUGG4l32zvmg7NTtZ8
WOs+vt0qEDXyE9txsuhZqZevraJ6mBbXBNHi8yG+uTKM6pJY4ANfT7F2QwPd1Ulz
dJPunwGejKhFvCriYSTpRymLoyiuXdWEZpm9iBM0mGvje9327CJSSQbJbpyeWHlL
7g2/V08S9vIFfG5h9IdFElpUsf5LnmzCQblZoahs3lC70zeUXIWespt057ydQegd
16ctQVcOKrQIEm4jOgGbuJXuewWhxGMLHIiZyVgKOX/tWI91QJJsdMldQQxjikjV
PWVqos2DgxTFtLqzrWk6fpHVgTzJ/KqRESXbRrgEkSNXBT5KrWu5YllcBuCXqjhz
iBab6+mDjhT4t8FToTuZS0IktVDegnpHvy2eydhR+31clBc2i0sTDUyOCet6AkSR
GbR3Zc7VuyE1MFwgf/4pU09ArkwGIg3qYffWh2km+yXq7btBHu8cIkXyozIzZUoZ
m12lDPmJ8QmG5neNvAwEMDX43O15ES2y4duJoo/AlBGoKPnQBzfv486I3Inp/x7e
hDNj1TP05JMPRd63+goOGk3HhaxrY/yh50oBicZFLncja8Zcjkf5hFlh9LhD0Hke
K6cFst9Q6PT2gAuOiZVjkowfH19p0tlX53n2NWpI0iGqZkVoBUGskUP073+L1Ced
F0gPO751cmp7iRnD16uLbkUrVRwZXC+S+joXVwFGMHxHNVyLFldbG02mPSCpTty0
zc3r340qskxKql9IKAbPTAsvwqSuJ2zDMKigdF1jV9tfmLnlD1Iuu2HLopV6OXey
XkIhemHHXi7bik7T0Mi4hhH86ibyrrtU5eZ5+tR6lLhG8HPu9aSHjamWG2aH/HzC
Zgi0piTGiLtT6vdU8oSzTyMAvCMfONFW+4Akjkr4fpBb8ItuvHZh9Ie6C+w/4tfQ
P3qkNn8vIMLYVf9Ddr6AqaFB1Q7z+0RZwet5cdgU2GYjf7Wq3JZMXeJbEZjvMecK
9gzNlTvWJSjMR7zOK0Txc4OV55i5gmj+zD1U5gAT1ketCyuwcuQAebQvHYkqMWfI
+nkwoMpJFlD2fVKCxxGjvZs97JMGh4hd53Y/FWvbwf1DmFoFlARDh7g+PAdx3cAj
uS7+eA6f9oubp+te4cifoLEQd+rsvR2KrABzfdMo4dh/2C9zAW6Fr2wUXHaM2+Pf
VbtTSzr3YSqA5PoxCZqW3p8e5aOCup2gm5DMtO5xrbKr1EsarS1Oj54xfv6M0bd/
OuJN7H6IdQoXOtCAkx10Cl74+oHAKwWNt5US0D3yyvaWQM1stWBebp0nW08OIXAg
2qh3jXxEhWHMK03tTEL05S/1Nwe6adMd+bgW+k62Ay5NcmMR9NV319eu3y15bAyX
gdYZyS7Gaa6kN2QFDBGjNod0KfzS60rNtBLQmKBnSrdP6ze52KZc6v2ddrjrIh5M
wLPGTeOC+bXhyjpE19y7Dgp4Rp72YIwOpzuHqkHQ9OfrMKrXKjmlv0GX5f4ksxAj
ys89nwr85M9lnt9i5ODGUN+WJmjtBa3hxq/qIohJptAPB5m+IEdhDgHO5BZOG/Uz
1j+6xQIcxW0a8aHwZlZMcOwkhdw8cYOJXLozoYFPy2BixPthNeBcW+eOEx2TMqLu
NLHtr1V58dfCJ1519m4ct0Fve7eId9dxxYyOjVSKi0qT4yKzVVVqQf2EJqCWJB/c
pIKyaklFomvmcs8rMtTDMc/uty6emVkfZLmR/OW0J6ddWz8MdAJM+nfnuoIDBHBj
uiayJuxW9ImhSIVO469QFsdsJW/IdnN/wzCJ30GYONJUCgunpMd7V6L6uhbAjYwl
fPznLbOLFNX9Bw/zSvoUfgUJoemwO83EGppZxPdrOflF0yVy7vM6+/wz2qyr9P2J
NpAzjJ8RPdXAIrsiTPsN4i8Ah+PhoBL44QI37QcOTb/7wWVPvN0Vjs9Ew3eMZGwa
XwbMmB6+dBW8sbSckbxrGrATatlZuep2YjA0H5H2o5eogd8A3HNUyNTHGk/hXlsY
9qhHcJTWSiPDlIOPedTUqDZvGajsTGc01MhnIK2xyLF61S3osrm5Q9BKuLZw5oX8
gstrE5rezJJITwYBoss5QgZ3KLzGBCPJv0JRVin7a5yG5eZzyMl8dIlrViPxSCY6
4he3pApwBXqygvaWqP+Q/1mgDMoRacXjcCu9uuRxQTpt839m/J02BVPiCHWCr/Js
pCSB/9/R8oMqQ+kakmlrjYAS+0CDnfkCXgGX21LgGG6s/UfyEmaB7DTCoECwu5Rt
+GyUpAO4GqpEXRv+FjDMI1XujDisqRhbsBuXVCwEA5MdfRFIVg0cSlPngS+Pq1UQ
nJC86NTdTvWBfuaoIVf6sViQzzNeJmcE5fsfyQm06sHObCJUW6IwA3e8OndUZafr
EghMual+NWcXxxlB46peEkQGKVK8AlaYOlsbk0p0dlZY6SP+xx3NHm7mq0zcStc+
WyMRfRwSJC3IfwHlPpGtpKCpWk34H5QShwIdTcx8QwiTLw+fEK767mJuJcd/DO1b
E+6igEgcC7YWY8RnscQInKtDvbLGX0nExAKw3PplgHEtHX+ecSHGFwbfoYh9ivzq
LZNebusbDvzsvbC5sADCrln5L5zOqkaW3ivmbjnJQgcZ2ls/l3OfByQuvX1eKJw0
xCDsuK7T4jYymTkUzm0pFo7/kQ9OAOhplPhj6ZCjjuy6ZBAFmPv8hrM/L9PFRFr+
wuRH5EUPansvl2JkP1yh//c1chN/4qHxXbFg2TjRhYeBTWv04zFKVnxX/fDJfyj4
tBdtMz5Wy31YAVzj7EftTQBbZ/8T6Ts0rT7cvzgxfVsUKL/lqEkCpZPG9a9fbDi8
2Avyv7HeWc6Hl3z7OGrF5oed3opw2wRPiWSlQxg1nZKu3rq5xYcdWOu7Apc1buG4
eERHk24GClrJWD2xrJaj/KcQfhqWpsRS1E3/9Ospb+asPfe+LJ79XT+pTQGBE4dg
Jrwa7QlLbLZnf6vjDVYQkL/bZDv7vnMwaaGyqfy0uMlVKzDPa1PG2r/wDeonqZBi
1VxdugLHs/2OCH1gn1J5qy5RT7cFiNh3dV8zKG+Azrjjn2BnQ+iowv+yDbGt5tJV
zrxERr+lYhYoGbAhigds3QvwiUJ8HSM/4ZP+S7t1HVpK+8KZrdec9namjLWsv6zY
N+uzAltrKD9Y+oGbykw5oH14h6xCeOj/5wnRWBgqAYhJJiDCxvkbWWELQorEWEq9
tLGFCCPcDKQ4j8TDIB877fFhlxzClMf3Ug+BCMM5e3+irKxFTV68KCGu4L71Hetq
q2Hlge7J45UrgMLVEOmD3NtzBN4VxBZIe89o0M2mRAUXvEfiUpoMUDXrUYUNzeEf
OiMgLnCRP7k9QYPt5O+MZ4aCXLx59tVaLKpPfjQldTwV8tWHuzyqCQR6r3N1itFl
4gC56xs7HqkDLju+I4MzPVgGdYPJ88jJn9WPkg2lS/Dv1ljBTlGRiKVBB2Oyov/X
zeoJgO3EsSxmpNbC+8P/zitQRbSeP9rn/T6Tjr6zVwl9G6L24KAkfM5nsE30aG7L
oUCcmAzRlTiFpvjrEfyoP8h34XK/fKNKJyND5aY5EP3n2osHFq2pMdo0Sy4e9PaQ
MxBQB3PwndrUVreiIEn3CyGL1bUXvc6QRGn6Emd/K7iL6xj7Z22qKTt7TGWon3TL
69qLBMmnyj1ZqnvZQhnZK2tIidjbuoxOlcbDQs9g8kVP315xPPGgrKN4C8UOLcBH
yH2dfkqNRTGC6qszsOhehPbGmNFx2WJG1hZAOLYjqwsDlx07B8/uPlY0BBiD/Egb
Gs49YAKzqDN8xSwqwKRICfa6cqNhlmwkbhCxCizmqzXkHlHfx0NkD5Bwrg7BVrjs
Rkws+8CQqeGGGHLxtau+IclYN8qczla/6RYV3k/GszR2SX136LfJuu+7MxdutqfI
gD4sqBA7WQETnW1Qsx7ZXPVzkld77Q5Yt78Ymae062HuzCsmeNwL3HzTT8Xuw89Q
B3AH/DIgc4EoxzYmLPkhJ10pdV+YWcNrl+jq9dqszQEMfFOMoj1VTQsmMp06Hpma
YibLVuzRUjeMGLZ1KzjkX7uLyCNojTFLVVFkqutnJOaFQTjUXflEn4e2P6lu8WEb
TKO27nfikrGVg0koUcuRBjUfJgS0A9tvct8/jqUpLr8x7kbtQlK4bZaz0dzlCbD1
+n94urDFqyLR1UFGN/CObZhyP0fgN5hTG/lXhOWA6QnLOpbgLy4MMN7y2+ZvFnvg
AE5pKoox1ZVfJi8kGxWDyMprgpw/1kSNzE8B9Mf1El6HtIcxM+bqSFpj2+5tdh7J
59gzsMcbR/B7iPq7OKnAtFHXtF7PwbknPoalECjTFldKMBI8Oj4UvIF/08JAHOl0
HJr2a+fxIv9TzywxeIcb83rS9GxeW/f7JIuen4MHje2SG5LdBJ0MCEc7kEKIXnNn
8SAg/pw9oFKGM0CJQikFWn3fo+aNCUexKbvs1GUWGt1BS68mHdpVu6jDT3FxwOCS
s0rlwCfvmfZz/WvikWhZ0YruWHm+5JMFIUlcHbyMp3KJV8rC7MT4/cxBBvWCmczv
bjl7N/ZEuCb/WZKb/HXOr2s4Gzwefu1Yl5JaIzw/f5tk9wEyYwz00XFGthOToMTK
S3PvQLf/Cglu5kTtrR29ibz6Q0HRkBQnD4lZbbCWQRSEsHp01Gn98IZMX4U0wvx+
DIxE/hoGDzfyn0TTBZ40/SSV1NOPe7EurYE7PmzeD3iWYuHCyB2NoSHD2TsI/xV0
sNxoBIsvVniPnHDEEBNbrkbOlo6yRn3/L63HbfGi/dUIe4JD2j6/Fbifd41qBbBF
nwjviMBO+KCtyKxW0S21CYVP8IMt+lw1MZrC5fCxDNeRrfTuBbvXppQw4BBwt7Wk
icBINMNVs5xFliEeoLfLtSiOVuOf0LpDi4WYZO/CCkDQzjR+zY2k3dA3Ptp9Vsg2
Mm+qD+gDWSbu4Xuf4xpOsSE+QsqGhWNs4l5/C4FLup875cAyW6apg8j7NZYZHbSA
j4zsRPfDa9dLj1ehCCsV6/yeXuEyDAU5u8Xrf4sQq4jv/YZnelFb1eXdUWh9Y8Wn
MDQstSrJQO+oflYJL8zZG2+Gh/+0PoJXYk3QI9oYU2mxFnEfseJ37popgagc4sj5
R3SkTMVfHNmAVePE+kOsoue6rjd+CgYBaiZqmUMoYCRhHowE5hu+U0jlpaFBgIQO
WINSx2YI+Nvj7Yb6g8oKL8QIkvkKI4bv87w2U1FPihsmi4nuumSME4l+p64CZ9a9
JdpYO4QgI/LTv/qHLX7ZDyrRK78GxLvBnhKQ9PddumtjOtLnjWRSYRfdDRkgVfkR
XLAO3WRURC9rR+bYkafhCbZQDubDvuA9pS724wKtMFAxNpIGk/TAQOCphQQWxv9f
s/J8H6jabLa1JRophcruD0SHLPmfLPdMOJQXrfMM87GAKB2J2q+FcyPcKoMYVblF
qBn8keeomfxSyvsFZ1gJnle7Xh3rOeNC2vrR7YG5t7TuYo7mnZRMLBcDq2SLjOIQ
OsNDiYTstHYLV5VtxEf6BKF5NHzyNZW5Bmn4Co2jzmeCMnNvhFS3lkgZ8v868mK/
Dr505BFcXUxGQLCaobfEwyWTH4ayuc//Y51OCmx7I2eiyLiShZ1V+EiJMc3WcEZD
/e1sQLjAcQ7SCQpOrEOgf1H2qvI2VhEVOHWefDfoq8XkZO+ij9XuCZ8ChS7nq0TK
6g+EVq+KDcsZq1OYzqp5VuOnRp9g3lijs3lGcl5rzRryF6nXXLlscOY+Vx/oNTaI
NK/U8oXdYI4OS/PM4zyjMoPmpZiGtXkHF0DdiqJswgFiVyWtEu+af9I7UgYTBO9E
EyC2pwzOBYVHkmq5AObk5S3J7H202bu3Zi7U3YrBdhl7ET0XfcnddDRh29343kQc
GcfIMb/5V9MFagcZPdWC/Ik4Hu4DOWm2HhOGvusigEulRC288S2jh1vLMcsCY4Q7
9/FTSQ/6xoVWukWwat0dezne2LRW+YSQvT/2yRgYcvOqGONGU0VdO2bWhXXvmLjn
GeKhS3HqvI9deM76Dn6UENyN3V6UOgRRl4qB81PyJvcjc2xsAKf5/X7mqpTVQ3d8
EXZ2E4uu2eYbGG6XUkcpwcRUqjcVhoSOIvcMsxc0MFKSOAvlh5OAh3GHuErA81rS
f/vre02SZaHZqgq064Y5kWu9z4FoACqBpfOqxDxu5RHwdKcNCZGKiB2X/UdcF8Nh
TxPs9VtN4K6tMSvaKYcVZbFK4ViODG7zcqUwmmXiPGT3E3JCQI5cOMsrfyH2y6nb
k8dtekwC6l9coomEKdMuCY96ouBF2orRIZhWT45BpUP0C0/cifwRUIygcLAVQFsV
gUMRiOovAAB/uVLbTWUKUufjngYjmp9VZl0Gpbz+GUQf/X/fvFcB/nF9QaPyCxDV
ii9s2F/i7cXkrK/6XMsv5VJDWoyilexHaiyjOKVeRhl2mC32WZmAAHjqbnnSSpgz
IytJJYztXSLZzeN+oG+vmrisXr2g382YR5RGkBGwi8R4XVuZh+NnzYla9OmxtQ89
j4WYWWm/USIDnbQT5uMLGorodpSXD0/WzkKdiMA6q9f52FUELM1727S3jdu3d4qO
eDuiSM+/2H7jfDLoHpwZ1XK9jU/2qfTGEX3g4TfGq+ys1sU3wK997/a8ZzQ8EmI1
YYH1fh85TBnVGGneIejSjuYBn+MVGSegYPoFFrhFX3yss0YByNKnuPgn3Sx5Tz3M
2XiakYZYf7MlTyDvSWDqDB0uQzGjBMOqS2sULAtLt97nn3xaHdPnJ41RhK/CcQW5
ciEED4gOM8BjOTXs5p6A0jNkOaRFBCvPsI7Ff6qRQ0AjUlb9iF8WxRzWXNiqFXL5
GIcQUxrIyBzRN+LwmUVcIZq8YmmctdlJofsCjFsyV2+kjDZwc6cd4tfB7xJ/A9hS
kU1fHtBBM4ry2DepU7Rfs9gKN8MA1SUffY7iJ/kzDz6PI6dnMUn5ASTIoZBc3AwA
SKbmsguHqGinS/ioLQw9clmD9K4ELRAwyXdmDguacoo7Z5b5/32IdMfeDG9pkron
v4aOiqa24djlZtDQtdKQmVYMJKzsT1Kbaf2LIOTimqu31ZuzVgzQwSGU5qZydRY0
vk1J7QKi7JrVOROGro0rUXeE0R5FLg3qiEv2ZZvdJUN/tvSR7FYyMn3YaFsuyiLZ
Di5S0WNzdG3zi7yN5JZ0/7eGW2UzD1euHyt/PB8w8kr51H6Xa3hYwJ2+3G2YPGFQ
7Uham+NttQgpGRwmxNEyw/w2BrXqPV50b/GEFlsU+1En9n9mhLF10p6sqTReLrbT
TSubH+3dPwSSzpNEUkzIucTXrNQxUzr7tWF8ifuHvkVtqsp8ogU00wxckKBkaU/5
z29C+Sc14S71xzvr1EkeG3kXiAzQPOz8iVOJwe/3k0IPDXkizD0MR1EJ3aYSGVw9
PyMD7++PSHd2ejlc41xVv1ayHhgr+q3B6m7QrZxxbKuLgaLBM6zmOyl74Bo6ahlb
INzfI1ZEJIWB/8f9yeFtQlMzCH66+c0kVe3BmJR+OQRB9tVlxFSwEClnVs54dUmy
fzituMLgsdSJB1226mL1/Nvq/JbTvv4h2mN0b6Gere3sFuM0aSgeotN+1LRk3/iG
IWVkIaZlw0x08sjoTU4pXFp2eO4ydZhHVLv2Qqm+MAqEQt8hFmqwRI1JyjStMxB0
fCbpyQiN+y9L5zkwPLuiJQ105K6a+tNhcTr7g1iXz17wDwuamuoPypgJfPeOHfpt
PVUha/NFTXVhm32ApKJfECUvkefdxMVQpLNIdObpdpPj6atbrRhEOBQtR3/isO3p
gbEAoPk5rBbfC2QmBKaZCm9PUh1TKEKa4dFQrc0xWkYqBeet2/On+fHPMjjFB1sp
KNMcF08e4/I37cNJXoiZH+57ZOVKlY/8YNF2JQUG6+YMc43FqAFuMBfmGYMJj8/B
y65FuX3I//617LQEP0QGenW5q1WEEmQ+whoGBnhbO3SguE9FKnFzdinu890C8VZJ
XmZRtLl7wgb8K95jkKdIf71W5EONSWOjkrZAf9JfUH44tWdYLhACIVCLoct7BooA
yHReyDLtSqS0s3wfIT+NqkDCHH2ut1/bS4FEkyCAhyje420umBF52P5HO49/nfTu
RdGVX7psCY8TOZfYCbdUVSdclpdAWzxgT3iLOA5zfKqv9c0lWaaCfhYy6/2bM2aJ
wjbhmfD3zsd0K/OxIQjwXVXy6aYZg01aVtEJ8cGywCKD44Q3kfDOpF0FgEdVPc5N
o6oK6OO4PqFbzDPTwr+fZWj+HZd6cjBaeTZGaE6fED6ny4UOM9/gILB+9o7jshya
AH+MFBL3sC4YpR7blDG1e8edrfSr+0sbFmgMrj8hJgBQVCa2688bdKgD3NjN34pK
4DIuTyJhNQ9GoixEIlN/WdE6B01UP1OkXbZIL8xsLKD7t/4utTulNylVJVp6H4LE
8pi6ZJ5uelBRmdC1kOjxFogl4d9CJ4sZLJbt90IIeaufBS255ehhLk7BDRZweUYg
mgPrKifXUXH7D0CZkvTxs2WMx8vpv0n7EfXnQVuBTVuyr4MsMCDg88QsjjSWYbUt
3Yoth+EywqBqgj6ILlQsTqvvn5ySW0tRClZT/tNDCKoAcG+5P1/nW4vpQ+Y68B12
w/6Cre11DmEItqSMDRtllmaBwRBOvzQMPhauli/yHaCcNxM+TI4fyXQcEfWTYR15
MHEf6yLJe1IMGaLtT6XLLlIzVxE7/I1vDN5I07IyDe9+tREiH59zX9YZ/4Z8qIq3
gxNoHYykBuRKsVWLrRXelXKOgEmITvSnYc9TMMf9iTwux8w7wmp+FR/uH5jQcx1N
ZWsLFElhmlgBKgHPax1xjT3x0b9wdfxb8S5aHJCTE/rg1625cJpiGgbUsU1AL764
xUPbhDteByxUV4w7IV4bwicVKFPIfTU/GOjD7nXYsUFY9PhCtjpvxq4HsBuZirL8
/iSlsRtQkGF+c6tqrZWmRD+Wz9lWG9XTbujYGCR+R+xpNEo26xFUUbt9SJ1kWqX5
7cO7iVL70TVSNqxJvWyKS3/fjsNV78MBdcIS1nSCziGSyeCp4/zRZW/hTokTFL8u
k2x0ncIHHJXzqJPhNPjuBBrdX9MG/QAKa3TlEMsBobgK3wr9UogC3YEMra53nZHC
/mUttdEpVwhefFoli9G78SVUlgYaDYwhWv6oFRestRqDNbpsZPj+kmeImrNTSDLV
R7KPdWQKx5EsCQ/YFzEMTGC41K2KMTc7/DLjajQ+lgU1YduuhCfSiz3YZsAtreZ5
+bz8yTpLqwiNFOkFjbPvdMfx4CZCshYX0ivsIf8QbQkk6R1eLO8aX0TWDpmAYEyX
ZoLYn8qXcfGmHZniYEn3qODpUnr3g4Gjn3y5Vf5ezgcejrrbgItiaRHJ9hVPlmka
6RZ0D8Xhpxvq7SEKT8qoMEV3scF1ArJSNKRhhhaTlSMdx/QD7FefxU+RPrZSibvd
IGoG3oMFXF81JOBvtOdUUWdSE9EdMs2fKxQLkzTIqy8Qy5FmgGurbnNigK/U5lsa
j+qHkflUSDzH8xPPRilF1nemfqWLhqw3uCJOn339r2Ss4ttGa8o9W20ZUuUGJyWG
5ogBBgodNDX9qhCxziMwvVMGZ6CFoiudrozJsuPxvoeOdeyZk5cMlwlKPwl0JniL
o/mp5TNUtiedMa3L5dKhBXFnFuZoOWjCzzqatDQb7Rl0md4w+5HhF5Ga7pOTDdRw
5I7O1o2UpU6wYZMgMvCGHQ4BEhnCPpImYZ71h5DhvvBqJK4iW0IkbxGTvGZEpRKY
2lH1oXaFrbyMeLd4gfsCSG9738PmiDEeKllb/ptSkvQKZBVz2MNSy7sTks4eh4Lu
fR8DFh6F8nxrUXREqp+Qm0QZ/t6znZLcdscQfPSeaPOTd0csYaNR9LlHlpC1M1h0
Y5gOFNiOv110/h0GlxGKJHxJYx0Yl3nrIytYJ9TI6bdOx95JpAG/ONVPo8I+pyxj
srsIe3VtFvEoCYQAByMFqAeJ9219u/zieDI9Zy+3RrsGxUv/Zrl91DyMeKrXI4dN
r1OgnlBdVhndoN68S2g0od2P87+51HdyxdqX0eOd4FklHbUS+XAAPPwLbrPnuFl6
jxtVMII+nCfeaWgYLW6MP+3JCWx4nBvqfPctTBgqvoKFGYUMKIbXs9NTQgL4mQiZ
Eyl18X7JoTOxe95xdHgi02CuOGK5KSteERpQIPrawy5oIHYfXw/LPO4aYCoU+SMV
yFL2yqhLnYR11xKM3W+J5eQTYopqtGtVaAmr+FcSbbf8WqPzPQ1070ONK/z//TRX
NGh1xebKo/x/NlTkP6UflYmD0jfx7DnZlM4J+24iP0up7GXEHWWwZdw1SZ0W2lVV
HlGvw/RajjTBwOwYP1qCpddxm12+S+5XkW6OYCM9tH/NRG5dmeZavp2E+Idu0YQU
3pqDnTJdtfHyzUtpcSGup6Dl14WOP5KgEezuczZU6Urc08R072ihBR/qAQC1ltcg
3B0rxsTCDpJtdIZIzhUOfJA7Vn9ndBu95zpRioC4ezt0CH8FsPybzB2OoisW9wyr
5JC8cRiHVaJ5Di++iBtdY0qs8aRe5Vc4lswqveH6BG2CSN6SuN1SMtrztSZMGDMa
Mh+aM70lNfq0RDlbAbxmjHUMgg7vXg7qA3w9WmAEx5gkRxffVi2C0tq+l7GzCiAW
Ygoj5xgsoLl8rxwYodyD0h+9LPraJ3SSP8bZLlME1+/pTY+sQ1e8q/pDSxtYSUzw
EYE8BA1GFdgP6hVSoJNaSF7t9cUcIRYjg3e8fDqJJjUZzhDm8jDVO3zPbkbV0nHs
dF9nNu7aMUmrkyiDBL1wwlI97MdYWPB61fqvgTWeZR+qOET1SdomJB4fzIUnpwym
OUk4CIZ7YepZQ1sn/IV2+vq0LhWB2t6oPsYfc1W5gAzFOUQ20vn9EtIXPCL3WYeF
NwL/N36S3SfqSFKI3jXtl9kTpeU0NMaiUzSKa0R8G8CfV0g/DVf+SDnuoBYn1+uM
hVAIc4SPU/7+/e1gg05+l/5682pDEh5+IIUn2GKGMkHYYZUZeLvSL2Neu/1QmZwp
ConpVypCJ87AmKZX12/dZWGqUnOOC3Drg2r2BPYNxWzuWd1lAHZxrf8ea7Yg4ST7
DO90RFGQ5Exw0Kxg9FTtn3qilpMjHFN9ytm06Uxfwe5ojRtnxKNZ1jkyB2RYSA2p
t7HqszUhVDTMZOdjuk/NsNY/6HCFkM/r4pidwu3xkY9NxxztLpHRXQkEF2XJWhHI
ScxDcq5FgHbvaaMv7uaeA5ZkC0mvlzOwkla2r81xZ1EcYXOfi8NKfOkI+8ahYYFO
q0flKjjgzICvUUKUOnuPgWCZ0scITvFj5jX95gLtS2HI7huu/Zz9LBft2qzwua+v
f8WZfmMLLtxjg7BjmLurI6J2+42c9oGJbW8CcbMOySxPCaLx1kApbeA8raUxMLTQ
VmR1q9rnK94t0sm3Ma/RTUvcdSo6sMzO1WB9q+nnwDgUtkZaMqpK3FGC+WmtDl+g
fM+Um19Y5J3D/YnyuVwvH5OVGBeZTCxg6316UnR6USk1d5Zj6sNTAYjHGVWTQfao
7JEKScozA4gaoBnAYgH4NnESEf7iQiblAJF2sl/cmtk6SeUVJSopls77FdSsuBEK
Xxd83jOEYZb0F+TQlPyox+7nmFsiPbwdxgvLAc0BzQd8ANAlwWTXddfm5QvQ2W4B
T0e4wWIVY5c1hc8ci7gwP494qg2Uj2zN92vQmg1hZ/hyfpepApSepmIPZ6kAeSUN
enbv7ZaPdGJncLt0KuuEXGHbfpoEapC13orUToeZiZcTnS5O1ha7STpab39GQGl1
AokkHkAoNyaqfsxoJqBylezXgAH5Y5BhgN1IjkPdK8xWYf5CavFNX5afsgP/WU01
yDy/a8ctDK0reDeHeDNdblm6J/YXwUO7+sY/4gHImfP4UxCkKBxg08S40Gca9bIn
KICIsvKxToMcKiVnyNf4QcsOeDQK5wmW8M2yPdkVdS2eFZ+GeQA8VBDd+mGj2lAJ
zNuGGdS7OYE7PrPI19Oc/j7yGKzkio7F3+qYmlDenS6b0Ir60iOVacA1dqY7SZph
GPuI2Qi8frM6FMhOI6xZ1UKfGnjscQTIxrdP+lzri2YCrrSUcKZbLBXjFh3YVyjk
qvAeD4zoAWebEcy5Lpwb57TUEps5VFRudojDRJzq3O6OxUorW9JOx4pqZS8CVqTZ
ZnKdmStq533d9D7nKuODJ/1ehe6ZjFWMptBjdOYXCYSLpp7tXReJRgbXG8mIuRyq
jiPM+CaZxZSC9hhnz0PpPIK+vNOU0Ek4wLX5EVV4WtvmkKwDGwtehJUtrYkkYN9f
HCKCwkjiO3cL+2uTAy6x7VpxoCaALqTnt0yhys5Ny2QYGRs4ASectJ3H/3ncGZi0
OktI0JTEgj2bXGxKtdnhojeC3pxm8kd//NMVLI3luXVckNGckbXZzzSB5duBXono
ra3XhhsIr5vDJH9lNCPkIcZwJPp32HUB9TFyqqjH4jsEzR1mKBqFQnTmXZpgoerv
fQkkLcvf2OrKLpUcQaidhNToXJoeZ2BEzhG4qja53u4NqaMv3Pos0PyiMxtNUnTf
4qR3/Lv5Kq2aNo5KYxvD0W1fW63f8ifjX4SMGZVXNlEN6gzmp4FhUcPkmar9L2Nl
1QFLml+T46T7Pq/hwCrqLoa5BjVPqHu3H6JtgazvNYJX388XsCVZP8PL9ZSdbHB0
iwBBB/MLVEQBSIkEsB3qzrpPpuPII4ihmXRVDrFOtxg1GG0iL6JrEhVByyavu6Hl
J4mXL+btHVQe/R7TgOmmDQL1lkP3YE1eqib73AlfWmQuoJEqnxzGCPbaBKOFCGI3
CEJQuothVXbZ8EBBouyyt8xeCOZsYC6MNx6J1hT7DPfFC0gws5WvlE4geLEiBxYC
uIThLVlglYPXUZEUljiQat1j2RfLrOj2fPogSb8Pvu+z65GW8ilrMCAhE+9ILtU7
gEwlfC9ze/Flk/TT5q/qEz9ZT7tG0pM5/kSPjx644/NxFgD0frD5umnKKtjMz4PU
KodrxHTqqP0IRVL9dqhkoDZ+5aemqT7BUGCOG+Vz6DCE7Ue+MxHk99PiT/vMRzxX
OlEWB7SgZ6lQt/0gkvD147nrcrX5Wx3xVVH9EMndhkm7hwrA3ZQ8C2DJtYlg7ViX
3CC3cr92xA2+nVWiI/Yjo4j/oIMtnx+a5DQ7MNao5u4FTscNXBPcNGeAV4xGEGSI
y6NQJpxnwvqwJzkpyB4kgSp4gQWVE8k0XXvJEt634xdM87zFrNFIbvcaPUGXqLpk
w3nEc78s/07dvuOH8oh66JtYmDdbJPYbEYGmbAHIeG1EjTapbv8ZjMkb61FF2sOE
3pB8nlJWXHc9WXeH9UgVUGji3ofJD333PGWtMhnBhgp4LI7kCK5xeFrcG9uoQK7U
8JqACcvhI1UqaYhF4R+QlQ0AzMygWZT43BeB0+KBc8sp8sPf7gctFEAnnBSDXR5T
0U1VzOXd2M12RmiArv6yoBKh2cGFLvgs38fQsroofcNgi5e39h/r0WqiLVOYfWuR
141YFxGjEl1+mzOUMXm09y9K8HghcKW01XB3kTPZbyRFlM7/s62OHU1zNH+rLYDB
WWi/ZPLKLPV/OqfGoIUd9n3hjCG0i3KfGS8b+f51WfQZKw5NDlh0EdjZNAwLpgpZ
pBGVF6Clbp20qHagRraBbVc4ZNRmFLv/p6styvumzJygoMaO/6qQhSR17eUtQDdJ
mAppyfftpsC1qVhtXNm4wwiBzQocQXAlh1TK12+GGLA6sfN2FwInNiJoEckTdKgB
DWK5cSv3Bt2ONj+GcaL0PakJuf4cEc5mhp+PrBwNUu3L4cAzoWIo6XPVQC8ykBxv
N6DE2Buf+zqG7oc2bI6ouNUDDAA9tddF/SKaRKrotmfScGco8BuevQ0SYVKJHpvR
kAVVRF9g7+azmOdCJKDqgcupfHjAN/jaJkOyxOmV1uxVEPiuC/K9HwXfP1Vuktf4
UlF4mq8qovwpJ/BJdWtC38OP+Lq0jmITCKmxT9kdtd8Ox4X5KWxZhMCzqdxN46Tz
Y2N3phpZ7DRHSSTMYzQ6DNJwbgFJbsGc8h1xLib2VhNAtY12bDcH+OIID2yzSJnE
M6pLYMccRZZIPYHTyyMztgpIS+2F7o4HDuh8S4r4JcwuqcgCQxZmhlSm93TKCYBx
HoX4W80w69kM9NwpT35sEx2Gj0xoBEjTf0zB/oMfJpGW6XmhebJtORlXhkE88GU8
RuXGBpZWJGGWhexBqAUowubWgniTOS/hwMrzJD+BFPuGXJJPPDsfBF7qGLXY61fL
02ZjUP+2zzTSb4BFsMpgbjcM5ny9GP5UE+3+cG3nDvC9i54RH9BDJFIAdqQhYOnn
WdUM/h2VPreL9WXSHQUgfoANOLmE4DPAxhJbM1n1ua6qUzyx70wMFhhtJB4vccJb
ZJr5od5yVBsrT3JwyJOY/GBLdyuYvKwOOnMbbDdNF84/1xs/M6r1OW3XPRrXV2EF
nNS5j2XIKHj2qnj8uy6odG/CfSm3n3kPJUcdLMZoIa9YDm8qDd3LGSr3vRXaQLS6
E7qK6dNvM8NM3EMcDl0TZlIulg6eViu2A6k7mbZpIQFTs+HU5LBvR7GY61QKmqD8
mQdZ23qhmFoftJLCviM7FF2RHp1CP06iB0p8ZUV6dXe1SBsbM+ZjKLqQDXQWadRE
QDdY6b5vJePRbR1fMCNkYgEjBTZbyIYwGic2MgVSXlsE6f9XK+Yfb4K1NeGK/G7S
IgY/giKz+U5+m58HUtoXAPr66MEV5cS5PZTC3DooAwngpW1a5asm8V8HOTKqNJus
mH7ehC98nyDZCx8+8IKpi4zoL9jC7160Ki5LPNFSzFCfQQ5hoJhrSiGM5zHO7zUf
L9i8+2vx6XqzTizGNdsUfEjqsgdEiuNhn6DARbg3OpDKBGWwY2fzw12UFhevnaGB
tCbSLWCzscm6MES5b9bVAls0mvJWIpZE5Oy7ob4uc33AqEKPkwLYmrAg/g0JE7YS
QakHh83bAMYsd7ClKk3JeTAfA+85siw+ffwM0kO4xqEgLPDBT9qzLLi99tFjqAha
uBLARzSYa8hlFfZ58CpD2wg0gEC04MUrGIFztcWYvbUj4LcjbJrucpsen9GAe5DF
NSIH7RKpdO6wtldCaAGM0gZO73QKYUsQKZyUYrHCYiVBwMo97u64JC3LzV/e8/K+
FP163zWGplG0yp0cdcZBuvtfoF8J1S+vL02yMroiq5UMiw9YeTArEUUTVkHwNYwD
ZLJ2oGVKPbTPAMZpxmAcU/qUf16jv2dN1k5euoJY2fqc1oqJ3RAmi4mZvrxA2Dyt
cmuK1FuBFP/lVTFEZbpmW4lTDzgyrx08KkVwPt+5vZOsX5WoA08K2EvmANuaNu5a
BCHtZ0EjWPEZSNnuMW9w8gKdMpF8SzVejlZ9a4Xa+2AIBhAjfF410MxwOxiDgySx
0DV/TiTuEYesoDNGVKsh/HWO/bOjPxLSDYOCMzGYchTjbKgvDeJc6JLDUKbT+UIS
nuuyCHSP1lHdy74hP+q5YYGkNOZoxM2GkZ+OYcMjIQ/1invRjbLdlUw2J80npoZk
pJFbS0rjkJOqC3yVgwel4yAXClrG8/irkiL4BiUoV6tZr2sgmkKzezsJ5gMaourp
RNtxHRpfPgibbqbQEthQM2RnjWrMkQpisJQFa0JLoL8+Edb6MMz5h6P1ylzGY0BL
/loW/RAfZxGT5tgFPMfU/vDowKLl9DJ3f+hvONI+1lx8xDIXymY9jDvvIJeo6lvX
R5Ci+QBc6o8X3TmPp/wGVa+bbZIcgS48sFfTPuA5UajzpYLBCOkecm/hNjoZUbG7
DJ8JYWvjjEtOtfKcrDrWKBntwlIPnfBIxqtk7HLP5ymYh10YFRjtpROMz1hVCmVu
amaWIAmlANECoEh8Q3oreAFM/9Y1m0I8OZeCIWU0uHIM/mlt8+vRkLnE/UkOmd7M
Ii5fHpCD7ES94UMmHiyAVjR/ePtdLD4fEoxojkk88bsnUlqBhYTr3uOPb8HQW8PA
JBdz0lgiqptqGFX+U13POlPvRK79ae7SFNGR7tUa40sAHJKiJ3iG70UJoO66dAv4
9YV+JDALH7zcWt6AYYYpaes0OEzwSDqvtl2Q8vddfvzpq3AI6LulhCp/kOt1iPhf
atOf9aO5aev1QQ1QFNPtqQeHkUxKqBmSMmRWbSxl9XUCV15x6ldmDQcCkji2zdyy
cuim+tXVGfQ+lHNjNmZAPNw1SDjbuyp/sOjkh1cjbmrEC2dGIc9drm3p4GFxOOFZ
5Q51cpwvL9WHIFuh7AT8ikHlk2oteu1Q1BKJT6L8ePQbgPRqe1JtYovXkY+ik9rf
a+XQ512Pfi7zFg0IyixeL74rugl1wgg801osExrfmmLsgeWXBhEJdF/HeGPOKabC
HsbOzswXjde+GvoiiMc8y7ZM+cu/oPJDnhnh+ay7RkqYUfXlvoXWtMpSWHgFbeXm
kS31aK8vosDN7J3ElcdGVtZtj9MB8dco3SoqcSBGEz5hGr+6T7YYzLQNXwhXxj/W
h9wVGdh6bxpwxDXmt+96rhxJwZyW0ypwDBDJwS9+/Vi36BT1fTYIeJM/t7Ni9yOd
GVp/Y+VyiI2Q20KNGjEjZdHyfz94wGjdy5QF7LBaW5VcqhxwWk8vgslAnNOcfjSa
iFeyKhQJakeIW6roJkEDC1APJYdBREP+JHc1JNrHTgsvvbHEqGVzMcGSf2F6jA/c
rgwRw/XK65fizfnYzFHFtJm1FWRs91pQj8Um18UFZmq/uWwETKm4TGlB9lbV7aKd
4vaqbgGLzeMfmYpYVIQ70hsGuX+yWvyP2vM/DhJ5Y53Eazq+veocfWOG2v6NATtW
EUoq8O6YQie5HUIQxc+27ioz1PoWb3ERyBwicnJoSaUJl/6LQoeToSg9DDwmiYx1
a+8/UpsXWnvf4MfQvQxekniKwLTjjjzCyxMeZdHn7I2QMcH1U5NLBQuby+SidwsY
qPPhDf/JRfND94/XAq1ZvQSnFhVTeWjtGY0KBa/DlLY/4Xu+hIydWUpWivf+g9En
lAKWAV7i20NjVhSkI0rbLT6YaEopRVdaRf/QROd6bkGZupCG28BysYQdFJilxTOr
RhYERg+4UfdH7tIxMeclWwy/1FRxppJQ+r5VwkFhUdGQ4f+E/4PRaEGQJw/2aH9+
Z6ibKqZhoRMqV2VuA/4XkbbRf1zVPgMd4uJzuNJBIThOScZCPc2cbOtrgAaaRa1u
k+n+zkQeLljFopBwkk3K0mKaH6XkhvKE7cWwQww+Ai50+iAuHtCIlCkxodS7DBDO
wJ/x8d8Bcic+N+t2n7okdkEup+CvaZ5pJ/PEU7sX+9o5Lb1KuehmDZb5/KGN40Dh
hWznFY1xKdTzgH0nzPwwq9SpCdwdgBrmioms2wJoUS+FFrtcmR/0zREmljqmsukn
UelmxS8ZqXYI5wa9pgNffUpRALYm7/OVqEcanFUSD6gRwNJdTi8Q5U+0hOnhSok9
uYGCuKiohkvAjJe3ygbMVvnAegbOcShSJlkUk5nJhjocpBwlobj0fWyEYYLqpqj4
x1E2+/60hGOKD9IKaz2ybA3w/xlS6OY3DW/zYm2BBzH4FxMJKPWBq9qluFOMlPAL
iNPl46tzLNjWssGVCqQ9eTwn1XvY8ZDifAqx0PLkXe1g9C6DvLDgCxuMbsXFQJxI
CMNgqZynbEjW4O0cE7OXnnJAh1sdZH6v3kxYJNAH/99Y9PkchTskFkdyF5i6mId5
XsI4oasSgWHQUCmBBThpaqTPY/zYJHdGfjWS+Xat1T2vRV5Eu0BOPPWVOaezT8hv
ck+nTjBhmC3dKIcRQn9r5984OfhiJNltWm0TUf3b/MhSyL+VLdzj94XD0+9J5H8l
qIOksfunhtu/DkEwvdS1AsFDmfcg3ne5S3vPbyMu1Yu/n0Xu3NxpiB61VXds3L8A
6rjzLXGbhStvb6nOlfOTtYZH7qm8AzxT04AG7wMJAN5VBkrNiprvwu1J8ptrlz63
zzwRY5VqjgLQ/mKlHfVudeyi6Gh8kk/yy2G5MRVBNN5MDNgoVIPkAWEPnQQkyeHn
ZW5wb4CBkNetHNarBKT9oU1zhApxLlAV8BrLzZd8pVZdFvrcU4YbNJR3aYS57abt
hvUgNifEhayxJZijmuxZ/HMGZsJuHmduoP3CviYPIMeAOK5/GueuA0jhABnJLCHS
0beT/id5qi7DVuVjYOx6dMZ03/dJmt766bfd9chepiMCf5R4ygY47hyPcpEFpPF9
R4sD213inqwv5KTeHk24d9xfI8TTz3ftry9XHtgoAvgP7u0LzMrTe2/GB7JsHiJT
EIA3jedSw6dDxPNOXX/ZuzhwzizHZdbTAVF3RZqD7m1S3bg7PGjJ4puZcL1fy0du
nqSdcSobcAYRxa/MIBYrFNxy7XUVxF4mbeu1B8SmTa38cotsK28cq6zud+GeT+Gq
qTX72bQb3SE8BidrZO+sxTlJSgtcXOzgU8QbSZh4r1Ten4viM7T+UoL8kRTxTQfJ
bpOLz4zf1E8HA0rmyv71/3telY8oJPLKBxWbAoT4O9xV7DmIsUD4kuTU1bwAgDGt
5t3ZnJHdFA5wAGjZr64Haiu+46wzKiMiWhGu7aNhBPauQ8cWyb5KowarNMVyv9PL
j7MjlP5C4dJZB36w+xOn2wei3RZS6FEIbEt+GQbWK91iU66ltaR19hpyY/2dE8Wb
EIO8JAxhPYwImisMFnALML59drypBfajiD9PMA/HcJ1gTok1JC8S0Qh7gQBtCPcC
zjGkpFMQ2EB9SBCzZRIIEs1GRdcDpl5l1RAznftiwYZOIqxbiy+t9fA/ZrCmyeIO
VEFGBWZUHHF2wwy8pJjrH9/q6hybhLlylzk5w9RSajqq82ccArtGCg/v6e5dOqFR
oGsuTDMtrXF6JfS6a+ug+HTevmu0PHUaHnbbTl4jIMgfqgB4aEoqHilf4kBDS8t8
wuNQvIeWNjZzTBjcZUBSDglKswOyO1zBNKJkLvudx3Qp3NimMW/cl1XmLXpvMkwJ
NhZMgMONppzgvSLZiBwLel00w3kqHFP0oelyM3qPg/l4gRDY6jHg1xVz/zS3qUbT
eoAhN2Yci4rPwqa/JgqKdj6LSBLtTEnYYydqnKGK7kQ7LCFNDbVtPLx6+bJZcGr2
JdFpI6P0NrZfCFAqsNwB6BvdGAqi9FmBzEcULqPmPyPpagd4eUVlzC0i0Z0cpxPu
1Wgd6D/BQ4QA7/MhQYO7fBuSp2/xSQVVf+Ua/NVVVKXOrjHiXOSEDegzIv0QWb2W
kenOBv9NI2iv11RQaWVMitKEG5UIjlDuw5FJorr3GYp2hYA2ZGKybSwsSHmYAWhM
0NK/FHeDn/n5iUJSjgDiKZNTOXYJbfrtSTif//wmi+NW2Fippmd69kjN1HL3C8lN
/6tClg3HOZML9Sz7Ysip+7yoUHIZQAJVWnTYaASHWRlVa2MFjteyKdj3JPtOFflH
F4ODngzjd4nDZIeTs5WlMcPfC2DRAl1Z/IidYqnqSfTg+RpvQ2dU7OCLZPn/wd1t
PfqVlSF2KwxjsqdE2HANxbpmYGFwTiRGsbGqVhFx0cf+x6QXoAaKEErDUzPfp+KP
MXouq3hjhLJQmb/Auprx8xc2kDzKN134cKxpfdTAAQEvZ+bofeNlEMeU+zULQrcC
0SMfLlBhcUSVdw+35uTajS/tmzuYDV7DH2fColIKTiE670B9rrTOae3RnIHt9jX7
hFEJ8Mq+ZrhI43KIXgVvVeYoukHDYzbeRtQgbSVKxGHKOWxq+b9vDetQseJvzmHf
pGtMsqA7YhwDKP+/s0XYpcaG5+LMX6VkBnDogswPwKHN6Vk2sr2ryn9q1MJIeXzG
kmoSpQ3XUCEzB5YGVJWqOixN2OPcC616ti/9YpUAPt53Bn8X9wTT+OpPtP7kqdDY
Djhh0YvEewF2mjjK3kg3O8PeP4eJN+3P01l2woc+kyBYWNranIJi2celDlYY1Lla
bl4QOZ/gH2S3BCj0ZHAquOkjyLU9kcH77RthiO/mx+8ulzwqro2+M3YvUSKoER+B
kCC/8U4x1wL9FE4vgJ01l4qOBKsdzV/w7eo4uWLibotyJGQXR6OZ73LKKjBzC4IC
i2iJ3QrqQxuw3lRTsBOi9JA5g4B2btQka7idYUMwqRPPq14vl2OMtT69QfJhS+bx
sKGSW+UszfpY8gPqMJASMPcRQxr58updGhAltbLbDDHcSy16tlaXqyp/M924hCXP
ep6f4JFZmAcSmfpOsiGfmqOeT9tGwm0gsGX3PP/J2ZOEzmdiIxwr+iR4+t2uBKiE
wwg6BQqQdingJxtTOZfae6smxnSuPzWNN8Cr3fjG5XuIAbWJv4XImYB2H4MISxkx
XjNDk18h0lMFpARdpaubbyYDP3MsjzrR3ybA+GspJOyywUqXIyOpq8x0ms3TLCyK
t5u1c9XsHNmDdQ+UsuRztBM9CUfQMD0J7wJc8nfCssdAqm/4E1Lj7R/3p0B+qE0V
RhnBesVrjrZZ+H87/CrebO2GFweHkn2WOu18RZmPkZR0d3KbWaa/nIcq2dXxNN6X
jMStXKmwBnA6CARSkwmlVU75SdiMWiC+92fntgvxRic+17ZA8GtS3RfptFAq60f0
uIZS2KcNDHYH9H/mozltldLkX5gsnqDGpagf8XdFwIeoxIBEA+P3D9wV+Nxlun2l
wTzL/9NJSRDHuA3EXSAXiD5xD2aWfJalnEUnJUCK+5n7jsqKX41535gXG2bQL7UD
qcWg3XfEXIiLHNFdPtiWDEVk8ycFF4H9pChsjQAZf1jAR6bDgzeWVcijpm6JhF92
nYijI2U91onaqFGt+2TpRIlkCOApouAVoATdaIgD5C1EHycxvhyQz6xrP9QK4kDT
27DGCitfo1sum2sSEgk8q3E2GkJJ87Ip443kTF5JsJIGAGXnWPsuRiGjWVifpHDQ
FigDw3EiE8IAaH4F+8pLe1ZEIUPhBN2NFzWZX5RSBOKivRWJDdNBQaj9Q+wWQNEF
cC9HTzKv37m+os9KJs6lsg0L9DleLNJkIJ5v+AqESsmegkH3O7J6WEOXLe6fEtcC
hIKy27IUbEGKiM/sFx+HOVjfT+U1dJBbLVvKQAVj/kGCKbbiMkv9t1Etpcuf2hKu
Q95rreOR5T1d4MC+HuxushIoDDzPmgXudq13kb6rHC++LZxbVy1Q/ZGmbofzfluq
goVwtRTZrhQrQ6fR65tcTJb4f06kSjw2gJ//Dc/55uSUg56pTbrANTtV4BeeMVNE
Aceu+pkzOjQbsXYknU0dWq7r4wggj+IbXAVdiMH3puY+lcnHTZenAJ31X6ANNu1f
YULcWyCWxCttRD7VDde/o8OoU7essJbvtf2Kyl3ZLvO/qMLFq3h7cJVlywjd1d2+
EUazDKoy1jYRJ/lUXVZsu9lMBcOBGf4dBaaQ7uvSKP2uigNplxgGhhQH5TNFdgC2
ddVByNwC0zq6MQMboBYdChs5v0Nj47ck5rVzpVfyPIXoSe/0cjQKqfHxlNYlT8a0
s15U0sZ//8IWrm0ibZuveQy0QDt0fV3lXsztHpV7PmPBrBmNeoKtpeumuQr5Tr4/
+CeRTRRgvLkFlDdsNeF3ftGSV8DVgcB6WjFk1n3nqfZtvxz8zTQWSgPUROmG5/bJ
hGyFo4WH86DB9agcRmbdz/iyboILAr/h2r+Wvf7VvRPL5XQpEE3eoJ/jb5NOuhUu
jgAnm2Trg0/d5EReV3qogae1Mh+cSShK81QG7LAuJsgfHv8a4VINCskHl9zvq+9D
xvLLLpgu+7yASCUJeZmn0dsDppax1Wcq0Kw5y3UvnrjpbdMf3tytnKGJO+TUcCla
I+n/MHRxwBFdW/t/mkN96WHJfQNTECNmAyakHBD2YkFPos1CWXHau7zOqY2L3k7U
YCuQXDWDbXCWK4LRUxIqCxT+LVRG7FAWXP2LhtD6zheLa+iS8UivLIRCwg0icZS7
azlLvoK6+8uhtQLAurgzA9G16MDe9MtEV+tXzQQxfsERqNg1PaCFiSHC8QeVBs2Y
+7ICw7V0hTuheNDSLX7MRUV0anaL145YmFOhyNUkb3Uf2AIyypjfd/OnYt+BRLmF
zmp93LyNQH5f4TWK/Qwias6nXTS3TVlCgMn981CgS4w91XLMmavWKqQNlYvA1IAn
wAPSHDGO1fOQV7Pi+kP/CLzQ2plz9kYhruaiQmKjDXq5i1/w5N+dLdgmGzPBlfI1
7ns8AEdG2nfv3rvggf7lOKlPbfiHiUykQZuYhrSyNpJXhgcm5xvprIiwHmI0EdxO
j8kHt+AdHByOqmBsQc7DQB1V6cjQrCuNRHQ2UuDlLxfvMQoC0ESJFhE6+xXCi0FR
TeYH9wF/S7vVVIXXo76OYvyhBMJwtoIQiZHY8/awsosvmddDPPMy+rcdNp+yuliC
Wnu/LWLTA8UvRPT1+agN4Zg/MPSeaLY1OHOOLqu8bXJ3oroKtYpbBLeEvobCSVzz
R0VjNcAbKicnqBxmwjmXUTYaAvudymJ0Q4Rh5OM1f/G9LPifpgzmOj/d2Qt9w9eN
pMSgwhxuf56Qga8V+6VB8I9fot0Iuz15xaWE2aelwHOVtPAsXjGHTc9buBWMv16t
0Ob7zB4CDUP0uvwX83q2c8rTav5mpL1O0anftvoEizP5RGPeamgnxOJxm3Ppb6N8
xFaehLM1C04d13URVEZbRZIF32eHxdbC4RCBJUTl6+2kyooca/VC25n1mxsbCc4V
jIVr41jGpze/pFw/WtXICe3SdlKpnm+vGekHszUaeqkUoJnS0OPJp7C3Y1u4ibXw
wPJntWJJ1xqZKyKxQu8PDwGry4c0bq35gng1N5wOS1BmFb8Z/skTQY0ea7ubpyWz
MUfRWfAuouxycY5eDsZLcRRNhoZNt4rndUpH30H+lS4hpFjM0NKjBzq66W7O85pP
6oBbBWTBfIDwdXZHrMTTF14ae4QlEsbWaPApbuI4xVM4wvIsAfQyAvc+wXWp+uYn
LYXUxGi99YwRxbPY6K7wzC1d6hBdtG9r6jCqfDA/KxLd9oblPDhUZM3s/u1bxh7O
RnQA/ZA+t1EaYzrv8I9MPEUbdFl/KMoccvlIbH4LyaaYxezLw209hmV6tHUEyb9j
VFPPwvQO44KUA3A5R1LCAhnSu1Z29gdCQ0tYE85sRL5il+E3FesZ+N62Ryi6RsOU
jBd0nslVu8E7abbYSfjPbTdVQHr1fePQeTAJ2jlhY8Rn4Ap68+e0Zo3rSM16qUdF
EWdGAxMAj9wz1wFFK0UZCMK71ut3/v4PXJwM+L7we3ThGHLyx8QmOifN1c6qnuTt
T0ro7PLNqUfBDwWkwNzhSipAanUhfTJjfpRoV2BIMvZtraepfHXF1oaqudMmaDP7
1Y0f8WjlnEl6SU4Ztq1wuooTcBMxNJgNaPUcO02mNpGx44oIEYYaF/mk3PHmK2sD
aYWjdNST36P5AxHCejgOkkPbL2odVsyaitQpJYBshmNtI43upV/2vGzx0RwqBZ59
Jgbu6XLr/NT2mRzkorfyIAIVngvd4exJR5W8+YiGn/InFJ5UJG1ldFmVMT5SO6Gb
CODV3pc35rY0rfa9TMv0LPjkSYX1X+7tThOcr/YvJmYi38i5iQFyRhuk7aAls57P
G3WUIMmCw0L8B5VvybQ5FmTYJfZA0qJ1Wiy82S2ES0Vr9wRpo5E6dHIooMnGH/0o
7MdTSH7klmp5YQb/H+5dkaboct13jOGH4mvY0uwQf2cGI28q4cjl6e5Lr0Od/NWf
EAsvS8QNnVVyb8eUbbZtGdjLVqTrgDjZRJsSiPk59l2b5zgxdSw4oWVU3/JUukpQ
DiqaqYhrOCYmsrj0/N9CBowRSzECZuX94WYM668jCxeOffy6ZNCxGic2bAfiC7Tm
aA2SQGKDxOucJ3E3htiNlcIuFXFKiBbAUTMsjiAZQqBMH7oM8pkXujurz8GJYSvt
SZ+5CsZdQzRVLElpnxDZxpSCCvyKF0Vz10G09uidrnz28j+Jb8qoVmQmkQIFKEA0
t1s1p6qZv1jDvHz5R/Y2dGsYbZUMkUeSOYgudO+EARc56JGUBmUOf7G9sPBMvHEU
JP/wXP0jREhFEOh1VFH88Jz4VNNlGZn3NWdSK2e42MH3RdBBK1ryv28GFbHdOD1A
oPXOEYK1rdT97/fJZXSTMPwe+WRpT1iTb5OESmDXToBPL9I3ZpMk1mjwMi1/IKgn
+RgsBJ3FzRQQeFRpmFmID4sdF4KnO/AIkg3tNlBx9MclKu/mxm3n69qligU0OAOK
iJkt05JooTXeakNpRh8arKU1Kk/poc4jnwWegzpfTeqNEGWJQUch+unREJZ52ARc
FzjYtS5zoYWh3Jfsagwpj+cPZCPThsSgbVPDDXyXAZRxoM7oJjAFrb4XoeuCeJ/q
mm/okzwn6/Wyh0g0pcCAGOXudFpqXzPcLcwRe5Jd88Y4pb9IrkGnxquFMtkTWzgG
1krMP6ZFTVQ0zJWrl/fmSe/I9wTW42uqVI7A76dX2i/2kl8DNVFxQgVLj8PmIDRR
CAaq44OcU/UoinuBD/139JAa0iw//pG9yCHjb6/zYArMLmwyFHfPYql7Q8Q7Y7YW
hDILcfDgYhtPbgZhkTGJDlP8nNM8kTd04/xAR8+yh4FRgwt7ztiUlkFowGk6ham+
hK/UzR7mwAYIX8KHyJ/oYjSgYoy4FQ6PMKmss9vuJ04tahohAPbCUJyukUZSIEHU
OPP9ebfky811OJWUwBm6io+kqXO2EAq4HZfx/6lnDofJW8mRens9BTHHH0ySTnXZ
HrWu3agGnu5b19ijGV4ehaSrat1B7Nvxy1qUeXSBHt9Lm6cbMBYByd4TBOXGhYaB
Bv39D7kRJpg20VT2QVLVBlzxZA/1d1u5XMTsqLVaNuwvMeoaoB9cRz1mtowkm7Nm
cUdNf3Zf5zGA7whKKMLVz3kn2uTD4izYUzjmv9VC5OQZpTojEshyNLh6qM0AjbsV
a7+txVkcgPmofmO/HtmC6sIGFGoJDLdUtolv4VjlbwOdBxO+M8l+ZBUufmCq0Dsn
lxLle61ldi1fm28lSRr/cZdm6GYbFTtf23hm5Xnoh8Y81zVOWTZ7ObrCGpPk2kB+
TTE7mHTjDBImC94+02fvrnCpA0t+Mv9lpiQM/+GAZvD3FyESwVCZa5GQ6+uiOIha
hfDIZ2B80ieRJmD0hkX10COrF/G0rgk+2hhy1qKnmMs5fRgQKDwmMAuE5GjKQqG9
A+cbc1JUbSPFIAPcqcgsEbFOgCg21OiFLpLCt5mLucdE8bkK7j8slWmoN+rkjq9l
l48xePMUi2HZXwDilViLZuHNCvviamtUIygHf0EPFMGUwgkLkFKCwMRI9QkYQ0eK
Jxb1qj8FJeDGxIRg+XtTTN68a+fJRLPsR0Y4EjQn/wLrjLPICY2JroE67MLkmcEi
Fs86v8ouGrN10OfoOsuHmeLKUZnVjk2nOf9nPIPVOed0OzU2lnKDGcQet9PCsJL8
yogaMOysz/NuOD5PELFXCWXVy8hSylP2kzLkOD5ZWSdud+DOfCBR0jPZxXeAy9jN
nOoJmprxmUgp2Byl9KrG0/VFGv8RQWTQRAIoTToU0dLxBATTFl/gyZmtQPcwNuas
zijHWWUO3e38duCnGXWP8bsDBiJ/t76VmgA82/bt87ePBeYWcQ2KU8d/Hp5HcjRK
/HbSQqtzpIPNrYQtIOLk6fyqcSPiwsY/tRTVPUZL7yenokQDGXruDIo9/TfSqOFc
NBkychNylxAqji9aCGcYmDnkTRdmPEb2kJasrHEDvU180QPNxNnSVZlsggFnnJtY
qxXqm6Ms1Iguc3b1X0MijtqcMT55SpQ/f53FanhMuazQULXS0amrIUc5C4mG7cha
7T+guxar8PILoj3NHoWezHpgzM0cx5Sk9V5mqlGZhYoSwzTiILa/XExZun6RaC0h
VsuBVHzq8Cn0BtdVQxdKGqzB2XOe+fafC6FXSrSuU+dTyZd8Tj8O4zJljiMfOp7D
m4EfsWUE6jUJDMZRMcJ16usfM7YhPa4bdvRVpTs5xV9EKDVJs85y9uUq2/nNCmDG
KvIseVX4hhmVxzxSpxDEk51wF9bMe2AiYAUuUQO5LKvK6D+STVqMKYok4TiUZ/Uz
bOVXmkybN+RqEYajHVC/yzmPmpCf0Cl7JfBjXtGb+ftUEbCbFuXusZhgAR8qw/od
ucuW3U1R1a+LOCSw+unoiCM6+6/ZKcy6XrFI+DQT8FhA8UHZJWoZDKXoBUnf0+3Z
5dGBdUVH4NUHGBpfQj3Pvon9W4Itd+5efqzIMm4P8KTJ8LI3q+mrizOEx7f/6McZ
CWDOGSvhmKeymLqh9p9LbqfZfXStkAR8FUFyl3SMVAzM9IC4wQmhO/3yh6hSFZXt
niNTguZKKLkiBnVxHRxtjze2EjUSnJs7x3DJPTWRvvaErvSHQYC/tMdTzbTPO4MN
7UzHYmbCv3JwSQxAABFHzWjk/9SlFOB4iNWTcuY4xjYzQx7F7j0eL43NYG/Ox9Fc
zfsqjDszvUJo8N9N1BUzfVlwLOG4SLSCFlqaZ7OOxbbnIdmfpZOHJdu9RHt6vrLF
rEAK305JNkbnLNwKag8RQFvL0oIOL3WPJiWxerjgwwXR5FwaRUfrnGnaq2A3SNuY
YnZn/IsCCpveAyQrtV2LYl6DtOq6nmpXPKeq+67q8O5UIpINt7j/lVduaAL7zFU1
bnhaB8XtaQoKHsg2DAENbC+WDSDZTFg8xztWI77ZXkw3TIMhw+usVaGaHhakKlnd
wXrIa8diXPavQ9Bk+mhIrQMCy8EU32Mfk/bCXR1remLxlKE3q/WapprRS/8rKsm+
540Q6ELL1xFkSiwQkpOcGwHi8rHgGxwUUxPbG13vSz0sTHjreI2xogNeQoVJ+usg
hFYQoSnXpMcbUNFLsppkR+/fiyupYw3eUk38WyB6f4GWa1uoY3c2fMzZHdjfIDd2
S71LX/fwl1yrrpeyWpL7vtxALIJF3c3b832fv7V5FpBBCcm/Z7rfu4tGJ8Z3tEOJ
Io99VRD7m7iOrs101+cgcLGzrb2fROxKUA/r2rNBFJIIhGwfmNWiexAwlgr+lHtP
RHXmvG65L1LJGrFNKhMidqD2BRq8IRzqtI/BBORuaN78eaPw9faAFB2eXQPXLW4+
xsz//3xQQ808XaEBW9r5EfWUpt5uqGEO8QhRhWYUfhyd8bAUz49j8FMko0bZjLlT
Cz/qdA86wksCm/3Y3PQdDOWFCNWGVf6kdDdwjtD+TGD9Xz/Y4RD/jROd27ikpKTm
FbwpRhFfowWsuTupfzxJkujtCAp4jos6tfNHk1tec/vfVBnn0fbWDruwb6RGpSkl
ExlrxpqM067XsyZ2hI9RKxISdm9X9C3Df+If8layFn4O3D4vh39mIcue8c9QbeBc
3VoVnZt1IGRXcQyqAsuzBTy5QFzVsH4BvR95vlaGdxOZRzg8f2kOBm3i6mFkGFGo
6JkjOdWmtLtq643Pw9xRC8mN2R5bpau3F8n4zyzefk4i0V5IaYXl3r60AOkbuJn+
FnNp9kUJ1owZGIfhFrUhIIX4AvMW2qbSnIi3XTFsx+iqTi4JHlwZU3astu9b+l+Z
A9zbm/ehitK6eftef7lmzN8E+8ycWEj939MHdk7caDPiDTCSqMB8B+9bGzwt73TK
3B1PpB90DdBzcouRoNDWEXsEeKf44g08yv967swMPF3YVPZn896ugcmkPQLNYeb5
rx4a2VnXzY2fINAhgAjeZF7dWQwGwezsCHqmUS3HaXnpDysxqXCHh4ttFG0ByqhG
IiaRiCV7fbNo09Q7f0AxnX8ImM1yGxDq+SAsKgW7Bt2/bwGrYq8RxHfXE3qAYepp
AZcIUq1zoIqmPPqcfzbvsTeQZLtPakWlBaEh5iVM6aKWwrwskgg8zLgTFZBlsJz6
eZOSgw/Q3ROciT8E9Fi0yV5gsvh/il2Jcspl79e4oT84RddgI++9egssYOS5D9b+
Ut0OmDMq1INrmfYAiKQ9ay30q2ClZVXnix++Y26ZbMZJKQmbB7qDYXxWdlfCYFjT
gDcrh9FU0MMCf6Id79BVx7mDvKkkooBs1iWg6jk4EEqtb54h71mmKt9JJC5663yd
XBFmBE2dF9MjuI6NAlGf3RgV3I1MNZa+QW5UvdfIK0WcxWCkyhYp8A36NLwsV+65
OINJuSNRpTllliW4sLaToQ7BsqY5/BSPZOsMIVcVriew8V4FGaN2CBK25/E5O0eK
RDRtHWEAVEPxsidYhpTFR69Ut9udQ5jWN8rXZaW4DqT5RH7jhYhakgZ1eRBeG8fT
A3pcH9VTc/T7l2L3Iji4GrcZTwLpOdxI8D6b/f24Yr2S2syW5OVO+nwq0WFXG9Rh
GSkAJO3SA28jjsbyRDjIrxDUdnPLPACsRLGvzGp07bpSEX80SltPBu+h3pT7LH0U
6fRyJNkNv9WIuSnvJXtwRl7Gn+PUmNrd/RnFppHRmUbpkykdJA85tPnc40J4sYme
shYMmFvHLDdezytOMeR794re/lTa0pB5yf1gOTPmVl90H9x0KNF6zRpPNmx7Lktl
2ng3Nzge5x8lH7lxRS3D9XXyVtudLuVL3lcGPYB9DoIWt9Ob551sSuLBWzXooqyv
5Z3mcyH3FvztbZYixQJMhBh+BPdYjSEHfm7Ko/LkuTirEuQxUHKL274FaGWyN6eE
WCi5YmMDon0Nt53Fmd5AGnuZzhzpk93ujDMyo1axZ0VX+3MK2Y/J7iHtTUBOMJkM
6v91l/ce3DEDOXbvO2FTxAeGSWtaQOEiSazbOFH1doFwXa5Oz56mWYXrgH87YMwp
1u2VSroJMph76bZSmHsi2TvVqCGNSTC8PcYCVLrLQzgjBdBdaJdzOiSTPsEeEYW/
6i2uAfRBnE+H/S0NnQjYIY0Jv4e4QqXdb3owQqULp+wc/RDsT0G6QlLWm5HneRzk
mknISffhzJH7vsc5UPRXcRmNRlzMRc+RtWOYsh2X6r3kcpmgqNLpsMmqxgyPyQ/s
JG7BJMIQ15JuJtOxKWczTfQWOmiZ2aGCf144vCcashRDVEGzJezYjWFuoF2uBIQO
SUAkVIpwB2Z52829L85+DKIgfehiUk3rQnLTvRnSRJv+anfTSIuZBsmmRFJaCDFj
8QQAp8i9hl+6CiX/xdFkl3xs/F3ZGZmt+wF4wr2Fb8ct928xIRBtO0k+bjo6NTL1
tCcq5wqUKBj8kpIWiI7OyRZHoVJwSVy4EF1hz0TYINC9Bpv/WC9qv2A7wRt219aU
dyAGwUtK3y0aIZf/doEJ1e4fIsy2/PEkQHBCeeWnloGBoZ/OnbgKaoO5qC8go9EH
DDV650Zf6RSgOgSV/8aK9MflZoG/Or79Zbmm4t8t97yhVGWMLUOGWpZvwYdgcxK/
yw6y8TRm+dK/P9VC5j+zs+iETLf2SMQLcRI/BMgXkAO2GxHBwJ8vtv0kv/R3w8+I
YbmytbLKv7APoNq2nwl2bp9E76g/LKLddpLjhkxrGWSG1cgC0U7NLhBuZ3I/mSDg
iqbFya+XQbBWtl3Kiytv75BOyyTJVCeMDQL5bZJv1v2VN2QOFd1VY/lcBH1z/8aT
aMZB1HNJNIqVe1739wC6BMIJc+fR9gvGt56oLSqXj5iL72sefx9vxKlJwSyk6Pqv
CvLGFsrTDP1fruqU935Ub3gLS+Md4o5r4+8ojY5mCdAvsCFbCJgRBYK1O9qkA+m+
HCQGGYmC4UBA6dXaTrBgpUTuE+OjhNEG5HXimSUOQ2TGvH9XIgjna4Vm3pKvtG64
QvQDgvZL/9/fA89nmdXS1YBQmeIyj9m6Rx2/NFvlmoPmVfW/KKZPenahAKQvA3yW
iPWrX0nYVoeEeF1YNRY9aEFp/TK/Vv0bnyMfvQmC85rasViVbVjBlb45eQOocKAP
eAfzA6sGlPU7HqzK3eqTMWJiH6YWKQJJdqZuU+mO9CHSaNyF8EfR2hbakVgXBu/m
fRdVhNH7VhAm1pUk0eNwV8ieXzgTuzWwAZFWEv9t3X+fpAm/M80dXbvW9m3RoPBp
xHMYRe737GGfeiE+flyBCmot8fRbFb/ff3sHKmTEqyOcrr6afWy94fz83L//mW1Z
Uj/BRFebIIxbKfha5FK9q4PWCbD30tVKcSDOsTZjBhGQY2oSzgMzmmlpMGXLL+Bu
0RdUU2ZrA8W4L3nTkL78srdizDvhBQFUFMQx/qqoNZjNcXbXdk5fNdMO2LmcSuGt
uxjzL0QOZjW8nR1UuYiz0vcGVsYz9G9SkSiT29mtXkWZIe8q5qDydlhacCRPuT/x
FUbr1o2Y8dDKfXosMc5QUHqZTR0AkzMy4YaAxQ5AUChNIDi2hojbSN1T0mtNC/Pf
qI7FfG08YBUOjF8MgKDmr/UCbz/SlGx+3AEotFK4Ht2wBBU8fGFGCV7+nUJ+jnFQ
1Tc0vLvxPSQ3PPqBBJ62aHUlb8Y/6mQeWcD1Hqx9B0bskof2EpJERdgRxdqhmGaJ
n4GbXaI+f2FKkVA8VupmnTeaU5Olbz1EodSB9i0GNg1gWTopyiCgTsrmBNV04a+g
sDSVWYUfdd7twUSElfQw4/gsmT/K+XgUu9W31KPBLvgyf0sCd7usvVbYau9HADwM
X8LJJJFx7D0hJvgyXceZpPS11R6lL2/lpi0wqhPkNJK2vkr23Qdlfisu6M06R+8G
CCFFkgqlBj+Gz5AkS5/cSX9BKMkC+fq0jhyIg0G+wIETu6hf8g0QklFPh4IA+ciX
v1Nb/W/dBD122brIl/DWThFFynJIqV9nvnUuw1cz0EqQvihThIAJgVhx/SbNMyFE
K0sMT86xf1rmZrNIVDrcDOEQ/1qNgk8/TOTlvsUT1RKq/UTKrlIk6A9MftPfZsat
zu4h8HRgDxWGMhk61vGMG0x4mzYWgwAWqCM5iobVIu5ExqEgR1VJ1PXLdKA7k5R7
uO9OZ6uSfJ5q/i+7+hhlzvhdvBGGA30iXExsZsXg0bHw52JjqGKTy9gzG6LncoCy
L/3TQvEwktSUsiAhy6xjLWCoMfA8eRcy/C8+KvbywyHN419yc2a5VAN0B1h2oNpj
y5zJ88ZJmm0PF5M46l60AqSNgLvCyKeZBFLuD35mUxshJWJ6Rk/Zqm/iUJw+Y7ey
UToUn+JhTpqSzMqPNz59o2FJ02G+FW/wtv2D1KzJr+Ty7H+/Z7+GiJUgr52atGqO
StmhOVuVPaWsE8ZJAj6UUhXYD1ViAaipzSwViJP5IKDieq5eFYxF5Rs2xVGJtfOW
p2APbUp5jcDj2NPTcA3d8iFuqahIHndqRpy0xSM2zOOZNpy7WLopnQziOmcKSg8t
v98Ddu23ij3Bcz6azzsOI0MrH5W00dJhBkQ2Fz2OePDjmsaLwDbKsVcdbJChxSYm
fymNV5pGgUUJEFfKuDS2kltpVQwhm/zi26n6SYgdw/FMUqcVhiyFDTsa4cc1kbyp
SdcT7/4NS0eAp3O/5SXsmgJI1oe8yuGodz7gwcwYX8B6VPUlWehaK8nZ76dd5rkX
FHGx/xrSCBOqlmIzBXIW9UqzUqCjbPwbHqD6aud9eBjyq6aL5k0ZxDil7MzkIOsI
C/bLo2Q5/74KJeLGUE+tgUfG168/E+cqR394NluoHVq/RCDNOGLiBQW5T6WhFo7o
uT9yz55WMIC+PHDT1jI0jTBfWGxt73CYddXwoBNv+GN0NhhXTjU2g8zNIcElGXzN
dxvjbe1+XBOfZaaaSLMENGK/OO7yjkrW8F2fDOYEnfw225Wo2CH7pepRAQ4cIkLF
X5+YyphZSR4RkauJSE67US/XCNS++cf4Nv9ErX69vGNL9nrn8HTD3bVEg1OglSzl
PpAJhcjtFeGTru1NcwhPVyQyoutr11LUiydG9YFfXzz1Bhpx6dPzRZVfecJGIMYT
ezMSURr7uGhTFackE3xfxfvDkS37PMzCcvckCe6NubKmXksu/h7n1r04nwTixuia
9LRv6BmxJkoAJhXgjXotma2k4X1hH0MV0stWGX+T+7FuwvYjXMDzqhznBaSJ4PKQ
yfENJ/vCnRpMdQRe5UIXkKbAMkqCdicBmFGw5Wt7sfktQfAPJztLE3VvM2BICW0l
qdVSvJ25EgfhRa7SJvhXpEBRpdIaL4uMyw9CtqYV6FDXvM4JLLbGx+17pA5Cu4mN
IWgAnXgnVJCA01ZTXbWSHQtH4rqGuIPW/tJKkqdLAC9Cu6WCYNrPoSEkM9bJ/Re4
jr8sAK6Ck94Ts7sPrelKZQKG2+EMGc5ksBeNCPY+M0e9d1sULytb1BzJGFqiRTP2
CNXFJPmEyRqp1LiYBeSGeRAStWJ9H2dBrubxTeLDAPUV+QMhRWbFk1TEG5UtO0Kt
82D2sMM4NXu/zWXFufNz30ytKsPNKLxdpr+4yTEzwJcmZZ+j5i6bMp7qcyV8xDDR
Eb+nDXwmUd9fVLoSacLdBeVcOJIjZckKczK5LOeHIJaCvLXB91LPg0qiVF9flTQi
rLb2YdWP1tp8keB4CDFHpv+Jkc/47qPw8nVjM8Ae6FoAhE+W2FMwo6wt3y29q1k1
dqJCLqQvByxguSdfatkY1r7H6EgYSOPxNONRT4IEM+SM/Dqbh6ginOGmaBfSHoJo
T3LwWznbUMh0fFHeurhvl9xtGA9MuYojFSjE9niHtFBZVw0TPc2U2uPVVma8sdHq
bgFPUQdHCqUhEElQMPxYtIUw2KSj+QbA310EBIw8OT/kV2TgeHHltkNDYQJ2jMmo
BEeHndN9QlynGqecoXQfMfAoFp11715eZR/Axb8ii76eHDQiKhKR9FnhMHA/Ga+5
SXFhFb7RhrqAAt+wHFxsGTDHljqTHg2aWTywqwLWOq9xg3xfQLqCbfphCxaFsQUi
Gy0Kba9+hraFHP9POTnWiOJnxGl1Ft4YaHBlovOsJdYpGUzY9aPbDJZFqLMj/L84
YHvZovDLMp+8I3bVEwT6vXsHCYc2GZsYzLoiaLn95011gqH6NekpXoHzCT4eB+1P
yhyQhD0lfxLkR6CAicdJNBFhE7IHRMPmc5UEADYWorjgciOPHTSU4FxGt1ox981W
YQ9RHG+q/IaDDmnitaoEPJgePF+ickOyp7FfaheffPQ6fu+rNi2c4DOyKuh8lD0X
QhVWPQ3YN8TWLxY99ujV+r13y2l35TXx7u0x+rXRnTwAAqq/C6MRqevBy2nSmQS6
gjaXhk2JEkEUUkiAj5scOkrUBW1jG8aRV9EEu71Eip/3+V+ctidgF2oyDo5Dxexh
Fo6lToMQENpg4smX+Lm1Gp28p5ckdpIlaQ07KmLwTZ45AokWekSbEewh1jTGIe1G
8VEmj6lBiGtJxZFl8kqgJU0rP1szTpS6DH8iNeF/k/GAePgFZdKo/uSrRTBC/9pQ
CVHzxLBj+qQa6msnL2v0GHDVo/veG0x9tINYL9AWtwSvNW/exv+W4w2locxOb7Tw
6Cuvo3DCYqyX+B3gGSquClS8P/v+dBNTnCsR8GfdkLIMb830/qkaYjf54J3MM7Uz
iqiT3gQE9cZ0DOjT2/L8YJChlEqu1YeTSWF/mT4+a5fffD+upJAGVcrffu2lfp6O
NQMLrujrHBqRkjz0+9UP85gJ5+CKlv5s9VFDp3Chf1laznebFl+gGH8B+DN/nBcm
dNZB6nDhDtY/Tshjjk8+L0cRAI+YFEIMR1UhX0fsaBGILAJ9NmDdCiO/yQvMOUPS
DcSXsSW81S0gwnEva7jHZ1TSi9/bYPznOzUYh3hJQdLf7W10UdJdmFDtewDSpJXd
RBHtPhtW5ENqvVYHRDbcw6FF9ycYiGPrdyflhmpFiRfcClss+HUdahAkRQFR2ZMt
3KPJRIUDaEGtj0foVrAObqphFHyny6lVHt8OEfOIXXFQq2yelpm1/ZSU4Dw8q7e2
xFjlei0teDGq/+G9dpsi6Xgdmsx5CfDnKYQgtdEb6q6LTo+KGi7t/i88Qh5GFGPX
OVL48jj/+yfCDWDGCO4bHMlBvj49RrkzvEaUTdO7eRt14iM/nD0V9+gNP2Sqmkx9
2ugGU2RWTIA8RzXOMOGUNYxIUvKh2xmCPXghSQDIS0ZB0FuOA8yJZA8QW7Y4hOwE
Ib16AglK3Tp/knpYfexsyhle0577ZDh/tTHPvhLI5ntLOvHNDO1i09ieP2qv6ed7
F3U/gqxJJc18l/77H72s1lOecfy3u2am8gNaAR1n7oNpCdS7I0L0b+R36X3S89HT
SMNyuzjGbjyR8CTvrHVyUS31jYspyWrm3X2//otCNE3PvXtCBuFznSjjxMP7obxR
ZbcQVvlS+ftbUo0RtKXr6l628eGNnzBezPb+2puUrc3tHEywh1fS5G9Heglf7IBQ
OLE2rFxtsqovjw9bqBP64tt6MYY61t9cPCaE3cJega1peC6zQ851HC2Edinhm207
5TMWY7KyHm0TRYqwNtgv1tYA6nPdZCnoDifGTBgH3otubpnInPF8mEGyxb8+k4fY
xYYLuPzCYpfUV782HgNzzTGyEINapZ43nCoPILClAdKwh8oSOIVcsUN9v2Q2sr1z
PGpbxxN+jAocBJANDnrx0LUVmfsMRkt4+kr3aGMaJUE5EERJVEjVqmgco5cx6TL8
w3uz7iHbpHJgLs4LOtEsZolYdGGDLoqH+ekfxEWn4FclXWSMMorQXqlHVNp5Wd5N
qVpDh+QT504M/G/Dx9TcfWuPP0bmY6qY00I4PxlW8iS4i+8yr5++vlbUE57bDIUH
gc2aluWIPQDqq5zo+lerhDDSC74+IzXqxPGxUg3UbwgRbcjR+i6NobEpt35SZaFo
8dF8Wj5vzU25kfIzztne7bwNdsysokp0Q9zd9TYTOgjlxKX03iBjPOs+An9xUwJj
Kpg4br3Ez/IIWGyRckTHBG3x5rUsoRGJYH5YbfRfvH4PnZDwPhKn4V/ExhNh4HTn
PP3KNmWu4MLtZnV+/NVxlXWkkYXJy3AXfBbA6wy/o2SfOEv+YMrU1DRHX+Zp/19Y
mvVqVV7gABMlOsJQEsjjvmxIUK1Qwc9ju/BA8d4n8BrI6xz4tqgUdmab3wXuKa5R
XBdlEI3VMKW8LFbIFk9HiGfiJzMyCojnrCLrpDN8ajlx0YQ/3JqTw8Y2wU8SSIgu
jK8qR9+0vlJCCVPySaKyIFPrHxqhZOpsOYk5geIrJl0g0dUYjnPGo1SY0AOm1u7h
/00wjRi9SLz8Ta/+XQTL0wWH9C9j2BQWHpoYCOy/PmuiMGvS4Dh3MlESoTwua7Le
tcy6ydd4yyJFaex3x6mB74V8sSLBEXe8AQa4RVt/7HAs+GIvIKEpzalbNXwpKf1B
7+T83itnPbh61mZXPKt9/RwtgMpc4qkL+vZ4WZgFO6/V+bPez3DbweNu2gcvJDMh
1bzzjFc3dOnQfVIsmqURZRotpZq2qt0LiatLTsKDEm46W2DmMgH9b3IxXHZKcLLS
VrGtehkun5fu6BEg281b5HWsAHdxnfyYdfENP6IWQxmAQHfN2KY7DHhl+VGKVmfp
Ua1uyaoN1XlKKETkXWUG+kH436H3r/qJIuUkOidOWfpIr1df0Cf1JonaXKWjOD+F
TmfcDYf/6IORFuQBXKqMaOloSb0Vbo/TcJFv8zucx5JLJDDswYpW/hnevaG+oamS
ZUNCr8aS+JvtXYhA7rKDXc7cuv5tkn0nK6dynG+xzeyClZqTFmo+DmXS4kj6ryJQ
1WwDuHq+1oYBj7mBLLYauNNLPnKRR1cb0nlmnoR+YbwzxqfE6E6yKQZjF6gg6/Z2
UIYozPTE2IgzfM63h7eNPDq1xlxKAmaGCiT3bJLZ4wlnVXFtY0Jvw2qxRBu6FSXD
F2UPCWklFMNwC2Ar3XKzt4a3XKpyHI2e76XTC0epr9KavXiA7ENYgOVM3FPLEEFF
XhTEJT6s1u95LYhIUbyMhz7X1EOxFnBAQE5PYx8Deb/7BckpklP/+X5K4R0YlnV0
E2P8/pMX0/Lb+lZapcR2/gzmhpRwv4O+IxSI0Mh6PSljAZsGcrKTzLu7lrnJNXO2
KGPnnG4MlZN5v2ZWxlkzwiTSk1Z9CBq7xM9x0nidtohekFREBj6r8EDwNro3cuV8
dHoRUarDimX1r8rH/bOMnWbktjgRsAI1XV3Dpew1/MjnLM2R3GTwWZiD4WXkrx0o
AWpVrSyELeK5NKlHAUGdb/e1fySASkJp3rtBItl6hw+YJdS3I7Tp116y6VhMXUZP
aHN/hW111NIbtIpFiCF7w7kvTYFIQNjzc0RIquN0q9ePR6C0aMSTJdpqQsi0HHp2
Idz2SkPt5btAoG1dtT3QpOzZ3sLfDCDszHpROnVbaV0+OK8RzxNzGr9mAtAy517Q
ye/C3bybtTBhgFZCaUGOz3wd+aMQyRUIQ41FgPYOBvIFpfSrx+/d9oDod3zP81I1
fRcbz0cOe7Pup3nD++HMLz+QWzSMrG8Ix5wWPBipL8GRAP2U9iosZcY5NJCI0wzC
ch40CfgSPueZWrqx99NpeNed39nQCV1pxBiZVM1hbI5LiZ2zMmmWwe8EQt2FodcZ
Yk/5JlU7xWsyxkFYSvoVtCGt/2xgdCxhkQ7yW2o57MRShAqHBdeO9uV5cy0vJVbW
kjQ/RMcpXwQH31LZ1fLcCP9yYf0iPA3oBXQD2+CskleFzlmtq6ZfxO5yjb88rhZD
2F9WzzUFnotfGD24lHBU3WdinvIkEqa2Ln0BScA1LWFaTelSvOf1S1D/61Kffrjt
yv/WnkoM7U5q5PTZCemtKLNW7zGBrBuV+X0cTcjAX6sSVf824/R2QVGenhsI3er6
j36H5QSqTkexAYbymqf/9DsXkB02jVljequLhTNofoUXpJKTv/2LkI4n9TrNMPXP
6SxO348EcpWngT40X7eg0/THhx4Hf7J9LMYZEQ5uJWlaZSCP+85l0KUaHve/IGKn
2XvlB47FMliiW8WYr+YEDFI2V0ebHmJE7W0MbyvvYAT66zT1FsXErdAQmqJjuV41
n4i2bV14iG0Fi3g+uGU8wj7baZIRwZhRQnAsxdQ+WIQUxfaILlGqog5YrrLvJTYc
isjo7UrZpnWjAiNyQvCrcC5iUNtGfMb+gbX4cb6v3IXtJZmlCzOQJIZ9PAV4Xuru
votawK1Id/eFHy24sQShg2U9dXnJ8DmJiuXpM+T0ACsk+oRuaS7ROJOxm3qqNWWo
M068vB+l99PPo2egtC2AagiyktbiMh9XPHc+FpBiUQA8kzILkwvsMdUpgEJ7Dv6Y
on8Q3UlAI6wDks7pNz8KaKK2oR3FWRzfPoA4LILWW/m4YfMzNrdWQVSfUXjCaUZ+
2zZVMa85F4wgMfuFzhvtO1JCjzk3Sdx49mN12HCs7OHhgdmdl9+Bx1aLeuk7TuGn
jGX5Jwe1vry48lQYzsmTZ6V7GSZ3EIrVgJrdFficUftqhDq1Bj2DfHq0UFpGgmIs
uM3I8NSJN0n9qNHNBhYjyGf0IDXdxTtAaQUPLN2ZtVw/xRpwVscAXDcuaktp71kP
09a3bJlwLtvfprB+SyH7Hh3zsVgWysLi3aDKp+giDmHQS76sISLesKGM6MZgvibj
LL+7hMMDTK3dVXuMYg/TttWWCc9Rilvs1klVlYVwNPdsCWM0qzAOTzFAxcBjKt8m
lY+odccJvQLURCNElAE8m2Am1CH3DVJ8tctwtvFtfui0iXDnYicfApeV0Xc4ylb0
U1QYfmIifpac3buN7B96GHM53ZcS79NSleQjzNlk/7tLfyOnpP5H4PyessSGKaJP
Q4GZEhOud0xZeB4RNoee2geopLb8MSN5ZIkwuLKt47nCK5guRvcUBRs/L2VrPDVD
ObwAV1VdQ6BqHNOo4mRTqDlEMXcwrEQDBZ6SwksXJwscwZHSZ4OlXwosaqo7VlqF
qQEAVOJZTb91DL60L+71J8L+azEevkNLZFbT6dPpOJmzwPkj+rKuSc6sHmZe7Kyq
5nA/mcGv/Eu58TpXQfm+SrsEehYR7z9vQytUK8fJUEBWxUFyJcqu3/nbFBnWRPkd
MC0cRUZtM/6J1Ld7C5Pw2bY0+jvpjmxZF8DbhKsFejmW0PqWIF84xfWgcKzWiQpT
RKWLd8Yukqp/MdIezXWwrdq0KbmfBgNHVrv2skut1GlTQVzBkGVhijbEnnoRi5yS
GyiihdUYG6SPfOAEO5pJJHMs7opp3GYulr6avRzMZqe0X+agMdMrqUwzMWBDz5Uv
4tifPzrtIz8GbL4MdXSHRqvq8DD9kLZA3Q3gUG8VeiECYJd5twXNouh9rTf003HH
x+JYLt7fNgFjWCkiDXCeKgXsJKGvW4VGtQC6/ow72azsmK8q5y6VPBSTm2L9qSEQ
FpgCHLHBRU0dzqyf1BB9F91UWtevBYb0zvPJFbhSjgvkwxYxkp8j8UHI64oyZOQy
hXJqTlcMn3Vtz2V7E3TIPZV88ftJmg2IoUtgg1iJKWmJpcJT1dSPtQOKFyYavKES
8EC2pkz1dqQrR7NhbIAScJKQyUe8RxiDD66UUqVAQKSmcu7zJRF21gmJj125VBJL
cNnb4krsAK1bdra/D76nKbEmVQv9qsP8aTrL9QCnD7YDregEeHH5jz7fDr7S6gP1
ZeG/TQkixsz99EuTSm4hHy+8yGxa89xG35uFD8LnyISmHOII12P+Fm4XAr3XvuXN
zfmzHiELtaN9UoqOlOgH1cTRI9uK1u/9pf7xJJhfI3SOTaQmfrbigG152XmjkjNm
uNqE64+TmiqIoWV29t5zC31V0MK9Wc8wB0c8eKgyu/ikIpaFqDNkhre2OrHzgDbX
xfUVb9DKwS23P/dib524ZgneaDBiBJrEgnaacEqHY63c2B9uO7QlPHdFHMCxQili
7kiiqt+2ecoQbQcRVPnPSJVbMFiPyCOKCcUZUtOpVUGP05pk8Kul4giLrQi+F4ex
BObUkwbthH2nQJFS+bYilBgZfYGn3LxvVVKcj3nig3rjDb3pF0nqLl8gzT4E3/7v
EV1JV4eEQK15WusdKf9uVx3tt8t5sUY3KbmEbdzCIDyWZRVXEYO2gflc6TyR5qKF
bc4SpD22/FlPhLQzNUGaXwt2idoRnhYW9brnjUihzLBakRr5eA3T8A4uTjyTHCe1
1mc4h2gCGdZxawCauKIxg2TPqkMhgTQK1dL8smHVDi/TpqS0xuNoUkvJpRh/ym17
TobNSsYOUjuBU5u3kTr44v1/fs9gMbLs+qHURjR4bK+R1pXWa9RzFdc+oX/3EhZ5
ugmV8T6pJG0xeqCzNEpSVRobGcufMAY1PbyibWUjclpBcN9edS0jSvYW0NnxGxfH
9pgsvTKcxLZApXRLP2XLw2/d4Rfh9B4Pb/G45c3mnHw5NIi5BYb9YGOeP2bUhZ/B
p930SJDAiJtnsEAgZBzr8nIhYjHHyj9sN/Z8jQAnlHQnJEbyw29+xjbUzA6rav0W
Tyeha+XiWYvUbo6prjkAC+igP46j8tAu6RxbvgmwjwfEIOvMyTc4CbXmA/J7kX4O
Ja/iFCHl8Y4EUN0mkgV5UoXgoHdIxYQcvBzUAeRh7ekLfq6UFg/1L5t9lJkxMtoM
AtQ7bdSzDWmQazKayT1YiCm/HAhvkmscsNSCZX9t13GU8o0GWPLGlWHsH5ayY86n
wA6W1HjNETkYmsTUoFYeo1MvLbHnGiquEg7OZEcVeT+2xJBQILvkfLmbmMWb7Cvq
tKzHcjl4T2y1Bdp+PapDskeulNmuBQgDpS5jvkJQZF+PofkrnZFxAlbuYe03BMtK
yIYqXAzbX5AS0Vtvtg4C17oB7RT5N0Eu00wivo915xtds2aqiprLz37kMT132/gX
beDubz7NF3P7SkMva26ckffRcfgLYPctO9BLMI8CTs8mSY3pSAMor5iVBWeSc+wj
FnN4WKZ072GyIuqB+3Iz+Gb8Ml6/JHbfrE/qMpj07Zqvr0nmflqD93SM5K4Mbt4q
B/xv1Ua9K7FWcl7CHGHb155Ew5zkZzXN7a36bygLbspztskv9Q2x2UA6x4m88l0t
OCoh41ew7NxoTYFDQ4LCgIdcXTnr31fEpy0SCngqGM4NGlD5v/lmQtywF6r3KRkt
Ov/QBtfO0v4Zbn0i3HhumJ79BRSPI5Sw731HMiXAKlhQedhBbmgshNGzXY/Lt5jM
YY6px3BTtHqAc8Va4eR7EAgqbJsKbM6oDHcVWV6+C0kxjovDRbEhWDLkltOYH6rw
yMzBJSqq3M2efPR+CakiblBs5dFuuzaw+o0lCgEOnRun5atxPytaj4Socw9QkZPl
fWwhHpWaO28Q1t7wSc1WlpRm0hbOACcBJ3NHhfEussdsgJVMuR5DdXj+/hcRE3DH
Hz5J2NJLQFIDCTJVyFcSggDUHcmgcdmdcpokteC14WRlJLsxx4f4Ko1hgaxLTfBY
3m9TPMo+CzzMYj3sGnWqC7bweHVX6/VDwRGi6Y/+MSTEyGOpT5ZjXet/YG4Kh901
8Anz7KCP1ndQguOLmZw2dWVfduRb+13vHwsI+lO/EeD4tbQ0gM4qq20g+wIKZifO
ffQgUlAP75xkH4iyQrPqGHgksrEszif5+7TYm+gpCVREpx0D5oRW0DubAJdm85y6
bcg1E49mRU6Y79XIIgTfBTcEg9SM5PFtwZWxt+N1AL5n88rME03H7kF6Pn2BnNNl
7GkCrrbuAuFwhDBhif6ctmwLACo31xZytepITUzVEMOxTHu3EhH6JJmd6/jcUGNI
PfZugdYsmRhMiUCfDVih9U/2OUS/gEW6XYe5IgTSH72eiQ2my/QD4QLMNM9Q8Ppl
qpyIkdyRxzH/n70tzFX6hzf8wyhJU1StUIgldJVQVM8Fuuv4rOcKTFHV8AP+NVrU
7JIZoM/64Eakj1cr5ZlhDvOHxKcEGfKUeENZS60rmhwmaXE5iamkM3jBb+2QNQ8h
H9xLXJb7tsvI3fKndLYzES21Y8IEKe15tTrOi3vfqxL5lf1qtJk/aZjTF/WogFWB
b+vxcFvnkz6+N0kINylAWiAgS45oQNARrN9f2dYTHUsRGUxFwtU1lcdjyYFUdgDP
zTyaqKfSIpQSuMNGandqYBdsoMIaca63Ec8s3t8UFovBXn9ySxVtjTMecviKWor/
wBeDoDgDe12poroSg1CWmcfL7DHDu0SeALGxLE3V/FNPu7fgIJReAXw7eLkGB52K
CCijnmNmetrR1+BlwM0LvwiwtYS6ehkKCQGr8KOiG0flcEWsJbo8+J2L4cWLrzrY
iGI6FU9MiLyyDfyWmbP33dN+iSYdf66Ph7fLwOBQsEohzw/CECn5vfUcTd02T+wa
vnvgNiIl0inNEiMD2ulr5mFJRyBlIt8c/93uYPYSsmP7c1xXmzKk9DBPtvJMlcyT
DKA+7B3P1+GirPlAK6A0IYrRr2eoKx1+CL093X42B0CsykmnongM+ByeUTn/VhEZ
IyO01qa1kQdna9eebog2YDdIM4GY4bk6H134jZUeg/ESnEnO0GukIkeJhiMmygt9
BABTBE7vRd2ptj9jzc64EAHawiwL4xF/8zTFbxxKBRVh/1t60GyMMfhCKPRbRKNz
MlE1oZXCBrtmCgmlxg5oWONguRJU9SD2816YBAGzhq79rQ+Nsfm+IWOb2WIBWA5x
RtNQGzzbxKgwj7KZQepTpev3yC6vhDhimhNgzGoHPI7FSjwYekq5PyhBxvlIR6Ti
bcQQOgEoEA/fRBnLmuh8Q7LSOIQYnX4B3C2vcN4/eIYNOILTT6HkO+bM5kkV5TnU
42UMTkMEmNNq0nFQjh9DDk5uT68xYgTCPkg9tgtxXZ4k92VtTbBe8NgDMgVlY25i
j2nx6kXOoLs9YOqhkoG38i73hYqRZGFMLYBfzREFw396IoWrbkp+kpyuvHIcbCfe
EZv4QWfU5OgtDar3v9YGy1rE4OEWsl9VkQD61twZ3oIdpCDcBtDTGWA33Dtpr8+9
XWb3x6HtFUjgHdYbL08hUOS1vdlwJE5NAfqdb5HsNIqkc1aI1y4u68KTJytUUC8i
TiOjAQ96Nnxo0v0NATILEQfNbVGt6ceYmA3cBYlq+nXd7twSnYjjDTPPx/6lsuP4
xWmfK9IbMpKY5jmf0xnHwOZi28Ik6/awLAl68ylN+v41dpuorKVJhB8u59qpHLBn
5DuJsYzRH+S/PDatD1xIN+1dp+lY6FXXt1MtiMz8HtUl4Gv+z1uQGxp2O1h+2yBw
4FxA16cN6hwMkqlRJPeDXcLyZOv5wP5o1Fj498pbH+r7jNpZcwlpc0bZtZBrgj/4
3I/vqs6oXJobZcQT+RQWFJbFeQ477sWsJSP7C3tubDx8KdtFiIoh0arYzacXHD4S
WahdBplAmsspNzY96RqI/CaNgtVtDEDq9waqfLf1bBi3fijBpCUBoZjq0paT3Dq6
4K827iLVeK9fAKIeBkfEkBnyEBubAIySXsfgIgKaL7Q336RiYJzED76F2DRI+5yn
4OiM0eVY4Q8RUj0QHsrABXKZmPWQpsouMIQAoDMaX3B5OpSpIFpVJFF55woqm3lM
UsT/BazNIoMeZG2yhYtVSBX5NRd4+EevVxxOY6ukhBrA6JbjkEtrEFE85oNFsIGa
awygxHRNgxBmqHqKEAozXiSWQA61XIsIM6tja/HemvdAucNDuxojSWGEVuM5pi9h
z+4rI1hN4q86+QkNXPfP3Zj3ol5ZGFk4kdwD7OhnxPfqbfmYC6HyycQ0j4/Mst7f
a8QAJkqn3kKt4IchAIBNTgn/Hq3X0TCSdd4arV+iVpFuOYErn6JpZNsZp+gOABKw
9e19323ZydznjDxEwM9Hjq710UFrQddGUMQaIT+iboRppUgkjnOFPybgzcIDz0ZA
oNWGB36y1HIrcdh980gljDvQpqj5cfDP2bK8TFDtsQaeRUBStyG5KsjDJXaeL9w7
O7dvuR0BMl/7M84dY3Ce+kYOOmMdAYrM+UePGwsFcdIXcr/N0Ufk0aGAry4XyhBt
/vPLazL23AMv9qw7JTsfK3s4+P7bAn2KJhd9XISlRxAR0ki3Bmj7cMXRJSLvgFkK
mXId8lrgnY0SiXlWHmS4ecsMMb1b5HdimUKn0oP28cdMRXNrnHCj3+ki07PCLL+5
xhbtBxkCMGr/SteeAkF7upf0s2Vsj/ctMaUHNM3pYF/nR1LRrGMVmz45Ga2fMGW4
EOJqSQyGIYQIh1VrbJTctppCGOmlQip67bAj0etqLCPZDZayCEFsYtEGjB5tPkL7
mbMHE64NhCxK5KLc3E/XVq7qoDHH83eSvjEYXl0UlX4a1qmVjZB2yLZzsSelxYSJ
ENmGIgr0ctqpX4/JAKHNAS5tlDMWu0YHDricW7UphCCs3fc4JISLrSCUuswtrjX8
BxsWooHMUxLSapiIdItvxjP/8Q9jm7CnJ/1BOKsOgtUdbo/ovrE4ZqsRTgw8PREI
T6kQ9ahcTBMcmQMW3NAx6VKSjQ+wWrxv6/LhAFcjHO3qmNPU5kWwfWpd4farRB7C
VxZm1Cha1SqGrFmSagBBVZvIsALyUFgRhOYvTMP9nA3hML8D1+56U242dD1ua8wH
AxWB/xWXc/YtNeO8FWkUXkT+GWEsJuFqGA5oOxDq+Pv5VqJ52Wp4xri+fyox3Sd/
2gISRKtjeKtQ+moH8mQfAViF0lB831iiAiHXkLsB5Q8ih1pr/RbVLloxiEtk5kTG
2AG4KoJ9O5+h61yxnZt8hNdium6k3tAae/qcdOrUr9CMnetzusDhVbTZYjDLXmuI
3MyKfigqsMs3ylnRpWSpUe/sGUN7ZTEQHdYDwAtRsCyecMu9KdSsIjDkenl7pA8h
DxhpoTLTthvrokW1kPdmlct86bndEY8hONp9B3wBc93smKI9pFY9L3pkiTcYdcf8
jnBIndYPa4sFaBpy2eWtJyYttj9BWerC6SIHsQyiDZD41YfLL3ZSbKUnvGrvwCFV
V34itJmJ9sBqMbUohHTlhE/fagbAd9b9rfDGK42T7YYmlLNnky+xzGEac4HdUx4T
qmRBEKExmcFi4pVUjB7cI+hx0afHFPIy5/hh4uzALx2gI9pRYIzoGGPBH2oduZ2P
TiRAG877oAbgYhpqcwC/Gkl3IhqUBnaINYsKzVKLaUUdsdr9P+pT6IzHFadDujP+
COlxOelcEVQsON/nJadsj4iPmczSq8p6EEUpNsFUl2nkuvhZfS99nlXjJl61l72t
l8DqixfJFsWhrrVgWP+NiOFDqBgurz6nO1QWmU2xijShhYgJXn+9T8jbq0AEzXI/
elgqb2G8bL8HI0F0iZUx5/1qGj8oA5dSb/B9Tul/cDqNAzXcapRXCfyDlK9Z2BNs
OdJaz3R3Mr7jBnactSkUWNLSN4R9VdZMlI0Boy00lm8dxzD4HZ4SGNANdZvtdc6v
XpgqFE5vgtLXJ5E2vNUkCx2w0x+mme3ddOi+6Gq+dM29OiF7i3ZDBofBK4IFNSU+
xCtDbBgnCcQSWfuhL7njxlmW6VXpBBfjTDyC4+DaKtqTgH36EiB/4QcSESRAHxFz
Sb2va1N8QxPbGYEROVlGhq8pxbdt7r+9wu1/15kqkLd4GABMicdc8XFj1Q/GP89x
xOnNvMAGNymm8PZbzpkJBoebwcEeXupSBNZs3nDn2tRc45p8LIb1OrZRsvkngXpX
4DnbK8MkOp913FI0VlahGrheHi+qja8vWqm8Xu4xJiBISOMlgqoVr2KpAbk//JXY
20DJ9SsGQtT4rT9p7+P00r2dDB4TCg8WSEtqow48YzoFNqoixSJTTZiC0WDhyRUb
wH19ikrRvEUlO0GX7IGZgh8+SDv/qdrZplJYm8dCzjgqTNcKgRr7sZKUeOsz+NVL
4kXKGDKeuMFw67V6ahaLC6cAyBjfyr/vyk2hbN8NC30uT7EeTmkMkWNhXzbF3/y2
CaccwrwFBlPgBbcyCo+gxI+68LtY5Ey2dXvNkJp0vPSpwuHph0Vf/4dLj/IzUMTy
NCQYhktWpcl7I5Om6YrCDTtYBVaTygAI3yJ2jRkir3fQhjv9p1L9SVU1nyLeTqEi
oYNoAUdVn84zuKflygNDPmYuNE/BpCXK9uFxOwVoATs6toU9a9ai+a5fAWS0jKm2
ptsgB3K+yImWrYteZNy7LIOiCwqH/9cPAAI+8IflI26GBoqSfVtKMxwasZBE23oE
80Qgsgbeb9Fr9pWVQvtsZWRW4hc0ZB0xxfI70tVkZagqdY4Ez6GeYfyqOFjGcW86
SJ5YuFv35CXnt8nU/OPXSgt157sQCdWyQDlcHCVokLdeUcFqWYnUGmWgog11B0Eg
wI7BC23RXgvQszyt12CK2tVQxn8Et1tAQ85vPRWXg6AHaXHIDah/eTjfgv3cgxo5
Jk/HZoqkvZXzsehbFNcKtl+bCrNR6c+G0s71Pzfa8wSlCAKTH1EokjckZWG3UCy5
N0e3OHx09Y221VItq1vmd7nL4xzs3F/bsnma+Kh4F/Ol6zMdKeBcfsTHGHgFQC3I
2CsXduEnJA0+/invxBmPOIb8puhIy75sEiNXq6ipFbwORZzMqWeZo0A0vugJ91+6
rOfzwY4MEyPL2cFxAvcEofpHjOYro1PxvZg/bJHIAQ+H0XVNUqPlp3H/48X3Jey/
nnMHQnpMYZX9UGorOfyP8thW89Sd7DJ8l92tlPOYSZ4tHyEdTDxQwXqWy/+bGU5b
OewA3cW+S7Pl4wwYYQc5jjlnHljCGuQRC6ehhUIDCWajsdZYoOs6vphP+cVFNLf5
1sV9dvcB1vrD2+I0L60jefkMynfZbrdw3OHWG/dGkUI/ihAR9Jg0KBw7+CSHCnMK
vKkPpaiX7uLg1dZ1RAwgRw8v+1tHMwaEl9AIrRv8jMVrlVKChFk2J1iJbUrkc6jt
wEdVlwmQY+M+vF3ZWghLyZbuPDw45gGZrOhdRqAO7X+g4xeL0auj0V5n1uI7Njbd
l+15+VRbqWiv5Ma1yp4Nd/1qr7crv+lK020W9cp7kznVcqHIlNC0T4GD6xI825sy
Xzth1sTyygMBsbk5n6saYjHs0cM54taRvDNEjSNnFO71botx0OL42brbx9pHnUiT
WbAT4LnGstQznYfX2cyxlPd8YeVxFQ1oIJ0BSLKouLsOWls9Um7JVZmxoZtPiDWZ
WTFXtLPn1ezjdW1/+PKFYyKdk1hPqxtAq6OxxPFMpPI7B1bLfyYsFzSL1l18/Q9N
RfMej5TTEcpFfQd/kvpaVtbyI/nbbze3EwSJ57P8bwXGjQQbO0KXvsVWTpQ3MkHb
ahTk0Fg5rH9IykPsLtJZJDmNS9n0yv4GIGZO0dfWYvXj9N1Z6Yl2c9AM1ChDfBQk
ReLi9vkgKkVty7eybDkCEZ4l9x4Fina9pvfp0aND68UJpQm5EjFUfOAEW48h74U9
ixqU7nPbARv8zUJZWu8jki6bBHLpMHVnTjhrYo3ObBnyMSo46x/SNbUrtD4QNBcO
UCI49++YjjoDP52yChKOxsM/DhvNWJx2Tp0Rc323f/WfXsPSomTu/D3jrBprvNIn
iTLdQrHs5DxuzYIKcyTBbJfBwUUUpuIIV7BDP+sajFeRH9Nhq/k8aKflzlJaF8mU
O44KRPkC57h8i0onDp9uha5399V0Pfcuwpq2EeqpvaK25L9oy4dpzLlZUWnO4NTu
sWTOyaNOTSqSEjxW+zmyOfs+EI2oV/wfHE5qdNVCabPPDMxxgQ+wkIeu6uJQhCiq
cR0Lx83IQJtZaLvKppNTOQK7W27BAjvCOJBGHQDrbBGh8nSCJfvYejHqHW8R0I5/
cx5U6GS/1XvhorjXzgKXiSohI5J+PjUD5YMrY2TwMKONEJsBlyz9+HOfzdVg1fzp
rLF05nLtS5drhsoPY+rxQR7JrIYvBPGzJg49rltJli3rvWv4R85iy+Bw5g7Shec8
8Z8I1MbrR8BaY4QZteaIh8NpmwCCtbHyKJm7ZZvCoz87iePBiWy55CmKFLXPrk2t
vHEwIRVq500MJ311oQ61Wy5R4urrPZPmchnMzEblhDgfdziMHgrRUMCYAyahgYFl
OwbYg+qYTdyRnHfIgSKLtVRhDpbBsmSqnM1Eu+NQxbQwRT5JfgxQo+uQ/WiePvZT
mgKD/jewEThOd8NqaoaTMP4CejG9ZolMyM4D3tpnIfv1UEFzjHp08qCyVvtPDQgN
NFVuvwjDbjf1CNO1K+Zsp75l+nRluuXUgvvrejAr7EaRfSIVdnNfjMsJ+A3jNa5L
AHg9jwySAYZ1yuN+DoZM4zLB4bMwoV1FmRKCzpO8oi9rt2Dj21mYcUKWhOyC6e6+
3Skqvv7gsAuMa4DiXVBzfwLr2rydsATDMBG4bdUpzodPOCzw6YxSEAYEqar/NalL
aTTB0LJEqA7Kzdxw5443PcvWqmPkrx79QFOma0t1bUNbPHDfmizfmHtG60AFUlNu
xJqqvOOSJ9Bsk882eexIxwAtRbR3Uziq0dSteFgmoxeza/IfRlydD+R85nMUAPmi
yUfwQNhIFVo6nbusY4+xQmy0NsxfF8H4QNlkKxzbeJlo3nGLNqzHe6ShQ/PHC3kq
C/B5YG3Sodpg8ErfYOCK6qmkmrbXs3B9jozYpphnYXn4j6dGTq/SK5prkwoEqtYD
1wEKdMJnvH8OjShYU58Pp/OvHpkpYd+qakJvDGV37MPHgUfMhXIKo8wpxnGuRyUt
SLme30MjqIkGN4EQpkJFyZyplXxrzy+w6BoDT5qS+opgRh4k+/mb0vJq1LggeM63
zxxWuRAG1TqhaFTk2FuJQghR2DwxWuLXzadVMFfVjyI5uWkDwRv+c/H3uiu/A6hK
W2D3k+YLx8kGCPaHH2vHHRpsyTugcBGPqhVYwRgTdu8iEmX8R3JaJbJliTOBWSoC
WHRemzwu/amMxsqKP4DtVKwLO3fhe9yjXfcUlFgGHSR743jNI9RmWhU2YtoMdJPM
06uEF8TLqt7LZOHHy6IYr4OTgwGqzSc7CJzGsbZkLvkIA5ey67/q57VHUezTh84v
lSKU4wIDxx8FS4jPl7LRTYKnUbyQNDau/4SUvutrEw+bhg9KASpMb9JwmOvoPB0f
RjYE/QsJiDCc8fni+Ardo6AdHvIR77mBAfxkSJ656bHV6VtgebgrP0GfP/QCWi4a
HbOZVj4KidNQ3S/5d1FfYfYLBNMt+PIqOYPaoReUyHrqbjPN5jhfB3hlMW92Lfd4
iriLgVCSomg3RMINxDT39Z0yT+M5fqT6DvpyjBypuK/e930eCYRSX4fYEuvJqypq
zGfjNKsJB4MPCwGpx/INN1HncTGSSD1PcCBMGACe39K2NAASqIB0h+5l0TFFE8LY
TxEHPh31IjXokBZ1Ui+qcE5LSfIbFu0aCn+kA6ysGmrYO+bNytpICE53IRxAumw3
3Rt4Z+iWnTUSuQtgtenSWRidVP/XlsdDea2rBGdBjvm3OJqFSZc54ZAZra7t5pgI
hei3hAFHtDtKseUtie62WMtnJQIwDXbw6uZl6X3+8oP/Vmh3UdO2zwEZ0WF8Rf72
1BCtdQYk71l5zIBySUqUyH/9GoUf6Kwe9x9lZjVzAr4KNe/fvLfIINPzkMouSN84
/2NWrekirVUCpRi8vJSMf7qAR7CKT320mQYY9mtC7eRTIOREoEOFVo9Oe1UtwgTm
Lwxquyrr8Mwv7D1eU8udyhpmpErHdw0OGL9KhEDMp/6bRhjkKW/S6ZyvgX9XtPBd
ZfLRDTBjViw1B1X7qx2GUC7BFLazUXcO4kfx/FZaOsYkLkLiuVJe99T8ZMeRKDAN
BBmPZ/gVRJm1tgsUyFet80dnmH4HZfSaBx8l7FXsdW6wR9mxr1IN8A82cKzgyUAc
aVkO9oOP+VYhOOb2ZCkEIUnokwMost92O2gne1lgvB4zgTK+3fHix7sD7KC1d3Hz
zDyYsl35RjtT9nTat3IkFkG3FQSgCL1xtSRwOu942l4RgNcY8gR2XSkkgsVTLNRr
VOIsY18KsxSae4nIqEf7edWA90b6smffLmbQBAAze9lJp5CU8Q1m0UDyfI7RnCeR
1S/QLuQd47Fy5gN5wsdZWh682l3dpsJokwpmViqXTz1PbXAx1TPEKYcptt27Nh+G
TB4uymg8aCYIVP/zXV2KOV9JKMgzqfBaaeJT9SjjaaarMbdQ1cX1D4KAr7h0R8fm
eV6x/zPvl0ITRJFeynblwWl+RmEbiSzirwOUrxoSSgd0DaT9qjnb6fjQO4eBS6Bq
OsxLQ4F4aa/KltPB1phiZzJ79ynZsnoAKXmL9b/KotgrzoDSUzzV4lnU9HVaBs+s
sxZdYwZjPTFNFuo9yDRLfstP4zddOa06q1yK5A52tcQLCu1GiDhO5J8nOWmPk+nL
9fuzDi2jqRF1QwNstJ4Zdm9m94UD01UPmqtJCmUaSfskvzGEEXmytGr5ABo5qpo0
IK2Ib4bw0DcTsTqoerWUOTko4rDSnxwUKg6SScKiup3bkTnkeA6xUZnG6f8WfiBv
MBxm7sF//U8bzk9j1ymG3yXF7BfXmPR2EKXD/O1b44wvZjrpdLn19iD3+CC1mxR5
qhqLHPsSIbGFo8cevfslSQjxyvDrb3Lp1sQlr2prP7YR0e4nt1akKtDvgMHpI3Ud
0cf07MseFVO6vNzObwpX3wj1GxoQAchxDWnG1My0RYuXpbC/g92HP5kru9VGVz4o
u1vZDBIaoGoWYUHMYgCZfjqLmFc/MjguxA0Tv6k9QB6X+AuKxrVD1YFjhVB8Irec
umVQJn7PfX4Ey1RoT6QVPtGnJ6zRFQFmDuiNTZhPFcaAQSsHr9WuE0uYgB7/EMHc
51tdwkDnURwo/sXtKB2fOSuTTAC6y6A3jkgLCfDzRbm9ldgOHbPXCdZrMclbtM68
H18o8qTvLE8DQoy3/E77puKm7vLR7tBc2Df1B2Bf+7jYfc85ykwialXYW9PwHHpM
OLezBNgcUaAClKJ3nF2E/PZ052OAkE+FYl+JvV7xlaXFe8Y5GC8USS6VxQ0oOKSE
IkyGOJJkQIx5R5K7YVrZrUQEeMIRc5xz93FRU8f2n91k1Eb5tevmumxCD1uTP84c
94ddY6RqV7ofNFaTM6up29w4QdlFtGuG3aieLaFeAB3shpWWZwOlC183+N6qTRCo
ZULu621M9FCfK8sfbV+knTP2bLup0YPoCOhg9xkkFt2ra0FMKN7mBXW4sUMrb72X
50c9t6XtVq/Bw+rHdzIssBzLd9KS7g0cR6nZo2yZasm9L1lcRCR075aRL8gX9mrp
IcAHIAR4Ke8Tx1V63qihyAFfDcgw5reRnGMYXeXRfZEsxrQ4oa6lls1Gg8+xwqg8
SKFnaOHpKqQS8pywN1ynd9k17JgE3qzw6OtU7stghGf/zPJFmNVpRqZtQUz7qRs0
V1hri/ph5pGOvBUto4QnRbU+C3Jvaawid62Rx1apbuWU45c9gjoFLtiSr2Xr4F4l
R7uKR68/RukzCC6l/s/swVDt+jRVuNLnMtmUOTU5T03PXQvNhnqZL9vGdgyPU0XC
LxtqyoLjNmIDlPnG4obD/1zdVCM0TE5MsFMX31kgXD5uzxqiUo2nSlF8zWa5lVM1
OXmsx75icd/WFF59/vngVrUUPuMxSVFfZ93jXeK/Gs1YfnPqqW4Bck1mdKJixxl2
PIFbR8mbNnB3nUDVPoydF0CjLjbFRp7xlI2xsgDDUPzk+YdkYc77vP1ISeeK8Vrg
I5eWpTKhjc7XyNmCAnyObQhDfVTqGr6FAkc/H2794SFP1C5Vg935DcP51dN4boKU
xdja16QHOOTBVc/Gm8SBlWRkdHpx7PfO7NuCnogBSr66djJQkrpxHQCHl+7b+Ik6
bdXurp+yRTvpZcY29cpQuuWI300Hy7ylhWtWwWnIT+YU1du7cDeZt3XDHEZdRmHm
h9afjeTxdhlGHKTLJWYD9VJ0YNJEsjbFzd+yB6UPOglO+Rcbphtxng7jagGIz2TZ
rfJvc7FuUi6CEfz5/aHC8NADR8UwzVtphBhFUC+MpLIhHkj7uVSFwpMDPG+RA9Jz
FW/tUnN0PXAwNXVXy8Nk2jduAiDgih6Vc+O55o6n0tiiya+mT7NJIvLhfV1D1F8H
PdUPFyQFteThxrbDWTAPd0TpwuwVkyVbfxba9o7nc5U83K0JVP2hhymVpxaEJLI8
qwY4rK09lCDrpVoKl2aNf6euu8dmFpkcslsHJtMGJMklr139Xs21Ci3ckTwKv/f3
Uln+EJcUlikZK0+pn2stFSNuQjO0XfrgyJvFfnZhRpa8ycnLpmB3KLOmRSPrzlAC
gXfrTSqhUOecgzwMG8w2unsLZuNLgye6OLzBJhpdOtapI3CtWTIofhtHaEVm60iz
9fQ0335J6z5PAZgxaBPy4iLISomvXh/ME5/2FVD8n1jIJ4XNuR6J/p8UWJbSDFPk
KAWthi2JIipH31OndSTIx3yCg4EblKCGJ2j/mROPobKOUSF4lgYZbbfrRteKcIqL
DoI4x2M8s4T32xEzvAQKhl7WzYizu6PW/x8iLQ9MIFrTnmFpvBc9G9VbZnrecy/j
qeCi//V7C+0ip9u0ubZK/6zuRU9mwcit1d5dse5EgB8I76+K93dI3nKpkon690Tg
hyHqAPiTHHm+odD+qOS5nWSjZkuLMIgE08VGU3452Lqr0gb9CZmFHaymmwmaVCp8
w++3cWrjCbv3tvmy8ociaWx74C6K8IxKjtxl+jlyQ7nhJbG9U0v9M0QupYrIznNK
PYR6AgETlVQvgquQNg57KTB7C1dbm5dvu/RDqEwuYJWVBbMpz9Tgx4jsfy38v46r
RIczpxP74woOGuE1tbwAjws0DcPNYszXLna2jL4eATw6s3dlYaXmX5zr+RnKEcZn
Akvjw5A6HR3zkhtkJeAWdsQsDocNwv8TvP3bsCI6tp5q7NZGe+X+pwQ73zBsT5jf
YDPT7sYPQNR2ifKYkOu3rkHh0EXt6QoXWdhhucERI3KEUWN8cBHJOHFAz+7ZVVPU
rjdpsCxz44r77yO26Ahx1nInobhALNtWniRJUTTwIHb8SjxAtu+ymlj5OoQuehF5
FIHcRNPCCkT9NqEUdTj7N3fPCobLkknYucCCmKqovn5Jb8ISQ+W/bZcdxtg00alK
rd6UXWHI2u9nuPMNIEbMWKQCzJBx9RioOKqQGRtmAOYh7YyQowAb2Ix8uOqJwIpx
LmJojdtXE7IekYifL/ElSeKz4ArmgiK2Sixbed3+OllatjP0AlpPx6LvAOdZJNrH
KQi54n7d0CUGBNesd0ANHhYIz2PR+suW4yYRACAhbOgltN0flmTwplBPyQl/T9g9
EQDz3P9E2sbbotasmZcswTNykgCmNrirJKrWDA60pUvU56fKlv7F9RhE9U3ZzC3u
GuditWHAbBdavM/Y8UdjBxtNRjjuJI1A//DXQCyVveAw3CCuo8KeaAGLGmwf7xg+
5BhbY4nsaJNNJOq5p+oGkopvdLztUd9RLvqks6QcyxS25fVFqXqjl4tI0yUdONoV
yohZKyD+R9OKZpH2t6alCAA6PcZfG8EnsYOOWycVmHbs/7IP4UcISbXPZThTBwiu
1/DHbTr0FQvBi/83VjEy/8RG7uIt3kllv+5UnarHJtNM+1XQUeKPIHbsFIQHH4lO
Z8iovC7DMXqH+2B56IwW7AcSQKZBWCFbwhhbGibCrh4DER1wbmEBGQA6npTrNBQX
c4jCvSrhZfPzYNHIPpvZ2xg3cEln0D+jx5V6H5m8mh5peh5Ngzdn/DlumiD1ijLn
0aeEgklnv4ldFW5mg4ZLKbGGjAaxLfr+svmamCi4+zbe2v4N+ns+X6xGFFLaVSfx
1jiyDy59GkIbUVhZobU8pZ2pVEPQp0Sk0YAJ+cxKZhZhLsaS8Hl3bIzS6gHEqoPH
2F+fx5I+1hc6LPC7hcFdBVeWj3116OO4xkON6pQh/Mu8/CsoN07lPIqPIWxboKoV
fkipKfj1IT9QPAJcSNWr7tcSfD50fjcHTPGQ/P7c/y7/vxySfQslq5ebGjo98cCL
8UwWJ4dYqDxknCUVXpZ/CAZJMfgSRYxdNQeRkB950bMv0b2bIamTsXfySJBcVj44
TJABzVclcQx4O4EZUZ7FhzQY9Om9T1ZHC4COdR4cApTkFbYIkDLRasHkg6wJsTTJ
vFJ+rRxeP+lkRtgT5Z/GGfUdtGEB4HnDC9X6b2dOOTLS6OTIcvdpWwt1xCFOCaGi
yI2gclo0kcIryWcgerL/g5sm+pqsew3QkuEKTREm1D097hDh3hj90o5wYNryvZoy
HoNaxi7IdoQzVi44CxGEY3VdmcJmm89BCYn5SlRm7TTqfqaWJEBl/qeAOHEh15pw
h3vJoTSLu6LBEoS6m/VeuVN5WsHmA7SswuMYib9VeGMp8zEOobHfGQn0mV0vivbt
DsIvakSPJNTgjHN33nRTCWh/cosJ55aWv/RjWjbXFNni20uYpfs4E1Dyo2q75uGE
dm6U9r2bH3fkwGtxwql6Gn+9m6DdPCDV/xtMuDck6bmsgsP1epxzESl7aMmI+E3t
UkBMxUlqokYZB/QLxXQ++iUYVKhR30sZpU046dFjuH67kUZFgkzlbNy51XJ94BGp
gnCFxIFrgdJBiJeyTGJHdtpSFUcrrtyIvs0AQqVKF1mD01gvg8ZBBqHTETOz53ac
Ji78W6ZdOOiQxALyJvCSOeyiKSTcmd/XjGGVUg3HejyjAFriplVD7v0FthpPYj8X
hk/m0/SzQqbD3siw7hZp+GuHY8vevFN7h4nGbFKY1fMaOkGs6sS9BbbCf+oZnwsE
Qfz9BDaJgrs38AjRSoD3mI+9TUHkorCFBJjYkuJdhASlRFB4UC9QXRhLhlWV6W4Q
yUBSIpfxAEWDGptalBTV02Buuf0BX+K6gFkmCvmPwGqSfmq6h3h0j6Ase9I5dK+D
3S+DWbO44ed8bD32W0lv9CahzjZK+n4iPrXkFGnYTofkcElkAb1CJ+X7ETpdbVyN
KGAqiUTuNlVJheW+g0dyKvsCn3JnWNdYcH0fnzlDgXB5hEvDJ2VyBNnxn961kTuS
CGZjDlBJBKco8Vnj5VTrNJcCRA/HVCBJ51UrF9+YCjVAGkHcBG+2nHoyR08KHgrC
IiE+KgIVZ7aSghY8P1bnGB+EZE+3cQSOZTzAzV7kLNsRSwi7WLNtij4j0/MgCn/p
t5MOtggjnHNsDDI67qXiU5wEk2HNye7feftW/xDAZ1JQ3AHE/nKAvyUJXgh2X2m9
aqJcY1JstLwnGe/Lm9USwgw6UT2pXAsao5FUB1AmyiAW9Ff6LYlprFKR19a0lLyL
h04m+m37w00CukezVwyhzQCa/F6oyk26G0O0QNSkTTNSFmkKSSzz+pzfevIywb3a
78O8SIMtoqIxD+YpyOGGZ4pVEyP5BG6gcMWbmCLosf0EkAY87iy4iB/aWXUi607n
YVcBwIjlxBTzyvQHHgdo/5NhKfkVmAcMCjfaVUPpR2mo5XNzhv3eXhxh6l9jfAIc
IBVIxzYBwkeylDe88/0ewMLCrQChkw7sFQnOoBjLvrZbWkDIefe+Uc3lh89hLikN
+0on+80Zc4FXjIjB3wM2fyb12MabXVp83+Gf2VZAdQXLyw+vLyYEewJHr85H0qBf
pFmyAqojTvNvdE9dN/qWiYSAog22UzdjEBMrmgg82tWfVbVHwyTC7ne32iv+HNUg
1NcJFo6rjQs96UTHwPI7OZfhZ1S4Z2eRaeigzIMqBZqIM0WttN8/u3bCrtkLwlw5
9IT2GGVrf3XObYrTLTetVyM72ZmG/sNVXrPdE4gerM67qXKGI0QnQ+3nS4DNiBWS
KG7zXIZDxWVELM0uhazbmaT9E13IR3j5AG8ZkfgaIcYPICQeyqXBXp0XbIHWY5RD
i+Sl3Jsk9PFGdE+mpP5nDI9DAkwTU1JWOVufYbqwQtir6xr86OoAfcI1z/Rn75+S
cFptjRU8ssJJVNrr7g5IN1Gim4zdWiI7+OCiKB8dRK0OzvKC3EgEUeCW7noFfaRp
PagGwXK8gOG58Cu1jSIaj2qnNTJ+9MP0GZExlhxqyL2TY8PVMQbmWyXnsd2+tr7x
6/vUvBAPQsotEcnDSicQb36ot3sr8NIKCHTxmXHe+n6UjcCB7/ocQEi1iMZ1x6dF
4M2XOjv9CpE9dFyaZwpD+nxajZ9+aIV2+B3c8BEvZHaFZJo7bjEUikjbDpGzE7VB
XbSoW+mFlolx3lmXlKPs3NIAx+OUTE8Q6fLGGC6v3zoRsnrh/l6Fd6g2ks+mdbR6
vNg8mNtXfhU/4RZ2U0uHGSl8yh10TDBDCxvkMnEdj6fdxOVsUpYm/uGQ3O14T2Zj
Ojcnvfs5fv4FzoWqZ88QwymprXu59FacgEkUXh4dvFN6r/cqz9+9L+tb2XheYjYg
UKOtEUbU1vMdMHnRxxLdp6GNPE6+le7gSpIMbtroV4ut6Nz17f+9BwJTi/lZyaWn
v+5oyxpfZIOb1DBFKKWKkwjr+xLvBsnTaxf5s9OJyUZ7yUWDEMmJNtGdbAKSFLsh
O6u1W57GpoHOXeFxfMpTWWavPbMZ05KJEYwOlYzBegpQZ7feVtb9Qn0/Of6vXuTl
XcyKzEI87f/DgFUCZ1epcHPbThOdUkt+SfaS95pTfvuY2MMXWVjkkQCAP6Epfag0
RKaUrnWfGuSbnFciVrwcIVvNK2fQjnqtV9u2o2UVeziRa/XHFzq7xDlnyVdAvEW/
cDiEBjcKZwT3CDkzPj6t+2diFi3JCPFK0fVpzoEaA7yJoOuDkpXOV51elRbFmDUC
WTWnM0Sh3mp9ynjG71p22P98pXYyHvNgTJTuCfdnkfEzCPYTVBYx4XlzRXOqgbdv
JwQk5qdEyLG/dMSUQNVPS56ce5rzR4aF5pBVlOAKCLZOp32+EzZM7NtzOmZ7+05+
mCBGCGzPu47AWTolNAa15JgGhA12ZcE0+RcR+Duv+a3IrhUQdHYg6r2KyC6WIv5E
kSbGhi/6ar6ekn3/clRV8sbzFd9LcxBGBHswiQGA9SaZEzdl9CBarT6KWs75S0tS
IrEQ1hcUpWhZMFVEokb6vBJ9HiVAadoHE1niEBC6VjY6vPYr49LSf2wZbvHzrTwf
/2m8695JSKPJcA5Ic3Zcs20LKBfE6f/WZLuCcKvHgGI10j4hQYHGI++mbghuZEPj
Voefo/HuMsrMaf7VUzl4Y0h63V6E4orLofRZGpEq5yMFNxYDqKBuNrHvFTQ/QJxB
Me65vE3I4QNSeH7jYCE+SopNTDyXfN47xvzAqgYNwd/R0PpfnBovLwRXNRjVCRKo
HQSiFXeDjSypvReJG8JrZzHiyDdOr0A8uCewsS+NVamde2JXuH3a1Dicy94zDq+S
fpR4Mk6MjV41ptv04fgv1eEdnPEnULjIjUe8oVYxW7dSTUyrR60NeksvdBpDZmdG
DLslrNm14WM/CGoWQgo4zdZJbt2H7tRrzK2EvlIt2Y0m7AmREZjuQNfEYHmLBMHM
LIeLQgAR8O7ZNCLpM+4JHShSk9tDxa8CdzvSP9cUJkA9GZsn8I1L1ez+gUjbtlsB
sPXnOH7XOOeoE/ItD2U1KXZ7xE+D7Z8X4jsXy0/EIZ/pOvBw7sq2ummO/fZ9+t4X
vTTn9XkUV1dVnj22NOGlCBW6/5gqyP4tLYGIf/LDqGAki6xVh4h5zI7RJfDb8hnP
gPKN9CZxdmxqYl3AyRlzRH8xWhQ+j5+MqFfSpaGWR8xj2dPpRFapnwR+669KDTcH
a5apbtZGRtkGKVPqFDRb4mxVgAZutQWm1I/BQs0RD4kosBUuLrqFi8EGSZqqdMaE
Y5p91mEKwDxcmTrXXz/bY07N8WEBSR/XL99z5qGUIfZb0pLBdxdaTuEkgTEk5Zrq
7thOyl9MQZoLwrmG7gcGytp//ek36cHpCH3Wb8olU1Bpj5+kp6dsDpXenqpE46Rd
vdU8Xw3vKM2VdbaXG7NHh+zWqFKS5fYYZf1jyAaEVdsdZ6m7q+hlwC34c8cK8y8F
QV/7HOc6L7kz1OVrdY/p+nHRGL1QqNAmHqD4b/Ej6OYBwSYI1F/f1d2hXeUiB9pw
9uScTw4HdT0krxfQ1HbCdUHRrdMMqByoP8HBuIjJQmSiH7STaBkGNcQmYN7rZ+N3
1JK4S2Tss8YNyhuikjKC9DLsK2OBs98qbEksZubohtNK1GNKFe0S0JwOo5hvYnuB
qFWvEF3Uo2Po4mDcZts2/iHTHteIceyXTkp3iUXh33fa+Y1RLcxVA5SU9cEXrK+y
zyoCt6xoSPMrxW8JV80O+ZTbGVTGaEdrSFwId0y42uahKbAcwemwkUYupJVZQi+I
CQXLndZewx1LCLRkeYuuJNxAzkmAYaA4+YIPAF/iBYHTQmQ1TqkpsEJaZaAOW5lq
Hpro4f2O/Bj6pSdRWjTml9rM8Z9HXVstsvMOdfOZWmTlKVRUrl03J+Wd4zts7rr1
txw29ACzYMkdkszo6M2mWDEtJEpsuRl1YWoJrJhSxl2ESDKbTEya3fElRFMnivdZ
urd6QVa5MsVAOHrOzSxIMRSxgBhmWX59pCJyRUnt11uBpnHDA5NpDPlC+kc34wUD
7Uq6mtKTGnJ/eDRgzlC41cupAfYdYyNrowXOBWj89kYHf+++GPp9tnHr3lsqXdRd
npzqFYGSsJod2elx0v66FWvqqDXNpm1ECb15693li1Kwt9FFcR41QucFc9uiDM4R
6UX3KV1AzfOP+kfVNC5tWEyEE2I7G8dmie5ijLXcXNVnB3UwWf8cV/58EnICdgef
2aKQATRiMthKHUUU/VmbvrxpLiqRQx6V0YXQJBrDeyWSe+YgKpRKY0PsUBZl1msL
ESzA/1rwFczJ8GCMelHNJO/vJi0XK0A9RcJhtqBINpDvqXEWsMG/Rid/I/V4nDMS
Ypv5fN4ux/QfWgE4R899f7/ePs0bwKxMVh8kFivnvyaf3BpO9pkUI8cyrHGROmYu
dKp1neDkM6RB6tdNYtFRV5qt+tjphK9jsTHUvghq5lot64Y7mKn6SHNm8FfBYnA1
DQ8S2XFB1azTYGAhLCcEg10isevUxeGFaCUHb48s6Tc49ceMbyQxjqYhhB8CmMJp
/t7c6oSr/vqbeF9fxCw5v0WzHKT+MK1ej7Uh/YL+2Nb93QKLz4BCPx1Khn51Lupk
EhIp0+eo+NmzlARNh7N6cqs8S6dzl+zma+lM/Q5MlXSc/zaKClrhaW5l7JVNGtf2
cISWL7UeaC4yQIb5TRoEafTJBDW+VJiIsO3P4q1Ky1RSl41BfEn2NWU9poCw+0SB
74dQSrgLmhA1+CRxn3vLqIsI4g5rAfWQ33Foaq2P0+nXQNXYo9u5OGDF6phUd22Y
YtGIrJ/tslAXLfVhg5Uflyp0+KB1KxxluJsZZztdTCZp97nnq05NxCOdnXZiarE8
73c/Y426fYwNQ1whiwuJzwWYImDU+DHETEkLJjvpV3x+T8Egr84LYsA06/WThCEL
Idxfwg7kXWtBNAv9fgDvxsIYl8H3wITW5YlgcewXizDFEFv7eKuuzG4MQ+ms5VJj
9151nJ8Xiprb1x2soO6c3HORqCYeYZUpSCjobZTy+x9OQiruKdJ94OLaTaJuHbuJ
5Dsd/M+LsL4KwjKmHhpZG9SckKo+fPWHCvxyS5Lxg6sdb+msB9to7opvlmA1E9ip
ZF6CekKpcNAHgx6v77m0yDX/zfN210twKHBi4O4Hdr+fkKhBEhylgUniLyy9zBxf
S3C0Y819bVWogygNR6YAopJPSO63IrNe8zUtkQrzY/8Ic0HVoQpbaZ9D3oZiPY5j
E6jDMpVj9pt+QzAfRXlfXFuIDaC+tmlC3zs9JC4NITUiqvNa55vImFMq/oQD1o7B
E/5yPZG9nliM8lD6rmnCOhhFdVXomMKZhzCnkGQ/8OuYTgR8REcHDkW5nKWii9xb
yWcmYkofXhV7embtm8UqZDoP1sSFZn3kyNdceYTxlUk3+zUi8EwzCu/+11rnS1yM
Fy5N1eD9GBYEKd+w9UfdN5tpu554eWH52bI8PKJx8qiwg7t8od5f/e3GYDY7b5kK
x6dGehSvutKGgnUzc94MF65faZwpJtt+EMlb6TGq9/ojEhvMusONJ/u2HIXSFoyg
5dwM1oYYGv5hlRw2ApkdJY4xI3Wl+MWtHGjP38qXDZIqctqE+dXIk9o9j/QbUnMy
BJVbfGSvngXdVPpUzqgxPFFhYJhF7d086WCwZHTz7MptDorY0UpiYZ7Kj7pfocAt
VRDIDlr0uCH69FkLRQVnkJkee7ZlQxSnX7Maw2/JU/nhZDuTduLzew4K+9A+ybKe
hnIJ0Or2+dPxzFVY3/x/tupk/JChluv1s2vFlY9uPZKN9OTI0J1g3NqWWy57qrzb
UgOUQIxIHP2IYshLbJmK7hLJHlPwcLleOdKqCsI85WOB/jFAUEQOYej6P9tchRRg
BqDlutDh8F6GjUh9dJGMiQ4F7KsKl1qpPe579+Kq1L5XED26ANUsQr+ej6CuWpYA
9/jqBcEXwqDP2yCu1elamnBdSzIAsBQ1DmXne7r3o0RdiBZvlb74yC8MxrpI04mP
zbfvYZg8PJMmZnWj9VwVs92VCELCnT4wmbA4hFXuIha28XI9+W3GhyizS1rgtezW
Bk94UBZvwkUPMlcvEQ/zwHghOQM2y4FnpC3z35AfqJAd8PJ3qIerp08kOIBuYtMW
fkfg4msTbcg2uGY53RxuzFYdhz6nyubRlKj/Is6bzoCAxRAC+/BmUOTvrF+i3lGQ
WSCFiNN7vxMn8iXMIcWP+tQOqCD2x78spI9gLFh1swoBYh952cYIQMXHaOuigz7u
l0TGSxpVXmIv6fUSG/teWQGKSQmNba3gTDxJ8w9v7axDdgrTH80x0cdz66RDnvzi
zo15q1EDFo0nb3l8/lHh6U2FXr3GZmkMVgrWQ9/LgDTFZAjAy6VAMdFnK6ZUn1/E
aniLBhdfqq8sAzaC38wj5vYIIwehHVsDVSRDnaK2Enr6IihcGe+YBK/tRJZKQscE
hvhHnX9nqm8LXQsTOzvIz6HXR83+qCC9jRsKvPJDi1Oq4Uk+2ATNKCOCqn6fNj6P
8ntlQhzq4f8th7phwFMPmdytg5TiAtiC157ITESpGbuypnq0piMXQB0HTyse83TE
8XNNkaEY4A1SvGlPmx+y2uWOo4kIa6VqVIrwdrqclNaZeLRkIHGsZlsrYB/MUS45
vs0KjKWzRxW5BNYMCrP17DuxljmswtDuVpGRqgQ+IcXpBtEc9rMxfd5V3fhjGJ9n
JK7T1A/sY6zxnWtkWJ6yIv7WxLOqvSyJ7GLpd5/+xBFrakjxvzhLzOLmK0Kyubzh
EkcfB+5lJYsjeipuCKZTBHpmp1KYBky7ziDbWTUTPtbLFSZK/pR8dLti6wuc1ZEt
vlhX9ppZ72if5akhHehoDfggwhy5E1COmtGV/At3y3hpOLlDqFKuCXGko2RTK61e
okj0HkesM/ypvyCpREe+/X+mw43fncgAcUSfaa+MgnPMr6Wz8pCUMbVVSq8f5Iw8
jkX17JZRFxoejROtt4RKdKUI7QPhfa8WdPWWAtr0/gNuU88EL2v+p9BqkECqU3IP
/sySdu31rw7LpJgwKWEkQ+4hqgYFgTSODiHTxMq6KH8o79jyTZ2Zc+MCtdWQ/xVn
hdfNQoxqQSJjmsu3e90Jo8IuAqCI3ncvJjkhGGnN7cw+KeE/z7noH9/mAJmXecG9
zGEDrwD7d4M8GqKJcZK/QxJPGDSm3MzOOTNLTVfxw5ZoPVPU/hzOmUuqJHyBcduN
Y3RqwsevafpxUJGKpjuhK0qY4vq9nTh4VrLljvrEbiev8yEWwNCrEvrwO4TrG8iI
G26555+ln2uRjjKP0ocVCQ04i8Z2MhsU6j4R6wpRmX+cd/yfmRN4ztOdtgdk+stH
bmiXD+TfSxGSnFMi/yq27fKcmmbdPmIEpash8AbK2AxgUUMqDUkkBqMboWMoKyRI
26ePbap5iCD2oFXRf8nOlVu7LdERipp2IaxnyrE4TFSh4Rb0tqQUFYi9hpgYOS5O
Fd52U7zbOyg+mSLNtmbFfZgq5WpYy7vw4sPOl5xdjsCW51Db3wpTfEP2yVTTGL1e
fwfvYEMDfMe2dy4hN3swJxsRxQBrY5wJ417dBjpdJA+I20WMrV1pgdNdNj9D0ZoF
Acddk92R5Z4kFmYYvZF9CUJH2DjVDhHMKzvgx2O1Kwtm0L6eZ3Cw+ui/j0rI3NQ5
5tbwnuMQeIOj7KsX3Q0tTXoVZR9EodcUoVAFrNbcfhVSo8V9AEwhmL7GIGf7bzr8
3kVe9zoL+3jvzE7Zkgngrq2RawC4qwIBtaE+UqXrwVPiQDPpgIbSSqAops9zqnPZ
quyKG89HOtsPLI2+72J5uWCknxbbcg54fX9CbF65RG5rjpXBdOa1ham9atcunqxp
0HpyKuT1deIc2tqtMA490euCeRWklRuDh2kxO6cbnCoSqHoxEjdYpsDE8GkE1vbf
DrsmUvE6N3c6XE+fM2kQpn1Ho7Y33E+9/jnyMn0amE07MqMDJk3G7ZKqUwBUL11K
YH1PCdGUXyFD6wMY9mD2uFWufItOJOttya0v6h1Wv01I7vwKSgXFrsBSCvH15x/0
tfNbo58fStMacO6ViTEKzjFTLYAA6QvQZf8OtFIG0GSJcpWdMo5UXPU3vA9aFRRq
xRb9knzSrbUomRcKjbP3AjQ1ruzeWibVbNm73LJceD2wFpAEi4ZOTNMA+ia5RnmX
5jR8N4dist0PaGaNb9eclVv4wPFp5QBt/QF4lBIFru8rlVxCqC5LS0HH7nDt3FsU
wp9jK6paUPphskfxS9cLk3QcNPOnHiGZJ+NesgRKtb1bBOqd4LZKz4p4atZR9EHv
YIQsqz8y6Oh7+Ulcz8GfJMMFoipGDRzBhWVtt5sxoZMRZjVeYesMhDmvtZxRg3ib
2bvC5zzd6yBt2XKOWsboaQyT4ktl+vfaMi4eP10J4kti2RawJWkBMLbAL3ScuRB3
icIT72GUhp5aMdLQBTFOaKgmtR9Ryr6oj0HkGm13Z+O6Opoh8FV3YHUD5+qQ7qas
sr9hGI9DNPdzVTdDkH34OaQVBSWP0M8djDQO7e+rl3T5VcbBYWpcnB6p4IWA5Hzx
FIVr9GZjKAFhhzh+K9Z2m89jYbQIsVrrUDP70JOqn+ivLgarRijriYcvd3oY1Sz9
KriqyRySNW5ulPFrA0tQRa8EAsJYfEUOpC/2IqufzkEo8B3mLCDVNfZ85TOUzxib
z8tHDqDHpEythGP0QJcg/p89yHHwxxlgB2k2Ijh3xi9agem7yLdRkYKuEftc4F4V
CGadHxut55FP9hpliBOBHKFqnYYJJ93G7nZJ3UYq8VYdEDVOAEGa/CJ/9O+1jX+v
9X8Ci0zVKyEXMmHgezgIAh7HEeqmLnTyD0svVtqXATLWW9rSLWWn79tCpgQOYkGi
kYAUO6TLFgeSkYO/9xqkdTUXna8rGU6Q+bsoYnbWDCgc1untWlj0naF3/JK0u7CW
NQkfw6+B++XbwX1cKrNzA4+A5imJLScVmRSZzKsS9vo2tVdNNw+ELqcI5uLQUn/8
vwscMLJwLJqhJdqztzTYTz80WxFBRHwtsIf5/UkpbBjHqhXVxwLTjK6m9ZkvOLo6
RAXD/fBWzwwZzogcmFlVvPiMKYwucgikbgcdzB+oMcyAKEhr59XDv76yn5G4hGNU
4vfcIpYdaoOn9UTxFIJ9JFg1mFMiDIqGEayowOegk0MaCg3KEaFLvYeM3Nwv4dG3
/THttBzB43ImRYPlHnNPWoRu8JxEp78pkMJTlFz1ilpv6uAw/zEwSoxr7a+zzZdm
iXPkJUifrBkbnej3jEyXsJPl/YUAFVYCX/9Uu0uw/4KpeyJcIq8jnkv43ib1sNGE
qD9ozKRhaVzCZ+vjvqrMevAnCOl2BXs+SxxlcxQ7B2qI4PLZl97gSnC5ucZVOfOw
KV6+YMauWb/4XW5UNWnz6p3u3gBCvshJ2TGlCSKgrYnOlGeh4w+EITdKNSbV6DlS
nQqqxIM/MYFugolWbmgeyV/6Vt7qtnJgLQYYcLrceiHnuhFa9Os9/r1prUkIv6Xi
JYahBzme3IPMRomGi9pycEjgsZM9f4Qfqz1QhBUt+I0JXBcVPkIhqi8HFb5Gj6iB
ziDiN+QhczZvgvqazTj8biWHbwVhIHLIcBkUbCP61klQa3b4T32KzuRt40xPp1aH
qNk7kOgzM7GfGH9ROdpXO1iBnGeoFQ06XdWPzWVwmaTkaSqsgSRhRfNakywKT+8M
ZbAR5wERXtKeIZJlO8Awd4vPjNfFvxuKKoh7GSJ7+ZoxLqVRJExi5vGTYSgmEwaQ
tuNhLN0yQgjci7wNHdZhxo+mV5n0c08e56KQiFWY+xOUPRdKpnXH5W6gdPYWktq8
m0XfUPO/Qn2fExukRXJAWC5XxBeERW/IOIzIPTapg5H0nqBNpYCK1uTJPbrqIDpr
mZJZn1pt2fLF4fjx8Gy7MgvBIBJvIsFYvYTdW960wWWv0UtqnMIjI4suEICSQSym
f0I5bE/feYgiDwEiYXgD9tpW3Xj/TbR/rS0qk0sUZ2w030jiW3OntewuO0Jsdqst
NGcsNzgPufi47MxF8NijvT0coxPJ+FyGj61pQ30W7u6G5zPzU5wD2KN9nvdPluhi
8ySDuNRvZASfjMQSBQ3jRvOszQCvD4SadEXZSgEkS4KVn9ZDEzrKKDDiATEud2Q/
RiKb7gkJk8EE1NLqpQgfDSOQnrbCE58um8j/l1p7F8enTU4A0DyQg3cxXA3WU3sv
q+Qul3zwu5lGFg0FLVTxwpk4exaMp3gIvo3CvsrYUCZn586vY5yHKCBS2IerlH/9
dnA+ZT/pPKTyr2rWo43ILp7BHyQWUUh+eoIFepH9yz/0OcVGw5XsEhjz1IHP4Y1z
c0JvH9dAeceqO08b90ipTRSiw8BPCU6UTX2DcnMsWNvDRGxo5901nJQ0apRXclgX
lKKXfeWST6ezUqY+yZZRqHXevaUnhulJQAojhhH0DlAJkfSSCjSDEeA+ie0A4QVR
IOBRBvIcosdBgUPg8kjQz2bnRHLKE4lwWixLydEcvPKXtey5rijj2fM8Ss2dSTaX
PJCm4yMHcHdTeVr/HFoyaULXoupopAgj4Gw1CGjiy/FiQbz0n3XGBjtIaBXUtSa3
O8e+GmG3kNoywWJsriTZKWd80jpRwq+3dzJWM3jbpWN4XB2qxTyH0EGQ93iVuwCo
236TKc6Tf5I/wTUh0xa+9y7U9OCPbslwp5rHv5IC1Uh1aAwlVCYhntk8EneG6oMh
Us8bEaDqeAFPxvlwkkReUrZ5Gz+b7k5IVkTCzZFaAf0DbeKQD4FSfGT1K4zidzLZ
gbr5jILO7OiL+rHbee0M5kELmkauV7MC4kaAIQJnjLHIVbZ7ngAikmWvjor7Ampi
Ehr7jwKrfSNemSVVmaRnMWssM7wwAT8vwdrR0Xz7wm8M8OLTGaZGQm77GyEARlXA
BGf4UhTtzIbeik8/0tBVTbfn3nPL8PpxBDPu20+qNaNmJIACbL9mGZ8ObfZ1LdYP
dHVe3sXpai4ODZIt36vz5lqfQcW8FfEuQ5AT+lc6Wb3SuWCce2J7Jlicqg4FjrDs
fqWdSVtSvA7re/8/JgmRd+7CCBTdkMhpNCGR7eywUjNj2JyhiwKzrav/zC0QEQ8z
1FY7FAcqDcUe1x6RInkKO8P9HPjb1swTncnvLOKWQ1cEL8YdCVEB1oRgZO9QqzIZ
z+VJBUYioSsxXekke+AlnPThjXENM+P0MtcdMQ3O5NbVAjtvv4QCelk1lDTpcVWw
0/cPYMLHeBCxGYLXhrjAxLYrnASBIkvK5KhG25ra0Wh5HG6+RDC/mKnhzTa/hc43
5WhdXKpNQouY+gRpF6yuv+mXGMQyGkZh+et+NpTMF6BccfwwF/8j+sBHhv4PuM4o
Ohc6GCJCEv9q5vkuKinZA962P2oA1ckXoe+heiwuhpj+DB71CHoEvU/ZrS3k6MIa
MoAmulJ5UKPkwrpmHzgeDz/s80tQPXAzUzfI3qgyuPY1vkoc42Xa5QTwOmEXscdV
y3uPcJYvJA/M6EA71oi3pjWdm8sq3oS1poAtLevYAwNB3WddDDsNLKvVueOmSBt7
HDqSSqFkZ0xpKjzvdtwvxANQHbKGNhcL90uO5OVM7t17dady49FFTneQvKGUtu9g
wntg62TcVuG5tnSTeVR6K75tpKofRLMIqArEyrthgKk9Wd/UrB8s58CRUaHEgdHW
TkJ7joX7AuYqd4m79NBp8D6uCgEvDRw3ENAyY63gER5YiU1LWBRHRyGAUSo4iM6U
1asCB9KY9Ts40/KSS45d6gaASi9vv+V9oqvKvb4aQzWDeI1rgSu5lxHxyWU4l2c7
+QBIK5VVem8UtYBFoTCP587i84I+yBV9ui6IYNp5xlM24NwM5HZBEKaH8us4otIP
pVook9wwzCQWwSbWFan9DTiCoMr9++rQ46Ag/Hc4I93PhsSNdVUk5RnyBsqknnmh
p+sc4ap36eFasK2bPKlUGvUmIvDdep+9n6NDt4LfXfvrAv7zoHpO8njb53K7mW5E
qgXoR4I+QhaeYGPSoNcT1ZK3zxVzVNrBDrSyD4MuY/M7lkD3nPdaArzkp5GZPxHT
mtGvc3Li7ye5E2kyERkhNyLvKYqw040puHiY6ewoy+HG+XyBi9e+iGMO5V4eaks0
Oe2FQz0fch1N4Rh06rnm/5ToV6NsUbg72ujzX1K8OVijS/00IfZHphxDW0MNgiwN
eoCG6ptOKBzqjzwP3iPlIttp7NFsXjoO9+nU8XyrUjr/v0SbaXzCCO3PQ3DZAW0e
QoIu1TKF+VIUUkGxdMhZO2bulGNfpv624dIHtOqHVNMRnCs7JqjBQ6Q++eqRVrcZ
grdg+1/3bMIlkNrPmYhxtdciDB8yVSrT3ZNUaqqAqzPocSbULM1HNlPVPYrBsceG
4hkErf6pyEg5EV8rFmHZZ8LiSBxmHr/HsvjQqxpPHiP8Gx06tZuHj2QnwVYxgr1K
AmQoxgtdUXOU4bI5HRphiuV8QPvOeqnrvIlqx86Ahi3ICGUnJxW8lIGzEJYaGSqQ
ZnGc2zk/4HWCB9hAUiCxUrjxkxnOMcsL6zkBXNLIMWoP3jIDpo1nn9mS25ms/w+Z
7dJN9HaSi+Yo+3wUZRP/vZmZLUQIKHRFnZwCZPJXsCtMNnCLF+a7h+yra6ND4AGr
rUDZ5nZaWDiGjeP35Ji1LSxdtHfFoIP8X2UdH7UhI1kRsWh3p82mghPoVpI7NrK1
aklBm6TXvCuE+HjVcDkdJmpiAdUFMu5Trt/X7CHxTnA7vgMZkmryHxRxqDmUjU7V
gUWdTi8Znixhfxw5JMqK0DWQu6GmtE57NMYZIBLPvyEgJ6yqnQndZfGNjaXLnyxy
T95dDYPdRulLQWSZiHhInsDv8LceklLN5OzAdx5jQ2qoQfj2jF4WCICXmHJhXQip
zIlTLFuuLMrb8M9+tJcGIZjvJTqvEoQ5b1Ta6HCCi8pwMXvtJq6QvBbwdSykHxgF
8votyAfu9TJVGnzxCjtrEUPICSrvFZGK/CVS0MhuEHmt3tJ5N2VXxjufQPAkEW5y
Sn6sKcijkdVDrL7wYEAdciE2/4Es728nyWmrE31blxzG4X1mXfFIwtjJfs5LRUbz
pE+MZrPAT8A6FLkxNTXr9F7hMJYwDNYcqeG0KWpJujIh2V92pnp/ZXPlCbVY0HnH
HTbv6cud2VgwLbqaGt9piFqbtkWKsDLXgW2lXq6zsQLi7vLmmqwTDMln99OX9iRa
MqM49xrXvhb6q0yyS6jmdofcRXnYOVAeB3Ys/ySPYDeUVmxZQfI5/C5SZb6Eaexw
eylW/USM0YTylIlP1aAV4cFmgnTVccISDKaYpkfVFDhFIrq7bC9CRHHLLcTbfT2S
/4OV+GkRcptI6uBVCJCUiWKLMvvmaf/a50k7CHYUpVF8LBlhdQUwW03eNnDR5owN
wZe7tXPMiFkZdq8kXtQA3aCSnpJ8ACTj93IuO46bk/44wGATh9xxu+QoXejWUx/q
cHLEd/kLLAT2s3hFMRzhUS9gbCUs+zRSZhX4nurv8Nlp4OVICNL3So+kbNBo1SiO
fSreHWxhqMW4LPThsPau/V8aTqF8ZtijIImgOk4owydur3k9yhUQ+KVcpKFhL2fG
g9+q8uJ+nvtnQtMVYBWglcCFhfUHLBV65sgRGCtdS6DSLHJ+NM1/GYuWzdLzwW0e
lKjt3ax2t2pwR84KkVfX9hNycHspmao7Q8RsTcfrsbIWwqD45QDO4mp4su+hSTkn
5Vm4X03vwab6m4V21efXopOKXYDW4sWmRRFaQXVzV17odUHR3cBtsKWOTjKf9BRn
irXOr/nO9Vvq1wlyWibQ+Iffyeux2RHHTJNnP1eSpilo1kzXZFbHG336NiUq3lLV
HGXE200WvXA+p/lkADGUGAGU8Ik9tILy6NWLGVOtbq8MwRpeDLWri5QfJytrFAOO
vW9UR7tU8dabUwVmM0kxxhMCJ0ei5jkxMZyeTtLoMdB5oWeeBl6bVds25u3sBaLw
W22UMQ5tn4jNtsw+OepRjLElho6bQZnMyArd0U6b3cSq2Z9tWLS+2x51EJalCNQE
Ff8zU8nZb9dPViqgbQ3nVylZZSnnmQYiXLU4kKrysSPpWzGBCmRCin7uD+aNg7He
MIBlryPJbFuCi3O6kuxQS6e5iYdzX3i/OmMjW7Rz02g3QKxzt7Kc46nj5Hx8c2Q6
4b0iRaQjUi2TYfN+itf3STYzDh/YkqbOLH579SvJDmV9ZERY+dbZrCt01CRrSx/u
mbjWVQRpjkXaJQX5dGwpMypmvbEKxR02nAcaBuCP0AQvSejUYyPIs9s4AyRHCMN8
L0f10KE/OWYEnH6eq1n3NQQirrnAG5x6AV1kFjZGSKCKVxq+7Dikqw9LBLFmweUc
j08idbJaI/g/qQROjKW/+KsDOnaIPJgdyOztiVgvkFqXzT7IWRlerN3ak12NvGuc
DWamEF1kAvurJDTEnlTFD7ef7XBkKo6c4Me1erIv04DtV2Yi66x7hm/GUzNJ7Dh9
fjUZgoW/2YyUspos8SxmXMdMPAd/+c2syjG0q6HE3lIfEJRx6vmmTglRpDPcYmCt
Kb1vIOecMuXdiLvFnMGyT0jL+eqCZt3J/KFFADS7wNTwBn70+qiimZpp6UyXVkDO
K1G3FvTLnENDi6y3Slbzgi+i63Cdnip3IBR5k6V0RCF1nKAmRu0j6Hc73sgIRYWm
1N9sHGVZs6lxK4Jr5Gc6RLDVLh4MKMpcgwz2nmhEn5K9ErzVrzMlK+0WouoaH6xO
xTRTzca2o+tN2uF4QQJ9yEzAsrhZl6bJf9/NyD0ne9u4JrQyeT/k92cKZNC5Korj
7yJnFJeOPvyC0rMegHWRO+8QzQcQ66rzyJdC3mnJuQaDvU/Oz8OP7B9wcEZH2YDg
dJ2X57Dpw0c6ezlBWNWzBS+SYSa4QTMhrW/kCUGpQJwJIfwTAnqPUg2Iv2kDGogW
frKQOO2RZuDCqq/lMRgqylPqP8/U8NduJC3oPqst5JCmf+IpTcKSylpIJOwA4P+F
6WXWL/VO3EH41ByTU6kSdHvC7XgAJXUU/g5ZqokEorFuEYWAZyqlSh2ULvwanLl6
ozxw6dAwsDQuUZr5ewDAm+4SBMa66fXuROsIoo2DQ9uTFtPPbu2NHzba9ZK8lN0d
yKUE61X8wwXfNzNNpQnqnEh344ULh9L3xI+ZZqZEoCJEtrUhtBSBWsQH3Bxn8nNI
TZ3ZqkNTF3LXD92R+zRZ4cOoaLlI/11LZi5IfqfIgGeUqoqhveS9apPxOK3YWsmO
3fbxrM/xv6CzyQGg/4enbfGGQoLYWqgxMvNYgxuUTxo3uQeItEcCzW6kRa087fr0
Cw2iFUBrSIwiZ3/CwKn9PFIRyFvINhA9JDKiampvpUGjvhVJTF4iXcUcKndWF+Ng
LbYv238vvih6qQnA8FO1BVqRrOedMKON6H23uuOGfo6xMNpnr05XGVgUkaUdbDTw
Y7hXizrL9xl4BkadiUSiI9T3o8TG/mkw6hWiuCvPIGxg8W8FU9lcbCzh3tPX6B3b
o7t6vbu1NX+b56U7ra8sVjsVZSDwTzmXKVnKfISvIxrEWJRwG6f5Y5R+TAj3xxK/
EfcLheSwkUYOQIITP6pkVXNfEn9AoKWEA8jbVktkH4vmc9wgRfsIJA09b9RWSxzz
JAZX+jJzUBASq5UiZpIEcfZH3NS6pa1e3/8MAEU/APyGO+66zViTzNAwDCUjAG0n
UXqJYDShaL0pU1GoqDj/sYubRY8HkNGNT6/b1Vx2xvcRyuQFPJqzhIey7g5V8HBd
zQwQSEvYO8BLDBZ7WbtnGZAaaA1qyMetPD4sbsjWsdpylqK0KHTdycn1+ra5miVo
LZ3gowc8L3fnuU/GkMyDLZ6vq5isxlCZPppz33D3YdgeqWnq2DJ4oXxY3a+sU93C
PUSjNdf7R/qGRn/G5qcV4cI1YZ1BLnolpSA1wSHmt4xZmi5YzbFG7w9SGOEy5RRf
Y1Qdq0A2yl27k+d7vqA/MrAelY9vB99aHiO4wnfEnayHVj2lMbLX54s8hp8xrXl8
ovX0GU8QwXP9C556MobC5lef14ZjmXVV4F4jvu8yQEnCfwLIeXZhHcaqeyQmz0bw
zpFzhAFn3UT+8F31eqZBG2kH6guM0vtqFTUjhtyDRzmV+U/LLcDA620w8H+mr1rI
lJXF8uBdqppPGxTeaDU3kxrIO2ZxhfyidXZo98qZWCqytfmCOIl1HAJtvQ/kumXk
u/yOQitnBdLiLLbt5B6hpOOijt0Sf0iXgGNVdxvI+QR9v7H1apg5nHP/x4nury5A
M7LeEQ5XqyEfEcqprqKB7FB/QH/2TJHajJYpoDaCC4Sd2oUR7I4J9DIl7pbzHOCO
jobA8NwRBnTzYqqUPMvOzYT2ZHfKE807QckegFHjgxb3bpZZeC8pcWAE6tAjd94x
+5u3yEYclbkItVeBVCaUKx6fAsU9P64R4NnEJFAYrguBuHt8rnZ7tPwd2gsPgtO6
MR6EBVGbsy+ynrZNYZZtXa2MfXUeeGBQ8428Gck/Io0WzK4erDsv8xo0iSHNItsk
l7FgkxFoonys/U7mpD+tAGm4ooPw3GSg3LBxOkuhpU/AmOJ7tkTetSUhvNJYuNNY
y6AefYJCiISc06a0pW1WrBfOvj9ep32ZoYSkRPA1c/bZ64baSvl6mbXsMRYqBmnk
Rm3Es4y3anK5GIcp2NtvD8Lp2arsrHlBciwD0PQEh9QsTof0ZWfQgsEnQfzT8/7I
Bow+KLDkrmbG9Q3oyvavDSfcWaBCV1uevoMayDXaUEBRqKXvHh12JW8OQZqBg8mt
Towg7KXbgzqyN1yRbkiIi84O4taeQMJRTu9B6QadATL3GdoNubAbCaUTNWcCuRt+
7kgfi+MhXvf5jtWvcWoovqFUuM2JeqcUFVmzFo2c+yhERAOYVtgE1Bkd8HmJZv1h
QfmpWgu5PGm5xqYEr8E6hm7Ids7Y0+8nUDf1xcUuc/me+0ACMjZ2+5BK9IatdD9a
o+PPeoWnLF5V5cdCNWdil4k42mNeRvQj8qbn/Ly26NBJ+dPs4SOEE1USMrbinqrR
7wS4Ny3p59THERPsItRiIx95c9g3uXuQePhYcF7jTZ+HNESwK0tDkNnXfW9C+I1Q
kXaVzXuknlpfptCKDDUG1DLU/+EVJVuWwZj7m8ibBOZvyZfGtl2IT2kPEwfpDHAN
C4fxJrWcmT9nGue02aH8qtfpiCHZJ2rAjDroIf84jcZh2Cz+kT9Rjc1g8GQc3HKd
9UYDroiLrMmhIOXfqaA3g47sVS6cHBCy3KuZdL5vtyONtzeOejxbahx0iiUJQAtd
dnJypa2eCX4W4WiGttp2v/2p2RySxIT3vP41h36FHMe/tGuFyGbI17xEhU1CkEBO
l5s48IJRaX7RviMlblSaEFAz1/AOajk3u4WJm/C/fxfHW+yPcxr1uwdfXb8kedQw
idfhlXMP/AqeYMZ3ujwo7fT85E4s5DciJg8iwfSo1byLXPy5QXMLIvn5xCbn7gnw
fT0A/QUMypFAxkJngS01gWMRC28TM3NCu8P983qPpEtcIUZfAP5n4p/v5RXFS8cW
yEIhgl+0JArQNFG8vfqGD6fqfIksIxFZ7FXMhkMfdeIjo9IJDBg06sSvTz6wlBDs
HMcQwsBoTleZYgZwRmEl+++HSNNXQhP54jLjevs5pwV/qCEej+SLB7hn+qrHDfFE
LSkfyIPJLcANPlvlIyzVnY+Gcw5tVgix+rTH56FRhhc+0BsKlmCZ0tiUDq/urfhs
m4+87LxJY0Est/zQAN8UZPHinyYOYuyYd0itgPCvTeHdPENws/hT3glElj0x4Cb0
q9xX08/h+/oQg7B962tSqru74UTZO9qcbmdXk5jbIqaCzf1wLphZOWlmmmi5DHeG
PkVrcSNjzX3wSqZJV2OLmFRhOApcfgJhjWk546MhfR7Tm4L4tS78F/H1zMrDdtbg
+0E6kV51OL/aqjuKeP8LKp8nw6++jNTxMXjNSRSEL2lBBlxSswQqkHiey13lCXCh
RYfE3GQ5C2J678xsVNtIjBVcC5sCp/qx96CUXwKCvIh+TTQYvISVy59wu0t92840
Ltq6+eh/qQ78idy5R/hlq8wfUk9XCA8i8kQD03ieKE1RGbaXBbNrD9MjcHyoE1q/
4oagkecwtx/je4Y0A8SMoJVjDMTWYbckU87W8DpoDvKTCb3wqMZl2F5okXQ/ycct
BOzAy8afLcss3fO9Gk9z+f2Yyog4olvfAYz0kKhNfcqfXPBOtDPlPzaL6i0C0qJf
ZxOG3sVJtTRCDAl4V2b09Tt9p/ABvjHxOPUH1w80PweKR7Cu+cebtr0++SYhmZt5
gafUhjalXjpGXUmuvXne7of5kVwSHWBlbd3tv+uFW7WL72mGtw+uQujBzmHWFhkr
VnhCf1kBWhtIu19hMEV5OJy0rX25wc+JxBWOQZYGNZaBl8MuZPcVk1cF94GVPyfy
vj8tesXKejRwcpwFSlyGjMBCCWJdZmgbiXlvjZmIN8IRB5RPSDNnqZ9MxUD+PKvQ
znG4/uy0YmjSNyzZuN71I2Yduj9kYVEP4bdutF3D5Uj/MFI3Oz3nyKGXQhuhexJG
8d2SiS4v9bL2h7K7J/MF/Vq9XMHWzlktgbdZK3y8aCkZyQ9TaGYKU5u7HRSltJmm
cQs/xTyYBLnYsmSl9Vzto2U4O1HPCRMIQLNV+m6OBTkGO0H/7GuIg6odIJ/+POh7
kNd41ycbnlhbGcNTdogVw/aJL71+yHw5J4/YOY5sK3v3t6aYhqNmbCE/u3fLjsI9
4KWmClOur4KoexAcZWp95iJ7//gD0lB/KafvHu0/J2gDCwTg10PSe/64+pq98QRQ
xuv1DgCYdOsq/3ntjtwWy25uoln/eVFPw+VyuxpW7JhHBxOOdtSH9c/gKZUSIe3j
DTOFN7+M4J4Nc65yudGfRnRyKEJviLxy3ECVRvW3biKM0c/zSpmXcPSsKIj7IkuJ
PW1AkL1Nm7+3rbyiqQtBCVxyiQtQNcT7JWfx2MB4nDFPkdz9nydpd04woHbq5VIF
r13wl5mQWuTxSXDUnqgVy0PoOD9GtKXTSS022B5ytJqeGg4Eh84kcNBjplv/qLZM
lkS8ff32IF/oOXFQBr+e7F+4bHptLoDxL/gD5RR+d5akLv5uAtQmampIOqOX6TE5
fUSAWsWHNdA9BWVdAf8qO5HJiT9qkDrqKWJe6SOEdMmLXUJS139Gg+7cHN7CeXns
VMSqcKP3eopuYsOlqblnVeIRMIDT7NleNrMwbaINjP+yFBcvhlguHiLt59KD9Anl
Q7aSDNGVrEBfJAaUGHxFQos/PPrft0zAM0p28sSncf2m+7Z5/Zi8Bqx9aiXOel/l
SScbaSiWuDJDkpZ11JT0QNJSR68eBV6sWAAv4Gq8dIGAkNm/jrA28qIYbrAAAhKk
QPB20gMR0k6lGsnigcWSmrOe3Mlq630tz1q1V61XYXp7/6tTieUFAypngmjrjM0Z
HpCeCTgnQ2vE/wELiNx9lRzt8HfBARQE7xK/I73yZqjIIHl1KlOwW2UELyPljKsu
K3PdZvjMPPstuKnP7RoRhmuDK4YXlW7S6pVTT10OVhyles8MfWoT0uDAo/uNkBMk
SmGzWONkLCvBbf0Y3WTDNAhkeIen78HV4FPit7Wfp2C43HJM9n6ZZudjk6CbJgJR
YqG7CX/w7ek5ugXC/zSDSqSstnzSAnve7o365ftqzgcNhRxZfZGoe9vAfgz1a/qB
iXcTg140Zzlf6BDJKkE01ZLrZp89Fd/nZzF6/x68pggPnNyt8KeEr05S1maoQlco
D6FduvQMtbMyYn2zu00SRhZQVtGMYjiadH20ul6R1pFoXI6C4a/TpbQgjrUoqDua
DTrY7y3o0PHlGJs+XajAx4IgPOUY+rC4BesbGAi18IUz8LFMQm1eIxdhRl9kQ0JX
Gb3zdiVVBnEVu2eNOE/1s21oQKvNAXT0nW2FG0sOYDMDqiTBlwexJ9ybV3HraP7B
xGGbdOPCMwyh8H6WMsDOzz54xN36OYSqvxZ/TJiapZxTaKxn9xERO0fD6ct0vM9R
yJY0kgx/Qa1w/X+qd2LB4u8YWfgOPhx1X+ow8cDrsjqTqr+Elfgx20U56kqWkCZf
RU9Zfopm6kBcMejrRrmHsWOByz8lkc3PWRAWVTfkR+u0vOlacJbjtMMTLelpQroh
xF63GJHg4BGZg1UyBDYaE5k6SEUuBXycq1NrgPW5f+B/ExE4aj4lvBh0HBUiweIv
n89CePSVUI38tWD80BQKRjYCfhi72re5Ofzv4vGu9WZNmh1nE3oz34oRcfs51aRs
tYw2DwOTe85qcYqzAeksL968w8Gr676zumgb4itCpjieQly7UysEpWC+rUy6dNHZ
Xdqll2jquI4RLcSnAC/jRIfLtAExKcd8mnntNWzxdG1Q/ryGk73kaoN8swR03A0c
1QSlqhJdpc7I30jYSnOAvRGHHkogaKHyNI+VvrPkNyC+yaZCUkE6t1YwdB1SAJ/N
9WG7ZRwpTRYZBG6WW0GiagcT9MhyC+GOO/0D8Ek3YyjEJ3F5tA92DxCjF9ovIioA
YP+iixqmYz5U1FJnN/3kj17Ro0vCkOn3oaU4ccSdgeoqviAAmU3NK2RhNawmXh0G
wA2mTm3C7ZChGb4rxQYD/zf8wdMq9LnkBAh2lqdC85SX2mNnDVjUsN/7HhgQ9dF4
jwWqRraxSi0dL19+kPxPGx2NoW2RTHMjIknaEPQozkZn0ut7Tu6vuBVmj9SoPtAJ
HOQq7m0MR13mw5ua4lKQVDsUY/M1IQpuwtREMGgDzScZJ3OzU84a30Pat5XoUPQz
6O0SY1pFgOJVWhqQE7l/ooNIR8ix+3Ci6I3nIItRu8Q+P4ulFypJFHSBU/eW8x0C
HfKVxt4niGEQHbxZYvznfxOvf0IMIqwHj6bHiLw9hu5cF5o2Ac7D3qbGMPsvv3nA
9jwpf/gWLAPO6cPjz1cxFCemwSU2C/vTvUox4PACb+N1wqA6VlNN5/BWnvCyt8oi
E4FujPw38d4kldUfRjeoNJP9YDLsyJt8N8uiYdSQnG09w4B5lfiXD7bB7K6UxKcU
dg2pPrjeP+J8rrvjrrEeHnQzDnUoBDZWkaSSDWl9r1kSJVDNnn7JdA/PnNwbFYni
/7ALNyJOYnzoWih56qd8q0QY5u75GkOnLH4hbG2m0TOPGjPV83xsIkZ5rvUFOU66
PfWjkzVOyTIuonPx4H/r9hPV3ntZeTDZSHelqqYra08Gwpq9TljwU/IR62s3A/8D
9jgbkMn6bQvz6PcaUE349paMsrJ7KjTfgACTLPRT+vtcQnoorMEN6vCIsrc9i5XH
nlehZMHLnWA82cNEfGCuqX3SqAfFojN/utLqPUneqdKgNHfBs24EmkPJHG6hSCr+
tikGFhjlv3i+XnXDEyRPVQt5k1M7e3k10dSPm4maKqgWbb3X7UUUTdFLUmif1Jsv
Onli5h030Gh6E/L15/nUQk92+FBiNgsev9jzftzxX7eONhGaLDPncmjZHMJm4tyK
nt8lIKFOhzwt2lFF0HPkh7fY0nIb1Fx/6mllYLazRlWyDQp9OhocGP9usXRozgzn
KJWV8frrDn6eGcXt9i4C6bdI0mxgSOXTlGz+0wVf7DedxQff4GycY0z/kaWh2FUu
9BKeKiRi+eTbVZpqaJQGIe1uy/TTjTy+DDHSPMFW61C0tgNirik4DnQ/V+qiZShQ
/gRkhxS9mqOPbbb69jcvYhlgjjgKX0uarF1Odk4SdMglsJz6c57GQBeTc59YBhbM
YSM4pvYi0b6hGfG/iOZNqA4Y11ctP/vC/2aaigF8hkxaUzSm+ebI/iYrY0k+0mc5
mo8E3qIgLtFhwx5VZMPIYR7uiw3LyL8OKs4+fm6h9jWdm1YJ0/HZXZzNJVERP2i/
i3geAmqJDvXSg4DblGGEYyAnjy8LoaD/9oCyIouG33z5C5KIWaeOQHIvIPxHOb7B
CDJTKoXtYJ1c5zMqxDThoUNwYWgIT4wg7eBwT8e8oOUncgaR4Ee7ZInOLtmfMw6W
6IEx3P2OLqx9MUkh5XgP/CXO3N/avcF8CGNfFgiG+ZjUwR6fga6WdZ/AGrPJRa12
+sdKnLEU+BtcZj/zs1SqQ74Nsi229zyAUhNUYK5zRBum3vnSVtcd42ZV36ECZaoM
G1eop9hurM1pJ/tvWnDf9QN20ThGR8pubaCZ7zz/fy+h0c7USxoYX44S72ccVb9L
zXwZI/6FrjvKcIRNFBtIuDXNYpDLE8P1zZIXnS5sgnDAXp6qvyJy/QmlAva62kwH
Y3T6ZtnJbH62fytHiNhYT6rP9A6fUs+PypTPI/yeMoiEW/YnHXKNM8/4zkUhf/kt
/CfQ9Jiu/+XNrtqpycPQ3kCvTTdW/k4O27A2nIbJat+PBGMV4gmzjN+Aqt+0ICWf
Z5SWhg/I00hp7Nol88Uf1+iNJ+pUv90n0URdLjhdMWs6hiYNDwU6AchOHEU+PXsU
d8aGhm8MpAC9pgLghjPCNgt1cIS8xJt0toP0n3t6KBPq3874DYT38F8RD7FDNq9u
0AbGNbGlTISDh2CF5DCrVbwaG7xQsb8I6S9S6NtCn8QHFuXxqbx7T5lvYYdq+3p6
1QlYX7ybkABoF4yohJw4FJrChbNOYzgHO1WtBuoNTU0DkJ002SABfBdxlZw4hSt3
pXjkHOopRJ9WbvydANTuXwm+2xGkGql3kM4GjhZ3gS0BrYlDzX9WnUK0yr1/2Ing
3pxysHrm92+1PJ9d8j/IklVAXzTolTCdbwu4cGT2MITVEpb10OD/OlCdjdTQCaD0
LsA30WSOzXfqgmiN9DIoV7pCAjZS9I/rbzF7u4c6Nilrwy+7BSqfBFfkYqzag6jy
QPEiIF0Fil9HnOAFrPInhf0mCR/DaBAvy/drZvOJnys5GZsyZKQvDBEOuUNFnyAc
9CrOI52E2vpeFLtvVE3uaJqfZsUcJ4+vq5s1qwW3hRwoBUKJPXAtQTwnO4MIC/CM
50kOl+L2q+ThVRfEAzh/2G2qSZHa91mpTxdL1RnpWOVo3RWw2mJWolW/hBYCyhS1
XuxskZ0tuPVlGhFAewR4OX1ipQAU0h0TDt3p4xXp+8RrNJs0oUFHQZgMg7OZEORa
Q0Xy/rQCT2iaDuZFIlx6vkcWuhjtWuUqcHgfBl2lT80s8g5pG17sl6SSv60wbP3C
4LJodhOiyP1k4z3lLeNwktNoemQ/b6Ch9qhHVH06vsUHiDSCLK3MpjklmpQgLnY9
qBZgfs4VBLoEzb3DDEadTuRHDp2elZqKC84b7GNi4HrUY+ut+m/REyrsgXWApm5U
S4KuZ6GZQeGXz432sXk8GW+ROw3EMO0HsiqlT9Ige07eWPzYrGG/JEfO36ny52Sl
24ch94TonlcBfV8g0v39NbCe/721c4FvY8yVLSstrCX9+2TEuoQHpByz3fVa7k5f
Jr6tZvB/lQHq07hcUvwEDGgrXi1a4AP1DsWa6dajVAy+jwzBYL7mls0QLLDe4wPO
95LvzExFeOeAVpdT2h24+32ZigUx3rHNq5Vua1T6YymnVrjPfqzj3I3YEj81l4Oi
hyVOAu4v2kM7fJhI5t6rU67Wxxv39LzuhguEr5ol96PzTzIWQcf8+NssehPDlETC
VTiE1V/b4I0CZPPUdZbiSsvCyOUkSN1+uDf619n/UhdbAkHM2RoRanxoRSqWErMe
mGza709Vfn2JV9I40ulL2FvmNUc+KBfQ/1Jc2Nxh5ThiJHb4hVkSpyI9IjnffvGU
BEQIyTKV4kY5Ky2VKvZ7SlivkrUWoJWP8Bemc4AzX9EOMCE0JLqd2mpFFcCq+0Wq
AeA0lZ3RLbvkeYcUYvJhN8scxaO5Lp+TOAU/5MU1yTlQKfoVFDS/78oNPpseIzTH
h5+zDG3S5wQA6rmNPK0o55CZzLHEWb+00EBbj7L2cGiCwtSkTiSrd2Oa004bfvX4
iEt03fu7sU0sV/VutgjaUQhj6lOd9HNIjOLSYZZEBnjnW4cSPnLfaYtStgoiJsBS
UUWN/8FzxcuP0hL/8dpXiQ7psrnJSnq2x6CvETvb4q2vjJqiItGFuHh67NHJp5wY
NnMLxqAl54tjilCTWuTjn62vH4GQrXQEqjMbLBK+1iWB4OzR8LNAgf2/6xa4ppF4
rQyZngpgnmO3r00WlTh04HL9OXPa47DilqDIPbosLMQsjw40og3u7m55P4zUjUge
V9sLX+JgbNb+0xtbNASVT6K7C5YbACrdtdj0h9P0d2BilVq2FEOjq2BZYv1oJoyn
aqwOLuY1H7Ul+8nc8vwHQ4Dr2/dDpiNiMEq+VBxDgjYyj3/QBFbFVlZQrmjwomp0
4AVMgwtGC5clC/EIwjTrjxU4bcjE4X3s/tkdwBfOFobDPxj/44JBnZaqKQuatrsL
2V55muEmaCV5CBRshT8AzG3Z6uomHzH1U69t3k2JsQ0gbcbO4L2zQKje/BZLKSbl
lt4xFjcyROPU78J2MR97riXYdFHAEakCCC7KCnZfPKSVBVb6kIh94UeryQiDuwkf
u9NzqvKnWHKXUuT++BIfQYQTd3FizXFIV5QaY4iudk4a+EpQbnpoHz8ZEE7M8mtb
B/6JIPsTHTu6UimZKruH9bbOABX4xynLwIiaeK+BVQ2uyynhRwnjspqc9EBFN23Y
98PoS8jqfSTX0hrTXQk1riwotAzL7ji0eTJdv7npvyuvnWNn180Rozd3qTJ/RPvJ
i/0ZZFmmdFLeSznfwYti63gm4v8plFYjEbdnxSJedOdvXtgYu8ygP/hU51KKsaNp
ODKMQh0WBT2lECy33sNlYxhIKME1qwJFONPYKPPOI4rw2C+SCCPwvR1Iw0Fn6ZO8
/3BDWk+Uzbhl9PLOH+Xe3ztnMmRdPJQu67MmcEHKde/Gbth4uWuE+usnzy885apE
q7yNxmIEEOxrWnOjvlg1ZOXR3XHK91JvNG/2dUcxB+bdY1cL3qgEy/Ra8xtp4AjD
YAzoXg4twUpxjVU7DA5t+gHps1hKcuBmeh1g+JeZO+uNJzAsdZDK1iBQmhFA8GqJ
sy2ioN50JKZHFkX+OECwkeQ0yK3sJ9/5oLdvK6x8jer7soU2OLXfJucKwlKJh1oR
BYsB6M6cpRrTnol+uTx9VwjvmsPhXMpWS/cWajwt+CFrC+K/kqvo3DbwyD4RV0Gt
5bZ5495mLClM8iQcpAHs8Ze5BFtSt5oSd4dnh4sNGeqmb0Oa1wR9N9OnS4oQUvX0
psrtpngLCYyX/U1QcXqXalmQJ2fXPE8edD3rWYAQWH6re8DVkmSmbcttN9n9pnJz
qDSaFbtvvcVPM/3mHIJcRL8YUBTqWkM+vbgMjvzEKQS8Z9rgTAcK9OAJAbqWrltH
tif497VokVa25WSxuSFNoB1D6RqzDNbNzvp3/IwDgzT4TBYdu3w8Nt9yMJEjb0Zc
7usLPJCVelPTpjEX532QXy6KtOBLng+7OPMPJz/y0QnSM7GAeOcHp+iQkhW6Xc0b
9uqdUPJw9ctR7xoQ1EdTZLr6AP+HhtDoahZRzmE3g6IBu1ziqe2VE9HU2hRtF52n
3MsqJ2BmrUrahENrVMn4NZoFGRBE33CHqtYSsnGSksMIk0zpu27yFm4N+2QGEE6u
J1Vo4Gs1pVe904RO/nJSFbaaRuA/Wzhr883zbOuk+i7I9yCs9G75ObhJYCSMO/4Q
0a18dr/TGCzdyzsXjfUrGv8NZadj9ZC9rBV6fZ1pnFQE5ngO1LsBatj0xRZ0Slkf
0X9XQjXGCzGkwTQdnT2JS+R97tfJUb84hCXWo/Eac4fiVuMqcywMLg4rwEHbxvC6
LuW9HJ2Ir+Y0w0CNpOYZ9v3a3p2yV1UV/Y1ghPE3uYk8kIlIrJV/rd975GzU7zhF
XyI1sPgh3lqv/Yu5BT7FBkQFrLsW6mTVdHVnGNu1s8I6SQhjAWJ1o4sE0x5VhYXa
eNA+pyPONVLbqAqQWHZOOQMWdEgvjChG3N2WoiIC+XHMWAI1P4SAobf/O+7DLhEJ
cIiBEhZpnN3WPwP6XTOv7NXo28lZ9l4IHcaABaOFG5W5vSFf/+HGvRFEfxdQR7MJ
cc51BIU6c1Us2JHaVVjN9z533aea1TP8tfB7O/7RQr1mvlfq/eAD1f6RvUGt7HQg
SPznWCDhoiE8ngkWDz/MdL2JGUWOIuy+TMqsMHmVvqmr4jRPUqm2CpcBo/nuHfHQ
T661XKccnY7GRS3zSl97fz1wyPYOq21bD4r2lxQDSARml2qTHCtlD/moG5gB6eFb
V47cCKmaVLLimG7nu6LhcC39xTufW0DbePWHNyhDB3kdEaO2epSYVFBubLYr5jjP
C4NkSVhWF/v7axU6vaAcOdELG+7/JhkNijUJWEdGzIfdm1dwAcncPSSZ11Y/C8B8
/9nhdzkSkBfNjbZ1uCuJeh3YEovhPfKmtNdbx1lJwrrgTOPPR2LNW2fE1sxWp+rK
cpiqxaHDT5l6tkCY3ffWycE1Amb3LBU+7W6xVNGn9sl0cl9CosR3UHukKaTisWSm
AZSWyI9CGaqjCONDuilkOZtfYDweYFoC32bCvDcexZnl23MoWogVhxNSvz00tUyo
ImdaASyEaq+m1YmIfqOoFP4OA2w1RkCAsOf9kh4SoJXMoJyKZpdY7f8m1UUSUzOH
EHidObjklKOBKbgnyuyFwEkkEVUBdZquOBbwVcMa8alGP9R+N5CukEiI4icpL1Ux
vOHnlluk5ZfDW+Ar2DllmP2+8izxgIsulipd9mJrTXVSuAnI9qX410LLKaqAHIMc
wzn8ptA/+v3z+3a2St3zN0R3/8c9c9doPZu9v4QJSySFCsmW/Z7lLZb8pX4JBfU2
fLKnCQ7vekM+csrhJkKyE4C4ZeipQNZEL7wy4jhWH7cOASaGcihG4CGEsaiiyz3N
0nLiJZzZEHkwT2vtbXDLwWVn72ts9GFEbCIlcT0Aydzfjz88jcGUgTdQ9jDgVTWm
0we8TAiYFmOEOIE61fbAKFIDbNMYwWfuFWhsYuvPnoeogFb3cep4en4nF5g3cVN+
4Fgppx8CWJ3E8d1kT2N+pLKXTY11maPkOJS80mG630hPBb4gBFkqNd/NN8cHan3y
3JevMWk6YzjpraUJpwXrDB8YgQK75UFSvXD8sP9357v8/o1x3nSrWN8DXIkYy8j3
cjrMEepKNaWz93nQ+1rcM096iul6HERMVNi31GwuaqCR9TQ43XfUK3gokfpfe/Tr
/sIuFqi2xMOY/sVKbt3kdeZUQnajLWYN9iqWCy6daWFG7yQtPvyo9GlLy5Qxyvjj
EjfJ2DlL7SqQAmJSLGWSBzLTNasvqt9cGo1hM/jrEWj7YPZC3+3iA11m6Tzz7Ny/
ryWJ9hqR7kfxGkZjq7nSQMd/36dSgQT/I30DBVqOdfYEJT82UWVCDa1ETijcld5M
pQ7KHRibqfO5CUw4eZzJ2A11r2EbzRNHO8rfJ6AwTKH+HQHqb+72RBtEIOBHTX/N
Y+5O5qqRT7BR2Vg1WpF8P+Ae5m1mkCqzBtH6M6j0sX6wXKLqj3JhdsDEtZxIhGf3
j2UyptPu+Vf0JxJOLoJF3Ne2U4S2d9FP+ezJEdBux2/DtvpkKAkzoRCPEWX+8ARO
MlKbpycI8fDt8uhI6Hz8eT8mvCnzwOS0erjCbQoU89fDM3PfeIn2sIRVPdpRuxHU
AGC2peFvtE/EFCWjwajjWLMtiSR5+GZD8Aakunn9edXdS2+iFP1ghJ8s+2tyL1uT
BEMBRj0HAyNkWXImatzEGpp+dZTgaX5z/kIIMktq5GDeLFZlCKjf87mzSV8WfV2j
yowfU3omm7RlJydHgq2JiME7GB2QvTVOgGnTG7oPdMgUBTga/mTxA/e8AfeUAoSx
Ca6DVi0DrIaUN4gntxisehI8YdsRxGihzoP7xAFNFIA5/IzLUPZ6km9irZjm5R/A
tXJnRPsom9g0OX0mzGsMhN/osmllDUJPn9FkqoJT6DJV62qz91Wp1SSIZOWr9DX1
EwXraE0uJh5g6MpzM/b5WPB9hIqEJnZrHesnudLMdv5Q4yuvTK1XYqFddSCQ2jqD
5b3oltEUn2ou+qFEpb3WCoQHuxjPuCFM8+/LsQ6NhodPhLsXA4yKlUL1g7H2lJWA
FfWT4Np+eZ/SFHqdYxTgeTRhJo33rUAgeJ8VRArWmfg3yeiyGNZC0JfDP4wj2RVY
92jTrktfm5xH/WClbDCX3Z59L2XgvYAaETM5wMmXqNZuKCR6bchpDBYjDcxish2x
WMfSaY6PIdFVCJMUOHqs2Oir5/cHufh9ZxWQ1vCBKFU3ZWtGULmR52llYOylo2Dw
ty2VPY39cnR2PRrgrZpDnJ0cCrI/cvxxXUj+KMqO2z+aW7zXC7yYMIHXyQ9899zm
xs9XOomzNZOAZw7RDMSAViOZ8bqDflnDvH/po4LT4A+4OnH/TQBgFc4p3bWnXjQP
M+ebkhu0fq7Cu1XwIdiU7RpTUmU7VnrcmdtnT3hLvQwDIuv58H/PM96mPgRcM8Rs
3qJyvddl1mwSilbDFPmS53OjNkGqhDaseUzhiRm9kavXuIHkcm751wpG3a3D+Nho
CjPZNx6+Mfya6ysQ4XgMGxVOtZOro8lRvSbZS/8iWANb28Af/KNCarhtsuhBMA3N
yTN6R+uCmgsFyeHBeS9JfDKpqozquC8c2GoW1OeMB6iLy7VAqDqatFmALnEKvR+X
CSxaIEyohD4GZbwmebwO2Rwj6H4sr+guR/aqpkil72+jVs0hHDJbj0xYJpItlU84
njcRh4SgnNxQ90qPt5VumlXOd47zdWN9eV+f8viKTjTqw13WTdY6fqniMjwIaWAL
n8eSxl5oxoKez3dvAlUanq1q708DBqXGA/9YBYzif0/azRvNFLUMvKHmnOxIPFU5
cqWJasTnXvEPYKMKuTwiO4XgXFyuXFvpyAIjJ++WIMYoc9bgYJerRPrOqW/v2uxl
XMf32zSOckUE0uB1lMFRkQQJIfVBU60HiGGZfT1WkdePv6p1X6dRJStE96qebdKh
5XpUz/1jEMAhzy4e4FMNi4T3JX7Nh0zbysABPxrVQyCr3Y5y2BO8eJ624UL8er8r
5RivXRM1n7KCqomUh1pt1HMJPba0zcDQO+iwHIh4j/HA+HqzB82i9BaYJXMQneMs
IEj4dPoELfUibz3lp0JZvP+jCzsWc9w03ZgrNffyoi6FhE1VijIU1RU46dx+TxBL
ZGMjSGLotWyofduS9Fk9/yZA81tRV4GYFoKXLIopMTrMERuc1xVwSsmP0/i1QNQX
/VAx4yw4in7LWVqAO5Iz91fnjPVs9As29gKMo+dYpG+oVOrlHM9f9oBpkHYWfAIX
rBrpERC70F5CdV0EmQwYsaDxmI3aAKiWfwFVlPF6tX/WndSnleJ/jW6ghhPCZE/D
smMI4HXyCbf5UUPqmHzXdxiogm+egmC7zXFXZRx2tfvksuZCIDCfEGB1mvhH1zCe
hwRO6bJrJEKeDMGbTANH3pqwbTB3dgCC2ccK95M59Gzo2WwZONs5RxJlMg5OCqOu
dVWuvKq15DhdtVZVb/36pan60w0asKlsYmSFGKxhCuuKi2DjhQpNEOT3Yl6SexuA
/9vLcTQWaLfu6ecM6C9ZfmdD5LxS/VMB9Yp4ZYdO66RRTPp2ow+GWT51yakNPT+c
0CjmD8qF6U6BPVP75f6NAQCJ9dfwkA7YTrwt3vLexW2mNC38QwqJuX9Uk8zUT9hZ
3g+yhUfoYzqnX1p1b79DkV/UcjHGdOUGVPEKINFFF0lFSW/AsOD5OdB1bZZSMAq+
sF73y2WH0sqLQWIb37bjZ0tj3/CaDPoT1Uevy8cKRHYeazqZiBPKBEFzTGeDCtVU
ZnRBLzOO+btTvwAfsOe3gWXm2M4jle9LjIojzNWm/jx8cIOiSyT+lL5zg/RfbQuU
v0k7qfro+IqWT8EDvD2IZwp5N5NYvgIoWyRENM1OTUSnW5q7zKTM3USP66/IW5pg
nS9iUFOzzeOaIruLliUJd6fIOactyEjv40jhpobvPROSIyw05d/Tz/jQsWfTr5wP
6TciZyhTNbTMbaeh50DOAok4PlHvqv/BE09OXtKR6i9ETZBroJeFcGUksPfqtsjg
OkXiSPMGY4yUWJT80OqEswnoX/bNU+/v3tNH3BeQ219iuf+kZabdYJQJoAibv34o
r8c2KovUMEe+3WAf5XYC87BBuTt+3R5Urcj7ERXqC7uKLmmXUi+QPTvuuZofqmiN
iRxR9EGNrWdowuWdVIoaSJP1NSqEMVOVOzJRfgM7nRoJAHy9HzdI9tNef2HUiWvJ
XqqUOnf1RFV5iJVbKNdwlD9bBPBpwGzLxj/Y1V9GFJsL7HK9g3TrUAxoxCvV8hmK
oSflz83GzPLcQAal9/+laZyDe9NzA/j7f5WzbtmP6CNYUyEPSCo3I6hY/VsJ2p4T
cr5Vss9WBVzuo4Bx3Po+93S38VnctxACUYycUv1m/O+qWv9MUfSd0dyzWJcBsyx7
2jPDyHJ1FikBE7eriAo9xbe+EjrAvL3STVBTlqb0mPnHMXGFcIX2dtxRoTX4JbvQ
AkWW/3wGOToMgb/XhGE/1IXjWzahvm++xLDv7BxquXMKtdiDnlCnsmYhcReJurXu
Ykgxnjuj6Gw1lBkAtnoEFbW02FYthGxLIY8wGhGbdCELtv4yT2nvj7GrvFFy6oVo
uLYxsHjFR3pwf9lulE0N8CUDNkEyrMQvXbgWSFQ9OHPgvU5yt95AgzblDX9Cd4hU
+DW1vV0co8077qJPhVB2+w8JU8zsv1mYA6teBZUMkQO1v42RdeCsl3xZRc1qvV1m
nxSqxWJdbWBKR1lq9p4qrRm/zsIv+reFEHSqHLVyfa/nmkihsk5VhT567D/lXkyd
Ho+DMgW5VwOn6Bg3AF0shb46FRdHqf1AZCyf/JvOkJguOGi8aaoPj24Tlb2Pn09c
dnYOJHtQrvfiX/M64LLcaw+QIfo9O574BttNV6vDyRvvrzwsAFyaPF5W7eLPJhTe
4mKE6Kqg2Q7Cn+cHcm3+YQocdCcnlv1MoHHeD0lWH4Xzg9vArex39BFMZuAKT/GA
wKP014k0GKRoa8Jsf41+c6OyuUw7W/5xPYSelBJj+HwPAdRJOKUcUtj0ROsgHr1D
kopFxhoMbZ2zQtQ1QAfcvmTv+cyjD25BzMiBL3hdsyO65f2985bu9a8JWNcL324c
mynJqWVUfNarWQF/95LqgWWypTyj/xsgyKkrybrEU8j/EGhUZy0SWqBy8NwdqWTT
xetGNJfa7fRNaQRX9DZbirIMyQxS2w5Cq4o1ImQBa13y9MOnQVDD1lJjBHAsYp+M
q3rQZm8+yPGPiV3rnl231DUfNVvnrrs1Q36477/GE7xbTrii5bIc1vGjGM3f825C
6XT92KbWTXHdeRwVUw/yxz5yDl115BcdqL1kiS4vzGyUCdnXTz2ZTO9Cnt52tEMO
kpNbs2AD3xCAEuKzz7paOigZYIHincceV/WncM3q6GnOT6hySc7uwNn6ivvQWNxQ
u+zuZVZ4WLkMEexaIAyqVf6YS0lVJUs9XKz/jNyuYzDL/5gl2sU27o7jbp/PPqyz
IxlmYUysQ8eEwp1hJAT1sevY2PGJLL6E8/hN8vrxrEtpoRhjNGlAcd93XX0z1gcS
JzBgjVy6BUE9wPBzylV4Fuy9D4+dL7k3FMqzgUsjOK3R+vkxB8VsRudYebzEr4EZ
NB5+jHy1+FcCOQrK/w1aKNc+FmD4HTC9RsZ95Z8xvPPXqSnCibvn1jT9WsFyVHxQ
qsW5Un5rG7/6sXHReRjhcIvV36alm830GuWomToNINBKdz6FymmVT4WU72kZYwwb
8bdyBqXSSCmcnRuxaF4dzFvfnZh6Qu2MsD+0sAaAnrMFCv/3s62ONPoWaQdSPVzw
WRdjwd8whTu6TmjZJfcD0u8kVtNTfZt3w815TyyBGSrqdg8eufFHWiSNdZFzhJXC
wne8pKl35MZ2iKJhL6eDxZXSJLhZwLD2Sch+/bbggUB3fZlnXS9aNgNXeaUophN9
Wvuyvhd2rJQs78HsrHkH3xwqVDJaSnDThE5by7lfZfXNXIiFa/xKaPmmP8Lwo6UN
3Qb9BidM9tzLgTqsO06h3mvf/8h1yll0QjWlIq3V/Tp9dwYsMym0x/IyTzaNOAmJ
SxDAJ8POQqjJoOBaRi35hsX/VL8QX7jdaZiNI3I8mQtk1qRkkaInmE/4QuzDw8FF
Ey2QcAOW+lRYNuFjlKmmI+Vcz0Z1wCG8/oM/mVF8Th1RSuub+0XjpCZY4xkG92cv
lPf9AeGjOzHJMJb24OUBemR3rF8knFna6KGfOiCOHQ93LAMgI6vT+wAjNb0+jKd5
+jJGOTHfENFVDpzXOVQtz4enm7omYCl+P1YGovWMM3EJULxRKuWeBmyAeLE7Rawm
mMt2fj/J3+A91rg/IJ1hoqekln2RhjQjUf/ANX3Q25dkuD0SFg9kF/gMYtzxk/x1
1HDkNx57olgpGk/I6hwDaNR0J2QHWReNjS7z50Hz88CQeLUZC2chgcmrUdNw1aEl
xejIAwoC4wtlG+wjYqEyea+pspN+cbYkbSG/JxOhpvSFqNbtABR33OVhN4wyoXtf
70si0I3EmTreepo1EMxR7Qo7FeoF8ncZpzKbRz4bOc4YkPLF844sJGMuV3b0QU2O
ZXBl1YytqaOnKNFATp3XAfQ9d3JguS1U/1lQDpm1rZQ6Ghxz3UnZbYZyQJTd6EjM
TTy9sIsAZ1oO150mjbJmx6LW+oKoBuLcFZ0rLgOnennWGBNZVsBEXeKbxRUhyuEx
eemc33L/0S2IKjCuEXdUqhEW+aLYPypEOFelgEaLUTTcnqbjT9BGb/wzPPFvl19Y
M1GYQb3E339ivUJRRVGfzSDHHozxrY782TpcYlpK5PSET6/GjbPQtKOrlQD6j0N7
vqjY159Li7FF5TbJmrQ6uQwj7weuBEXM/OdR5CXpzeDb0C+LVCb1YyTAS+FMlWdH
re8hAE7CBfaZa+IpQyfFGNsaPZCXQ/9rbQX0Jgb2mjFSTh2cg0pys4WWbOFoM5RP
nXut0zez+htqkmly9Db1nrUUidKEsgXGoNiOgnoyAHQHPpFToAxS0EngGbMbjq6o
fbTKyfS3PW/QIj2FrMNBxncqWXyWLBuMxIoR2B7XRqYir1/fjjFJFIdzvojhF8NO
c96Rn03hCEvFJhvgvm7fW4G6u9bBRMVw20WqTMkwMCEGSu2DuetbyjKbbqA+6+hb
+AChiERjDu6E94gEXJCzz6h+WUaF1aAcotpZp7ERIUCD0WobXZt7m6T25WISC0uB
A6/iAgqtWYTbdUnqW7YmpNo3WW3ZUxRx3mGFYs5/ygph0LmLuB+OKQDPBa/YGqUF
cV+73P/rTaI0rvRGuuICHFHqiT5Ju1Wk5tUvTtMBMlE8hjgYOIh83xkFrBfSpdQV
QY727quAlbWyHWsMU8w0yT85JblPfJgykqU+nzZKnxbogy2lIn2H5rJAOSgw4F1C
FI7Z/hpsKbv8uOLUjRo7CaJyB4jQdwHOJcS0RTkddpihba7bC7UpJmlCR8mUgepu
vMOE9+eq78xDpUZ6S5EE56/BkzbIEo4yNxbB12x7jkuSj6CVU4Z4giuyTAkaP9hH
9a3Trx77PyumiFq1FRdRLGMPkGuMiOgi+5PJN1jqLglbyxmzgGaEfxzzvIRe79le
XzUvrzf84G4vrEl6/0SshcC//GAHZVFfKAPzNtibgS9lW+LVBR6AJvuVoXl/ISwh
inCXUGlmqG2F6Lhwy050YXO/KxpBytj6xw/WYrnMFuKawiQ86B8XC+O9WhgPc+J+
kf1BeqlAaUgsKnYSLsOXHVLdQ9shefrQwGSd9IlGTz7ym1jG/zt2GH9DuxRYygDJ
AzHtYQm0INnSB2iNabge6PAhfnyvSJ/vobHnrlosWMSlmy2oM2TjKRLWMODm+7ZC
8gPCt0KcO1UIYuhzpiXU+hDxdNSqRXCYXrj6+jODx/o0Al6JnQoVUdfId7IEx61Z
rVoBwdjpbOwfqlyzMT0SBKTfCyM2zE25dbZH9iACuIidtRMuEcYYcLtHf57TfnAe
JX84UmUvT73Lwyj34Fq6qXpAgQ80wYDo/4s3/7CejK9zGJ+vK0Bn72f6JNSgn1Er
Yre/CefRot5ZL92bvWo0X+lVHSmqP9Kx9Af4Xb7zirVOsGgL2t2zUobZMNqfstN+
p9L/QZ1UVmekhZ7XLr4qB4mhoYtmmRwmeYTNVBnshn2GE5NcPQhrLQfWWExPpeq4
Mf7rBs31luWByoeRYKDP567P/VOhPZ10fDVBKupK+tILiWgaCQo4qHJ3W9ExeCJc
Bwj5mwAqMEN2bnWX0SvU0Emp+iMd0Nxfh7NAo0KkR6lXPb/736HhiOD0wmn4GAfy
ZLwkxI7s9UYvVii/cDMAJRKT8OCn0urYk7i2uDImzlMFiHNB6yr+4Af+4TPUcU/s
aiJ2aJd/JOZLQsgYzyHKvhEbAYwDYMwm5vp85M2pQFVZOZ61mhVJLWB9uTHJugQc
6HyhZLjh7yPkOI1AZno5akYMOEMUxZBQzj+NGgBg48Jiu7TFtm+3kIqUvYwgQsOk
8GcIKyTVtMjg0KF2nKDTHqSdtnMTMF/5c2iLvCiumG1KtKzrhB2q8M4tEbU8whDJ
p5U1Cco1tV7k+8TqFbrl7pheXDsjhDTH1EEE1MVE9Z7dQWmMwkEHol2iVm1ZOIe2
Rb+D8T98+bpwo+2kpLNoQcBSOJaXHFZsCYUbtNJ3RqSwj5ck1LYFqhOowS/r6cHc
fH8PBCx547STIpnUxegGclynhwckGJrInwyPY6to6PnTEd8bkrRH0n9whZaru3oW
Kc3HB0hb1cGGwIyuVKQkmbPQ/y3gmmjAkYm+Vy8VYJp3Q+5tzM9Ls5XGxk3WOtXx
1gg7RsTDiO3zDTPmWO35aONgepVgQqUDpSV8PiiS+INM3cY8G+Jh69mGlpn9At23
hn0RDw221wou9umpxhYKMlueGTcX6Z47NDRwNqJFJJdB+47cSjSyXEfudSaQBdPa
oPdt77CJDxjjs57nKUA+Z4iZtxPdVQiN+ZRTZhnugMcbU/H8nRDCGM9WMNYZBLFg
QzCFPxJJiIfpzNxJ1e8OC7F4rGLTlEppi47Qw3cw9O1HD0mbaGk8NKgXvnzoa6r3
U2U4cAq9QO6hMNlVYW3gzjeF47LUwiznrjc5eqQFTftQN6bl9yIOlgLyDD4W7LPv
v2FrdNQRX+9gSWd94b5uOESsJ47C3ZWfByZ89OSYvr1eogbCScSsbYKGM2upGI+2
sHN/XOAPgRx0cBPTNfhM6Xsnkygp7/N0XQnjX0hUlOS8dSTKOubRhZVRVl7NnADN
Zl7dNU036PBeFP/wy/ftPo5q2t3tQiMansG3rVNyA4c9d8GLEnk9e/v7IuohJE+H
fOmbrYZYVEoRYc8tKKCZ2J7zYExuqpCnPtEmWmw5rKMJYgAcgg01fftAJkvwKKRi
gppwOhMzYgfSbj1+aml8guHCqIy4iU2nS5jzF45nYO6Zzn+icVu4tkWwbrm6bez/
850M8+0U6SeYVY1tLLk5in1BjhSoEvnkU3vDrvERI2zafRLtcWQ9gO8kHmn1swdx
TYzhLsru+K1iYJwNwrobl1/dE6rVu39DwaNrbKUGlVZgcUUgW/4uxXfPQzLXC7u2
CKrst2/bDduL/juMKmvrPXAo5pzxOK1/2VbBtKkMBKykQVzL9KgkXoWSA0ouiro9
sm2ghVs0gz7OLTMQtZtLxHj2ThDYT+4pjzvF/p8k3y/5QZT3HK0OSIbct4shjHQ5
GGihkJmb4grKHkUkWIVxrbbyDG+NnmJdYaZ/wHwjaqAAJrkFcjRAXuGWQopzx+Jm
24k9knF9ns/y4Uo/8l5HtBM+gYQS3DBkmQE/Cze5yh05W66ztts2v1J6U3hGqQjc
NaHCOPKbQWMXiYLQcqHHbvzN3G9XRwMcIpSY0hZEMrnfbSJaAROZVIt5iF6fIH2T
m1/zI8Xs8LM2CkpHPCmrkS873kpyIcL7ogHq2GTBsjgaK3pXwYO5KlyrcGctBEoo
b8SFdqDhuTXP7WJCv0NTHIEniDRb3VL+whAn90c38qa3ITxtUZPGQtvYlNbHvcbA
61UhGawqbFsxnXvnGAuHQC1GIdzV7Z004n7oDqDYNVyj5NRhFzB8l0On0c3qaHW2
j/vlKYncSzuNOnbWk/6QOU2s5awkNHPvaCRE8BewAwVrB/b+KIA40yL8/kSsl8bZ
/MUqQxaxiUvh3hH7OtbDH5oByiZ7olQKrCQJuf8UhfM6tySgR0FP6mBHgM6Qg9EF
RosJYwSSPk5jXgTp70h4LCzVEQ+RPo3lnFo5beUCpb9cDEBXopq0wnqeIdTjTV6f
dtjvBQZzUgDXcbZLPoeDPisILSiuiyeS1R28E+gwzrs3+kQPT+DJdWjcDozaiBef
wsfwUWCuEZPuspPFiUViwxN1DqkDs5gwScr0oNVbsKLYR9UUZSDizI1aNz3f/KbL
lv35wLwmKhtTv+st/ae/6iUOl83vP0n+hh2WYRJDRGsRSDQrJyw0w0A1z34LKhtZ
DFFLJJqmt8PR6m8EB6cfeNlQUCoiE1yofknvGrGImQFIeOXtg2Kps9bvI+9tqXgl
B/C/qelI9++9/cQiJeYz911mR2qoIDpCLFWD1fg7p+1VyeapqWC6DofkIPi5z+EF
v19Zmq1TgrakKfRbdzP0ZpnIaNQ3wAu6KDIjpLRNA4dSA5PrTee7J4IXlkGsnsvZ
G6CAMexQqcOobl8ws/z4NxUBw2ArJ+W7rwKf5FXktc2Lx7ZVzDiOtrwuhWN/KY78
KMHmcgGrJdZtLa/ix/gDqwaShCZiQJXFoPYDP3sfPHUEeUP55oEthJ2XS2NulXDS
v+tPhwjic/ak4sUPN2GIn3Qp9K0eMzoAUvAjxw80yZvZOeGayNbrjRF9qqC2ueTC
IMFsyPuJAJfZfRpsvwAugIqsECNfz6qi7N6IaJ2/ZGZdxD9rLlBrs9g/CgO0COip
oH91m6jZJ3FyVRoMi5+8j/OeSsVDxj5FPUBgA0SyNUfPLk7p6V9iUgmTXP+5LE+8
AIX1QWqe1Ja0jZuX+TEM+7z0YhbGAPhqtjJd4DnK0gQCMm7V+5OKRba+pV266IeG
HG35BpPuZzRsAz6VwX70mEWTZBv7qxvqQTbAg5h5rFQzqS/7kZvGOjATRRUfNY+R
4P67G/UbvKE1f4L1iGNqEss4Ai/WupUHx63z8Biy4et9Q3Q7zyed/ZhT3XqlSsz1
NkSdTF6e0xBL1fAKHOTeYQ2GzQn5XxG8bTMczn4MXwuAAVvy70T0NxWwVz0ebc4n
4iL26YR2wCYhD9xGE36ofJ3kAr2MZasPcOQzHV8yA8nhuIlzaH/IdzxjTOsF+FWJ
yfUvHD/NSJIWnpf3Rc59/gOUXgVvIRYo8HZ2yAgwqcAuGx7pJuxVfaw/NEEM/Rgy
x/6NYuK19dtLH+WUsusNlYLrUD3QLkEi5eVx8fSW/6tWpZ11t4LJ+FiRFjzraNT/
qVP9S9SjLf5p1Ip4TI5AhCbQyVrTtc185mG6+bGATocXTZrKZNrU64zaAX/H4Umh
M/Y344dh0sK8pTuBDIL9BYa42EyATrgxXh9YChL5Whz+3CCZevstzuyFyLZaB5uB
I9oljGxNt7D1C2bpDhY1KiI7Y5KkkDR6FgdEN1HNSGkz+vXSJGZRAE6KVgJ0cZiH
n1Z4NDdLdFJKB7iCtf2dO2uGvMGKVe9GYXTaU/9biySkpmUYoAQtsRC5qsuNZ5GJ
ygklqF8om3eQ8PVGlIdCX553nrkzP0l3lZ8i8O2qGTMFn7hlZ1CCnVnWLZ/nIJkh
2ZKJ1wIxSj16aQeaRbb5dgB2TcB+p0XxGEEObzPqUKiXp56Rgoa7NmVIAoZhf8EM
6U7FSN97r+1gE92RD+zt1oJ2O5817zljEa2eZ7vG/wRySfaLMkdcvEK8TPV9Ne/h
uhYVurbqCb50BWBajXs8LGIMIbB/RtNCAB3BgvRqwe78j00W+4e98yuyAuLA/sfs
mzb/kTQYDn4pTg1/XVz5/7VYILZFbceeTNilDzbQXlrWf3c6DvlvYaJbE24hCBKQ
fvvAMgsuoJBTXEX0m6qo2hxt2xSVS2WZFt4+tudOhXoCsap7Wq6VS+oWwy6V6wtJ
XH5ZB0j3d4ZZCLy8I9ym5DlzBz/k72N5pMrvEKkq7Y2ePw51ffzgwt5+v7cp7S6e
onBTiYwmbD07pqET3l+uo33YntVPc2fr91hzYESW7us95dhhlfrVe7peGoFdjFIj
n2cKL5BVWIzT4HmMUzyKzYyDhYW5sHrhi6B0jfuHS/mqvPNkCoGtoGw1wFR3rBBe
ItZcU9SXgMjvjuBYrqjnJobV7GYRmyWx/WL1Eld0yVTBoKrd5Kiuu5o5nhobTpxs
0tJflzKIq0xS86f8nqrotpvMn8FQ76TSyklLZfj5lnbVX0+pZAddwuhUwZXEHBgG
lkkP0zy0xAK2kksUPD1hrgsQtqWq9/HN9r8uAn3PlpWVJtAuGyFOUKEmAdgJtenL
/XUZnhmuBlCm4EvgE1e9YZK3+hDhMQNzwUOFS7UXHqE8Z2rvlq3czdl6naXEgzY6
bTsHbHVs45Qm1fCBevfREUmsAn6kXuL2H+sLY1lBes9TyRqQN7xUdps/yaZloAna
nGYJOacyZ+pt9GJP/zit2RwggGLSNEb+NNkoI0OvQ4kUvoL7W2els3ybRJ+D69wL
wZnYZWeuOUAXSLkQup+tQTg0DA91sfzo5L+Ha53cdHg+Ri0v2jNNTdAtcTkGYFVf
SlUPloCWIHUP3WXKZ9on/gtkWiU+EFOkoEcs/ht0IHB91BG6FTfSTmlM2aV9z9Vv
EvyXZU5TOSMHO3cm/PkoTmZpgtqDaxdLS6STl4VH57nxU2wsjcSHehzHbFBrMS1i
+k2fJ/h0O9rv5YSADQDAX7AoO4RLdu1XOaNkzf1SCikzGEt7kzZBLG4zsUhogMtt
yCAzE8S/xVqQQpRUWxMIlKiAiZVRTydtBCd0893wY0CM9lE8ZQsvnMMlE/VbPkUq
ekDFVeOSHYoFCap8yPsJPkdWIv+3+RJRy7zhlUCS8Rzuzq4Wb+YcW/fDLWjtLHBK
ydJUho2k6HJFn+veBfwGsyXVFQEXJ077ug/tXKOjYBjoP8+yz6R5GmlEsaYf3Ff0
H+Z4CshSDgvh0QE+OBbbU+uGX8WUU7dVFckXHX5wULYWSxPpFM2EsDhUQ365T7x0
nDvjJa+f7RcBJoFXC/pIBlYwvPm4tvSjzV9c26Xk32jGi48jD8dDNOA4DTRsQzoc
r+V17YbDR4IeWr7X8oVaYBMr7z10f+dbzkH2UNJiFfyPWDFHf6uphsp4Joa2Sx9X
/hUWj0MivmpXWrm5XtgvblF0ys5JTEdZwZJTcYswddjpJmQuBCKbV0Hm1HcFeR6+
f9CknlVcEaorpQ4u9f12FW7VMwx12JUBxB8FnqrHapslsTKxWb8vFoPH17GeQz3P
/yyzDoMcLCxBLqnFhp9EFGcqgSOkN7odpPfgflnQN3gJXaDKb1njXphAAkXyLOK3
X/kRDY5JIFA5GtLW5rozqhen3Y5JAkWDhjFceh8K/13nRbXG1OcaASdlykm9iGNZ
I7vmCUXf+/BVTEMu0pGXBBWCEEZj53hxg7dZVcLMPTjuLT16VAYCNkoC+S5uwlRx
V7Q3c0qqxq1ArZVUXJXozIawNZwqhIPKh2iNE+pbFwhwKw0PBTdj4qVAvGVVrorg
e4sn2a89wkkEPpBCNRYhF7aNypr1C68ir45DEBN41ypbDMbaMx+GQFRFZP/qX6uT
zbChaLbxXJZjLpmFARlj5UbRknnMGey4hexln53F999KnpTEDIoTMnZO3ixymDad
rqCMMQuEZVNnB+axq6wFzHes2yqt96wYKo0j9ALMv2u1oUUkKdoG7Ta34fkO6vy7
UALgyOqzuVVpH7yScTdtnLGpZpr7SFI+mWfyfgdbcqA3Gr3DYZLoCn1PTbZ5/oOQ
V35VGPnQfoaCEutb46nFker+MBpTCCrDCt2mMtj363FtNDjyX2b01L1ou4MlNRiy
9VLAzi7I1KvlWrv3wczWBrKtG3xrLWkNwn8KZ5vpvjghdRrq3Vi/t/lG60slraaV
ZK6Gnk6L9rXM63+h1+XVgoCrW8wqZLqkkRnWpzqMplG50fk55X6450DKDcOmUSLn
CnuOQ/V9m7ItCzBB9vrxhg4eeQbFMyhn0nIw7bI6EJC5+cbH+Z1lML9zFtoZv+ct
1EhcII5yEniWFoJQfeni8QMVZNF6APJbTUUpaCgF6G84FaS3qLvQAqqt/se00znf
3NbK54JSE0NB/wuc3vvkjZjo1CLLnqPJfYNGjdsqUde8yiCPdUqPOlBaxL9hA96X
v2q0SN/dHlfk8isTbCTq6eqC5uxcfFTw9z5OBZVzZZlxbR59TqB6yYmXhNdXjmsM
PRPgNJ/qmnNx9gGKAsXq7yVIMqtr6N5q0UiC5MMVDf8jLew2fB31ShrZJVAqompw
kq+amS+tG0vr1C4DhrFxB/UdOgSbVxyosVWZRnb97Zs2aTorZKJ437LeJYlFPV0w
yBz3AHwh2zW1i+EkvZ2biCb4qhlJR0FzrpO1UtunpbuDtyHmIfRZYeu+ty3MHtgK
FX33G17lQ66vDSpdDTAwNz2liaoVxSkPlZy1Rx8hueZdHLc8uy5mtpHXAUjVqVGo
TGkw/nlbpxwBZRkl0wbBIEZRwDdJFpVSf5uSfIADPOXe2KzPi7sAYsjdz8piqMcE
9ZsZGP9MfVR23AtNw/D7kfveHRRUPwTxtfhH6s7ozIWH+qyBxgIuaQWRDAyrpqdB
6VAF7i+GTfnrUJtwzaVXRf/txWEbRHEEgL9UhZpsN30PnLhUaMJ04Gv0RFvPiWIg
oRK3+dRd+k5/xUhzSd1eUBD/BxKFlCcEdiH6td4Y8dtkwjV6ruRrT0y7qMFReuzH
ExK1SWQcwuWH8AzVXK6hlUPNnZb6hVqH1iPlj5lMTlqbsh2ksYOl1KCeTXG4Sv9Y
kw3fXIrTG69eDm5npDXbtXXHOtxTvIIDv4P4HjSl7mMJCzhFvXyLHlbM39VEVaWc
jmncd2HDpnrPQDviPzGa90CyRRzq+LC944zL7kWgZPuQjMjY+uw3L1ABo9QdFx6X
Eck76U/8arpA51BvB3NNj0P6su30oHK7uP6Y1/VrmnA2yeszOEZMTNecHN9DGiov
3VTH2grSZv8vThGt1GpZ4T8abgG44rhTPgl7ikNaNGSqUB/UJJEHympQT/czjmYm
3G0fqXAe0J0O3NaG7w20Tuc5qPEGyLSYZrdHuxLAooYuS6pDReviTjI5NRYBrj/z
JOu3MCCZjHQpQzQcUCZ5geaNlJduAfzo5EkQVKbLKRpcX02QFNEd5EZDo4Y3Jd79
9aQu63KbuCQ5rXjjCVxu32RFjHu2H7h7s/VMdliuFhxO40bbBxffk26qoGwpQXsk
TN1/mFQuAaWKn1F64n1gzyFPWU4yLKhk2Z0w78Ptv6J7jaJJe/qk/43xNMo9vJH2
wrAf4JnW6tz2q3rqTFjVknISD6se6/jjetpibxe6TKCfE9XEtlXHhxbKxTmU1K0D
dBaXRTfCRoi/dvMQuE5HJDUV/oV/FTd9kuhD0sxwWv+t9NqZe//WEpbdRD/f4HKc
hN5T6X3JZVPV/wgsqyWUg4zp/DELTVSnFDqn4G3kqcLgSRRlBFeI5sCml5kHrcc+
FXzE1qeQXkFAP2+qUxjSYajXOTrjH0C6kaTZdPIlbClmF3hCTs9gjpnfX7lpi27R
ZYiQL6BXQ/8R5wyUV2/N7KvDQDtuMndmqtcUsHGs/Fs18nw/V7HNpK2hH1JfaAby
WGYulzHn4ke531mAQ3cnXeSsAY4hBv8GFdyy9ZhsFeUJSbmhlBiY6Kf4I9jnOXh+
9THtmv1r2dtQe8t6Zgxz8Lv6Ck5NWwRClEo4iVxqGzqYTmanEFadrfTw7n69j0Jr
t5GuiSZ9rW47M4bYvQ8wXMKzSKbR3UrF8GCkCSBv//hO45/CVz6SsuisbbUuoT9f
tYQNB9d8mU5tVRCmioVwhLpbZsY/v0sbXdmqCxtkb6zA98AU5Ix2EfAJ06cbbjoo
A8UZOheO7QddCSAUZ2NvwzvPCH9Hac20q2fPYkbS/Lc4ja46PYn6y1/XE0/db/6l
kt7UBFBOnH1EB9lC+D/I9bOr3K4jWhFuwrxzbvP8e+kuSE2tzL/Uag4FjHz14lRu
BIEENQ/azd4Xh4nShT7gYRRNAsLyU/lOaWHhkzGuHfjq8FhujmnbTbrSK+FamC25
hbbSLIlLyNgAxW6KJT53xXsApQjIuW3UmwpQzBbphG5cQ7pz19vIV81+nbEzquge
IKNTpeQp4AR72t1WxWKBP4ck0guKZb3zSBp2BsEYycUYA1uPo6qTFiX9/xnSG5Ny
zXdk9SIXzXLruRGvdfjgodI9wf9EydCyi/VXuHxD4QPxfnGucd0ra2f31Dtq3xyY
YPQO4vP1qghY0itqeLKoWVSjNYw7M/LuQdEqbbLDaPsNQEtTWqIPjIw+lB/P4Kaf
hfrKQXnl1RpdNQ0LBd4ELxghTHP33MzGuy2fKSeeZal8lNGh/Xp9cHwjDP/0VKof
MRo43Y1mNZFgNlfhtntgjr9lpt5l73noXt3SpbiqpIJxalkxD0weAiC6sEHMGTie
hFX1CwFY+ljRjY9su7thP7Es9HwLWnX76id0PjUksIbFQeiKLpr/K+Hpy0pjpcZU
vtNEusbQQogeFIqmcLvQnvFgWWjK2NdRoGQQfJVDr71aVMSc5OkDYRbbdeRm3g8n
5EDnzzQw5Gz5JfBHpbu5p5iQBgPqdAPOQ9ZLrpZqUerz7Png3qB/JLBKH4EO0DVR
1wxEAMcPJnhe8Mg2h0u9PfHn5AgrQMNabU0myHOCzFbaeJZ4Ly9dPV/bIvwRr7zt
OqxGufiIlirBhMnCCmYa9a3XP0SntaOKtt3I6b3RYJ/+cq2VmOu8UjSDHg1sFYVN
ViQmEkdRZY12xY5bAjWgpdCinQr43KWHo/R8Rkbx5qFgQL5a5ZSpgvk6U2ahhVXd
MxAsN5oJp6xQPTD6xPMfngWPYvKPwknF+nl68Z9yWMaugUJESP4KUsZkljYvOddo
3A5bnaaxigyMT9FFTJEw8slyo5EmUcgoon2/TxtP9iLU0V4cIHdn4hXN56WKH746
nxQ2ID938NIFHS3XzujtRmJ2nP6CAdEp+KW25Xpq3nao3OvFiv0zzzHuliOU6y9w
WXqA2x9wyfR/UgLyJmGL7/EuyVAc8grdcopn1YRxxmHjZ32kTTK5IkIjpS+1MTHO
R9dZA+trXpYK2QT8cRyVEudaA0tnUXaIrrPnojc3dzhzGxo8y7yrpVxeQxXSRerh
uj0dK8fQj2B0nJZqSk4iLnV31LJS+vtVTiPLKQXQLZ08YUapNph43upzqYWi5KmL
o5ksIHkYcY4Dxb760VYvj7Y46kjqiFf5lWjMo1CTW6r6Dv21dyS2aE17CtgObh5Z
Zf+3ioHSEWtKVjJ8ZbzhcxAkdYR+pnMEXEpZbFxWiRANM2c+KHbDzWt9HT2cCgU6
W391aZhCDZGKeShhqBempGvfgKbrJDecbHuAdHCov6rpqnE6Ee+MLiY4n44yVVw0
fNTdx2f1P2f3uHHfyQswiWqZykvwkkt2yWskA6oNHZyqZKzjHrPM0pIn2WqBXylm
Ca4RapSz2yb5JCb1KrdNAXxdeWwy3LgRvPItNKx18gJaRLufE/VpVnhJ4caVXcnm
8w9rXZHuUS7PRWuG+f3LG6LUy764vLA6KSeiiy008uooKcyAsZB9WxYptwYOW63p
nYovxP5Elq+ptKMuP5izr6Ax/GIMRjEoUI3d9Mmk46Xyvvn3oTnqXT2BHYESWvTZ
3cDQWsipGub1gKr5l4CBYzaeRLvJV5FB/g/a7QMLZWFQbIBxzUQjreRnDzcU4i44
tj8JJguiTibZXUoqwekmI7sRxlHsA9zkY/J89ePorXwnT5GUzXOlA/1+9ipLylaB
KEiwq8kf7uVsaj6/DP0MIvNH0uTC51/Sd1kYvT71gToqKvcxQwr0MOKaboP4kDcO
Ao1gwmmiJF+qntFt/zSu0VnGlnBk3wFb07zNSUxCpXOhwONtnUXr1U5sKR7BeGVU
2ffMgQQ+2M9mKaTuvPh2vR8JPO0QyjQz4xERwLDzb6pyjMv3ALQ4B8Eecd91NNYI
eIXtMEzdi0TQEqLsoq+TZIxOEs5A0bZCDIAdnq7HJ3vsac60eb8Ja/+eKxIZXRt4
0XTzmRBUot8cGmBJgMWupwJVoQszRYDkgyTB1rfrlL/0uIVTKG1IuykUDHwHQbgx
qovW+H5hGrYQfjoVBh8X0EZlBj9CaA92LSYJvi5fXqNuW/pusNCqSZbfaKimLVam
gS8XabllrUE8mct3e+XBJWKMnvu0ep7TDdKX58BBbTdzDvkKNY3/ucX8spz06giM
dzc5vgT7G533yWmFcv1MoQ8Ref643ZX0furXcw1KepJGrKz+zmSwWjjzlA2GAtCE
0xVZZmxwR2lL4IESXqJjapRCow0D6zJk/Y96CZXi+45DLlGReWWN7AyupK+NL73h
pLnfGjNM83JMFr9hbbo44QOUfeEh9N6AxLPErwmjy9b2yev6N6SCTvbt1Y8ep3ah
gVJFuKs6TZlNYEyntOJZbuHtwsPJpgp+5SSKxmaBq42tpWsk3wVA/MreWR0fUPD/
wnV7GpI86d/EcGLNCLiQxN2pRLnlTBNl47rQ56NvqjJShKqIs2q15ZbYuyNRcjPt
CRaamekgJw2KHY17fGwsXhaRTp1zvKdvaQUTFeTqpsKu1jEg1ZSv7LLC9A3JKwuL
u8vsSM7JBzqY28z8Qgjbhkpul/WD6ncAOzWGfZzOMtwvay78j5BlIACgBjIViyy2
MpHmBIpEnEMl9BOO5abkxGxlDkpssjOrm2aO5EgRjSTG2WMPHD9l03Xje+0xe/B6
wXPqC+BJF8tCJUGRLvKX2bXOw/Oo0ld9GMpEYMVSJd6nfH3DkVxfxSE7pTMhO18Y
JqsHNssUYvZctgQu6WyExYwoEHn4rII4H/iVVfHfzpRcY65+aVI9Lk+sXfvzPY0B
FAKKkf5NwncyKj0otp1pRjErlPNWLAgGoIdVO4PNnWnWJz7+GxNlaJRAonsuMOsD
CS6P7qc9PEkpdqFNzx+xZQpOEszJyHtJFhnOfBaabanGGe4RM9my8GTjmgJb8v6U
ZmrQ/vofUKrvFQyV7zDLa+irkOaRjyJdDeKxbgV21BuDn+5fQM8Vk5/XgpXy0SmS
ItduS1DL7x0xtKYaNFIwZWOdMlFdIiNaRO/hc8lxtzDOsffWzZVWBLKK1hKWl69S
ffEmZYOBUhIREJvQ+MHRQ2o6ckyBtUCUtMy4XWSoOyWrENu5bjDdwb2U6W1ee/2P
xx9poWCvHR+ca6LaYAmG5dAa1gUg9KLN5JPK0wJGG5Jc4/uYS/LNgUk2ib0gVTlQ
I+YLwfwr5iCXj/lFS5l3p7rBvVDL6koAMZkaYxBbF/8VoR5sux1DTR3D8m9TueoD
cYTkUlpv798J+w9jYQtjhgUsfUfW1rkJpGgpd0U7+/asFJ+hPqOaP+35QtZDQtJW
v+16wvc5MKR2/9lS2Tl7yrs1QPomPA/+oCukfaql2FpPKRY/44lgpNmflSAQ2ukT
3d0bhinNcqWa/elUcFWgMz+sqxt7qzQuI09qN+fXO2Y5fmNc2vbkgy3Eb2KqH6iT
nGiILHCspDIcTc21HCh/gMcYkSJTs80+1EaR1nmRkU/n17FqMdm8Ro4om4w8+02O
f9Dopmx53MD6guzt4TGWJVZydBo0KKvQvZBkMVr827/7Iw8l55ACEFEJkIrCKqyh
XO+vY9I/gYldL+/3vB6EvhobV4GAkzPUl2uuo9gPWEAiZiMuN01QVN7X36SU9IZV
YrbnOeIxVLrcQaNAMDtkTk0/G2NM+M4C1T5F1UGNqvu5YYAlWV7Xm5EtUMFDKQrN
ZYK9QiuL3eJgLAq36InNdMfUFdGkAJMZ/R5unAnNn6fcm444EjLm2ld1M1JQwddi
N2bGjXoKlmldqw1MmCky7k/4RKCxOoRYsNNEp8C/Nfz5woO+EZ666q7o3kb4Rc+2
zm3uyeyKARJlNvMEFwbrgvmAjEmgcXoJkT935zGc2+VV/HEVIQSPFWdKudsNpca8
5xdHAxaNCiaIXn2c7eeGlAMvEdpeOkaHjJLhKIMBVykIfGkKlxo4T2MIUagNQnE6
8Hi1YeAJBqNuaUi2KmlGQZjRPuRlgScT8oBOoKmDPb2Sbq3w6RlSw9+jJUo9+wpm
ckS2+PPFybEgAbs8Eiy8dfsjynwz5ta+UjbiZOPD7TZYlRR+PQnd3oyZ7yaHNvTm
ecCSMzjAbVLc8Ia1IOvrzlTPn9D9MgJS8HBCoTWhGqGSRahucwSKWnaq8j2iSAhQ
bo3r6gxBaqcWkcsJAdt0Js25C/cYrcHw4Ylf9cuWtTdKBlbV3ODMDHlPVaOWD7eG
eyGWgGe4aEiy/Djw0Mhx4fU5tvkrzpBBwTiT5ZunVj5i/fDWcy3hTVJ+hCcnjAkN
zIcC/skxCvEC5bG25iRfdH/Rt2TuUI6sw036skkG3CX0f7JQPZ0tAUvFjWKZwgJH
B4no7DGT2aYmbYIBNWrWxs+Ledz/+qh88zSsmlAqXADyYEBNqVFaFyGIBIqSvUuP
fqw9JMrMb79VTTaSw6jtb6PfKg7O6bLYSZkYcl7LrcpBz4O/KyKp6voW5EHJUZRp
TVu14vlr1yHsAdX/efkEOd4LGm94lNaNcfgJ+y/MD0HWPGJ2sZsX/EH6enY1Sh+j
bo2+XjIvgrWfc1sBRZHWXttYuCZpDzFVFkO8vJMgRwO6cpNtnAJ5tLBy6Zl1FVPl
yLBybiTWUb7Kns596McrYLuNo8utvHzYAY5mW/NTk2vmhHThwi00n6HdXgYbjpp8
fyI61SoWhXu8zeYquP5AK326D/NizVQmuou+nsqE90TOkFXNGFAzshQNPmcfbO0A
vNY8kqw7DndmTih5sooXKtQdnikcd+uOBrWoqadBrSXCIV6TI7X3eE5FrAJ5ZPnY
TAsfiyQ1I8joESeurAgXhFONvsMJtOy2M2geDuLThEaRvUvf/Aec4qI+zgKWwL+P
2I+OdNt1km+cFh4jZz/3wot9uejv3IQUO+16CnorOuPV0kxOQW9TkdZDkdGBLmfQ
UdDbt+jBg+/57Q1sLFpY1A4jFkOZTAXFg2n+ewc6JFeO4X5kBbAwzH27Tb9BqG+I
iHh5rxBlWopsmoWMVpLejStfmWQvKqBwODJmBULea72zhuw6N6l6KZ7A+TVbwTec
yUYoBb7TB2MM7xaYH3ZZpq7NGP+RuLckTzjfMccqFnm7LbzSdaJ2NM262stwpnHO
e2Kgor1q9u2ik7pfGwmx/bQADMClugGGocCkjqRiZsSpU3LpvqIusuuwS0J1vuO9
SBy6mjtdsx03IIfoXVdAaCibAvM4K+KRuswrgB5CQ4Krw0eqOTi64VNF2YG7rUTH
UUadaafrNljfGyACD+rTXFMJ2Ut/CKYs4UAZQDSKu7leuUYCrZR2XQsFqqp6CzXI
M+w3CxEYR8GqoHe9A9up2RVpGIIKhEi/N9mSQk24hAr63mly/j1DqAaYfMpBvXwx
tfLDJL2l1vE1rd7cw+09z+GP+UKoi8bCruLLC6u4BLXse4dYnEjMEE2fDxRQY6qU
7KAp+MK9Gr8bzVxXxpTRDgMHCVmem9hBEQLLUOSM8zWkHfUe2XJvefXH4ovXQGnh
V4BIL4PIgaUdn1mqk/QBwC6/g26BYZgxkozA8vCa79sZ5apFWtj0YlvQvc3pxtKQ
4yaieNljzaQBM/774NzoAHAtZxT63oDmbjUl4gb+k6YvD6bpLuP7e/uAjOlZhTtz
fmUkZx1FzDKR1PCMoIREYw5ivP1VIEhW+sxzq/wHUzLTG3bz2n5sRtOpH1pXv9oN
o6SExKBHltHRVPDkC+wtnZF1rOlnfAj0YHf+UWo0LYw8LezLjeVHz2r8y2qB7+9R
202ukkPK1CwAcPTLawVl2MfP8AmxlImmHK1JeT2UlgpsbHcMk34/PteXaMSzontm
SSVfzjzM0HSDH3CFsJR8Z0UWnKrQUgt5a/Pf95JdLQjWyt73lHgxCE9eDCUA6I/w
V7ckFYp2LwZroESShIbND//9Y6J1m6/CZONX5vh61uFP54TMpW0T/QEeJNG0IloX
nyu5cpar6/JWmLJBwImvFAJCygJd0oriwS+zIoLnSja1PAC/aL3yJgXbYBFzrrDC
wnZqwoYxHcvnuZFPvgMjJHbVTA52Hf6/uU6y2VA6IKXzKIN6ffdr3tUMcQFoLsDI
skfXYnQPTxx6QFdSGQ5oo8HM1F900VNCykO0q0zrULVvN7DOPWstxgEPJJYhMMR0
AMJODStagGGFNi+dnaHHY05WQM1/8Rj0p2wWY/nEVt8hoed36PRvfGnDz0mtnxuz
blR/gd+eHWoVTVudWTJE603ac4ytyjDPHeClvNTYO7s3bI5d6iIArTgYDTw52U9S
cJ+XmyIiKWm2Kx08woeqs2D1roSQeU/JthPJufELiVcN+s+1sP7PA9XnYAboQB2B
VGx8tU1iKcH4aYTkrqgyPvQ0cK+DrNKrX8GICI8XVS6va8rVNl4vHcqdR4mHB2uk
pTaALhQfRFI6Jjwt22oKeSKjv4xxVnng1SpTnExav2TWJ+pulKiuOColR1KalFKL
yUROt5ourOiQqj3Sh7ukk7nbfat8/tYsUks8VECmz8RqgkQrLpqnNnwB+gqOmJqI
yV3oPg/Iu/E0DFcKJ6Smrj53wneZS0dnogcDN2sbrQwhDA0Kl1iWG9smY04ifGM5
lzJ2BdlZ1nrz1gDcOlzlDxX2iuiRArXDs3IrniBS4RFbMhpABSgOtMBjPzFkk9H4
vBkUoJKyMzoAwio+JSfwRnqt3lBLDmm5hP/qXeuDfKw0evxxF/3INpZiLGIput4f
HskcqGsmIZiF8FHTZK0pdtHKU4Q23rOcG9A6oXrXyvsyVVLHSj/7cftKJrzHAjj0
ucduYYt+wQ7sNTsl1nN95+pkozYa7KNZjn2G+CYILgYRXIjksAQzhTgC3VB4a4aY
A0SZKt4jClO4PMT80yEgpklN+as4BJ2tAIRQKFPi1Tl9pQsjRcbFxPHE8A9adFgh
6qwwHymIr/ivbZFOlSPWcRKDenPoPn5jsTPDNVM8AIFbW+7MsdSWaKD+L/yHMWjx
mFm23X90lkklSEKuV3jf6jf4dAHs9T7zspaB/8EedUiVs/A5S/h4UzT0EXjcWYSj
62eN3umOVeaL7J/V7cTrbFFSn3+S4X6ZULXPnWCYeRO2W6baKsdjbmu+BT/cCyFo
BZSwReZ6ze9b/Rf9UJTZLkd13Yl2UszEyq3BJ0efBbjRgtRHJzEvC2hJzZq3PSgq
Xze6eahPtI8/niTCAQWlPrD1NVNfB9e2wuR0gu6ZOcaDaP8Bs3NYIdAfqTwCp46L
wK9BqN2/e6zHsbAWkqQlLa+A44esZ+SXLq8GSwrWWkVWuyh2ezTm36LQdUZFlwxM
ynZGp3jB9/eOVibV72JiI1b6mxrHH1/RxiyQOsFBxt2GZ5vgprKdPSaQscZHdnj+
TlwEOIH5tYT8nyQF53/jhL09EiBgiQ/c/sjTuZN3c/WPtrzTZuq177E8EkQtF6SH
XcpS4vFSz+vBzb0ZqLcJcgHao4OV++m+dD5O2FiDeb2trryDEHR1BZOEVb6/w6rY
v3RK1GjooJAZdzYV9XBON/LOt5/BOl6Sn2P4H5zd36Ol40YBBtI2Wd5f30ELzPjl
RbKYpczaj76sHmIMqDsEgyxMxS0+aJgt1SPGpPFfr3eZLpWNlC8l1BhgGiWeIC8u
JYcW4TPRRtmvyI5CTPeR8IOPwpq3le6fgLoW8gY0uVCSpks+rpJVL8GZ6GredeCl
2UPYVnprDRF0SfB1l1/ZNE/id5P4t6TdMFpru23xeJ86kKEP+Z1MX+hohlrxc9Qq
KtNl5nbot1KjcOHMEMX7+HjYGa3yVJEAio7dtmz8SAgnCQddSkJ4yaUijEnPkI2V
E9t5BQYJ7W6T2iI9kJuH3R/PeqKy8lg3PPQaTJBQE7qYP9oQklY7Dg1muCE3Vpil
A5TkX4jCp95ocHIE6aLFAGhx2EB5ZRhwvPgZbayPT9q1J9vJcE0ggVM6D13oK59w
CSw5TbbN64h6fckdhQCmP1nGvruK1nXsETLFdqsLMbYblFR5KMhkHdg+HZSv0TFh
b98NDNXduocwLmOU5maZRAgnGXKLOn2uqSNh780MDR0QrhAf5USfBeO/MZ02Ed8t
fsqhyBhmZYMNcY9IklLQJLumjVj02CC1OPVwbHtys9BishlNCzusaxJo0X+hAsbY
VOWWj4hlv1zJ2fVSX6nvjqfH2Q2BuihXoaldtwyWUOx4idYJWDWZmIl/qT1FCC0t
rAbMw4copitv1eOCrNrdfq2aaH/i54Jqme86AFbUBO+S9TkfDPaFVWAL5kZpzmtr
s7E7wIjeevHHez6TyDOMOXv1TVEC05QPXla0P66PamuaeSVpxtBJTjvfyl1ZH1TS
YvaVH0uZPAF5T5eMCaUSw1/fRS0kXcynlLc3luWkZIwtVJXPWKW+aDEvDUpRs/Gf
Oz8mTm5OnOeDORh/YVyDpmqHrbOvB5gI54Hy7icSS8D3VdhcpeW6FlASsdLWUHWk
3LUUUY6zvwmJyUOaUaokynR9srB1aXC52BOxfzx3Y7nCoxpWMGDsXFBjI+p8xdJq
V+5PnuVLvLt7KOXaRhhR+qXa7hT3GITxrbkrrVpYHlT9My3M3T9P3QtVzIpUxJfs
MRIAsQf5Whyvlc9XDt2ugx++gjtBYkL8vV+w+1TfYfIEOpEF8rb1tbVWCH3VxNtX
FMbFtePuawqnsM+mnNk8XcCOtWkckb9AALhLx+eUb6MdnZEtQmqPmTk33BozaA1s
1Vca2C7OSG4wyPOrF40X/DdVYVf5hbR23b5h3wl13Vu9h+AKr/Ef0ZIhNj0ud7dZ
fdRT1ed7bLrS4vPhLkVhUO7YRv74HkRXUbtMvf3CLGPPUlPST7gvzxt1aMrU2+M6
YLLS9V8LHVlSl1XzbqAJbH2EM1ocABL6P6DWb3JhUdN1McLeZSkcpeGkHkPJRA8k
Y2isLTyp19pBFou9p9/7ZonQUE1wkzcsNpZfwFCXFzvjMQHo07+wir44kQwaTpym
vn/7OK/Cmw0MItgC/coXb+kRQV1uZcmI+vkKPd1823IhIGjp7WUkqYr6fI/f4+Bi
ZMirwwLPsSz5a5llJU3TEKiIjcF73t/aUnmfm8FB3mKe6LzeZljjJKHDOeTkI0qJ
bzvDCx6MVR68heO4vP5FMyFghQLrab8Zo+fz/rMspTk+Ce4GU4sV5b7ahhQxMA3K
wuEgoh1BVg1xXw536Odmc0ksW0JskcqWZeFrIcyNb+l6wo6LKvFiJupT7X7xwUBt
mK8NvD8JeNbyUllM3+SEXaleo+C2c16SpfH2rZwZDnkG4dxyUsz3JtU4TTptGNWg
drVwEVH1z3fspdxdzzZc8/HKhNPtJUftmvbWNYAC7M+pg/ALnvwUcOwDTECfysqg
R0i4y4a306hn6f9/u2Q5ph5eFTmfEZi6pqFxygY3q+B3blJm97rdYmavcI0WnYzX
zWvcWkWqZ9pvL0ZbLtx9fLg3vo2jBvT1LQz4SlxdBHFmpyl9jZo8fdFjrHp9K4Xa
xvbTHXQH1ZurSr/2xnfgzSsQO3E6sLSH4QypuPrX3tXQNjo8XGyPagxjrhqavl7O
vxU2LU78YLmtAMrXdt2HTSwMTsDWS3EnefT54VJoL42MytXkaDo0cqTOVBUodi4K
0OyPdAJwq1ZHDNnUg6SZkqD8+e2CpS/evC/oGXa8KmJOO4WAG+jOk+A1VUKr3yAl
4dc6hQKHoTyHK2aJjViOvFahW2uy5hpFv3klGxee89hunhqOxaMuzPwEnrY3l/LF
ONDOZygKqaBLlE7N5SQDg1ziGhXpxJEMMxtjuZ4z7/GwAPFH8HNubAhR2673xLDd
HW0z1+Mwc6EftpI4M5plCGhi5PeVeBjxHlQ0kP6oROyF4InNMqJ10kFWzWOILjqh
XaIsN3AQ+7kLDd+YnI0T7/Y4ueYXXi/YmpPZQVpbssVhLvwzFe9AZe+pzj3MEAm+
tWbHBHzLl7uBL3gzJwgw7dSDJNeibvhfvPUzBUA20yL9gZmKYFaNwKJsr6iv8OfV
gt9+To/I1Sl0EIWxBx8cryTUKzBnjToLOgIYAOoqXKOatDGigggluXhIA469lxPb
9RIiBhKaVfX4ZRnRA5ADSpXEWsVifzWyyXElP3qWVYxmX1ZcHYzb7lAoWYAXdMJY
xGAW/rslo7z4xfoevZuAGOlj5FYhC6qmPfq+raCcFksH/5Ndm1lei7i7GAh+AwJV
N5Tvh3Oi+fEPSqySBqvcfMeHVM1dI8k3d7OmZKDDs+bIkP8b7RvPcjP4rmjr/WTK
DesMr3cxVIGNyK/ybRO3ymvV+wcfk+UduB5deMFICeS2Mpu2ALaOQjm6BkhlEovJ
hWEXzDRQ7yg1Ts/obvKZmaLGpFc3Q65NkEaEK0fkjw1mzoxosdclyTEQMXShKsmw
70Pt85yWQ4oZ0XYMiYHdSIGdJGOF7NxTH/PTfNHoXlX2whVt3rv3bKn2a8M+47S/
bLaqhrEj98RcmlWgKuB+z5O0Muj/mo8rDzNvT4dCp3VY6YGlUPaDflDNydq8Gft3
EFz/OjjRv2oyzbawIfYnsEU8uYMyHZ1+mpTYm+QetDsSff5K0x2nhbDbQiEb8BRE
Zulgdsy1iYmGuHmvFkATBV5YMfdXlyD5A5Ogt0fcciKJPv2B+6gD4+HfnQhRc0gp
Dn0Jr7nPP4wKMdbP3scaul/xOWN3+pN8ylJx1dl0Py832v9EAjA4ZF6zz0A/xAvJ
ogpbu3636wTRFJlPtoDGT18DifLrnog2kuAFXRM8xR6Y3I/FlWcZ7lTyByt2WGh9
2g8JfviAn7t8y6Gw18OVxkNlsb1NQXKdXQwoP0zpPbI7/qoU3CEzlNPr9htD531c
AsTigfFC4mt3JTuVPH0N8Vm6DsMqUtN99+O6KoBnTMXF0pdU9FhP+KHIfaFRsL6j
UE79gUhcKek3We+1NIRc7zYufZr8MG6NaEaaVO6X/gWaKCKMbE/rNbCaJjKvpUOW
1qs0fwQxAQJ7XipNMA4VCiA2kxJ2+WUUvhg0+7stLuyXpR7SqeLpo9se7rfwzGLG
PjMsiErXKK6zykbXjUqcV8szkhDhSxZAiI4IYbj/kakmRWr//w+ELHzX7WkYuq/A
syil80K0Uv+4oD5x9vukE1B+grVtWYuF7njgDty762AbNmzhZUhLWWJ39BXDp6lY
yVgaZcq+ZPkf1FyoxDDqUPuYxCXXOthzYVDg5qSgQIIo+UYQzyMTkzN9HA7VXDBZ
vhW8E6URl6FAWTzsh8+oTHJFLenMFyGzNq9W6O8kdyWV2lc5/Sg2hB/ER9YKr0Wi
scMR+bRthduKm+KKU9/QjsfQfAuiMLktXAn+dzs1cMCs9QXlUWChmlP6S+Tdzpp4
1F2c3IF7JiIrNrd1edJ8BdLf6qwCR8KbOfwNNcHSmG55MoApdNVH/aSjKvasMV2J
3dRhfRixECu4T8lQK/toAZooEsirfCFe/9ebfnvewVZkL7KX7lThQkZouqrO8dAp
6lkY5xzx9Rjcv0ndp3p//5wLxp+CpoOtKEv2YvdjYA8xW15dB1wrXIbz2w5TAm5o
J9nZTAx+lipInNQOi0Sul1RQ55qi18lhb8QpE1NPZOKbt0kc99p0PowovaXTZW6/
yhwB5fzoaQP4M5lcs6XsFuio2VlK6ys3I4v9HJRwcEDJ1mseY1Xn14E0xQgBc6Yu
/egwQTjsU+n9i5fmNWgxuKa+pzwvLvhNHe+zFq4SzaqcPO3FxMs2wpBBHbfkt1dF
sepLhMVpCp9em89eoO66MsWhJuI3xoEJ2IA5kxh1VO61S3XiAxRRsKi5S8INN2BS
xoQYix5a1X9QC9YNNHvBh+iNO1GYPhEin9DVJV4lz/ZdtdIe6R677rv4hHDj7+zQ
cZq7hDLx3YurBcAqn29GEqO15gyiKXGttmDmu52QGHOUhH2uq1EhHpF+3BVmPsLs
R41NVF6rNbQtaRSNRfoW82JKiUzwLFSaF0uxGVo++5d9TE3aB9ptb+fbNCQAeAFB
Qu5mspMU7MjILlr73UHcxQ9YAe2qFNC0/+5GLSAxf0rXNmmnAoXyYZqq9vN9gUi2
tGR/GRwHB4yGmyyXJxA4FEg96aMTOcuRw4/+TgePY8tkn6MSY1ddfl3vklXZ2d7H
ztUODmBDMlgTN9mqleLaHIeLbcL8S16Lg827sV6wN/oJyrdgYMRaUMoXDZPPx1yO
kjPgo0Pf5pmINgkXgI7S2iyMSbsjtMjbLKf6+w1EtqucU4xAL9Bp9mxAYk2/QOB6
GfBBa4LIRgRKFlb3UaC81DDLHHzYaJ8yeO8/tHV2vEZIzFoK3LglE+uFRgdZs2OZ
cgTTHPPGkKw/T89Np4dHm0PPkfVTu7VBPmgBGQqwWis3EWZ6nLBfl2+UEUynfrcl
vlRNzLtrRvqFFCrF240DlAC2Iu3CZx0Be5L4YApqmyDvPvp216WNNkLTRsQsjWPJ
EYicGiKtud2gBmfsh3NSZWhALMbE62W8dokyxw2WuA/maBIJnBtI3UlueA8l5ovO
udgoY/oF9HFelsOyeOak2SA+s+LbYv4b2K6kzlUKxnELscxPqSJ/tNdz1ipOKj6q
m+vuH/ZBR/iTCoQaPeyEQyRJ4JnxqDGbu0QGAJf9m7u2SVVrl6EybpkHFvo6bSC7
XOD/AEQRlQGWzA8wm7nZvx76xUkjyxQnkD6MD3ndQnvGqxPZ1KTDI0CuX4yrErFd
NkxCaF25+LIY7RyA5+vK4lvG0kiXCAJi9wH8eRaljluHUtvvFSYbWPQI+6HPz+Yq
5XeVdmN2RH0Q1T2xYdIHkRMN8S4mi79rOyiABKjLGIkkz7FF0/g/Ffaqyiy48WDN
GQdteg3m7j8DLsLvQLWeVlNxfhGG8pA105odUZmxrZ4izR5G0gjTgPPr4ZUrZ+LQ
8FqhuqjljPFVhO5XtD7bK1MrE5y1o1zTb6wzq5sNtG0u/wR3aer9qlpLA4P6+rrV
1rqR2QFQuyinF5XaWTjtVpZ91fJgjfaJU3T1QbRqB6ErDRbvvHzjhrcR8+jP27jC
X3zUticCgtmde0xbsrQg8IhhiihWc+/dFdKTOYV5lgC3o/1v2vjJYY8Ny+oOtGqG
w3SstnVes/rs/vAZ8QwC4+XWDIxHcETHH7YOkyRHARXX7FyT9Tw0Faw/qTCg0i9v
kxsosmEcMoojFY+zCM967wX2dCG5sJ/vY155cpTjrwagD55A7c+X0TG1+h9zZTkK
b9fYgvaqFN6cT8wNPen3AQRSiEdLqhPNckeqjVtVASF1ArVL/mXp+rUwVUfgmoGi
/AVEydB7jJyGuCP/deBwzZCVeMpB/IIFEPxeoZo4WhkeIaF5jpxWAenQW0vKfaO3
BgA7vnoslkyYv7pPlReiAU60h+satduw5rCqkpxQzEAqE7wQbaykMcEQd/SM3lIv
EqyLdB06eUz4qFUk5m0wAwuucsZoOmH0ro+tLWvqk6LcfaR/kKvIzk4Bz3GEeOCY
MnNPIw4FHIbnJ1EzAcN1jDF0e4n4hPtxpsali5GGutgDuvIE2ihUaRbqUEhhsrIn
4SZcgaZsThW/nsrXpl1A6D5R/0eUuq/+ifxqD7THRghre3zj+Tpw+rYyidhY3lZG
Y6AFfONB8Q3I0L1ZxVkxwbVGv+VaD7GiUrZc2M0UUb7p58cX/a/E6k2c8f2lXHJU
yilAL7oLx5XXL/BZpc2cLAhqsvF3f+Oxd4+P5WVQjR3V0vjfunapuSRxoZ0uW9nb
HN348lHCJj5zmi+igv0NZMWh0Uc0RIXwMlUM8DMFkQ5njiCChszuUc4alvoJdafY
h96Noq4KRW+/bZdgV9C/fegKzGb+ccrFDNB9hqkoDuh7NncaEm6Vf+1UBZHRNlqp
TgUrw2yjPzq2lVXnBEZa6Ru68d4mhL0YFxo4U67IWwdnAeaKcmIUHcU3dgT6nE9z
itq7gC7Rn2l4P9t6p+3MNHo+5TXRf1Qc44a0nwgolCvXamQy37uaPlzoc6rCBNlC
0eUJdmqGhhEOC1OgNLHKUv/gHKiOFEL9aUQITQOPQ+wUlKGfMgC9WpL2svrI4NjK
2Dil9DevZzS6xI0MOFBnX5UwIPdFh07qbrDHekhnJiBILD1oNADWzIJ80bDAHBgb
Tw1rXAUfXb3M09UUjG/dyGeugpzUEsvrE5ZuDVShqYbh9kPg8mvlOdCN40Ck963d
k9AznVaOmyQwicfssq2ysWyHo43TOeHrol2eMSgY4olXaG75Q5g9CXwy2TLpyBER
hizWOuZME2dcpOrUUPyAGfLaX7tLn1zCq2gDEyqJa+iPV0/rxaHRwr1QSx3w+cWo
SlH2REwr8mKVeo01pVxHeEcPL7ELdCTJyYkZ+ryLwkuYis8J15K5HdI07g+d9o/v
Yj8VvnXLoWQZlUzSVMEZfUv2BLEEOV1fRm7YeZ+bH6y6ZKS6o1v0E94t+1gWi66e
nK0ijAFoo0cxTQdjI87qk96Z9ok2GMDYbUl1F9UPnQ5WgnB1oDf61VTLnHhj1MGr
ClyFIkWSBjwcaR3oi0jG0UaC0b2C6QVVlRh3oeX7t9SkSwMCRbv1O+/ctpB4eM5M
BKpaezPmu0iUCopIp+3HbsiyeTD2wkMsDeIW/wrIbNGrxETI67flDr1WGh9sL0gw
NV7dG6LuqW3Np2bzNqKXNRAVkI6QBIT7aT4ZA4xmdZv/JkJHon72yqpsQDvYRdFc
PIesbbi5NG97/Xq4EmtfpYPTMX3QBW/Orieyu0FFdR8lY1PRhqv3/ZDIBe19KgOg
7i4nwVuVg8BQ+CsVVuOwxjdsjt/fbckkzKJ72SL6MQDURhkNKO3TvxvXou5xRQOt
eZRsDfARxRF1Fxt02lximnZDWcAj1crxAH8O66n8TFpEQY9k6bMKyf4gbwmTqZp5
P6eut6r89ThtPBYLN0vbupQiuKEr8HSCD955tXb4auERZGxXa67iQU/0R2w1eEx/
OLnARA5tYXMRiK7LhXugLOM8WfqpbhL3zaeHJcMtAorywYiL//y0TlHfF5v3Lq1M
HoRkKaNzJHJSxynSywOoa+rsVaNsX3y4I94Ct1BKotjKF9pvFdfqzNQBfpR+upzQ
/Fa/gxz6arW6+W5qFdyAL+r8YQ/xc/0BQlh2ttRzD9WxUBx/4vW/tjUbHzSKImOg
jOsKgyAZO8y9h3u94pmNXy+xJzTj51O75QpPKQ2fhXJrO+1HEq3nMrcTzr3nWm2V
+VU5iS4XeeGGjhdzCNW4bO+OplQ03SQiF8EhIYHmQn1VwflYvtM1+63pwjO/73oa
0x6fBCeIM3jYzWbN63L/M2d5QCrzdT5OpImmNaxj7YtArvu7b6cJKVHPjva3Hu+A
9NmRcS+2T8eHwe/g2kmQjmyi95jq2SzPj/QbLdvOHz6Y3veLqJQJASa/Wl3Z1yp0
qzmjJPAM7UsBGtErI0c7MwCFVp8BIZA2YBUKGguvWepStK4vMhtp1pH+IrgyBSH/
Ji8R3cvKS8+iK92+/sVGjjd8/i1QoUKeDFDtjgPE3liWMBnxVK7ZZUnbiiD3Zb9K
Sm/g3kU+JGgyfjFniKsHIwPoRr6j0j2IPQ1HE/gTGQt9NoOhEZyAgF5GWguETXXB
wCjH7NM0dkgp7lgbXdqBuYUjax9j/G7LmXrZu/U2cyUe0hoDviqtf5kZYVG58ZGU
dxVhzKgtn1lPpiEdce1Kvav3/IoPWKRGEuqCEFDI1dgaHSv9RGxOZu8AGugVcFOv
xphtnSLycP6QfFtURKAN054B+FbxweiI2HOh0uNXYviC2m18Mu+btT9XMikKpUrC
HpLo5DxTxD6mIAR+vhZUBNzEKcdp3lnXvWVdz3tQ2U92ddY5ZcQpMjrc9JGm1NSf
ejq3IBNRbkp8f7FgqxxC/wrX3xsc8rOwTeXJaRAt71WZuNWdI6BBFyXQBZpMKPhk
Y1ZN/+Ueg5mQ65wlSl6vcaEPPqAh8n5NeA3zAZ0P4f4JDIWszloRT7uLg7nj5Q+S
GsmTe0J4nXJpvIjolvIEZiyT7TQt4IP1CFzE8UkbIGaCreOZmhEMM7FTlPzlAiRV
3PFxAxTqEYQ6OLZizsizKYgBHqpVA1tZb6K/5G1eFOg+JhS5XI+XKSonamO2WfVd
rnzu/oaLNUDpDccphpwWJnYkKNpcPULezx5rJXjjcpWoaMi4T7u3mwGUYJHQE7qN
rmSWwzOBNukHPhWeAAVrEtdpzkDP75m6n9j0Cbp/43KCIKGhR/hIUgQ5T5gvpZRI
aw4IWWAkL7RJdjw1bqOySMjIfevnaTmAXmtrVqcYN5Ii0RBW0ri0QxTP3bJim5sk
Eto9L47NQKcdhlWjkG2J0Vd5vXucr2aBsyVrymjeDL7L1x2yGUAAUcCgqWuloaMB
sv5gMK60P5yqcbG+nLThBcEgabwvlHLVFQfjIvCAGgPnE0iI0b6HwryH/uukl8oK
FlbZxG6qrwUaFV0JtDZ41FXLbFf4x5PnBbzUAL4f0JeMAOdzhSsgvCusbTHy2FTS
GqHpxODdU+KF4agn78t80SJNQUR1no6cvmgg+UDf943QhBOib/+pzsMI33SZyXFS
QQ7g0BlKn6wT4eQj9WD3p+PEksvALVj2cFtW1nwh77eukvswl3se6woS8Gqm3/Q1
6rabsQLNfn3AfUM9HbDDAMayTpqh7m2c0bUcjUfI43L9pVKf3THeTNoEvKicXmVG
Wk8ecW0bJmBt2KahdYnVHc3LOmGEhn4LrcxQRCuvZvUz2A/a/ClOz+sGkzGokncM
xJ6qZuMwigG2gbg7OTpngEevK000N/V4dwr7zK/z0kVEsoju+itzxxignSrZsiNF
6P5goqUGlqhVw8f9Sey3+MOMccqsB4RkGNX2rLsbqhujuz4+wSHnQL9W559RR0NL
N1iBX/szAdMpTrNc/Sm8R9Oc8YROAtzw8FjXncfIBWxbtl6tDL3hvUUKa5f3reOw
fTJNz19ooZ1qU/WAvYsw/RABoduH0TpwqBTcCNiZOwldGMCo9UvOs+a9GQsjWFo1
rxKE2RKGEomqZmz5erbfjXKAmIs1oY7Iy1x7SO5VG8IALWYqiXCXM9/o6HGG6YVg
rEnAaPxPOI269WDarAfVJDwRhpTIvIBiQAaKSJkRLSUdC2qBXhcXC5HZJkqH6/81
xfQ1X7/IkF8lw8kL/X066+qTmpzkLDoorOhVDbLIWIJoIKDUw3b66GOcOwMKmNzO
MVG5ovnw76c8/f7iAAjcJkxI9EcOYzNjCQX8qHlZRyJ8SwMy3pB9i9IS4ClARGvN
PMb0/WgeqnAilfps4GdbRGzYzpy39rto+ZBFfuc6rMoaP63UXK75kBaLVX2aWYso
haUqnUPF38sYgDLKk0zOP4/WezBKBCGx7aITpmOHAuxjPQfG+UavIoX0mfTr09ak
Ormy3o8hxPXQTl0qsHgMt9dsm02BinWclnmjxhgraPsx1eP9K/c6H2ebFRK/16np
bm20a8lYRgK14P7WoFdJEIqbt5Q2Z67DG9nRJ9BlAUk1v1cahxYCPM80TM6rGZZd
Hllv5XqI9DnyRynJfd+OreLPFMlwf7YukdID0MBPKQDu3hqaTwyjY6LfYxueHeXR
UPq8NdmgiI6m8sF8gPYdfYwDuNXtK2euG1w2TfMynKlpFImKNPAgGd6mF/Sks8i7
W2Po0V/vFnJEW2zJybb7vXf+1kCcLTxgw5PeAVZponlRxHe3MIEBQ3obZrLfWbrh
exqKHR1zZMFTQh2MTmWjgyQ9hFaiNzLGl4ZSu/FtSvPXSLR3Y0qR2K2GMgnAfNLl
wC4ItvlMOkvpHYB3+x7yN+xEAjkfbm5z5OVjTyZtPZ3CRxLnET46bYnlFysUVtLJ
PR3NR+dZiF/nzyYBbgLKomNwroSBA5f384Uw8WVNS089r9NE9iecY/Xegvuo3a0h
TPyU0wOWEIjFVkaGvhOxAQWf3YsCRoetUgQFxYiGJHmzBB2QymEpe9qm3KIOvukF
1pfR9JYl+ozZyBWHaicD5R0iR/eotTUYH1+phWvV0Kd4/JmVueGnWys2HKuBtyqa
SzY7Rj/Dr5mWO6ugIuLfCnxPz6swbJDi+EhllVK8nDSTClvhz8PCaC/8A46RY6iN
nb5KW9CZmmHr0KtBSi86iqEppKNdrizIgrlJsM9CfUXhItxDBmHQuduMRahs/9lA
pcfUWCD+HLVWTiqGYn1NAZV5+5GuI5sD76C5/SZRYvxxrnId5wWlh43ANEfU5okz
G28CETusDxOLdnAleDGo8omiEtxNUDbN3DwHfX5jzm/izcyE/Hcaf4MDVsjuQRr/
kwmeI4mrYC/YTXpg/KbGS/PFiBCLGN0ZycPJjkuwbYeEpdeUuJuDV1IjmJcowEwB
HNjsSAEnvtIEt3XuqLlzCoFmwN4mSCafLUsI4P5gqKDcRtk8RPE5yzw2rwQmp6A6
CAAW3BT0avSW/9JpiGHVO9w2j8dbM53v48W0Vge7wdqAGBsDXeMxq/p/8FIrzwvc
AsVZraw6rUZtkYp/jnYG5qyfWLbtvvuvT+7liniIw2su31ilc3HNXxTuqFwTCTfV
rY8e4MoZ/RKsQnUMH9C3skaQqJim8rXhX9SIIyWlZGvangV1lwPQTOKiUvMUd+fC
bv67/xsF94uXguhfVUJdbb8DI3kybe2+mtfnbAPMuNd75mpL7tcEfuhhxpP6XaPj
HhJ7LvOuE4afbC1IJXCN9rh56pa+68OwsqSP+s7VQoIYUioMadldcz60fpTcor/i
c6kpYmIqX7xZKJlZvVIqgCciHMo9xmUB+PqWBxkekmz4ud/Z5lvh3mvdjnOf80i9
Q8lma9CdPn1j6Rl/ujflTolVmgETNcvkVMCz20i/kmzA+Trc/uciwzKDJdwBxNMH
JPeoQaOOakZ2N4hvcFr7T0RwoWsBuU8kP7X24+K7cU6kAelC9+h5blIkTsTSLwkH
DsPtEPZ868YDr1q5kNq8AQqtZNmcSEHjjrnIFeSkGyYrWJUgjqo7b/uY59Zfkp9v
7rf0gQV/kvbBOOD8wT7iuxjeICwSoHCbCZgqyfSuy65iqXZGt4cg/qp3MZb6rMvA
0bTDug9rN+k53cAplssijHCfbxrraqlUhEjStfZ1DZUABgost4s6QeVw0QMlmr4Z
Ppm4HfeLVx3OqQFJtAW1rcfXnw13Yi3hs4kas//d2e2tCk6NAn1QYMrt/ql9PJcB
phHGryfMEMoT9kd5tJ4HgN+omBCKZgfYg5RKXDNoV0yfLvj/GdxI5XhrqRLxiOzM
l9EFjD3ybhEyB6UkVlRS7bM+g4f0jZc6FdMkBZFZncGadLsbkd030Ddo72Mh6cnV
X9GWGf/HsP3zMId9WEFMbpFC1aKU3thjxlrWK1YjcwZ4GaVKdWWWznF6T0AnCHLv
WmvAbjguTpnHBW8sEKxufR94FWTJh+09fUgLA+HQ5bjEcg3IRCzJ9DLV3BOjkVF2
0yrNNrXkHAF5kMWeEjHlm9ifIisvPpGR0D0XduzkqnafWcdG+IyOx3GS1XoH9Azg
o8KS2S+AT+SqtJ9MLbCseoCC8WvPzIJPUjxCs3EkKV1cO2FjUWUq5QeXT0gGRQCf
y5Bq4O3UeLVr6PCqgmSWl76NoYJif7U2mWKvx2/9UglSHsDd9zeDWkYDVcrM301m
8jO+5a3XjqWDnpOWupHkSM4I8T8pHZNaetHi8D+nY7100vZs6J+ethOJMOqUfufg
mq1pQxj7AFLnapS83mS0mD8ARLGDHuOGL4UVHErkQ78341WLzsYfoZbRR1EOpWvR
jj/vNYt8SNYB1j/j81BVOwXRTZe/iFX4l/uaIj0Q9r+HZ7W69NMMW17odiMZZbei
Oao4pHbIjuFJ6+TAxY0qvMJjA3JlHQ6YTs3b0I3VkFixJfLmDb+Ds4Yj0C/g3Wor
uEhmV1fHl4aMIfobCmSa1eHJAyU2Q0oqAP69O2gLj4OXUxTKSTgWM56dWzMpU+aJ
0vJrhzNPw9iUDFnRuUJIUJqbGbtKjH0o3xiVCrKIcrSAz5hRY5pfZ4Z2MeQ/wlr7
+neliNLVXQJ7XQu0n/9txdwGEf9oY5f0CEZqsPTUi4BB1Rp+sjhzUB+2XLHdxq3i
yWyGPxkTLLCaPujskzp5Z2o9V/kuwKsGR9yHXyNUeMVFZKqbG1URAkYrfW76swzT
s+gNu5/dD46IE5BCgwZdye/TL8fkTaWAgPZ245vOpwcu2ipWfLRvGk4bODMq/qBN
j8195FtPV1DMOCVRV1VJYkNYpo59SX+4qTHhM1m9iGX1w2I/xuW7NmBURZHfWqme
Wptg/MMNuO8ngydfybLL24r471+NNPFukK55/LBhe2N7NGu+/pz7iW2xafHb6vzU
Jdwy7WTvc2B/udfaAI/oUqhfiVoUlJk+Ztx31LnVUmSOvj3bYUB/O8kYgPliWs9M
aPl0Hvvjs7knLQxYaHNDiFKSxSRHmJpAmsV876X/hrTUU/FxbZyJILSWTwH576vY
RCLC7W4upHmCWo+fhIPzCSxkCYL3AvwThmab8wABYEvvNv7nD5Ddjwj4n72wicCG
UHoXu7IR8dkmBc11ghR1gzZDIDs9vq+FpVN7vnUEVevtbSgjqBJokyDIBu8yg+HA
H2zTOfU8Lkjf2CJFR1+pkvkAd3zRAtu3T/sQgCq5ws9fLfTeXXXDIp35YmNtsPX7
vD7AmiIC3IMRCN0HdcwjUK/s2xoKzK5k+IwLjGZpEkmtvVSexyf/r5px1CVKznRf
x3UWz0lPeNGytBcy0a51QBqLgv7t0ZH0aDF1MFiq2if0SgFQeEuHZQ1mSlUMAFxi
FDAf5v3VN592YXBslZHZ8/cr/tA+13N6/+xF5jXStjDCj56r7DxBblWCsTsnJ7a9
vFvImcZwjzU/qXA4dvmKlUaLOsidCbE+O3iWb8K9z7CM4hu482KmMNs2hu0c6id7
8FmRCctRnXbEURdwZ+n29L80eSxfpxZ92AthP3VE6bZCPFuVpHCupz1nU0IgTKMV
BLbpiDQeRdj0C4Kk/4LBvvJ9elpMj7CDkPGV2b22l22w3hAC1LKGcU8nsjJRYgwc
1eRIJQXHQ9oBhJfRTUDyvuKCX3aeR1qBVlTcdFRMJXDpm0lQM1x2wiTp0B7hPZ1E
ULcg0RT828fUhD4w68Z8W0ft8h+B2B8DxjZtixH5iuQSKI1z/tSSPmQgbdbdBerr
8qEnI50FjOg87fuU+Vq9RxLJqF7FoTZcqeGpNM38jVaYKCKw1M7j8I+gSpFq5rXL
T3vY5wjWAxYJFZfL9Njzed4pZ1rfiybBCP8Qq5YlMPR0tH1BjAwvpjunIlZxugvE
3mbFeDXsU7AkhAHYTydt6PboajBZ9uJog+0brHuwvud9wYzt2BStlZ8pyZPcBKHQ
ruxPHy9rwJinFqnimrX4Z/ox0DDKSYdEkf2Qxx1gTzPV7HR779m2ofl5060f9KCd
qP1oUdH5KRuLhrAeZwa2L/Gd+/1Hqv7p2n3kWqhW5jC37bFX1+POop02/yBgmI4x
I34Xxk65ER3wfSgVvsD1xseW8FrDuA7vYhvQWgP82CDT252wBrUCPtXU3I6P7iRt
z4ethfhJFvFD4GYWUdqywxvlnf+fAsBC8TKZbO8QfwfV2mLRCIKwNTsTSbkG9ugd
WsnBxBQVWZOv/8E8Z4aQwmQ9wGsrHil6xGEsOwJH/26TGiQd+pOlv+6MvUry+/J5
tQ6A9xEGZtwXaw+J11BGRbB14QV/4Oc7QhWUfKezlZcrPdxlsIFe4RDNwuufKJqx
DMx58o+VNq4gQUGZxKJR89bE/tTjKUC0MSeK1Hj5tUoRtHoPTnm9Jl2yTVQryXH5
W8ol+22iWG9fJkvrkL44nwwtBXgaTJgVoQThJc4mmkpVryCtxodRBrqvLOe4LzDi
jCi4r5+W3axUE5Mqc96KYB2J+htYrAsaCqCDkf/2ISrN9luGCU1i6txe0xLs46sp
2U0rJX0+LYrz1dKQW3G5gFCdSPpQF8wnjZVFFV7NJYF3DATTUQmZUUF51oovFEh5
/mESt/rGkcYusPuQi8U9kwsuY6rFWIiyIn2e3qG57mmKHFLODUQoHdIKCUjtO8eO
xDbV20Tfu8EGE66TZoX4PCfP3EWv8jopbi2OVvQk3aexPklVFqrvFplE2gGPSFuh
8gP0sLukTEnRxj6Mkj8QZ5gQC8Eh29L3CW2CnmaY9nPVfqCiMMaSv96UvBvTfpwX
dx04Xs9rTWryarOuiYx/HP3s0jMjH1zK73hJSLqBfUg6XPV1KG3H9JHFMJDK5W42
iUQ3itrZ07rmnNgFeUgl+1gJ0/4QuHYNBUYo6Ic353Eb0BUqjQ1BHFl1vMEFVEes
Tx3poVcGBedLHKhD+PvBAoDAuP++GVtUj4+5+KQNr2pktFUxnT54LND/lguolgyQ
qzNqCvFP4P8lNDpEkrqrD/VGPhskkgZB4o1AspUoBPLZYfu/aYuWqLxwjp29qcvg
nzJUfj8vBG+/k5+bM+x7VFlsiPug7o7gIVB/dN0rz1EOthixMCaZmeJBwsZv7i/Z
1zErmDEYx75KvOzBl9S3Gr6KAd2vSDGP+4teZyr48f+fsd8+YNHiaUvUB6IeOX3q
1HqbQYgwK0hfeuzMNnqUjss446u90jfoH3ERsSnu1ggcfK8bnlpGgS51iHChvpvG
0N8gJ1yvKk6mJEWJD79wFVOLzYPxH8AIv2CszeNdg5CFWBRBCAqMrP45oHJy6GYy
VT4tZVVvzSv+9Sy/X6tNnOJI5jm5nFH6tpTpOchUujCr0DY8vjQDEsKf5mq1vuD2
alJW5Dg4GQWyQh9QOKcWX6oWJEMVwwKXe8VOsDImsPQ5uix7z+TtjpUK9uYuc9nN
SzMlGEXX0yZu9dnJi333+l5D4xWGqVmz3/znWYq1VnmlpTLoZJgL32UAyUEcjfkb
WNARIkIBiH4huECVc++wS7sfvw/cTBUxWXYww5dRV8xh/PLvoCeShJmYshlYKaao
VWL9wx6sLs9G5SLtVfj5So7grBz0VLoN8HpQTBY7noq64kNpQ77uCXeDssA2uE6K
tH0heCfKow0Ui4RefSG65qWbrPSGHSItLK5TM3MpQtz2vF9mddazmvete3Qlbed+
yFGqp5aAXlLCOhBK3AUzCfBFwUmjI2BBrcfDF0A8+QdILR7+pCgprdn8rG7QinbT
OqmHvOqiZXTBj1+nQFEp8zJMVmW40lFtyfgmGE3aUtCMEkjKqEK+Co8VHMgOKzfP
BYLQ4GGh1mOwmhNFQP4jQfDpqzI0TdT534qE18DON+CwhItBDf0wHR1UDpbTKwEs
oWWiu2lDbF4LZIkl6Hcvvo+QBTM8554LnEQtiGfYgsMmztBsjCmKmlmLsV6qfjPI
UoyhZffEIyAKIgcSv1n17d6vbMS/Xfs2lK5A7Y1HpoV01OYlXgI42g3z6W+86xBI
v8PQG7kWJcGsfjIyZxnC9CDrA6HvJ9w64VKyBktQc4Q+PSbDo65YpwcI7vQ0r4hg
xrUn9qOhNLh5WR8Ns57x6ZE/l9eyMMySTwv4UORngCk6nqpyc4RZevfFuCvQBIF2
CUB4U18qhXBLC/wGsWFCW3qJfEUQvVmVOtZeiO74o+Vd+cvcpd1uluPJcW++0sZq
KHKNxiJqUQB67E0Y2Du2VvKrkfTQC+yVIRQE4PpxawQVtjEQ8JW1j5yS8HBFys+z
WymeIWNfripX1iUXJ/Ho5ujo54G6tsLu9+flk8J5Hbte9I/fyvhw8ZD84dpOFmgQ
Hwr8UbqLWIP2PqiIVe8oGnNw7Ma3hWPgy9abbh5tG7T5pO9evpJJRaqZKTBBWyEh
NYgZz4CWygAaL3g3fdE38+SnilWGkwPiKGPi3I+/DMGnYv+j+L4xEgOv8sW9XwC+
s2kwqwIMcaBnOfhDz9nbd4UFVui0IxsmjocSGq3a7387QY/GfMUrZ3cnc27M5155
D0ourr/3s5kyzlvd+fsgl83DZOUaneefWn2qmBxICK2B/f+5C34CieyBFIWE8Lf5
Z9GVzSIio64dA67UAY5pwKivj8yb56zLFa4bqitbvLt43udV0ZqC86seK7Ybt5RC
LYdIFZHv9KD5nWmgY13CvGOd2xc12JxMC7Wzimmyotds+nBbZFo0hGfNy2UuvRel
tjYS4M4NdPA1FvpuuM6xgJdFG7CbJbKQZTgD9VZRHu5w71TzbJw3pyC7J2ZDqhGO
9a9AWERkCLF2ERvbb2qMCwe4fW5cOqI+tq1CmZHXAm6nXhqgFYTp1ZAn+Y+qVPvV
8Lyf4euSwHPRpX7guVFkREgC7NCg/zRdGQiIb7Qz1pzgeAKDFGUyFgVIAtKYoRJO
o+rzsbd4KU/qCvQ969vC7r9XJP/zNceuTf/pJJoHa6aR/zDwj3SWjRiRVsl58mud
17cVCQ77xj8ZdbwU4O9XgHz1hGc/xt85XRO/37PK6Kz/npxrsRCGxrzENgozxIbr
+tUanPhO3ASkF2V3AHYF61ZhBdPOCBT73AdAYKsWKjr5amHjyb2Hl+c704Gtothu
jdNNvgnTjWhOCnCpzLV132UfdaUbki0egE0ZuLaxcYKR4RapprQ8wsCvkB7SLg2j
CT9LnJrmF+euWb6EOXzyzUxgoKn1VmmD4ky+8jut2qNJ/AKj332DsOatxDFMR9U6
rX15+PpH67IF7arM6X7Yr/BgdzTBdE72xqxqtIwJ+BD86sx8t9fVchR04YOHlMaV
+vuccf4iQaRjr1ujUvEogxLMXIuuOilOwIH7X/6eAFeB3Ts93knm8DwN/AUmvEtJ
PwllWDIvSiM5xUGHCcumvRU5c1LncXk4VgmPWqrpAmNCclamFjHS+YyuPeDbFsjk
pGrEPI4g1k2Ffuc1hH69n2JA6E5nf7nS0pPfwFZw9qYvAMn/SBxAhRejW4yukS0Z
I9rMU2DpWIlEORqTaFj4WjbfLYHSfsDLG78Ru50vFTD2zyLATL5ewPom4TFfs1El
n+JzdynNW6K/b2WLY2maEZwPtrUxxNH3WTgowvtsUj4CQ+F3AHu0EHOKvgPYrdVp
tsHrpp+Zf7uhOeMG5SPvNHS71f6gpDpXWwwdUmGEfViV2eWc0axmKgmZkchjc5xM
mcU0vyqA9K2HK9b52d/CZQb5ZZQBfZWhuQviMKJ5eRWRRquckaNGNUP5TjeOWX8Q
GqLAmdC1c1KJ+IeqK+/tVpiOSRtiI+SgFJdVrekSBfTCZb7fZnZGc7IWcLucZjKB
i6+Z0VtSwSqBH3jtnu8jHDRi6OHt8swypv3r2eznJWEwaKI6h9EoT5IlMPjxCnFO
ruYurUyA/J+Rv5mt7CYBgj6PWZbDmEheBWgwINQQiwKESuu0ZIeWAuVBqENDF/b6
lmoPtawJIOpu+CN2ObEd4PvUVAMzD8aCeKOLup3EMawDvpQtnEmB+xoJnG8D/mRB
BAhozVmsmBjI1k+a8XHf63Dga6jLy4cUIo1Mr1jIeLU2Jct31+bfhotY26sVPQqP
K3MXf+WISGC6DJJYP58h++4LLqKvMb2+lYudf83pNOaXmY5Bzda02hNIF5h8vrG2
MR5T9v4v2QJkUI6g1v3/l97YxocYFn/4xpvYVKRoUbniRjS8zMEsJrFAzCFh6uXx
7/xs6o2yQgA5lkq6FWTrcVBcLXQ9urnUy2h0HYarZMobPQjVr9wXEzMlqxzq0XMf
BmnkKITesZ9xzM1ppRLhcyivfNnk34wS7dVGuuVUzxLM+DLAL6vmEoIiybQE5qE4
JY2kbKyBAXZkuvI1grgObJJDxggT9jJH5Fl892Loh/opQCENXZXMjK+b08TvjKyZ
h98R3P1VJqWjHxovV8gkZAt9gNarjgjL34wtPodm4qMaDulqusfTY00oiAM3gxo8
Jn9DXPjT7k1pJOm5+DP/x18hhDIsjSIMso9H1jXA/EeLhfncvG9FW9NBUdO/4pge
lHWTEZ4KEGOwuGa/kMSvURy5bpHEcdT3GcisSU6HGthIaQoBQDiRvljMov3NrCcl
P8RHsKAzmNvZf5l/PvzMThQQhNoUkdRomGNR+qFfyJr81njrlzpQwBjRGDyZGZRi
+xloWKVYpgLQsPFSU1drB60ufNgNeYvPYUgG5qH9AEfRCX6dCIc2BOpOcjEs/uMP
DupAw27nehb3Lp+/6+kcaIRuYhiEcezb+tYVQlIA4gGFSWb44YH8Rl0C565srRym
9vtFjXDWqkLcDKwfCcRrs0p2ww4Z6WGrXnzLPEBURdBD5UxLjnucyNPbdmktrI4A
NOBFrMVulFbPNWZHm3+Zmdxjmom8ZdmVojulOAHoLjmzDQ24xESrSopv1dJHIylb
JQvHUYQUl4ZXjbdkBOO8juMFmsC4in/yFIzHMwc5oFkmLTngTWG9iVD/LOfBzUit
CdFIiF0Y7UJNkEW2o27G7s1f64c3UEZDUj1wgl+OiS9uEqH6kzbAqILmOHy62ynJ
nS0uu4DULhvbwsK5zXeTXtcvJ4he4YKDjC1EO5RMiMEy682QgVrXXR1X2rMJ+VKX
sL3X6S66pqtLnDmJ7f3gSBPNenN1Cr+X+CpryJx4Of/PHgSyeUKXKpAp1hfCSjWc
z5+0ytTUZ8XXlCG03xyHCqhB/EKqjGopyej1IPQFU+SfPWCryisI/6ea9WAwFOVQ
o+hMdEqFZ5r3cnRE3X9at8QuqGBrjcmX7R8nLD5giDkenOMQ+6gff0MY43e3K/nv
5bKl7N56ctHua+flgeetLjnJHkw6fQarRB64tIfR1Ytju8J0ejTY/NO3xMj2fZDq
gZ2SMAD3VKGMLQ7ewoLcXpfpqf6swt+/s9HwXe6H64dtAtzNIivktj4u0LAU1fcG
cSqBzWC8YJr543vKPq1PwUmE/waKbTS1X/deuFzAlyYvAhBf8VkXkqTLP3b/iTZP
267nKnSuorggjJ8ZxFEqcokXEEHo5e4fQVYsHdVS5wtk//hlZCfaszg41m84c2Du
kQxSF5dGUUBg/5+63k/OLZYTWp0oXXLjmu/a1ARjA32YqIUY1hAMTbLz5fd1xJMf
Kmq190Eljzc+s0T7nzn7qB0NF4ZdUzjOjHPFIK28E77kM5m7WaddS/b4Osnr0vBj
839yHDz5BMuo6Z1NEwpssIcpO0tjPXxGEmxNSKxF9KC0EzsvBadH/39kgJIVp/wG
/dPEKkcNWaNyrXmzscfcy0mWgo7dN3b6iFnY0LLTQtGPglX7mJaEani5sucS1Iu4
OMhJNhZ9qRjkht3uHWqkfc1j0/b9VWJWJaUoZwBTsM7NMAHOsse7Plgh9RJu9oKd
ECDcuhq8VT/CLEaQ4H/cRB3J0An+5sZDCfGSwpLrIMiNyqAY5qkTOnDj2eAW0M7z
+kv/F/OveQq2f33r+E7QNyUVhh6Rx+lzHwZy6HC4i4Wue3RGz+TxEhjZgjhMy48j
dIyINK8abcCYii5Xv+Bi1RdeczNSg6QUU8OKADlF8psX+82P0YN5MaJnhVC0pi/I
+BhJBmt30CTJBSNxBEjHADHIQZ+Ka4yLo8Qoz+cvEw6UWwFeF9vcDcDM/bJL+FHB
7zjRvwxP1kdFsAAbCaQqEihi6K/8G44OclY0tKLfLa6LLX71Djjc5nKwGOYClkL5
95U0BzZRAcZA9anwTwBBb/QBxx4mWS9oOSFV64W2N1bHYt6zzaqpbJKmufz/dbnB
RnWpPZaXVR/HDyWGtpNYhUlhPlxFJi9FrzjBGhATSrF/zit9qa6JLgnUHEg9U4Ip
olT89aEYcgljtJrqi9b/f3XLyvn9ZkJRZPhlJzGcmcCPBvzahyk7ZZ9owdvc+oP5
7vWSKkbA0l8rSNv2Cf+1GdI4cd9XTJtFKGGBUpoKXpDyfA3fhu9wEZCfgK+qIUy2
95aLHdactsGDEnt8mJdK0LiFtNJVWpxMa5JybS9WMCrzmWm/h4NpbAAA3vojzNiR
l3gb0YcUM9a7wsfrqSZo4zAmhbI+QsK9tfKWRokgTYenvjSXlvpwawwW8G+e2JH1
GW63IVRBlsMlv+bczrkXBBO0+RdaBcQcJ7XQBWNO0dPdEvL3AC5qCVHX7qX8oFN7
y/2FRO3do6jNDWrv1F+AyO8QyTlum7YvEuJ/ygMIKHIYqt8it2YltvOKvN2IEfOs
ryavDhGlcgaBb8U0Q+ci7VHhRrEDRI1PQPzIksfTXGzd04P34HB9I2hkQS9CEE3w
n5ydprZvwGdaZyB+wK6q6gngiBci9aRKtPK1JN4mwEaL39WAlSNJO8aK1anOwutm
AlNsuoYyfsZXXTckn/gyF+DtLvdUiyBP+985iWrAsmcWlvel2LIvmrl0gynoc+wp
k/3aHm9yDGLhDkTnIbIGFYGoMFvzXomVBPiEhdvgpbbftv2QZK0mBMLbD793Iq/1
Yv56WTZd+13p+oJhgQrgefz3dZe1PvlqeRWQVmPiTZSo6sglGNiwdND64YrCY44G
zeXigXI2sVT0aSug7bJiZvvRB12Z2Zo5Emyz/yxrhcbMWbW7jNYWQ89H403dgECO
9RwcKCO2UwOSCN/tmr4D6QugbL0UbTADlK5D8oeHqNKbPE9isQSal7Kflee4sNLE
8e0wegi0Fcaq4/VTy1VNTNuLt6NoiPaBuW74gW8fNPnrDiSMl38x7+sJW3jDpcoN
WewO90g7TpRIdWNieTvXDeXVKnFvDs9A4Zuucd4DV0WNSItuS2HpU9xRPgO8uizw
jPC92L1YVlNX34hxUaELhHZmT96znTzlXd1ly0nubeTXgXvgeZKxNSxFC6b4B9k0
osCSODLcUXD33RlVVc10Hu3tueZ92jl9TncWpNI1Igq0q70ODTj88S0weAUqrA7t
ECAbGnMsXjC/yhUdIx2OUx3X1USMCD0aNExgSRf86iZrls7Xwcu3Ec2AKhUxA3N1
NWLLuQZM+cc3GFURbyYKyqtdftF9tFF2A27ei1JFs3g+4P7Z4CZrFiRdyi8f2lTU
Kajr/EaDr97MZyD0FY9z9qokACxH3RJeMFk0j+zwE6B4YW4L1R8EUHc2zok2rnrm
jOfj8/RyL4jj0ny9ZkC2W3btOmyQc3zBczgY6gf0JAsWOeypFdR9mQLegEBGqyP/
KWNFsaRvFLofmK8lYr1RqVZtBUn1cItVkQZ21JKUdtIQPkHHfPd4vKimrHEGmS62
pxT8PRAKluT+juVEzxU3w02OpE90ushtgl6fUch1z27ZVIvNsI7860RfpYP77mjz
Gw0R18vHKmKb+pHioxqELNkep/Tq1S4L4ZBELiEEdxpzbYkofIecxSD8UU1FWtkO
JH9N2pT5eggZyq9/fJ2izyOFthU19NwiiKD9f0y2ljEBFDi3xLTuO3knFa4GgrcN
UKJ2qc0WMFWD9DHowb6TfcR6vSp+IbpnrBb9wzeyJEaYk6C/Ke3PyUCFgzZ5s6z1
Ic8MqavVsLaXptiFbAufR45decTVgYDBcoSD6G8vNAOXZAnR4DoJ++9rsE/sRUkB
FLBg/EZK/zzAAVGBP0ari+rneyOeuiXZ8B1FhrhZ5tcogNOQmzG9VO2pDlWlvS7g
2XEYFAQ+n3oYlGnJF8MD2paBslqwQh7mY29XMPjcPVxqG1fJAckAZ6nRS0hkOotc
75Nw8asNBI4Qf/6QX+1PbyVWzjHojo1Jc5Mrtl4WAleUV2PgkTc92gOyrZbu1BLp
UYV1rPI5aU+ix8rXWRCrWA6UyK4xwatCtS/IHYqO32NXE5MW9I/LKfMRntwP82Ym
j9rQnl/k9T5WkFXsS8LOweHlp0v2MC7hPHBhaQhvn5Gx9v5yANqHGNxRD4ITm8HO
0LwtruXt+/YSUzrU5nQ+PEsswiGFPLGhg5b/tXM/kdXaBw7pbhkJc+mCGaQ+4uEl
+wlC2IB0MLdxLyjcEMig5X7Sen04fEAymDa6H+TxvXASR5v0XO7T68Kq0mhrXNAj
fh3fS1MWDgCLYvLmIJyPMGT2QkEynGJOEHxMgB3GLV+entAIuSRL0hBmgdyy6i7X
D89+gVgOOuAUALQjiwW/Z3iru1hmGA87ErNjvZiV3zuz8fhrwa1olSJjdMBBTfVN
JUEx/Z0uYZuSFJ82UcC7wq2VFnXqfFE1l5mA5yBlbRX8JrqbidX9qxdGd4Z3zPg4
jvML8oLLxNOp7l71FjQF+iQVEGgwckSesVtAycgF5g7tWSJ7j/+LrUqmrZfsU5I1
ZTHwB2WjsLca82cmmnYmOBlSJTR1crGiluy0tYE5vdTnHWi0PElENfGNhdjZ7ZQJ
PC6nQNulKO38I+OlXZy0RLSMsfzfkjND98RHJEzOyW6/qxXlvUJzYW3TIdnie2/l
Kbc2gXovv8ecUaH9i53l0Jh148TRcf2UTLCdKxsvLTOM4KFeTsbFw/uKtV8O3wz8
M3xYgnKJsnCjHEIgBVQ9Z3fTzrqE5/C9xTbiQ5zDTC9unZP4tW5WCdWZsg00ov2N
XSSucJw9+hMDV86Y342L3PFN8ujgaTQdlTqcQYU4XoOkP71EjSYI7NHQ6/ChJgbK
H0mDVstraJIQZh2GjOEIYzDsJwl89QXa1MT0wc0wdZw3kP3bIhJYTS+ekQB3c8L+
nmmSBG77EwUMS2ogl70zWOcmXtU2jd1Tc+2szBjnLZesCHoWeL/E/c3CFs4xQgdG
NShXHSbm/nI6M5epbMNjPa0nntS7sjCI9w2uj4D+YwZwpQbeSVRIbnqKwOVZxfK2
O2punZwoh4FSK08ImpgpPR/AI698hIMUQuVlHSVwvkHW/bgyPwf36lyAGqNgd2N+
yS+iSYnDY1i1ELbp4Gnmtv2KFwp4VUySbicrte1q8yNBtu+dntGE4sWCD23gv34s
ViUMWfj2b4u6/TZjk6C6ojmFbk++MXZoBvgP5nOHfFIff+mqx95qjJaMH726qa64
8M5Zd9xaokaFyZFAYJ6eFZ3otJo6zS+QVsaABEbVyNIs8JqujfD9crcMLG0Ih2L3
3RoGDcphJ07c7yX6/sfMDPThVV9BVYZMxmbHIF7Wez7X2LDUb9ByXBHdkcYzDtjx
uWFDYv993hpnXWL54gd7jTfIIvLooT7wSjLBbtWHy12u5DAGvG/bkPWAjbHiBrhC
cJsZWwSAii5bPy5K4nWUhAWSYfB3bPrBrE/1rNPFs2vfSRyt6/FIlxDuZk+81jNf
uCGtZ7gh9vBdghKvYpOqHEqDFDnCgKJrHFJibk43OQe0j4YOnRNnDVlCIkLiMsEd
s4k6OcUcjfbR6KJQrqFcWR04ng6t8UvCy671JdYUEU60LmxekNp8PV2NPTqX5PTx
REoAUHWwG2KdcJbdBc+mDmA34IZ0A3JpnTrCB8pcgV6+fGHSFuhYoknmDR3YKOT+
GCGn1WTwFHpg7Q1tixc4QNOd9WKmk4UOq0pYeFTfQmFVK6AKzGeC4LThVQS5u1ug
oZELbtY734fYIC/+nT0Spdjb2dLPolhtNv2Zo4bOEAZ/xSMuFyRPnWW9HQC/VNE3
DEysrjqu5P0DSBCO0qBClxJk4sWbz7B5jqYscvcbJIsBYWL2XQQ0IcPaEkCyjeJv
QP0XZkIcxZCBLpHSjd5Vv8ypa0OU+0k9ZLV8hXbT+FVdqsD2T82WIEYH1MAB72w3
+7O91MMxk0tEkONmzVhAL+4XyPulkcZdjw4TsL1DkSq6camjz9wg4eRvxBdcO1w5
TfG7VRk9pgm3209Sp+RpBikuGoMwkLpiwN8PGTZoexFmvFy6sPW4Te+zCeUalKAE
S5pIduzIjioRhNDdX+chgtleyLGDB4joce5PBQekZmr4d2Y7i/GPHO4xlbnJCYS4
7cznKzfqXzpJvF5M8U4Uor9gtWVlj7chvMrpoLEY2QrGjHjNFaylCVaEyFD1TObo
bPBgOn/yG3R6sCdVhodpg2OgQUzv1aYQYM7clTWRpHSGdN6YWc5x7RpnSw1XVEaC
fM5sOEZsyg7OQuqQC1DN/jd8XDYdkWAxMFAU+4JvuS0zCrPz8CzIqV1WarkUjEuu
zXfy3mUty2TwmTTayUHERHwwCWR0KwoD5+dOoYdnYqFI/n3KHQtYG6J6Q/+8bJPw
rsTMxqRDHpt97tf/KRjPdYmJL9ZNDgN2aodAR8oVr0Hpct/4gKjbVz+tuWacsIeR
kC4jJXYjSX1tpBbNWtypHnGxyZvfbWYN9PhO30gUteI6vfnmavtP0NCI+X8UQPs6
mQ2BcWmRdHN9ETcL2hqdueL8XfBKCCdP42HWmWs2aq77VPuqCIXX+ce4wjRFfZ7l
BhncZ0GVZx+vARIHxFdNUHYI8RkcCcBqvUyw/7JW8R7JpE5l0PvPtEXBqUTCuS/H
0/DDsNjbDnSTInapuXPrvp25GnkMjeQTfKS6kw648kav+I/4hqS+suG7gPp39080
ASgncQ0bH+OM2PwykpbMAyoXB5wTaoH3Im9YOn3r9Wtzpz0GjpHPFi0f1cskq+NS
ZQjG6T5byprwjsudOxpBHErBISVanLG7oTTL8iGgpDG8UgqcaqghZN6aa7vgzzpg
2xwnA1Tyi0cgWlSlH+X0A3OY4VHqijZLJWyW5lXk9MEnCP9C0jnsURstatFriY2y
OY7lL63g6PXd/HBFScDkW2nHsClmAo4oKKenCbWJdPSRRzcgyWNYM/kaKC+5jKKC
z3qvjesmZUU2YnEjs0JEjATLzf1AHijcOYKjoZV13GsNWDl/UpPf1FaVjxBqy9Q7
tABX8UPA3dzcCKQHKbqVAIA2WFGoF1WMUCllMdV4a39uueCLRZg6a5ZaoqyYBx9Y
mR8zVBATuviBL2/NL7205LeZALMN7W+NdNguamaoGFqxJylUaPnaEVWnhVK3vnCZ
snz+OfAaGiSC9609uYtNH63bppdZwR++eRorKV3muflXYHHjPjlzpRZFHu2qqZAt
w4TOEvPj5+u1ume5SWLvKrLH4v3W6Yw20FWigunGwJrU1WYZJvkPyEFNAdk7l0hd
tUoXduyUeu5URIm/uf5cHZ3U+T0JseqC9fntglD2wjSt3eUvI9BKu+yRAVeeq1dy
yf9h/BY5MW7foKWLOy3wETonKBsPL/Pr26lNgxUfd+TV9pmBDe4ssn8OnTQgdd5a
UyMsDPNofQ90fikv7zcXxqNUzHFMaB32UKE38/RTLzDfoPMhZ2QPefmZDUruwngH
hOtqUuUA+/JT3UhpXJEMyEEugtNCXDDxWuDhKlOcfe4bCX445RSJmBuw+biHnts0
YNU1ZnohfrVvhfylZwzTqXX7urymuLVUOYBDEcm6DXQm4S3T/SzVvi3yIEEVwmaf
LVHu80mLBwfAIANMEs8H3PUHzOqFwWCtwC2MssbFPDddrvaeHRU5Szvme+JaTKyQ
vEchZvZKOb7bjT3mgT0oKtfNX2nPi60XuyeFk1cRe88Tc6uunQqT314cM8GlWrhB
Mmk0o5V0wjgSsFSJ6G9S116XLouE46mHGfalb5VlnxLoJFqdtSDAPSycvZ/KSRYa
eD/z9v827vl8aj3T87XX1F7h26bXfeUvyOSK9nC7X+wobfv7C1CZ2dDWQDI/9Snk
AN9jAfBNl7cRi0flIJRimQ224bV7pvS+v+/JUMyxgMGUJThDoI59m0i685FCT8UA
fTkOtHEoS3wfADi5KFGCsNRZTsGk9jzCsPUn3P5RNOpuZ6wXAzro5+XkCI+6fBzi
60XZfkYiA3G8KliRK0OFth0DoM2lq1PbkHXeJt9pt8/4azlOhbEGGeoKVWCfA3dn
qdeTU8So+JXTQV+P1/asToxzqjKWrHEaeAcJCYyxOPt566DRY2kOtmR1gonk7DB1
z6HpFU0ArrUHxdJ+axvQ1DYR8wZWPpxLpgqpNuhQg4ZBiC39AWLYx9WWVAAM9VEr
KHzlM/PV7dv2q3yaGeutOLRgdDk//SKve9vAvDaF9Bnnvc8ajoLsak4UYh93wamy
vwspykGJ2ItdYBd+5sd9bORpTE09MpYKAOEnHd6FnTvief+Vi/93kKfYuoB+s1KN
yGSQetcEKpJt9AL1nKZBFzL4XWhMM7zIGL9ZV0OYLhPhNJdJ+EDoISZ8HWGLgki9
GzM62I8/XuJTnaE5rgAXQWI9rGLirqy7P7kJlypDmMBwIWrRf3lHciGOi1kk9jX1
bP3LH0CTaFlQNV/ijIbV43QG/+0Ucq+tnGAtKUVYub79CEY58UgTOYqqyL6Pd0Xj
N8ptfpgY9d+eu/0V5i56Alt6e/pQ0hTOkAVxmov75ALFbhQ2+T+w7n4g1gyAEotv
zcnP19QGbAQmDse4EaQgpCXZp8rhbYygBttvWDgdF0KZO0RkvDJ3OS8WdwYY2E4X
vFJ9bqsbg0NsXhQxJ0EtYvc9Yn4uTHl7UmHtCFTxmXxXaTcQCBm4e/ZWhmQK5lLY
lYg3m/3AVGKcNojFYQs1FWWm/4bvkkTWfVp9G7em8EwUQTMjepMOaVl+oV3kr2hD
HFar9EIFRysN/ZuxyOn+5HFyGzJuEKpOhs5ctRo6C/tAUFDfjwaG+vMjLg1rJ6Ko
0ENVU6yvtQON0ItwmdNDKmh1gyzorCqvHup0BLdAFAwsLQsGRpuOV3rzopvjaTvb
3F/9SXYKUUv3bXiirXutgLUChSjSATXmuAFp2XVMdGPuaTtuDOWxDHMyfV2jhTPQ
E5UXQlO6uxYzBalO6itTcqmRKjolWWpbWE0ZiJMllbPekEUm+SeYMDYmUQO0M9cJ
L7sk+ZjPXq8P85pFuYxnu4mn3YTO+rhhxoIwAEswPvVEinCCxL2Pj3V1JKDLJydh
RaSy78V/nY3ur7ZUE7vPtzyAedkOmUNHnNxkGUhabu9AJ6PTJ+zoiX6gDNfvH2S1
TbE6lQPRBQPvyH4DjU7O04PBTM578N1UDkleASyOeBVNmgUWOFzkzPXO2P/hdzDx
UzVcVVr35RYcwx4WBr5rwcqooeB+8XSgh1+T9V/vMWh5nqlTWvAlBvNDlC9IhZUu
gK63TilZpuQvrqZAwD7nPIrawngT3B9OLxh1tq6s/C8gSvHdzZ+EvG+HGLxw/6UB
Kjm5OYrd8Zq7EKdk9aWhf6IWV3jxpxovc39/igzdX/6M/EG5bEnowHY53xJDFmH9
CNUDvkluQDOarGZwE6r1BxNgcjDdjP7/T86XLGKiKDQNhjWpRweqewNfZateph20
maHyFrb1HzaaUx1VeJnR6vHoegjQZUFBiHxR8/u3k4wENZPLvLTm2arAFestTa8O
W5EfT0gYkNdbwYPpsRGP99WKVQqpLNQWgIo6Qj5OkH8UZCCO7cYxOIob6Cq2JJLn
gTxF3B3jWBWsVvSREsvFvSFK4bQE6aI5uW5+466V3liwW75Kxcwq1dsflwAoMnnk
MeTAMz8NMsWd7GBaqUp+H5rx//5CZ4LEu0yEwrcuF/ZRT7GWOUSygefNTPzW7J50
/tPZ2bCx3QnKlt9x4KpNPx8wVZ5l+8s6F6Q97OLWRh9CJrD+0+MgSwdO9CqfjiHD
mIjBu2s397oc4yjRo1VGLchlmdlKk7dGX34DITKFYN/bfxwWETIgSUBSbb4CBoEg
9Vx428oH/dFfCarQZWuyhyNT/FDddvkvUuRzSLLHmosW2wD43r1Y1fbijO4+66Zz
wDFeMiEF8FeY4OYCgc8vMHTBm25Ij8Y6n8ROeXnOEXNQN9pNfb612erEYUpZVDZF
C3ISmjFzv5o3v/W1eEmi8VBK4eFZX493NyqrvJ4Xf0q6NMDBGcsoazKEYYvM0GP6
wEYhsuHU2fiYkCZUv4WVQTSzNmmnCqwhYUX2owtQER/EC8s9bco0V1Q3Jq15L80k
SA7rXmNzd5cH4+T6bbFcc4/psphb8tf4iNagqtAOJie8DWrwvBkFPFlONdPdWTwU
1btpStAJX4J2Nlbpg+a4+kdJbHr5Kcb3fUjFD8vPWlEgjphan8BvlR4mHZjAj2M3
PA+jt6yi/BppH5NCjYU3gmk2xsjtFabjzJr/WkaUz7vvmioQwh2yJLykErg6je+S
w+GJlb2LvyO9n/0KIj8QqYhv6npCWKIv/QXX3sQHKOqfhQ+4n0f+of/t7zpTfUez
yWmmV5Vv/QOWKnJ52a2fwAwS76akTPLi8XWI6CTRAKRhOxnpv7gMUmvpsvUDpRzx
7+WW201CJ0bSN57rg4HrTmP3pwM6hs5TJjmRA0UNA6212yhO2MasQQqcvxGTpaIu
Z7As07HZtUxywUaOhaj43aH3BRI70/Gvbby48ajh1qsTC2RPCScVgUErYtImrlkP
fwCtk5TQqRMpOOna+jFlNS4NalsAf5Dgn6tY8fWtHki234NEQSmgALDJctKKr8AV
21f3KDPF9tzn0M5/yaEOBARlxNHAktWiqC3+Ct6lfefzhql7U3lAtjAEy4wcCRFT
F+NrwE4wg6Q9zYRodlsGXNHCIGULZT9YSNKTqkuhDVXVWB/7So7sQtiFNt074obW
TML8nIKL8zQxuW9DquRZ2jZJRvBdumdDeQzD8l3UUPjKpMWopBdPxJ/GJSjD7xhc
9Fd/patWpf5+6EAKaFfeQ2LW3tabu5U3LCiRKyMSgKR175sEL0WPurETnQbB++pC
bkRw5fvsg/Mkx38S3vrPmRQasDZnlPlaT0Ci9j+q+1kuCx4DEZqJo2we6WVMkv5V
ekHTOdSrlhfwgfs7i5D0wtLtfZzSR07OUILkD+ZjAtied36IIedLhLsmCRxrT7PP
wdciqliyqGF+vLVCEgMxQ5AIGxUKqaPbBdY7t8CnVaRlDsX8SvzvwCazfJp6WcII
73Qai3/nalK3NDoEXcec4+TvBy/5LZuqk8wWCWVMNkTRzwOIfie2O3P2Pjvw/cMG
YV/hQ+tjdFZjzW9lRPwTbRE/4Xwse3ELVEIHXaLNCI/a3o2dezvjMHZRjFNaIwv1
iIexP5BbkSyjjx9k12+ymK5ud5l+PmNUjH9ow/yeh5JIuyceI/hB3iu01kn+MsTo
cLkhzfzgJh6/FaaKmngIegJ4VQmyuDSlnB8YxBSmQDvVDdRsZhSpnjVua/R1ms8A
GFO6i1Mpn9DqkpjZsyrTOAQ2Pv617OzrnajUsc3Yb5RsQeiIZ3NqWsw3XFk2YW7E
X9Xanoe30/o3nznrFcCtZ+U8GsSHyNSHPdzhT+Jle0lnTGVcY4c26XVZS0JnIMS2
pLTo9kxdXjr14be6n5m8c3cykZwQkdfpV+lzWq96IRWgkD/bDZr8iyFM5l5nx4eK
Pn1AmliXR2XTvlAnFIFMaVP8GeneX2G10C0bO3/A1lRw6GCkWIW1rOvistlzQTOZ
AXETHJrzdiE537A1A95xzzxMyig1dtJ1K4QXImpkMJLym8k+h9OMgjplXwugdW5K
ZKoLhoz9AIbR2RJhcWMwXcAnqYVGDFdrRXMwnYj5SoPn+TFhVFL8MaMG+HxPPw5n
Z32JYY6DC2G42gVXVpDg9NUM/znvV3R9pAwkJOgl8QxPFY5oMpZjzi0JcjFcZXvX
MgjCWNixA7z9G34IzT5rglBvp1EU6tYy7EZvJUUjj7v0bknWt6VfLTSvZ9xXNTy0
L1f9FrF1ROunhKySmJfDEGZGolRqUEyv8lWFAxndifSkeQiW7jgn4i6LITx1MFm/
7j5BV1PfVGAsU8QrOIN3hCtMZ7jy8CYM/VNH/fzD41EE79YUo7WvE36mzCjL5YIn
MVNbgzAQIaxwvkVGLggoxbBcJQi6bHTqiQ8nKa1/jTYJIvLsRHraptQop9pLUryC
58nc3iCo+H8GiqPcXyId2E4+NIQZSRvBK882Y2WpELRP1ozMFfgNr1FFe3jK76Kf
x9TyOPft9AHB981XS8aN+iqBRj8FqqsqZWGecDhvC9wcWyvDB4RkZtDhkixuBcuL
J6gpqHblsof2+rOkbH1ZXdul1jq3VR890n63DIvxMBecRGngnlt/KYWdPBzlq81d
xiJ5ci/UeDCY63GjqK4tfHm3LHUVySZaR9OXvbuHrYw/hMFdePAq9gc895x6IgAh
ODYMIxe/ODPVLc0qcFwLld4w0TfH3HVGTHOznEdarwfAmAL2b/vYpjEkEjB6hhmT
l9qFlvzGOzsvty1hzOP9C4kol/0WJwVXNHO/ydb/o6sPUoelHduDeX1MBiTyNlML
SrXySVErw1xjSbgZw2oB2+ZNI1XgduCAdMMz/9ks4VqNm3W5QFA5pZP1xi+232Sn
vv5jHp0Hio3Z12tCqXUd5mUTnslkQAjoJHfrLBSp932R77uyPouoHhM/sAcpCcMH
NyAQZ2A71C3Q+32IEB+82kzKntVtxhSa8Lkq76dTC19n6F1VieHrkR30ffRkROsZ
q/DMDx5OVGXCKrHihT45NRU8RKkodg0IEI+6OvYlAd6aBKJ4qu2RvQSvcXTf4bLd
VwPUjl/UUf+QsgLlLWMcTu5OVBudE9fIiMiK7klmzFKDN59IGlMJUkTlau8r6csA
QcNxXEHJ6Vp31NZZ2rvFqJV17gdZSCOZ8zMJPrZgDDpOHYhwFUrydFRQ9i4bCWjX
Mb3vTCC97EMSOotpCGH1amVABnN4EwY3P1Bxmx9byjMAcWfRm2oV3bb6oFIY6lPM
8Rt5+RmykosIh0Y1BeqOFAmk+H+RGkRDd3lZSB71o7xHSKnGCkDv6NeVGYggViJ8
eZKhy6ErWvzYnypcjkx20KyI4/of2Kw0xJyG/vt20vXFWxjCZ3FsfLSN0gnDovC9
cvUjcfRX/cagLwVp4y4fDRCtK4fKtwjinOeTyBaCregF8WQ+zt88h68i1Ddw3gfb
C+ELJ5/lzPssAlNrfiJAIHUDLzD2SbYXKs6LmbNIMNcqWnHzAS/rc5ZC8IGcW8Dk
5zA7AujhtipEUhNvjd3qEXIw0zqbIotnkZmDGtpSBvMJaxg5skI/qyYNEI2OrkVJ
SQw84lNkk+o4lGccw0shhqKVVvLrISVZP9KL2eG7tf2YUEwzI0dq/mJzwvXfovw5
RcrWubxR+2sRYQy4XbHIMEOyCaiJsDbleKUuwjKoRzQ8NxAAeIjPbQtf+wY3LEOw
Yq1TMQn2jfvGc5pg90T/fwo30Ajqz9V5kjzL6WyDEwvgoZX5UVZd19nGGFFTWhc9
AaVTMM+OCbcLEhkUe/6l07Yc18EdJD66v6Ro30oD7Bzr1mB7fHyWfICSh/0R73UT
oNa+RYk+yk6IC2kjo55EbR4pKhZrrT5PECQ192PzIngtIdzYU86JfUHBLkX/woW1
9cKKFopPgsIUnlxZeGYAJf34xVr8Pc27oXdtQC42d6IyyCBil1QHfeswKyrPXonq
JUiS1tFObd1fbdTywO5JRH2XOBoCrHcHzp5Q5gTx4E//H3DyZu6KambEcEuYNiJc
CDz5l0d7CmD58Ib74anZ9cv7qePJtWytlg60rBKcUrFuMZJI1gNx5y2E6VzQI/sy
f2xT5O+qPSBEJX+kYMjcVdIm8exFZdJcm4If+iorP/jD0iuDio/2GUXbXeZy1Fch
8g90PdZhXj+4ABuaPvLIPslEhhrCYevmfby7dNXhi78UkAADtObhrZ3XbaeE4OEr
uY1SNBxq8zMg9vRL7ei1Zg9+ZYXbcNuBGbnQIlMnwsONeBWQt3NH53fxMcES16yr
MsR7DX4VxFN0dFt4R/cs5coDI0dqmX/cRT7rPT+Q9UJi4D+K2qSGhKqmXqHW/rAh
XsnxNp1vq6Rbef+9K4u3KkEojHk8QzRCp3zhneQII130NGHpOPWFjwIn6FlY8UkD
izCmbnJ4HS4UTXcMnZWsLbAZOiVTq7fxUt7SQ3XAbkInnB8uzqJ9pZUgQb+2tDjL
E+HPNXQZD0us5MouWbTRLY+FoL32veMCC0vhd4xXCX3lSHYh+CfKQ+h7xe+2Hmts
ODWoTxNUDlhkJCwvxAX3MFl+cmbaX8ClMzF1rqpjcmWg6F/ftmEhJgj1XJwkNmRI
t5ZrJFkUI6yJXiszMGpNgMYfSloab+0dKGwNw4+kbi15wmNiLBD9f3ZWCGK+ifWD
DgmFUKSGvDJJwlvjFemxZzu6MNhdhujp9xZAMV/wYF0WdkgbbrAjG+xBoma8OVzb
OVsXyZZZPZPpLEBEIEzv/JpIt8chplIHt6hQI2Wc+DVGDVo0CVK7vN9ZNbbUuMeQ
VhiRn4+ha5qGw5lbRFQ8vlWJNzdj+Mw3WsuRn6O1T5ixmsaRXaXWm8q7q3jiuWnw
BZKlR9DXIiuTCi/lt+tzVGS6uBvO7Dve81JKtejVM5C/CpNK+z5M6RQhikRZCnvF
8e7/AH57LwYR/hJn/wTfL+LkDqEl+BXuH7RbEfd50q1drSFGBGHIFoyrjUirYown
d+3Lxwo8eFQz8K3LemU05YUNQj9iN9mQaQYSw+3yunauGTVdxG1vkSQY3lPt2K1f
DYvJ7kaBbaBBmWWNn54whTmE8pNhHro04unscnCLRD0R7ELlFgPoFQZ0+2ejVOkw
W2XB5ZqiQfaVSEbt6liDjKo7wWcqylgL6bCTRLztnw1WeQ3LY9lfYDJZzDD/tsO4
DuNIliCzh+od7Yo9VhD2y/8DSRvpybBibutSE+W7GbBPnBd2CRZr8zd+me58bNWZ
2Nb8kWPU4tZ2VemNTgwl/e39m5m0lsmjinRGaRZG3a9RHQB2CGFIt/tocyfgOTjZ
Dr3ZzyiBQCft94wZajsYe3Ld5wSd818BBfn2a0ijtO/O1NYXQPKGIgpdpe+7q8//
zht5CDnSzNKL2gdaDtH4H8mmpkM2h6ns5sdNuiO1C/JeDdkKmtalR3XE76/PWOCJ
oDNRLXW19X4V8sinA1SY3sqbVCvpSnaj8j6/K7uacKsyGDzaWJQfuQgFAk2nAPD9
MjgCtosLfoFLbFAo/I7A/w96jQUjmK7M9Sk+He7rgUR2dmfTEAmfKVIamf3tGO/H
uESqiMm7dx0GNuQGmxTRtfPppDbJzsGF0UcxFKyyx88PBkkYj9u/Aiui1m+N5YG9
a88twxPNw5Iq5i1Qs3GyiGxgsvZUNZL2eh+sT+uxSiIidVOSLIHF9oenKU0Yq2Na
foJcb3eUhS1LGzaq0VPnPNE9jsOP8uwlCYonBuKOIiv6j0O9Uw37m8jAkrep/nJJ
xlqcFP5efNM+FmcYGAh3o8Q0LDjXWoFoKaQlb8Fab8Qsh5PD+dF5Qp3auPLIJ955
juOpFNehc8+hz3srZTutT4jYQ+IwYM1MluzQCBGpfWEePmr2IS3Rglv6Qz2htKR4
ljN2WSVueCxqXx8ufdMrm2m3Oa8OEpizHQOMP2yZFBH5yviggetxdgz9Su8RdMtX
dHdOjxgCXAtst5hJoXOkj1pkLCLpPlqs6r0LuHhb8r1EHAh/D/XlRG9K1lHSbGWW
SYxd2eqHkbje3amwBzH4NOThV7szidR+BlKMcUmxD8dHekwJ66qCOlDCY4zIEGz0
nocJTD4bfZndI/xmhWkN639aapj1RRbRt45oUR1n+fTzoc4c7OXjtP0AjMjS+ZPt
dgP0TefIZbPrhseKlmlT2RUA3XDPqNUtl4aj0SM0tY+g2W5RnkQIFe0JcJ55jPEX
nQLPeQ8JS+xVzp678abGnHPjBd7ZLGxP69e4xR+nus1k6vOY30mVpCTuCJ+4i/2X
bRxfRXeHdjRoE/RSw6gbYqP7msWx56s4cvPJSPz+rS7lA2Ty7HbASUyW/kBVCCkF
vACOmro70VJ8FYlezR3ww+ltDMP7iR6+dL8wMvIsHWuNx+dlXcOe0GySJ+eoplsV
6yZBjxpva7ADOvIjmzLLhGuWaMiAZdB5bIIitPDS/8YvbWu4Uov9NiFxT9WbWp6F
kgCDnPMbQOk4REcALbMtWVC/gjcE8wjDMT+8HldumhRAOF2niBIuXjAO0YsFK3y1
9GWKSHQiNBdfo5VlHbxQ9341kpp8srBjHRfqOFztLla6ffXDtKkfZJfQ6+/5fVSR
mX/Ptvfa/vAdyn5JfL2RT81vht9CMJ6WOCX41JHLyfdS1f4LjSjatQvZSMsVCtld
w54wHithl+v9wB05zua0I8ERJJ8IOkNp4TOWnHQ7FCjaFd5HAC3qxPFWx298avLo
MDy3AOuCuPsV9y/c7zRcpwoZUkSs08Jj6rwIPMS9b/SiDAeVdt92ZvZHHR83qWtG
OIl/gTcrVbHbzv6Fjf5JicPnA82MX1PEQFAzrND7JXn4CX9g3Ei0KiBcrBCwhc+L
9sisfmk21ETpHVthtjX+ICg0J4YBDZPYUFohdtzB+/h95pFEK1Q928Sw9NCZw1MB
pcuyAHpx8ocU4BVKmB/WL1UIPOpBOgA9gnXxUl+gw4EU2HS0EpeGN0Kg46Tc9d5P
LphkGWLi98xL5f5azh5bZBORszj47TMh0UAd4/rA/2EtfvkRfdWuZjsezJ8CyPrS
PnydhEK7UvLXSg4xSjJp5d1nsC8yJZgvJZ12KLAOwFDNU0ZNUx+7rVlSys1y8Us6
cAZM3vobCEsIgjtJAb0J+k97JyJtaper/uE/FinBmxMYJSOfgvFZdFDr4dZgEWWW
g9/RVNM7h4Q6P3qiURm/JbGMy2VB+ZVWAwjUuEVIbSQNGlL3fhu8FyTTvgvNgP9s
MAeCV/AtiUNTl9aN4twvdEdiJk/K2BbstJnpvdZ1IW6s/utTj7VYbFwyo9SDw2C+
P/zJ6BTEkdPbL/olFDIVbxhi7D/+FPErS2I+erfSof6ySaRmGcI5Cs3VANK9nBtp
5SFF4WQHi4CKrI+F+U59ZtVfym8ZwrQH6eAiQtquTuWV9/gt8PVpL1T1EFk2ZpK2
t41mqzi9IQggkHxSlYFfqtGumRpsyKH27v5uJnZYWy9YWPtG+8cZxnbjkndKeYfH
VuelrwhXON5xO+YAWAeqy/RkwlVjgXumw7cflgYKWb/IuCfdbbBZiHduLKJku9I8
mzNWgk44hTIR/I7C2QFLOm9n428nLzG+dQUdQ5bp5/HqHAJfpAgQOoS0/HBmoSDc
3Qp0QdHsWETvXltS8l0u46/sE5cpNyTvT1/iBA3YoLpgOAUvTmZeuHhUjJYm385d
vD4G74qFz2RusARzZYsgETrC3cdorkOal1nYd64nICAm6i2+e9Rt/j92BPGM7zCS
X/T/UVMc0+WuN5fdgrxEG/VUfnc6KASz4SP2nIlR3xK66buGTqXWGHmiq0Lc/bdw
kQ/gmZo8ubkY8LfJzPzXn43+D/o1G6UlBkIn/wh8Db2QZF/IzwTtRw9IeyntnAxz
galdd81uEfh50szCQBe/X04zVyZL56fRsYbgC+StDO3gMxh85+vhkdpcOXWTn6lk
1YJjPy9D7CyN1Vf2eL/4XHd7v3BkmBQA6WPysFLoPnq67gpckU7mC84eCkcAB86t
srlevG48EV8rWUyHin/dyvlK6PVR/I//YJqjExaPD1Ui+/vjLEREilPRNafCPH2z
sgUd4+4ss45PSmlD/0YYAhsaIiFPG44aPabz65c9x5pW/L7bGOOG/cn3O/z8qTtd
HvoLlusAHxq84TDJ+gRHsOwGlzgCrhjCsa4MCcKmluwibpoL/FwJaOyEvFtpbN7h
WajH9eZK3Hjn63+EgS84s3OBa8By+eVOuP31RI+auAWS9LNIbL4h9QQsYA+5FeKJ
fqItL93AmRD0iCYzrpU4vhH1SVzxIITwG8lCRKt4lAX1xHny+FrvFVsKDivHHCub
gicAjlXv67f7vdaCz7BOo/+SwsCjeIWqUNmh/QW9R21pJ37f/s9iWtRJe5tEb1t9
/FqKW8CdiswIgU07rPWbyZABiV1Fgiffo0x0CFo1DSe3ZBv3SbuWSj59isxsGQmS
Krydx43GV61CX4aXg5dvyBdIDpPgnv+NFkJgzWMmLg9IBwPB6MAwTt/gccTNAvjc
pcQ7EVaI0LGJgo/QuDf6TX6OmIPmE0Fs8Tc2NEhNP8bnkcomY86PKcO4+qWEmT4J
cq9mnzKjmAmS092Nwbb/LbWtYbn16F8ExUzp9z/ie3TQPQ7F/x0IRHqjKqQmk8Ax
xlA42omhE6mJagDbCM9wE3y9+FtaIdzaXQORoRDN3p5DQ/k4lIBnoMBNfaZXoL0Y
g7mXn+f/1vpAkhmnP3ztTjKljgjpveJjKtw7nwC62YCma2Hkdqdq4vUPvx7u7GEZ
tRCi13McqS5f20RZU46BSJxBEGbuu8umRh2gACn6vMlRHc2cRq2g+jyL84CryoPw
OZLMkniNundUPxr+u0xp/gzu3kspNznh2FSExQfEz8VQNeUMiOw/ezK5JfQfLDT+
Lo1AGlwJGKRTaE/2ILNH5b6LuDRUcwXQwmEyocLdDtqEBC+YTVa+ut0/WW9LIhKd
pP+PczPR8BXF7RSpgerE5aQ1oKK26Ts26T9eqBKSQ8i1QoStOCfGoNrvHaqheY8d
MaQX7QKvXgqObMHGB86DLS9wdlVmiSYBn+rid9ttmQnRCosEUy2neop4bhJu4Gnc
2iBGFDJNDlDQPJWr+PIEo1fa/eDN3iYe+eNf/psrI83dacclJQFEs/bNr8IUmmlU
JKLW/gtH//XYNCAktpmIxKeM0GXp3brxNDvMGzFF0yBfvFjNXpWRmYxcBuNhEP8A
7vaG6GaWsI3VhPQ+5Iagfz0Sulll+LaZgdlxnHo8AGkfgvBQchohmcB69yLget+Y
QCtxoPMMp1HNSvEc1GGU9A4q1AT7yERCMY4UVJ4ztrZ7a+7du+mm8cvFeYPCisv/
mDiYeYoA9nVfqU2pjl1AsipiAtM0OtWXAJGfs2PRLMzYDSHW25esifvX5eA5/+Bu
Tpa9vXRSJ3Ja3R6RCqDOi6wrAwPF41AlAuY3IVtG2VtKu4cU5okWd5uEfPJXOn8W
Zl8ukb2UXEI18pyppoaOzjnnvcQVvC3h0y34GQjYWq0GJMpFKN543eK+k/2TyfAd
EQESm32rgblf3vc9FhR891h1ZsH4Nc0gPzWoF98ckCTEWj4zt4jNOfE6jI2prNwa
Hrmc8vqvnzZZd98l3Ja8T7B6zsr6h28PoUHn7ajxRU/3hGYlxaP41ruqCG7RCTY1
SwTpP//QcPWJHqOjQSIT5xrHvS58vFVN/HokFjDHlOW/9Kj84BLIQIiSHC5+97AG
lLgSdl+aob3BCasE99Ml6Sc9LqysApCtIeMgpFrCfVxu6e2glqghnwWHivbaHP5v
FHBMjg61POYM+dfV9EaCFVvDhkld5rcP73LFedS+a9693CTxPW/c4iAufn0eR56K
7e1u+xlkwNzeR48++Hl9q98Dy+DzRgpkkV27fhjMT4kMIOmQU05VdEL93dydhbGw
iXUE2K1Fvdu6LD+V+AC6GmkrCjuW9o3EcWn92Gb/WYC7BThcZPCcZXS4AlRMCMdZ
MQVmFp/pRTgltty2eIW6yt6xxSE7NsLB3ctJ8H80s45gk69iQkVbtCQk5iDY/Cfz
q4hwANY+YEpLMxlFmB1T4m6CsTxG/07zcFmsa219w15z1Cimm85V1l1D2ac9kVkP
YkEN+yQ8HgS8mtJHnR/gFmmu0yCqJyJiwGalRk96UZ35btAEV1dvclQPDtEy7px0
B+ovqVj9IEoTeXeioNLrD8Dc6/QgytaVNvbidviezGM7i7CmCE0GNqt/WQ0XQ2Kb
lYltHA5+0pLQNcclxvPt/RDhJTS9FrjTVcYQRACC8yqZ1z8gvNeX9nYzs+NWizuj
m1NebMTMexGFy785NRDjshSAwu3NCWDhPCviVUBwI+YrNK+9GDrP/bLHzLpMYKWA
9Wgxh6kt7N/B1oxRfhXZxN6utXK1f5ANbdyXov2v1TtkUlDBCdbKfuVT30cEVvXJ
KqAXtzgz5Arj/+CmT1ZBGRGmDMwaqMwytiEJW2CySCfVMeptGkJVsQ2VmVMQHnyC
fcfC8aBuPVOZkcmnPGURCqM5vBSS+ugcN1P3Eo9HOghmHWaXDsfHnrTUT+7U2Gcs
k8/9Ub+FBBSMFopsCL0ZMKiNMS6oWHvu2juZSHuU1mc+n3f9ElzUItQD8jc2yu01
+8E6/uUtCPVQbXRtAdaP3v6qYsQf/i2Dvno+L/uHqf+B4y3L2e/ydVkiuO5/4QrM
dQknvoxDq/F4C2Z3x7wm2AJdc9MQSKovV1cupZuNGv8OijbJiR0PKuxii88gauAt
kgh9y0xrgF6txwuJCuJp8rqh5103dsyvfmxSFYDPwb6KAjD2XlmpToNX/4A5T0v0
0/ZxIOUPF1CG8JKczOfjRCAz9ocQi2ZiCfx96zihMvwfBeN2qqP3ugCIOqp1xjm2
UBcSI13NYjRT8tVXXoQSQFw2JU8iXeCNz5hS0k3w6xKMzx4rX+06H7GWkVWfWdC5
M+T1tHItyOU28EWxUiKsLJBzpCu5DtVz9icv+/LGz0wz3RrO0TundMz81LeRCiF+
hNYIOnUjutf2IF6MdR2yN5QYqhZYsIq0OacincFvAsZyWJ1iBfsYAZ6aWtj8be6o
4biAkgJuXJ7DnGJo3go9XFLx0qoePTYU/TNUhbOzkITlbSmh3mV2aZPLmN1vGWOT
Jfwj2YtF3OpwlCVTkTiMX+0n4Q/fjzIyj+CUlwiS0b5yga5Benpxe4sIMyubaIA4
glWsMx99FsTAWfFh0GV6ai4CfD1nDHyG/bHVLotuka0UF6PY3vHCicMkldMEYpVe
le69iTX7+jBeSji1rCpAAsHZIH3mvJ9cjk2JMIBlD+ZbnUgDZYZ6WlbmMoNgwNtC
u8EeEe+kE2DQywK3bW2m+WQvb4USEVZgf9YUsgdDkRSAjyDkh7+sHVMMSn0BtNB2
N2fk0MA/SIIIlBnDIvqxFx08GetP2k5xDnEgnt6/+EUgR5mxOQxPNSo1KBUusKzU
6YZPfPBLGc+5XP2+eWkzMjVXPzVfOnkk7IyfmCdxF1wIB2o1whFtl+yP39dUZ4Wt
J7A7ubgU6jqmX+NbKO0PM/Qlml9SbtYmGLI/0g3MDYza66o+VflwqpZTIdH5rYWw
I6F+R8AYp2nIE0NSNdf94Ew2OtZix/DoWmz3Lkq2AOjQVjhXbBFzGh8a2WGXNufZ
Bdk6z1pP9xFqZfv+jcd+n4qQawlAakbOdJcTgqLq275qJ2X36kgG70IX3vTH7ew9
TT+IrJ3JbOzI4cDWiHDDCyHXs/leCPKdIPjfjvJ0qQet54lWuEM3i1vu3iuD2w3Y
1qxC0+iM4P5yjdwFXrHPlW+pMhgqAPvJyFZjEKq+AFXxGHcymiddP7nwNpt8gtUt
MnaVjrcioSxXM7D+oDHtvsP1PZRGnLzFHSu5qSlcezaNWlZhBWYSFM2JRc3mhCS+
Jngn3aXHsAnMtut2aX81qYS+UKL/UWl1Lpwe7hKXREqgxsfyAGlLmZINwT6uNEwS
iFLJSWxdHs6ovitfnJqGS6ramV0bBHkzZPeWTl0TaYiN5qlTvooA9u/spaWUzTQe
fL+8M5U/LmuoGKLNTte1VcNUIJmP2sbwBRFA+FQh3DiRPsS6WXB+QPM1dabz+cJQ
OG2S75MpMVfaJENFUk2XnYuq8ym93m2DphM09kvhREQKCcavJuJFf+abbzKaAXxp
vEfqMmT2KrqY2+efz/RAQmv2GmUy/CkKNMRAwgKFL9Ka/vgtp2gWFqikzki9KVzJ
SYEDMziVfU8BVRK00pf0DJ8vubnynso0PE72e5b61OYboacHqfXBRtZmvbbJv98C
agHGRCeLcLdxMG9/vgXPDUG0gV3u7LZOkzAXYHG84MMh9H/+kfigtRj+fdQaSWKA
lHMxq1fxBLMksUiix7c5CQyEFR37u2xjvrkOS6wHMoUDrZY8R3qOI1ZjAaxBgzM0
M0uC0cfzYlyh0JJJDJiPytkR2E509GTV8T/6DB/UvPDpiMXiUmzj9RjjMqaoOGRU
8LQErUs0FDYVp+H8b+w4HwhDG/fXsyl4lGVTSuXcWCTMqMrtsMuvALhKysz8qKEE
553NafIHtamJOBqHv8xnTTJfOOoDc0Hmz+VWEL9cX3azGtULQMl8PRgJV1vPzjuh
Dnvo67QbvuVJycC96NPNn22yYPDBR2dOxL2aFW/ZCG2E6ivuToPwVfwr9A3aXEYp
HBguN5c4q/l6PAWXeino3Zp/3kVvM8LXVtKa7Er5zGtvS/6UQafqaG41rErwJnnq
hkj1fXbmxoYkzdDYz8BXg6c/7+fzup4X0MSNn4wRB3wbUaBi1gxi9XZVwhXOjxJu
NJupbkTR3jbiTaJ1GlFPDxOCbBapNENV3hOOdqVTX+jzXm98vWHzQMC1iQTIG9+C
GT1AZDN6AAN+es3qBTOy2SJQebVcYPjwgbEbvJ4iptumgYre9QX7depk162qUA01
4xIauwyQYSuB8I5Y0iNa3WpM7I//nLQwV1oNveMy6ymk5BZzESh9NdgXr1kMbafI
jAjrWtuIx42xQqXOok3Bc7VLWwygnG6WHgmji7weJNAYj0GzBxzZNLUdYBxFsxvV
t55+9piphUOHQ3r4JSag0fwJV+ukt0lnHLyVVMOdGw86UUetBf0hsYAPKIXr7VN9
j833sL76sB0eU9UozlaQeXBu1XzXJkArHCeDZq2To/J7pvvqylWS7azK4LZ30QDI
6hrTJZO9yo4/7uz/XrM0RFQbHg1QldI+9wz2CXxYeY0xt60/h3n+ggbDG7IACA8z
B+Bj5EwiFdEq774i5dvBJ59k9cfiLqsGAL6Y+TFj+5fLCGUsCtwo7h0gEAK7dnL0
1GrWWMVKfSSchEwEGmGjADvqiY1sCO0Hg9byDj1OW7yHYaqD62heacSmRryiBVgR
68ZWvIquuKJIlAJE3YJsGvs2fbpsXax9ar7AsU4XrepL1gUfBx4ggVqMR1Z2JXeM
4XrjFd2DXLgvw7x4iaiCLVR5joOxgj04mkI2NX0XfVHoFwhF0OttT1JCPW7+FaAG
ly3tb1iqeWdK0p8wqn9qkFxy9agCLR40Ar7IasjyqoGh93H25IXmRUTA12cnzCQE
JVJK3Hq5O4CxTYa6BIFLgEvxl2SrveB0TcT4rvr7WX29yRyeW9IHhuUB5MmFkNbT
lBaaKVxskgUtUACz62lURV768GZ3HEpoce+lFd+DYSEvEX5TFFJqMN8XTKIQyBJu
DNCmVr8WP3trI5z9OVDV+6HSwJ+PU6ZvnORF1TQ8QgL+xzTqANCfMMr0GHDTR/G7
2vWunv9NDD+ebY5uZtVQyiudScKBfCQNf1bgz+GE0/YBnhfCQfxfZiWDU8U1X6Mb
r1fY9Ecfxr0CCCqp2lSqjIlTcG3bwrqMrqOgNQktrrpeCrTFVN6Wv3859XOlOQV+
jm/P4ukFZwQJkiVXMwCKso393/5oUKeeNavoWQjV4QISsRQcTOxb+HQJRct+Fz9J
Ci0QQ0jISvtPxVcWNpbKQqkgN4AGFMTnCrtbZsRkvBSC1NXMqFyNFy8tSWyLqSBi
27YobrHZLFklmiBmZqjA2yHOdQ/p3SscGFjv7NDcE2oLjLVs6enKJvTUx2pbyAB4
m4tXlZkt4g9PTQK4ZC8KJqxEE2yExgIeJRCkiiQK/1ZRztj7gfwGuzfwnQnroYqx
qUAf6+EhqDBIuRxbOJpAqOcmhB9V8r7DYiP2YLFBMz5xc8hOewu2i/x2TP1bLbw6
Fm0/Po6lXbfkDf7cKlosSCjn67DEdqbUmhvVARI6fv9s+biyqnF9Eop/LaOA5Ad2
rTmvtMV/PrrjnyPFI5sXyRRj0pAjPyTGeUFkHoNHG1wyM5fgeqHDGh6SVhFRko5x
3BPS8YhSfiNbwrWVyfIRNzWLeBULlW+REUas768KWNEJsq4TYpVVDBolR7ysGHel
ibxnXD/8dgky4MWSGq3dSk1Z4ti66ZvvCgLffYj3GOLIkTFHupZDTx7ozZG8afXc
JMxG19WUV2nm9X1ATkfZssrvtv4kw4T2P4Qp4YbFvzGnP6f2pJbNy/BwRiYHKLut
ffFkwTDbg1qD/NewYn2UoqtEWf3YkegrpEuFZaPyFbCg1qHRaZyr2hTLm9GtvWTS
Zs8g0hOtN0mVFRx66kXW/pCy4+5H6QHGTM9Dkdmf3EiCwv+3ZfG0pAsUu0xvdPSW
ZIiqT1Ur2XC2JJyAw+/sXt0uAENORGiN6e7XxgJ9v8BvwcPbd48ETCY5SNhxl3CV
x0e0nSk2l7/l+S4HeAxniWmQk0Qz1r6S9qmXA/Aydm+MBXnQSi/YHUSZljQQXvYX
ahE8qLgF5kHfAZfICsoR8A/oI6SxbsBsnOyfe3KyIcglXZf9D8w51n1PhFF3G6I/
TOr0hVd5Z6v/voWK0jlsQfNh+S3+vUMZ5hAV9OhyyBau7/TkmtQzk9F+Mw/LDvUr
pMs5bZktIZqE3dlVaH2n16kf/Vow1JFtLPAlXQ7DIz/J1KCm33lE4iBkSk4wUUnr
7kmFitMiXyUpC90aK6ckhUXmqUhjsKqrtUGK4p0Fws8zBgxWhtnVWiPIEm5PDgIm
Vl+dUGJAtHFEBlrgxmfcm1lP6gQq3z3jZ/xsIDmFwI8wvxAxwxKjvVIwOALGWqQJ
qbWhpaP1IP3Rkd8KrcLYZiL5yNgYTKi0gOcwBv5v5VxPz/uYdiCTcmisU3zALM/f
J21hmzzEZ1PnLfcMy9XojCEEeMQ5CYDHAvGzd4TAzWBsdke8PImkOrammOM1AiR+
pUXQWA1om9Wquh6kZSd6QFCgdyvXvkHCSNLjPgxo2j7as38JdZXAT6PgmIrO+KVM
hTOxg7V318AUSQMfofacmhmzMDmhiUpeHKb6T86IUijJtkh7br8CYJ8N5XHcOgFT
H2PEjtvDDMD2dVctuOGB2WdafeCHR3CEtrZSRsBk6ECemcVcwUP9vBLqCkhOXIG5
y0A8srTU8q02K42sWFxlzsXtj6Aj+1JGqXSaSlkvtaP7vD2vc2E9x23s5DKoTeHK
08PELScxtKmgaNsqw+1LvbFh31Z83SaYZOiMuR2Eg6KybzivgrWMObRWoRydgqCR
5cNmVGAPwN7lUMs8vaRkGWQcA9l9mF8M9gcJFZsXbPZC0PzjjvoPtYmFBpQvi4wq
9Gr9ZLp4BOMqev9mLIgspeqOLv6JPVnenTcWe5/rNpwpZAdBK0msbzSC0LpbvdPv
IR7y5xJR7gHYMVWhyGBUc5FvWVVcRusk5/FnA0rRjlJyXd9hPTc7PiPuwrNC4zwG
vjeCEjmggXXjsWYcinE1wIh2ehxN5BFXbH3kgFhPOx1g5MQUjJkjT0j+ayVETnDF
NtVu7K3AqJEf53s0bgU6jenLNUS7NoC7hMCRbbntGtYVhiw53n0N8pWuqPx1CpCd
wP4lFFaz9sFZHnDC0vX3QxhXz4eE7MZ2KtAPwUGvmYbgjIvb06PaRE4dDQJImkGN
AroD+q1HVTFqRSVMBanaWIAahJeNGbEuEIpFvOW0D4lO5RzVO+9ZQOVonxYoruzC
IiPicHTXZrlXHf9hN/XyQxLX2hL/uC29ouN4BBdiegJDFfFWMeWuY5cC+RTNVrP1
fFM74aucOPhFr3OH9vqRqRHZg/QW1T2AKJs+Qe6OA0V4wSUFYANlnv/MMMY9xG9z
X80CL/GX5KUG/N8zrZwZ5QBrt8A0SOBnuiPDsK4kU8HVfltfeZ7e5ck1zTGcyQvR
MzYrNaorB9nEwTH8Ts2FhGXaedRkmd8Z9pb2hBtc5ObltlWD/X8M/iN3dhjhdGJG
YuQnk1m9gwIH3lQkQPwe1UAx5UD7Gt1tEKNP4NDL9JjnZ4km5Ly7fpsjnLQeCT9r
rxl0lRi5dQ/EdYaIEWYkfvoYSm9GwiB3gcEVWcKcGhizPZDMU3a+WX26kEM/46yn
S8sL7JEIQezY9fstMp+PFSa/IWV4QoErisbY11bYivXm2ysthAk6w2SFu50D/H9O
GiqVL3VdUvOGsOHA9LLmgrgO2u3QuYaG2NVA5CHhZdlMmKacawwdIPZq+KlGHoOg
8yPwzK2pib7rrRBy2gXGV6yj8XfcqoMGTfrJHkLADsEQAQ/ZhEcV/n8m2A6/Uexo
7ysm74Wh0Y2I17aAya5IdSAtHcwjRIObIZehKNLtzJ0pQzV2hzCMSipbZKukpt7a
GO38lQEZ8PtqVqMvAIEu2esOeltSyTUwaAIMSWQFkuiyjCf5m3KRF8SgT/7W+C/N
y/DwquSqEmRJQeG8sMoKKKKNiBixqlsUE9uBLzt6uMr6a5g/FcAp0eM1WJyhpEQ/
rpia3VpQ1BdNFlgdsUhqNoccB9dOZk4fBUVDCwmnOcW+CvPEduOdZYWTlmAJUzrz
rCvkGtYHNOjTX9W67pfLRHvYsufm80IaUzgQ7L9KtoOCs02P9Ko/HaDDzVkNnXh2
HchxuBMVxvxWv9SRHAifACaiHLdU58eeV48CBzepwbYMLHNoDtaG0W2liClGv1ap
LnoOts38QrD1pEUyiHh/R9EjgzN1kI+hf7tFzIK6qAFIyzmcgeAwgcP1xEzHZeBQ
Liw1FLTrHj1Rw4psjvdqNziURrrFOsOcI89MR+BTwvOwy3wzx0BfbuhQIiI8ykN7
teN/DsXK6Hv5OlCx+HoYbpd2ApmQ5Gji1d1e6YGsZkyA/Oj+4kYA4Fzty95LIB23
ArBKonYEf/T+tzxs5QYgGPMLfNbkKL06a/2z545eyRutNKMz/5bnoovkaqoYcBmh
pWRArO9ErMgLqQc5CiK1QSTpAmbFf9arI9r+MdF9nvD8gX+5dRBjsd4GagL9n63/
zvuUhXRf+lWjpEzAVW8rWx1ym301dG9Exczrd59Xfby11jrD6HoOLge9AxK599nL
yJctRxxo24VEaDgBIYQOC4BOq80K8CRLLmF6hcO7UfSL5lgbZ0aDLjg/zJ2vQort
XaRVgnSpvEVSYYOYXmYt2nCqLgfy0vDUV+Q6wYtXn3m28/QMvdnMtwk7SSf+VhTd
y+07fkgDtsk/Hy2JcFmUhZv6MtgUoVPQpAG3OcOLuKysPUFupND2d5xA6BF7E6b0
JyUJhk5aTF74XU9nplUyQC3l12Nj3MDc+ISY0r06Vjs98FJ/AzCe2Am3v2DwT2oU
X3/E2oKi7Y5Y3m/ndg2JVhwI7WlikCNv/4QP4n6tUj3vwlee7jrDQXLIkjuayqVR
hg/xqngYv70nRcRwclDZwlnPfnDVDV5w0yBv2TkK3VHsG/YV9fZo6is7HswblBnf
VPz3oKxu3etnj5Rw5xCCBINfg2EaQCZCPFZjE34bVlhFtKU13JzHmi0Z+EsH8CSx
psULvYwCJSK6EA7zJ3O3LXepBi8tt0XRHgMh+0qScrXqgBXx4pa4NR8u4MzaVZJD
MxoKJ0bBTM4Bk3cfCnVGE42fPuUEoeGw/9t2RUDmBu0yAogq8IDIYP9oQcN7KGOZ
FnFKFEbDIBGTOrcgEy1qShEFx7LrqxSbyqojwIwucgNCtKIhDH3s5t1f1QPPR8I+
xRDa9lkc2XsqLbrtyccGyT0gmjsTlS2HJ0dV0YnMsmgaDlU954mE99hUX2l8hyj/
Sn42JHK669/cNGZDlpiWTkFsld+9JMjMJYij6OtTN4uRTC1lNkJdtLeTV5L8NBBw
mzrv2y6nDXfOBV9Npq2Cag7v5EP9engIPBOoSsIEtG5agSHk9eyqsUuja83IWzRJ
aZLkm4xPTzC2/JmndRPREA3AvhlPPylYxDj0XTdZKzhk+0LkjK5OrZ5PO23joMYy
ZQFC0WgdYjbkhWEDbWxCFvorkyuxLC4fiak83m/YRCcpXZkmvdroWwOXuGNH0BMj
8El0EB7M9/pc90R5McWWEUD2+UyprdcNHnVQtgWwhlZPHsJAGUT49/NvqmwnMij1
k3zJ9kTLwXUhQUt1X3NVgirQBtR6K426k9cw5Rrb9RH2CQXvxEHqJ/+D8nJX/9qF
/D6cQ8zv1vLMhcr47i8H/OQIRAio/nrivuI7h+5apWuvxJ3ypEROdxu8AP4lTwCF
6fzSROaSCDxrIhEYQQnvLeoOczaHEtFYuZV9kz2klcybOiwKyzJAXiPi3i3ti/h/
mBFALl0mrc/0a1ttRmsOHG9LdQG1abizOfLGupygNSuIp7Ea39oiWoySafiE89/L
JOZ6nyXz3x/5IoO4bc9fJfHV0jXs7TIOThiuILbo9Ne6v9Pug+KY5AvfVoAGDlII
HZPSD/qzR6DUyoxiw29SlYGIOXfMi7IOzpEIiSYrPTkqgQ4gmRzOkVGsnuYGIhpp
VXU9ZOg8i1m6A2mUwLQ/LcG8izv9rfxpM/qFWNRCXqJ2KUJsPbsqi9mBUbp6PNi/
vxCDuTIsH8yuGPqY4H8VaDUfEogQ29yol2nu+bqdo9SZSOZa9kA1Nfgwf4NcxXEp
UdrkE/DuSwThyFPBu7wLp9DLMo7TNI8qHJgakDD8a2iBgjkJgG26Ev3XH8P74Ci+
0T4dT2uJoCezD4WK+vN1ZxOETw/StNkJELEf01xc8uQUQ3wfnTixAG01f1mT9ivN
7IJyvpHzo64KKAEZ7HDqONXcvqNaF+aUpW7L8C/ePdwPKz6paFbsQtGHwOl3k6OU
eecACkSjDP+f5S2Btgu1zVrOp41c/CC4S+G4AX6Db2vDi1yhwQBhNJmu/YWgVwDc
VXyCNDQjuPh17KHZjuRwutFd6Nt4USUuLoCKnDxHuMNjRnZfLi/OMs6TpGnuQEue
fY/ZnbNDutDqA4DovnTihTtHYuMfk1g2KNinQdrwk2hfVXXbGMGaQ5QPYRiIl5yG
88WOIjSCjoCkddwztzfFMYMJwBRCyPd9XKvQFq/yqLLdJgghfz7vadYF0XfZuE+f
2ZaV+eA3mxt5Mkrh1cbjEHr1Bd3YYziWrNO8uJOyHR4r+xD2+CmLp8g2ir57XoA0
A30Pf4ED7YecbYAmB1rcNi74PP+ck7Oc+0SOhoNBRm8YZNJyQihhzbEQy6kaJ++r
Cyr5m/9f4E23I3QBIyaLjUA0P8Z2frtWS/re6qab0POKb0T9UZ6VTjzRmUQdH2Bl
EB+IQaGeho2q0q5DsPBOntLiFRFYoy0Y3JsVAXwZYwnnqIBtkw2maYsjeIKl7pID
CcMFjDFqD+JlvTpbCnirA5xdDJk67T3I7CJMhe+BO17vWeG49ZON/knEM3Hk5egZ
WDnDlLc/6odOhO+zfysONH+oKLvEV1QtuzxKanB8/tYma1oQWEEYsIVByBdhqRyD
ee90s3ss19/6gCWAEUbE2DfkG8A07azNV6I2ucHRo9s5BMDZb3uELt6mWheb6QZ8
x+k3z11FOhvFIv8t2F8KER7p83YrN+d3lK9LSAN/SmLm2iyN9/qI1TWlgS7fJLa9
O50XNsniBI4DEW1NB3LJu7YSaHoGSb3RSJUNrUfnH79RXWE+Im500Aq5pVe0tC3s
a6XzTsNE/Y1vL+kDOIqi1ASunoCUKkGPVX/kYMXQQ8XaNSTtshkvAjaMp0eaQqXU
P9Tt6rMxajdjBD+jsnzQ6/A+X2vJoCTx/cWZv9DqeyVKX8Hij1PtdYWXSwCLGBG9
ybfllEnUfK1JT2nyOWYbqCYC8eXFk1jOOz/pawDd8srb7d2mKKkUKEc0Z/ggKvDR
bdCS6ID1/sTIxdYrP8ZQxygy2jtrqb8Ed0D736LGgbUFxHH9LnOMGI1DnP9jCcW8
wSmkfAVtdS08A0co3GBqDG+WVpsdrfojOUEm89JnNQZ3WFsB2f/JJZRz6G2l5Cge
eaW4HNIvvARmbTK4rpfsVL+xkWdtsuXnxorxuXCSu5I7c6OvWGVNpJJFjd13W+Ay
x+BmawCv3IFw7imjFhy7OTMsgonFbtHQuGwyydvg1JsPsCv0FF/gxY1+gz0GDS6i
59zBfARyUYpnQy4BgMzcpTCikSdxLmdg+lRVcVXPflVNiJvGQ9aVWpbQYkDqMHyj
c89oQr9uoV1lHo3L0e39EawdGQiVQVVXZ5GpQD928ThJu+fmLB7JeSkV7DtMT3XZ
wmpFlxt6wSDfr/Kk1urEDdi6vCLDfrUQseiGbfFg+wg9XyXBRaX13FISuFpUo+nh
2a6mzOG9viogR16OZCEW91nmRHtxugkC3k14ULO3Hf+tnNzFZf4dGQVDRPwop3NF
3kF/mQVABwRwQDEW3AgE8sODCDVGvz29vh6XBIuytr8sp0qRdeEZonyUdtTG6PbJ
RDnjLVAPSJ4pTfws11U6TBXbVQAQ6PxWXZ8ILD8s40nhz3FRbOftjvZaSV2uJ8F0
nqG8TbZyQdNHYemHeSgbhLNVgBoaKTBkw81F7/566DMpPMHayVC53xJF+w0z7dhH
6fwzBW3m/TmuwrY8lGDTLTGknVTi87cTpOXjVo3NoKmL705WVf/sadAbpEWFeUtk
UfaiTKcFbOOEkCbiB7EsaBFzR/l0nczVSvhHPpUW15CvfPCUpGMjPu7CP/eBZVl/
P3+XELT4FExzMG3hfoUND7TTStzyl7uS/V3DVs8cVBAGIZNkmQ69iHa1bBn7gmMd
U9AP0DKz1Kqdyn24o7HpZ6pKgJTFOvGGzORK5ZuVJBo/brloAIWIkf5/TDxyhpsH
Zbs6D2Q6NGn1lP5MiOC2Em6ghsRqzjr1ZTNhwNzL+EwggNZVvhHg6icTOb6v/73/
ZYOAxQoSXWqhs5zMzp93IoDaMVeNDf2C8Pt/AJYIXKgAmPCO5ZGfR8nxRZJYPpqZ
bej5zmphQs9d9+IIwEnmHP8BuQaoxO2crXepybwTlgrUEGDN7m/GvaZXyPAAMOLm
VykSqenw39RgR3hK+3kRAw1pkN67XvOhFTySOYSRGmfTuj6gNlpDfbgdntDxe7jV
uZk44ipz5Vth3vkM8E3S8Ym418ECn7QpqXeuuiFrfRbj1XjMfB7uriNOQ5e8rSrC
W7N0yzjqt/tFx9JKDrqt89A5gxfGHy17iuoUGQxvz3zaaMlG2M9embAB51m07g31
g05DseYzbP0Hz7wMyst4gH9vQ7ba32BSEQbGfbIGKKuws7VV53L+DA9koVx9aOFM
tMGuYor1DYfmhIXg31S72FQFeCaqLwRaIAP/8fX5FpgQYAyTyVtzZemS+51sVj/z
D0BnjCu8SPMTmITtiOnhtnYLoTajLItQzgySD+Tev+oBUHO2s0bF9EAEt/Di+iZo
u4ZvEFX7eqeilmneKb3Y+Ae03l84IVTPBDJrECcq5iRDpsPDrON4yq4vQaVMYYPB
JSEF6W7AzvM6wcZ2foNgIfmnbHgqFQRpWBf0p5xlJj0hLMFhhQP0/GUDmqwXFWsJ
3KljaAq/4uG9eGSLtwtSu3SwIrHC09FyC6mdduwdfoYCHLFYbxE+KSYpGPlpY2KV
Oj1mdtwyeAzfjp8onEeFN/koyi0c8QZdXdp7xiHd4ta/xPBkJRpXLHPqrYTlDD54
0714WyQb0XOD8q2YAanWuIFU/jpsAgy4xIIxL5nWCQue6AWDewL2rGJtdLS3841A
Tto0Hfl1PBtD0JHHvxcC9oK9q0x91FbHcepDdmUxsDIMZ8DAoQYEEX1w4iRohfkf
eEjE23EinIKpjKhlSamerzf3GwaI48DhIA7U/2Vo6aZENzdTEKSy1y0J9uzhsw8Z
WMWbc8qBs0S/1TFH0zvQFjstFWN3t7qyUSuwV7kQN94IMUPHUw00jXaIylPg1Kx6
LMqE80EI0hv1qecOmqGy2ivf8/oWOjT/I9sRaqIpuIvrIWOaaETnG3nvUVdxHv2m
JhyN2wLDRCOtpUoWb9M6IdKb17zqPQoiUqng4uvkriUjNyOPBxPRfB99ZIClJ9sn
fEB5BkYmFqcABYtUdkhgsP7+HbO8uswXrO6JlnfFghBfGjLJJKBORH7KS70MvUC/
XOW2jSCIAK9/2Dgq7/PgPUkrLtWo7Y29CbjaAJXPGUm4fJoKLoYqSFLiKyYDyTo7
ajPytSJMG0zI1nHeSyNwtYw5g3tNpe6T1IYYeU6mrUTQIVICfzZHf3GUaoHg7Kf0
ZFpNO2vR0jHLHRp2K0FO9nngQ6Eg3EZq/jjhVQHM36gBQp9gouk9uZB1gIlMRy4O
iwZ4oOWUMcOUxTycLwrayFFlM/BKW2PDuQF7/6X89fNVmYzfzWyNFGJi4/T/d1h2
oIIGBW6LH1NKnSET/KnNaagb/VYwzMOJ5KXtbubuWwJIm8qBqPMuA+4wU8OLbJ8v
FzmvV2O13kgajfmrDvgF3B3pF8obsAQqLKo240FJ3TN8K9Go9PkH6kDeqjHkbENr
9xZzRoiawawMzTAhNE0VFdCpoqUCvfKHyQP5fdMFdHE/N71ZiVCC0ETm3mwH05XR
jcm8Rxa+sG6sddOCg3lTG0SarobK82IL57GXYNnT2YWDufRjC4mW2uaOl3Hrg46V
GM0I/+D8/XwA1v6h6xKaHAsLJ5yz4MdlDpkBaQ+jOHRBtX6bu6L7AEgaJGOH78rl
jWxOPEQODNamNeacMB7TndEM08zy1tOTryqxcNA/l9xd/zbbz7k4+LxK0rNMK2Ij
J2cQ03Z45MX/xUvWaGrtsA2XnKtmKk99S1dvWnpFEzXWPxCpwGXPbvkInNG4EL5a
wfGTcMt1ThWUFDxjf5E5dgEPnzDh5P8MfxDNznGbFSJQUsRHl/8xn6g3CacMxU7n
c7TnjNBrIw29iwvj9VeniIJIHxqCyFIcfvRAz2rVN/ZRNpAort98CvdGYIlc33jx
M6RKVc3Ewxj7UiwnvTKWlPgv4XsmPZ9wXWK3b8scNWL/+QgLremGVSSiTckUZrn3
CmlnJpG9ZzAlqLysFqgMWmXD0cUgqhQJD5CDPGskkerVFkd5B23dMafOsFkSO/BK
WOxcsYm/yGOECLWoApnxTGgK0GY875E8gthOEdinaYl5ZwrmJO34pZ1ytAAu7JDu
LepXxE8HOoUEf3GMn3/GGxh0Khy0+Y+/b2R8O9eqGmslVLxtqGT/IJGe/5Cm4y7l
jHDJat1KozQSG7swF6O8hDAR+r9VpCYhCGwRJUYup5WsQ5igph6jSr0wixTHuq3i
QTUY69GSQOc9Dqnp5xTRzu4ffMcvSoKr08Y5BSHdLbu5u4tySIgADGVyFJvuBP2Z
Bpd/07TZC1Wa6WIWj41sODx7Crqiuku96hRnALRgJdCkKzzspA6BYYN8mEkqNuD9
ilO+bhRP1C3ih8BRvLdF5iX0ii7BG6Q2Vs4Y6bM1T7Zo82i43qbcm4t/z2q42VSL
Eo+2PYSCCNZwDfKcL8mIpQphQtBwm0k+IWaDv7EgxPt5BlDXvooMIzJUc832nE2u
9TyW4EdvEHdxqqc+5EgnZuSpkTKgnXKsDvo0GNTaaSVjG8EnTTGTqHonYJ7a1rba
JqxCuq0GEPvgAX9mZK2ZjIgLvqMQ5Fp3PO8n0t4EZr0DHja/vgckSVMi0/GBj4aU
A3Bijg9WZj142y69Rq43zUOoTqzVhcgeo0qVDR8qjNAG8aYuK2Zd7TodOOOZhHMd
alL79mPRGOnZ+ggDdfSu7Qp/EwOG0jMWkAeJd+ct+x5R3V9E24gfbhTc07w9/jeQ
IkTSRdYs4zcStaslGvgxCXDs1U9fOgY6M1KGb9SlUY4krXyasLHpuNnFPtkC2Pb/
G99A24cq9RKOTQPssC/38u3+9H39+9GoZ1j4MFM+crvWfrS9rp20IMBIy7oGeCrk
j0Ht9Jvf7yUoXEAu5uaD8CIniueenhPt0DIQOLGwNiczROm2waiVZmpvhzun5HN1
DX+2ZhhSUHVVr2QWSxCIbhR0fqzjxefnHq6ctmBGDoV0qn6jNPnYRgK1tGaiYTSK
YGNTqduhKB3bWnucR1ZPiUkiWOglieZEypCbH+Puc2V1AuPqg5D7tIaLhCilxQMY
mgB39kIkJf8VUDqXH8JAtCVl2Nw9PEtOjaN+yoFyKsVnyJCDsqUXSDfY0pxH+kKy
v4lN3XsWJHNIuLmG4O5dhWfq9O2uRtIrOF3yczQe1wT1oLirYn79Q+rfs39A0E8j
bdSNpCfLeIK2OQtM/VHjbdhYVM4Sr1W7aK5VKjFDPdyPIgrhzELdOCDAYLtLGC1N
T/r5nUU3EwoyMjVuL8KX/e39BPNH+qLx1P7ZJ2XT0eT3NXFN2UbPKlKBA3M7BE7W
tOhuaGMcqix7YNmSW51zzG+xR7He5/Ofz6jBSLQ+ap4wBMR2WWb4rE6PSwtxplGu
ElDiTDfh28ice3ME2vkC8+PM/M/ZTtD8ed+r3Bh5QwKNoFK5vho0BcKl1yg0ep6h
i9e3Ftxusd07pBzhk3qUQkMnCukeOxVFg1pi//+1UPKqx/z6JR2A8W5sh7nBLplr
NtQBwbjj48oady/p9CwSOEhKI5GLQmBmaloBhuEFp7g/YbE+a6ZTeUuK0SUGMT6V
jNfNtmN6PxVjhbzOPK8rApzMMsrpTXNGrSqnH+Dqc1wP58AeInos4VCKpEDkz76Z
Yy0TJo7dCH/GCi4zhecUc7L34l1CGaROgUoHC4slqY/U+1C8ir1utRncs+ktmDLN
5ykBVz/jIhuh/6tliTicy7JZPvcQqftgdKqTsX3OOMO5iSBuBftdpGBj9+SQXBg8
a58nCcwbpd5wjXozYupghXvoT1z7QxfSL7clBkqxFBUalzfyXdfjCdTrAcu0XxqQ
flUp50UzyOa6HuiZzM5z0Iion8XARdhzLqyWT3Ov0brlVijJZ813akN5+y6bpYun
WJOfAXQzJTJ2cn9iS1f9toROQF6O/pXGQTlp094Rx0nfutACKcvLd7aiVuKEBU4C
ozAmwWDnaKzFT85bT5StQbXl/hBFuiqZabGFQpYXqWXE/IeGjklnSO5MLgWVpD8v
naIhm/kGjJGVMWloV3Sb9T5MDf5bNysf68WF+uxdujmEgXRyjMCJeGmDzuNFRG7N
CTJDNFSK4S4Dc4Ldy3YBHHr+BPyihTzDhsOwgQReOcy76e0mO4YjJSxGxUZgbgTC
gc8o2e0YV2FYvCwz2ikretju6T6NKE1+lJ6VSNK3XJ6A6iwMbNfwgFOrY5OUJsAr
DUU3uGno8E4Mjw0ya5a3edgvzlFixLRyLo+cifUvqmzInESffZckfvpBYjiI4F8w
KDeHh3q/9Q/Dn0FjvlLjOrtbOPSLqAIbY3ly8UkiCGTRK9+pUuaXksz+KuA5vKsp
gqvWNeSfhUi0s+rLakAf6HVbLp1fLem7JtFRQT69QgvUJ1yfJ7DtqhCDBN99J+3w
aq1cltDQ5ISVg7ZK2/RbDfEG2ioOJs2Q6niEtlty0NHN3yCRyLE0B9r7xT9OPXAN
qKKL9YjayRbzf6DgmILprMosGuDjOGkLf3xSf0Gg6DmeTe5GkPRVGrLQHiNEZPCd
GEwW85KCqSa/fqcGc4ptCXi+GJUjehEW1qwKkXmQsgk4XU0Q+AmXtfhQJhIlcTi7
dOgNIwK2ErB8zRSexUTXVcWiTwa0nxbaj9yBJ6BqciQsWMwClglZFCJSDzQPqHhu
pWt/X08nBMc/Yo+HGqIPikpS42Q3FawaTKWV2D2UMYZLkqfBRdG+4Td7vt6xLia1
fFUsycxEqyMa5I0kDWopLotzuDgPziF3086TJkXE/1anPXaQIBDkMghFI0Sq8TpL
HMJuq8EQkBah7w0q5mG15ATPK31DXlCVSZ3ZFkvk22Opex4QQ4ehtOvZSs7AqXoN
k5YIRlIBoUB1l8X9aqoVO6eDvth3euUDZDxlGIjOwAKmgBotQ03Gsi4XcB3gVCBw
l+/q2byKoFq3ffJKRAmnECE84cb8FqXKXL/htpKa+T2c+mPSFex+rIDsxm7dPfWD
FI4Ly2t2d6U0V4aQmcD391+mDJqGZrlYSNjwKy9KEJR1thIYh/kmLuJGd8u2ecF8
bpoGI+MdRbAk3m2NVfm3bCxS6mThiE2MAxZHTobOpJWUfebr+AV5HF4fk7HBvtkG
S51/I9MBeMlUywY6bUNFzvOAgeJJQTpDggfMGSoeyIH8/ptndIxTRMhFim4klhPV
lz/2GL81RusGG16fpV9OC6btC1Hnn9mjw9ZmChXsVc5UtCo/0lWsJ3eNaPPLmlhi
Vg2CqpExaZgCF9KL4A7gCFtaAwONHMmfbgZzTiffCJp5mIv9+8NngHR2VQbc2MLE
Q/bDGeTTldp14Sft5AvQHNdznLkPzyq1Lv6MKMVX9AE3X0xf0lsXlUzTco2QMMHQ
6u13BYHR9olR30z58WMlXGzzYkk18JhLYkzBY7mnfwqOGPpjNGIygPJINubiWdkE
MNUrpYjv3nSswObMRbqeQnbCbV39RQhigjN/+gMGOXEvCS00EXNRwI6k2+CzcEu7
g0rFfPJZ0cEJtxMX5SwnbrSwft2T6pLbTu1XEQJfpnOaggOSySIxaYf+sjnXRTDV
rbmlwItBmO7O6mJBlqCiR4EPvtHGq2T7/3+KxGmU6Y5vICrTtatVhEqKO3hukRmB
WsfbEkOKYvSmH8exCjMw97uEm+z/sfPuxWBcU3QtupPtnwE8s+hQmcCH/Ti+DUl3
SS9sYoXQFV4HLYSm+h0sc4f/zbXQ5sudShLPto6OuonVbbhXr/cE67lNBTVZREXr
vDE5nDe3S34PExmQdzu6OTPnlio8KdOW/fHrZ9/L0j+uBhq02X150omDGkmXYfrg
ZExMx0U3abkTCWCc0/8Ceea+kyvEyV5PAo4rldJMDSNQKXt08w9k42DRgGHqT4Qb
xbD1X5hqMq7mBjvnHLr9taMNznflEvwaQVa+DyGFXGIuQStORZdIWJoH6NXLA1in
T4UuDqZW02CJCG03hL3FOH6YoylUQhjxCKpNZG0AJKZsFeOqW2ZDvj3CJ3uRyyqu
777W96AeGeL5NQg6fufrCSzcawwEEvQUqTnVei0VNsagzpC1i5yES9/opSGlQo0e
dSyTggzhfEO6A1rlKog2SvnPXSE+KYRrJwJR6gMotXeGW/Bl3SASnefMvfoMNl+S
KWo7vfy6oEcnUPAAbQ3ZfN1NO9ckFmKLLOnzmk/0ZFoVMwIDQsD3OV4bqMV0lyFC
8d0RyBoPksJGSW1Cnleq2kHXydnpsuvY872AhbfOlgXNnT0QgZGlesR3COfbd62z
s1/K6eJEj6sh/AAMUb6p1QNxhkGBdm2c9saC3r1fKfYsd4mEXnWebyIb3EBxjr6O
B+NHkhALF7ZjgdGaSm915UPFReupSifoc9yAl0uxMbYziNwhHLfh+6m8oLQy/5bK
y7OkW6uQFA7Uq4nh/I8/VeEubSjeg0ev7Pvdmv37jyYqtzpCB2sONlmmh4s0D1cw
6aZAmDxCRJGKIhVL6Rza6zEi8J51t6otHugE21azfK4GEXr7kmirPxmgVkG6SYmA
0ns9rokiVHceI068DjyqdQuBfU5KCQTvXzH/9oSH+H16MQxxzzr9J8e7oM+idqf7
XJnolcPL5ZDjtFWsKFTNYDEFq8ZygholcUbcywCFGZF6/tiIJIhtOCsgZo6ExGJb
bshIonjjV9PFA8sNYBni8Cq8ZgpC8yClutkbDWSBKjFA47zP+tTfTHfJTXzmwcGQ
hUu+tzgmrRv4UCnbNLOiPsp7Y3CK+rW7BERIiYkjfqG1lQiqZjtZR4ERykkPZli7
ZYgZgfHCaA27POzwzLj8wXpy3smlWPRims3dbND1kTSpIyoQQNbYxv4B9fNC8S2Z
tXW7v5UzsNnIIHkrKNCq3JTaZWhB8KSYQKbed7Bwga1LluhXVnggTgS7Ghnf8P2M
aoolOmE7/L/NvDySgsyZIcaQLjTE97J4qJt0mNItzwycH+59tvWpBYkhlpEc9/tp
zLoMvzcy8Xss/YfyF82jMV9Ebl/HoAGihgGPPax3CY6NPsnFo2xv7VZQlUYxf9HC
VusHEa7TjvSa5vUZ7jn+Wat+XnoJSoAHLElBXCOcIrR4A/x9/Cyn5UuKz1M9sq9Q
zPE2RQ7RN7OB6YLOmvu1WoYvbhfs7S8X0KtbsdWPEfuJOuhIbz0ppZbtgViNf3vE
EERwx/1Tj/ZUQOCar93B9mlIhijbfPWiYFxOzdTCdMtOZDaCVzrsKQGugZOTc69Y
BVh+srTFf4O1+UarMOVVeTC0SEMte03/i3+D1UK+2Ln9tVgWChJF5mKc9gm5R3sl
WgOod5ngpkEAkeLwxZv+PJUNgIHLhtJ6Ctvodltfdosw/wY7D4uZBH3ur6Eld3wc
4UFGpvhiFtlM8pfShn1mXV4HqXsJT9ayxbBfhC9o/TlFPtjufLFfQNFC6n6krjGS
GffChZUhGlQM9gFUhUYIvALro0jJbkmfJpPi4N3QHi80hi0WTNYqCvGuDDAliawd
2I2kF9aBoKWWE4mFywu2NTGwxAZkGwb9VT+WfFDSvvktUX1fu2CEsQMbtUsnyXXN
pINgIGaimyuEIh37KSdkqclWSB15vgNtrnB/asFMomV/OmE8RRv+89JLHA2SXwFC
WAWcLvCVetkQqcyM3p0vZfqkTxKs1HIc5e1rl8W+JyZKv9QyTKxk9dtCwL20+y/K
EDjo3VT74dv+iLYaILi+vwed6KZD1PYoFq306nefApVxNTYtsYFTGOusPuLNTIsd
XJ3bdISZhCXb9f4LOsrfPPXjOGTKA70xl9ZVZ+fWM7+LPqvuJy35TYpyTvOj35zw
np2dm3z4SewlPhI6OJv6cUk+dFeqGgM4lXnt2yl4U7fpkpLbAQL7DVc5KJbtZ/aY
GBelIVloFrsGhf9LdGeHRLttQ6EMin5SNHxFqnqhHFaIV6NhA+8eZRPW0hHiU4ZE
n3fKKRuqld56pobrVEYZUNZxrIXBA9BFy+wnvfmXlG8qnxcxbNB5HSTWNJc+nJaT
qjBdzcA83KlRf9VQwhQYxXLzy7brVhkdDVvLEmrygzL44oLVq1///c8P+kLFmsib
piFATMIrg5KsbSFQpLBtZItrRTR2QMF/tFS+lKgJ1v7fobSLxJijwePw4etIQc2h
A1HdhMpVfz/SPbw6UP8HE72/2oTlHIZV0VfFVscS73mlCnwMrqFgPkVTGAtHqtiU
Zuo9G6sdFQGSFNZYlBTWNB5DEOUN46yhoHtLbbbTGo0qnXiWhlkZDClRneM0Xgla
q3cUcfGtPdmbmf8VTJmGnrJ9uZSERJLxoh9ObPdsHdE4wlh8nC/urdknYOStjezE
mdvb1iEk8WOGzwBqncG0Se+gGHT1LZYmlvX1c2FYXsULIcjtHEH1RJ/wnBuZ7Y9C
e+0qpxK1R0avbbqSzkXlx0s+Z/l7iHWk05y3x94pH3Sgi+4rT7++rks+lrGXftnk
2nLPGoQTugParJeHUM6gIYLx6spUwPI6ccSLi2dvHZwDl5jZcJVIZsD5X2qEtFq3
N7zQVbqcRWw81BIvQ1iN/7mfr3AXM+04Fhjt2/zEQ3wQPXsc6tYmM7G4OE1Twsgt
EoCsO/AtbD8Nh6yVqDQFJR3qGK/zotYJZqbHMOvNtosODIbrQn8u+ss2nUPPjYHK
MZLB7tEFf1zba/+Ve9O3YYADV3s28tdul9terkZsYTNJ6wGCFfW6Sphzhbrqjob5
bRAZezJkA9UyLVTA+AAHmvvJppnJzHMmk3Rt+IsOcQf/r/dVAe6DzAjC75HWhBX+
TM+0dic6omvA+R7sbFhJ/rx5pZf/j1kl+o+xbPeuk9rpq2rN650x9PlHxCDnf+b6
DZOUUHv6TsUgHktSot2/Yc9vpRbDzN1mKFFmxsTJX0JufUxCObUTN82qPA/5Ozlv
/AAdJy06KHZyfhUq+ZLAmwPkx+iMpEbfuM7vHVJLwFfD5+RcNGzsF3AH1LDBD5cq
lh1WZK5WRwTSqkWPzbbcV69fIy7FZPRElBO8LDr+zBNOhfrLGhTm+gWX+ySmJ5XB
ZElFn9CLJUsPYJrPRayijSs5mAtbfAzxrNGi/BfHdSUt1Yy8ZtRMGEM8ndMdKLU1
Pw8VIiVE132Xs6AUNoZbj/5aPMU8hG91HNXVavyZgyWhmYb7ecV3gg6FGSmcrI0o
ghNb4kiSS079+A5+XoysfrILAnoowx5XG1zpcTVkKWAb//HZIPzKAxL3+5GcFhA4
/WbClDo2mHKTdbj1Uo8/Ye3sTyM6enLDxGYhE3aiVMtHvQtbhCYVTLDE6Gc9y1Dg
h8RcMUPNhXB/44xeir07SH2J/n0yRa3faYLRq7O07QUSDxAVEVFkzO3WTziYRcNd
MJUQur6LVnyXXrsB1vqFtBY+hEZMwgaw/hmz41SYt2hM9dsI6CmVYm0b5w6c9CoA
x1WfoQdIytg2hGl5xq6p+YxrE8WBcHuDeKN4DuYjCjef097Ls79B2YNN0hH1WB4g
0vDwWe05IR9IVfmgI43arLtuW6TrXiKvPIcOb/oII3bJ4XTOyP+oJfmtdXjde3+h
gaJLgFBWiKeeHJOx1uNClilESwqMI/KPfG7RaE5PHjZw2x30yJfUoTaY/dMPh70U
TdoVLZPoQHiJ+K3B6dOoB6+1L/XL41+b0EJLJ7IPU23p0ZtKD7aJat2llLVS/qWK
vbnaVe4BJhbUzd8+Ixm4IA5HEBmyNxuHD9ofYldpN9Xa/Jf2Z1BayIyGC3MTMJ0f
6ATp5uTV/jIOuqW8Ye8h9e995oSMAdvU9rKZu+F9ZxQmD0jwr5rmvl6Df1B7erWd
nGzJ2AcFrdBw2m4oUGRwe1WypmDOreLWKSJ54L3fL2kkMoGcdfGDoohUdLS+1wZW
c8hLIAyTnb4QBnAhCLZjI1Kw1OrzLWJIMQnGOWr2QhfeeAhJDnx0klqhiOw4MMeQ
A1ey9QZjPDZcIsQFAc93zlwkENwgh36Zp7q2tYFOfJV2vhbIh0hVZkoWJuSf0+oN
OSJK9lkjW3cKAN2D2KsqA4zwjKRRw4Lm7JM52UuAcNOHgUuVbnMV2XF3Rf5lEm0W
SnUoVDOVpyZ5eMCbrD2PoNCrofMHO+Ki0HQopKAbnI33wW8Aol7digh8KPLNg6Ud
Qql8pzcDHl3eN+JsJb38iZs2jZnMbVCYxB17Whj07CQWluSBM/+nwP+ooBvGRs19
iB2VlUV7X37jed7yiNU/GyEwp7QuDdU4VUm3qbd2bReDgg7Y2ootyuDnTkOeeygJ
N4fg7caZi4sYE7ZexPrkK0zdruZ7ajQnhHdHmL2GXYXHvwg9h8QmpQk4we4gZ5mp
g6DFw1bkR/YeHhFgdqMiHd/Q4Gdo2XFNxBOfcDa3C2+VX2PTBJnNrJyUesJvetOK
dwynfPD2VPfgiTvTw/XHr2K7v1T4b/fc0Y6STRkz9Ej1I+vHKQBG9k/G2Fzl/QJ8
XAPimOJmeBUufG3WEJRONdEFekmkRpqY7yiTYY3m/B9XFADeqLoqjfsmq0KVKAJ8
9aCFJ3Ay7je0/wCkA6l4NaoJ3jGxHeJQe9eL+STWehdnUdHldr/M9b7FwFyBMmR6
SswU4+pnJ3tVppjX05nNeJazzlLZogiY1q8x3pD9Td5/yDTqoiLeskOl0uHNDiqJ
AjFRp885gyoFe7arTDQR+KTbvwc64DRVJovKsg9XF9HgQ77bEgirhym3KYe+HjiC
X+ywIy/OH+YyXJNz0V/YBCXZeKn7EZGlzhD5vkTAz7mgU0PI17khVvrYOP3GhRhF
rYA0I0YywKrNMxHTgbKuE9uQyYn7+4Q/qODdrr9g332VvLrouSj/5XHPtAf8vyfn
gqh+UccCBVaROs4xe+b6McaQOJKhPazuKmo4fHBG3C6+E+H6GdDBaNGXaK1tC9wP
5F5I82gfvDcuMOQZtvCtC+uc3Dj1K+4Y158qqBLpQwvy+G+2TymWIwlS4XssEESS
V0nFL0pa/X0z2H7RZMrkPIx4lcl6zptiScMJg7LNPljaKqNyR7W6JA0qbl4oH+FX
4mEWNrAhI24+fDSS1RELWWQBhZgc6UrXUL1ILgEripKdv32K9TzzoT2XW+Q9mN4J
IxnB8T5iRk6wsUkoIXm/Z9iGWhYiRsufhHGWGdg4YRD08ps61pEwuRAnltugpPQo
wKfaSIOCviSP8GC88CF3wFRRivse/cSoVvqRkO7aazMJed652PWM5+9tLLmOtWRM
rmvDUFaun8AI9YjK+AS0aSCOowCHAmtTNxFIkb879ibdJHpWQJTvgXmN6GtvWTDz
FfzfmZ1nHbG3omd6OMK/tirWAEbI6d9MQBCqkS2ujsMnQxMGd9IzvgRU9LpZBM8+
9lf/yPqBHFD+zHUzavpXS/N8oqC5B3gISVsdBG3hX9NYmZ6E8QOy65TTDdgFYVHY
qjz5yEtcytkOoZCdV2iYnBra+/FRUWUUs+ik54AuZWPNzgYQlenrn+gGg3O7Mr9y
4RAqUff0jFiI6kCLegbjE7cHQbG6Rqejg/vVVgc5xmSUYBHFob8REvEHfXDeNuoS
88qorJpFy4ZFx+TTq2UDKE2ZzipAfAQpO6KplpZug2o6xpYLVJYTNrWdLmidZfQC
/9O6GsgnPbOSs5qExmnvhsEinJ+gKIYu0ePZaxiztrZVf7mOeCslln2MI3Q56svB
NxSbnIovsRqpm/pHredV0tVSofDHlX2owULDKLrfnIbjHtxXfgdMS7ib4gTB1H9s
1tnNsngB/W5AybLNDvP860MfKSt1KKv1+C9jZiGFRAD1VmkAOr3SbMxqXaMnZdl0
JRq1FuAXv6BDLXuBDC5WBkLTk6YuPZdlAYBKXaeEOw3mnj1rBor02D3S/+/KGxrT
1pIMHuTzkDvOC0PUD0JCKC7uKprpBoaAzkmHDuCxbNTiToDCv7qmrTa9OW4aWKck
e7Gko6Mpe7Dt7WdzdgfZ/rBGYCWTOjpKrpyWkbqlJhuksC0RRhbl1c28+Clh5+sx
12DCI4hQoJ7ReFCzAhjnNIhi8cBRJl98FOXdNx+cGttbBImBix9CeF256MRw9npY
gELsEwvOAPUBbVWEPfljWvftLqAgw1LoFgWmF3PRI5Lkwdi4tFbxUZpLJQVBzG8g
BVeopn1btV0gtNVxI6uNSxOzDJw1rYF2T7Cb2pW7Yq3+T24tvbe1N3SwNmRcgJJS
1t9aSdIn6r2sM83nkg1JVGvv9g5H2SqcMTkklF2sP5lECIjWBV0GJTStGLjxEJfC
8BL3WiQMQytPJE/6ngC3ausF8df/RFQRH/VUfibiQGTClpCQ5aoOspqBIhMB1HrV
jf8i5VdYKdipwTaYqNpnxw7nOr46SDDYOPevErDiRBYx+D57ov8mn8p0aB95cjEk
S8bqCJlJPLYWkei68Xe4rGwE7wu/0SfgTsfA98TlaQhZvSXetXvng59kFnlcrzkh
Rutr3js0X88P6q9FfexBzE46a0esBOuqKOR8Bhl5d05IgZPmvtmYwHgd1dpW0B9L
9b+Wuyh132IqNrTWO5+x/KxMaSowtmBpl5yUGY1A02xP2YhZ/AwXbU7OdyG9073h
KPL9ui0vHRMGXFpBmIultBQFwyelQ+SbhJOArjehfucWa57Dp1RI8ej/X4RC3lmO
RJpKw/Zc13URnU+ZiM7YefbuziFN8rr1oHgb/AnlKIez1u2BbKyAytbiuYwrfX5y
oz9o9jr9XSJGogljDD69wZnLM8g5wd+oXmDGFH56qCbjLyuRRd42ZL+fU5uRjYns
LTZzqZWL1OtXd+GmUXKJDBXZbSTlSeW/GBBj1Ymgd/nMG/IOlyvxi6UHK2QL1tTB
SVsjcVyEpjHx0r8m4Nnrw5oHjWV5lCAh5lhwQa1hcDNpcLybKyDPKGX1YiGOnJ2e
thE2K5kVm+C1i2bvpr9w0JVnCr5grE5lUUNo5RVPmygNAf7lTBdk7Y/CsrjCaktQ
LrWYjWzTpuV8UgqQ+GMfdbQK65O/l95Tn89VJ84tW5E4pSlKjp1SZfhhOszEGtgF
vwyhC/NyaB/5lDYyJYteRNkLl6YHA2NHf1mE8eJ0bsRkk/Bw9mKvjD2xbqyW6l5w
BcP7n3YRgtAAtDlf233VphoiwfnoIo+f2BNGXvkzYHZ9c1IJsQBR6Pp8UTSWxDNc
JepjPBcZWlC26y5bvhciG2ASqXvjQeuq/uocy/cQ2RIGTX2vto3tNjUEuBHuJZ8a
mkIvtQmANY1z3n93KiaiRJpL9CX1vDztSjhnyelDmoob1GqwTmsazVklXmBhD5XT
YG01EXXV5G8NdrheqKt2PJkFpEXC4xJojP6JgMpoP7ZlGKR7ZdcvY40ozWGzGpXS
aoN8PT7D+lEW7dOKxHl9FOh4jz1bY3nkqgnzhEO/yNvgEd+q8iFJWt63Z7oG1sNu
ph9tMuoGsuyEJsV72y5dg9ltDOLQAVA7TOaC9xLiF6pacuLOg7XADA1/UTeOK/TT
kYHpt3yPHpLoSu5hAloZy7W64xXf27tnrQAEZIFPQSSXkDCVOKQwuW+NK/s3nZog
KzMe0uf5RVM6uvN8vmjw0LW25Y2CqTFEUdWXIl1yydDka0tHHjn7cFPKlSvPaseL
htDj7gWeLJjw2rSduQ2igJyL5pjvyq38S2vtGsTcJ/al9RRpUCxNOXAhLeSl+7NE
BzK71113w0i8WwTsSUhVDR4ZD4Hu/l7YZH/xbu1R8c1BbvW6/v77oUIajjhbq8Kb
t7daRas197jeOe7O2bEWhiltphbI+P1zhGgoDECpELlc2w21Gxxl4G0mJySpaoS8
Id76EHjNeM068urQy1bGQFIew8zjH27w4Kq8ZUZy7o6aBhEQyflRavfLzCx5bTla
8CnHdydYbb1GB0YXuJET+Ii5cNI/Ov5GfsK4lFZTXx3yW5WRmlu1iNGwRxUBcWha
2dQK6hGDEmehfDnLw1Yuv5j+09tbURBgkZ35j3tGQpJSia3wKc97Cb7/EK+tN5Jw
NhtJJKvod08fGVQAk8hFozGp+ZXmUimsm6geU8Mt1xxzOgl5GBCnNvp3oUcdHVzh
CKFEHxtFsn2n2su8QGQJVt3kLU/ctP46qu4xkHa2/YBY5lm2vZ4ySGR3KZWGSpj7
CRx8oFWo79JhUwZuR/EyDf12UyTqLR4mXG2QGEO9mWSyqoi9zk3GPbV5MZ83C8V7
ZsPR1gobqLqw/eLENYhn4mONjjPrLpnUYdcT/ExrLGNBOfRhOW8yUzZWafZseMQS
YnlZjkFcvtL5iJnagnUF5hPGZvz+7oypk7xADBlEpwj4J0sP68cxo6c4H7tASs7K
KMpiPmV8wUCTE+SCAs4la1DHusIEWGg/mKJYjuLfK7PsvVz0p2W0nfv/kyxwK2xr
wXCFs4YItOmEuxQNchKsuZh6ERs/7ihZEre4IUmF9ZrkLVevydUXtZQJJKEOiewy
1/iBNb72tHykKNDI1KZgIJ/a/EW90vzuM68Jtnq8o62BsIeIDtnKdRpGq2iznTbY
R2FMTqU4+c1xDRhraIGqQSdQOa1KmsuH6rtZzGEOctaeDEPPqgd4cnrYk8sH1RIN
F8MaxIHPXmVNeWiRtHgU++m3HKw5U8NIU++8CGyo/OnFXd3a3pWcclh7eLBZZRHa
o2zYsc2ml0oPPJ8KoWCuVTZRvUtgEs74qs2dE9SYL5vpde+gtgPGL7b0K3E8mR6S
hY7URkwt8/HEQ5F19I+kwTCjfVFpYDvw39H2GPJPAVKeQLW83B9gesc6uSw1n6nB
/Ph+vH9ULEAWXLOku+97wzh1LJVA8RCvPkbTrHXTfsrqm8moI9FY3NMLWgbAlbgg
dalatNsu8klg0xqdPclR0HCUG/8mv9ryODGTHZ44zaITM+kXPhaqJozy0jdS1fZF
wkegg0tmwO4cctx4CKK8ZzOgw+2r1ALeVKQhcU6g6f9HwEZfsKDgys3QcyytSwPG
MYm2IiotK6n7kU5R2qeSahq8zwJCsQRyBSbFgahn3UafyutUOtvj2MgOuDrrQpTs
j+koexBupTquN0WAxnGTC7fDm0z8rh+F3cqYTmDayJK8YYt5ERWKoe8QBCFyb9od
zikfBmdkMB8a2fRk+C4SfXeWwTy2Wt5NCZh30oqXEk4dgSEyrqaIfF7Mk+dYzuRL
gxOrayFTfefguNeKQt+VmTFg3LBGJ39j3yNGx8IUifWtRzQtfijTKquLYfstnU6X
BYR/tB4MdsBtG10Exuc8PWVX9zckQD7k0P8tY+hyVPIHa3OYEpPHEL7K2cByepIp
N9Y4JH9+VXsRCdopHmSyMm2NQdOteEKTgOmdgpzlbPDkqoqzlpj6O2pV8pjnKQU3
esEyZ1M/wOcBM2By0AIwJvN5lq1LIclA0HjO5m8UKo7pHv8tQFIL9LvQ0Svu/qaB
XXV24aq6KQpf92vHDs3wrV4cxtBlJHu7glK4Ck/S9MEHS7M4ENBOC/ilnLfQFLia
QmhI6o1KNQX6J8M5G3SrwL8qkYdqx89AhpG0/Wn0b3Cbg2JI4ixjH4mJmu5Kvj+G
QQLoszUSjBH3beltUoxbgeo1/DCQXFvjSMWyO0JS9Q3arVd6yGMFjSHkkuoqd0HT
TX2k2KcER2DReFP6410POwho8rU++GhkhhaHL+e3/rWzC/tIum1eGbJhoZyRF+fZ
3NWfMtXDiTEMMidbRsodVgsvyy15isuCjIMmqz+L4sV+xCgniSRdA+uI61b4Fi5B
cjDCGqU+rr+P3s/b0Q2n+1ciuKDsOrfD4ksygivmfu5tLh2HpHAydruP9aKaN6Hc
QO4KBs2dB2a+ZMGJPGGCV6wKHOl2dzz3YHn3ZUEAJ6v6wxG0CKw6CSGIj66M8uCh
BACycwW5UopBK3fuWryF9BC78jKIlUeLwwV19WBPCgkbr8Ur6u2MAlKBPb1TfV79
dqPJ47UTB0w2af50LqetdgccbP2J2EaBEAtf2z9sYgCiBS5LkTqk9p2rKq/oFnx4
glzew5S+OHvM9gslMhxPzXQiBj5yNvbnt5xGFdZpgDEGut+lut/qgciNCKC7DhVK
E3JBk8DT49XSI6e63oRSRC4Dn48q+ryCB2HkuKzegov/EiWxInHUYMzmMuk793X8
fYKEAEAQRsBXnARzQi6Zw1TtKq4MxpRSyPBgWtBm5+UXEAiZkZ+Iw85cdbIaBzm4
twXF1R4NxfTFTxCzR+BdkhJZd61S2TjYI/tmbhRnBOPLYObGildf14Gq/TLsNpZj
cnD9Q23XskQKooWSE6rxaFygXWXDxr4MbzGrBO8tANVuZcM4cQZpOCp2iwhzxR5t
dBeupWMQ0o4BiEdQpVyTqpCImIveopCMmqzAlcgmFQEn90mJfR4w7+d7KCnKqpmV
/MF/O6cB/j/zkX9YIfcgN6VtkxBsLUJkwQG4gsEfvw4FZV+trIwdw1aBltqFsncg
/QSdERsBllVAeTCqqg+CkqWx5uLnnw7/+HS0TxNDAcVEXk4LINIfX2o93/RPgEPi
CUHF98olbDeOxMS+fwOCeyCYkN5nsfbl7pREKcR2D7FIaa2BVTGjJeVi7b6ThZDe
89Rqo5wQ0TDH/UF6Fi2MojdILNXijqChvLxn1Q8MWgRe+T4I9ji3+O5demI55S3E
Egfz7nWkSKTCycgdFRpb+8/MFn5EIku++sgl0BMfexVphyUNDLDzg0jrVmTEMTG3
NiqbbeGRLOcUhT7JkqZH8qKAlwjuAWE4Isaoal/c3lHMqfJP+g0KDm3rj8crhdJD
DNweDcUGKXCmCSlYFaCg0rt/aWPK+FG3n1fM8G0ww0+BIpSV/08G+cXcW9tnlqmZ
WxDWySjhk/pjHr5LEd4Vl5B+V8syAt3bVFHjOrnxz7uCLHEd8FMAX1EtcwKcu2af
QEMwsGQGBS+9JbiGk268keiaKN5Mi36TjUKA6zzTPOdQeb3CFt06pr8PfmAR+ptM
K/obBqbmPGrXv6VYs+H8mxQ3f0IoHSKTsCGIk8n8t7WPf1zOi5grxsvFDiDw2nzs
ltLt+R21DYpQ90rxk2/WTKRb70Ao+x3DjnDGaWO2OyWulLf/c1l8e6yTklttxknC
RZu9clv0+iJWcvDZTqXquMmb16VghX1UWW/DXlPJPfnvhxstiodUINzwnzTCqlKC
g3Ja0TRgemoR1SDtKULGxmqGhH6uhjgo1IAuk/gNIzfgNb5GL+J+o+zQY0UDoTcC
pCr+YZxfV0iC09j3gc5zPSfJjSbgBiAxrRCrSOrVkkfmDTkEdV9+PaXBHejQtpzW
hLyEGygixQhTqz024ucsgvYVcPHwdKuJ69203Scp8/voDEIQ+WttRHij1ab/VALx
YarXuxKei9z1J3MTlUWrJrKBQSD8ZavMTbYJRzMqbyEnBsV8pbeY25al6MPU2XLA
9AWoiythrxk6PTTTwlbrLIirUQ4Pao2imAUD7wTS5XQnFcKnfH8MKSd/WWkoNp/c
yAdBi4E1BwhLwKcWbxLQXMWBw+39R2BhGLJevmicpctSWCIceTedoUg2KX3hmMOZ
ZwRHWZ31VvPqmvz/A+jr55PXBg1LWNVMMySz45N8COeURHCKDfamjVgOQJRWvPsK
+0lx6UkMJBTbq0rLuBnjKwac3LBHIHj/th1DoXh3ZmOHkQuaOvEgkH/LxIaFS62q
ki6+xQ0p61Twjf8HzMkQ+q+nlwukcZ5Q4FkNo5WO0DO6aJ/p9ARanC+G8iNU9iii
HtlqqLO7k9tWpQ78Ka2fhh9FIQQW1YblrSQuRpY1cAEp1QehusPiGsuSyRYG6f/l
FAhF8nq8kCRGkfBBvna3CpJq8/lbrw6tO+JeVlfwJIrer/J+7sxKySP77N05xPF4
R1NLBEnAxhzkevgvlV4BZ5LWl9SHZu7/0xyR91FLuvm+WsPY6O/ynOq4152mQOJG
xoJNyFuORuAQAjzm0tDdYqrY3icXYwXLrg/CtGJ72YrhZeSIgtQAIzB9yKINC5jB
1BWNwlw4S0LhYhiGhj8y1cp5kccoQ7Wn3lwXJ7H2ewkeDnlZxsMd8imXECKUvRc1
UcpFuhV7fajgrAheV5IGDa3+W1ynk9AqBhwevOoVtsmWhr9J3vQUPpq3EI0deukw
LXavQAILSxt0LyXUqV0MRhKjqZn14Lb1yArdQ+De38FXI1/E13e6ufpkib1sxZ0t
mwMUcjAQXWzVKjoLxb/fzdMyFqmmoJHaPfYgq29ITNdIKZqudaPQf3MSzGeO7aG0
7KM2U80k0c1dOnzZsPPZ7sEzbHfmAABaUyqqbYwCBsY+vhOTS6RltHqMNgw9aPKY
oDhX87zsofcRN8eDc2UB/D2ODMIERxKzWA7fQoaY6O2gh8qrDsLeF9BSzsu3fphE
d8fRHO7csJ4LkU+1doBup6M4vyvZYXomiq9OEtLVDvEQZU59QNTdDqLkE838lXP6
aEwESi+sDTVfNXXSxxr/3+ltvUtgJ66CEmnSSuZyzP9CNu0eBJ7qesovd9k+lDw2
Rkxlw0yQyYrmdXuQkjY0rouKdLFyYiWxoWEwLVrndOyam0HSuLhwh71MsqLL/D3H
LGznb6NRMffcdxYFFtACwWqEvrs3POwJoYZiOjLKKMdDOW++GT18ArNZubLI5fT2
x2+XDBxNe7cM0CMcvSWqywXSE7pcKmuhXWRJRX64wQ6AIYjt1kzAEzBuuAKM4rz0
U+5iOGekylLCn2kL7E+GUTIjxL18G2JgIWNU18vhA/R+cCQDtGX8bdz/QZYyNtXN
FCDNEoXoZFM6oFj2MS2zY4t44O7lKLGCnkAEOo7U/OcSE9DxSPllFQSuQj02cK80
oisXbJUSW8p193RBAln6tsaFgTUcZoj7oXBMtKRuuIyp8nn+KmN4UxVb9tCprHyw
QMdeHCLs5pyco0812De9gQ3RYHwe/aTAZz1l7iUFxQjkHqa3TlWRH5lctUDnrq6D
+EE9tB52byYcT4GOTX3ygzz+09fzh+WOnPW4NOvHTcCbBDReGI4qcgq44ipSAMj1
glOY2ZX3Qzy0kcdQOj0BwGE3ahHsqWs+V5f1TEWKkcy2g5BzByFH1fNHg55buIiU
fdMlQSEBDC2JSwnFgKRwzKCKthm/k1ZVPwwG9Q6EYl5set4jF4AydIjRQtl1tx19
q+F9kfBVTzN+/lA3pIZnYlszr4t+9J0pClGse8eHT6PsCTbPMo3I6ZcrQx5QgPZV
TGEPS3/8BvIudmu/1JLajusYH/aEZKG/gNomFh62h0skOsxXv0zli+6yo+ygHagz
7vCJ1pnJItL7pu/Pr/5p2OIpj7pY+h/oDmKvKu3z3FbibqIgFBtCUmoY12K6OzKO
zngSEGeuofj5z6Z+9NFYLX+bdSlx+lAzvmXGQJkRMNyS7XaSjq7cS61fRsaiPuV2
7p4/BKQrkIojyA4r1XiYA26t+S5GdiAX2UhkgMldF7/sn8BkTCBH6QHC3fxlCr8D
3qjt+QDnv2zb5bvEM7y714kVhtT/gdSOtYfXKlPy90eXhh4RUfruuoxqc5WIJobJ
E37KzBIjPaMwDIi8khjQj/iz1BAwHc4SzILZqGMmSfdgUJdgmz3nQ49bwdDzbrJf
DgwKPeRl7kuHOS0iBrxeWZrW3ZQKWeE43NYCqU3j5F9MDOIEl4yBzCO747XN2Ehk
mYQ3DjVtpMNmKxJ7YO7Yt/duAFuETv/BSUcSc/HzAclZqBpjcJHq8pBclKHrm26P
4O6SKGdyS+rFB2QSMuIq2oFQOdv036KWBHdxF/7+QfKKqP1sjapF52De6xBUOsI8
x3RTONfevCaQASAb1Ui9GzrzxkJVKt58QlgR5Re1/21ELRl1GPHJt8phldR1ASHc
xZE2QOHXVhBaRPPfmRERxIXRKjQONlwq+BTx8YcqbXz2jAYigkLhnWtnDeMAYLww
jYQ3nR1/NT4kLNQwlo+0Lv6WZv2xVeltjVBGTrTE80ul2PqDOE3vwgbqKFvX4xGf
dhu4OzZ127lZ9Zd1wr8yC3dxrdG4MuUwplcQWCpKiutVRq8y8JejwVdlwF0aG0tz
kFiOvPC58zKQeUPV6BCndVAM/dCWZOnPK8Qf/JDWmwZpLkIxbQ8XTbs/2QlE415+
BVEJuYj5Mpd4vDQKw2TORcmx0a8gj4RTKCqflyT/bL82kPM5u3hfK9alK6qmqZjx
B3yU6ZPexA5kQ7G5Z/8FztjR/OuHyoR46IfdmPjcrmjqddHzF/Kzvt1VYomo2mFh
h2kp4PSb+ewq0OBO0m5goI/fcxmwqWSe5JDCZsnPmmWqdbGtcRsanOP0aVEEP3fl
rCTHRIDT2lMUUptnYi/h6Sx1YKbliXHwvvTbSD3P/2UJ4xVyCxkuI4YlbxK7zJ0l
3sTFW7fpBjzUZIrZGjhLjFeTTpKYupvb6M8qBIw9Bqf6mahbD9ZDUlL18Ags5t19
yCmeCjW9qw6+bpNrA1Jox+ets+7jWSDlm/XlSUl/q5JGfIfZCBxR/e1GUVhk9Nx4
Kt5oi/WGD3APL8vzNCd1ILSAsnFvGPKUXlNDy8xBwA63+H2LtFoSFnc6xzP0HtXg
EtmDwzcXIY6bNgJco/Sr7NnqUF3c2pdVSzwNmLWZ350E4G0LdlT8Cxkgl1qZKAM6
cphjs9Nu+ajYglh8z+z7eKdEZhev7ftfk3f/yim3Ktg2cjAAnQN3yEVecfsLIxHB
LE+7M6IKv6uNvLIRtDiwrGKkIx5Kvzwty0b7i/qhL/bZH6KGotmrEyyN9QZmyb06
3i8HbyrO6qrLqhAu1BmvmxeY1ej5/CcxlMcMKYGvgpuIdiG6IAcmkZv2Q3yuGY9h
gRGhP2TrlmuC8wwQQvktFMsv1RrNI4pW/wvOk96NSJEoQoFwk1lXPDzboUcTJ2iN
hfcGZcWQvImrq05KvsmcRBxpi+4Q6tTQhzs29nFwMG9A25zBM42/DtREJslG4nmf
DM7t0iYk92pPRjl+aX46uRNRkhDr4UA8Ctq0uXh8dmtTtEjkJp5/fUWAFacLH3j9
MJazSa+SXNHQBMufcYe0YZGxzPoarHg8fRm7AoPi4Vx5KVhMRuAXLejj/pfSaWrL
6hryYsX3ET7GFciPWlhz2AzRBIO88adA/DYx2dfYFVSCCzU/6up8IqQ/pP8UGazh
Twixu2OH9k7tolSS2SMqHGNq+1A0pENgU0WJ1yjXtoZaO7yKfOF30nmCaLvKuNxn
rafDLtPnjx9QhgMVd70LeoSjDD1+AwTTXk7Z22ogEYYQxtmqFtOohluObfkkoCGq
Rz6Ps/OKXA4123UWNBiUAYVT4Qxwrk9kO4x5CKDjfClN/j+YWhYyJtBj71EGuM1R
4tYyEJG6AxeOh9gmTBOkuHCelGxlhlaqb2kbu06kgRttqrkWF0+WO2IVRZ+foAUP
qgBuug61w6RrhR7Rx8DN+R2MOHg3dGBC5lGENFk+JUvRWyKiZuCMPnsIOQbZsSgm
ktEHJBVw1GDWtpFf/ZhjMu+uLamxNKDJKlp1YHsqOTcRuXPUFHOZo/wtb2Rgmt8H
P3FM0wRBqdaSIAYiiM7I0PVdxvyhzUP/4MdTgDkwTgioHiR/zUdLta8PoNs4R/zC
x104A3Ezo++wAkEG6jwzUb3UoAUHnJAnunQLXiSq47wuqu5PGpV1x0+sbmNh2r/z
LZMQ+zT3tPu1MktplLgVlrAG92a1ZmXTWN+oogd5NC7QPXmJBH8F8n2fWHjTOyQu
HBxBhSc08/mKCcAeqqJp7xpSACdP11pyvnPCGswjZp3gcLEUsX5xbjL8xizu4YDo
dtB/rYwyDVGWzBi3UWHcZsOH28hmoLj7f3H84uPcDPmB2C6/R7VAlVYweGrK9nBZ
5Pg26f+lCvziutjAwXzVi0LLBmMgNWQ1m5QxO9cy/LrK9cZqxPDcVFDq/IsTBNwR
X7KjScGDH6caCU7a4JH7K4t3h7R99Nf+Dq+VeRXRFVIsfmsCuY9+3BmpOpHUxEg/
o9Eum5tJXk5+Gc79TbPIkvvOpGb1MVPSSs66THNlf7qmjWJIwurYuxflKlMDl/E3
ICOKJlFn2PW9xUQ2bOJIY6mxF9shEnq40vMuC5EzFgkvyoJ2vQ9IBI055XqhNbmo
jlyxcPTGEyPRFXOonv1TZVoQfAvzhReQ1mxDsuNvkUWra7ogeDeKOYsLlw6IQ1It
CQAlUZ6u8MVjdbtICaD/9fU5hkWUghlEuiV6UWeXLLDTmyRls00LTyrkfcOtzkDw
rhWgeiA9FklQD9E2ZFHrfjEIQya+HN8YjF8AtcGX6tn+tvgXRT2hx16ZR2KwGFn7
J1Xc81c/BwGSa4g1RHS1mjNEw5cF5i0yDIWZ9I5q0QIi3Bqm55t7/Wb8AwmE0/Vt
6bWlZZie9R6WlvemUqEDrTNz4/aaPhiJ7jUKTAj2ZPTZDh5eQU1Adial4HQnIGNi
C6MFoSDhIP6Or5savetMA7LovXwlBjwWgO/+f9GkcGQQVOpdwy6ssFnHDHIDOQkt
6wN1psKF8okrHdvqwakG10nJdBDzZWEbdMGX2sovv84+EQsysl6DFs7ZlOCqkc3c
Y65eFO+LxaA+GHX+OkVs1n7R14Q2/iTK36dRxcsrxtgIUpXlm6MPB4TCXXp3IFWT
+jcbwJShFqj05ixv/j3jLyVrbW34uPCSrUFawTn77RoZL3NZkwXCtDXoqfU27giF
5LGsiSLh3MLud50vtSXCh62x9EthlkFmyaOfQwjciie35RjS34V/nJ/0hQKuRqMB
P6zw3/4G3RgDq8ADmj1x7RIrFxvvFOaPJqNW6YU4KVNKyOmzBoD9EtVsFcZLLhzM
/1xkZdDZO+e0dm72Mi6l+3UfwC/s+IHPeqhbAjIRE4PVe9qNE8KFJ53ZoRj5TOKE
B2D61NEsiCipEk1mCAoM3lr9Nsu3Ush572hR1KD7bjp+M4ZVbcZld3nnnPZb7HS+
PGW/qQeRPaXKdaxaqHR2GGv0BVerrOw/ta0Aim6RnSDe03e01Hih3vOn4qw3iy9X
J1mMXnvVxfqYxrO8ZOa0wULU/i5smoUsziL0fI4oKMtEC7KAaZD/ZxcKLn5eRvVC
3q6IUfizzgjYOM+JQhSdKxrb3kEvVnG51m48b3gMfVMOemjfriH5PtPyvkpOAMni
g7cUg/y3lLkYQ1TMBXfGUcjMyUVbcAzKv3VWhQywCof5moaA2aFBK+FwZBpSODN4
Sx7WJ0IF1nP171ENt6z5Dy8pQdX8dVRm0eZHY/Y3qVLGOW3jhKO9oXMzHRgfwHso
04yLBjncV8eX+ehvFnpy69mp33yyB5JNbwDZm6TeSIH/KVmSxANAdAY55dW8mtxp
e5G16hohV3fF999aEm7tUqh7eo8gWyEPcNUYKUC1NADFX4vNDDJTcpnmZivTVjP4
LBXGzDPh0l4QHgFzY1skShZ5qF1jR4B/PCC3DjyYPYJ4wedIufGEeDJyEcL97W4/
0CrmOd4HZheOSu1lDmmh2reuC3nlKul4dhRcT1yZVcE5hSoljz/yIFqLU7wFU85b
1vE4i+hjICPwx/TFVhrdvB0vV1wAnkcgwtGZwBZkYvioQilBcuMvn68QHh/WAku7
U6WETfJWiQKc/Jvmqg85XFlMVs+Ci9vtwFCTwj01bi/9ntdL+ysdxUuz4Xf+m/I6
DKkVXW5xrCpxzu2xUYtmg6RurVGxn0eF7EFCuS3gQqqbDuOcurmK6oWqJoolWqPE
8pQRpYidJYu4xeCJJkeG6Ox/fhRF0xbJrhnwfKNI/5fzT1pVfj+9/Ft8X15w7Eua
1eUhpf+6mzN4GjV83tWWXefu3q/jfcdmByodaBgv+R1wzdhEqukMxLIHaMzlX2Oy
6Sh1vBPPULaR+PVZxZyJku7xU7d9MNnIfkzljDowzfUteDmYyHHl74sW4P6vPoy/
+vJwLE/LUouqCqsea0D+u5zsbJrrHQ7ZRI6MSLV+xV1eOusHUT47RCB6Dq7IEVgW
BRgFW9DZzCX2FvowV8o0wxGubdfdkXhZmZZDSs5tLe6Rn6QBipvjdd3VUmxjTy/t
YkrI23cH9gMh2HRuS+8aYBEhszsOSLHbOX/2luHI3uBNkQv5KrM9TK1J+i6L8jU0
cj78c5QU5VCssA6yzeufojcvqhao6MYXeqlJ2Ma2X/ttWnQySSJ9XgM7xzuRxFLo
DAtcoazQpMK9Yo+WoTHYkCBo7H8N+GOAITT+VZFYHJedebUpxhMiXa8RjY2wqC2P
fkTJSTG7Ru6bjDG0xf33rEOcwVKAUae9HPzWB6Pv0Zq5vYrTq5nDmQ1JqvjHas7F
N2bchL1VmMJLfTBC6tKbON1CkM8cAJ2Ql78RYoPuaFUrXJPmg2rUg8Q5R22ykAX5
mH/6J02S8lwI+nP3RI12k97B6GwKaf5wFFvBQcf3zZt9CFTteuShzW+2L8c/+Lph
IPzGEXFg/8eOGumWmwEmpL0gyd8Tt6rNMmNx2TWfXPI4NimGu7IX10CVor+Fc/9O
nTGpnXyEN7/6PhzpHI7TVaqkQ0ypWp/vTPFLZfXL7OCvGXGzW64eQ7FPwmyzLklq
OE8XjjVP6pVS+9Wf2A7R+TW/EcvCPMpP9KWw942OVnbFLjDQb3m1DDJXU/2ZODEB
FoFmyQRE6MkorOmHH3KHS1QViqlx5IAZPRXNo6abP30+3RnqJ6LuZ+LHjWW6aY+M
FR9wpxwqY+FYSw3ycE17uf+bVg4j2n/WqDDa4WfxcN+oWeORYgAegin5zQUnPoqQ
8vBq11/7z50YEnasBEe+lpZGoXQUU/6C+WqKsv1qAtdRyzldpR4/Vy5N8enK79Py
H6J8M/ewtd+xk6FF/w9wjLArxyau4B4s9WrKFe3PIJQWH3wzUcmYlF4tSTJfou8P
bh5t9601N+TFPcAqVLmvGVQLfmgia2TVnbrRKQOAv+Kxmb59+83JFgxFw8Ih6gN/
yhCmSIeC7EtwaQIGc1HF652JlypfZ6hikXsMkTz1lUMSkTmRJzbStdnlfzleCcax
pYXPX6j0WCC1SZ90GkaApTNddTEy+CFmCUXAUHv7/cLF7P/i4y2zCx1sG6ZFcr49
6+/9vN2M2imDiXiEjTSLi6uRgyFErBi1cAEpSPvkQ0++5NrWZ482cugarzjXc4Ue
Ut1jGBValuqwSa5lCIsTekbngKcpIlkDpgUjHy4QEauzYw7jofcAThwkdpZFN40q
dyORKX30qJLr9PhLzRoGIJABJqbgm1apMFAJp3kUM3stBr+QoyR5jr3wlEYWfwpR
z6yt5gnwaK6PQnPl8dAH9SdNr/8Cs09rXQyKDtzupMRjoXrEtTX/tYW6Ma9qYUed
piTeUHEsKEE6iS6p5yfbB52xJrsRz3Y0PkIGmn/U8Wy15eLYfDis/7gq7M5d9LTW
vne+Yb9M78wEFAwLCSoH4k1IdyGmG1YmYK2YZpidy0m0jUU2ulhueU0i/14aHnRr
1AXPcr/OA+1OOcUylPR197Z168pTUhuETvx+Y/CNfE1sAEgtHwAPZaVBj1ryR1ze
82+Y2XUzzFvSJXu5p8qUkcGECV0hEa4yoSWpNUzi70QYcEhbGT82+RdOC7i979x9
qtHsqaldaEiM9KseehxiF8jbAP/Ug+9YwtrV+Mb0wR0pGPZQ9lA8Gg/e+1Ohg5Hk
qP5ZaFN2v2Bi41+F2SGpa7Fr/5FwwfbDzKmBlzhucE5PiyOLnX7Glo5R54P2rZs5
plPr2GxExU5rFt/aVpUiYNPSVrkf0mXORRJDi1XTgpC8CDxOeCYni+4WPaIcuv/C
vVzTFzriRWHbeiAUL7v5dHr+W46S6XzjmQA9+wCYu0NdwB7RY6QN+ku2RcdabePI
GolfyL/QLcc61J1K8/BJ0P2oXnU1TbhW5o8r4Q9H4cq2BxrtBp/5tCLcJnlFGkZ0
CpCuAhUmhZVRK19nPFcbFRX4eJk+eIFGIbaAZLXM0QGqjXLtJdS8gyvC+yoq2zct
znzrKgMyQHYxFEZxpj2vaSM/YbUbOLd183pd/RbkBXvC0jq0WtTyzWRZse6f0AQ+
E3H8Buq4CLU7HL/h/QclgSiSczUkmx1o0RZYGHgYFFA79yYE2bBkyoQdubGOv1BM
FVxV+WcjYLJQd5G9YFh+SCTE6AYeYgdYUsQnLfXoWySurOKjzlegpo7A9xQK0oFs
sReeEgqiKQfnAVqdxcvQJro3qv/6uO9PJhTyQ6vraMQbwT2Qw07XOk5hKewkBjR3
VUX+zSLWGYQFWZi+yyc3c5JVFyWmZercQ5tj8an9S15ZhpoK/icekucY6dzT7/VT
A5yLiK0ykNEZQtnbqZo5YK2x+FCTR69gpnsuY3v+GbF5MUgFGm7FyYId5Inz6raa
3tOIk/yeA5b/qtPpxbFovxIJEKRQ7/f5dPsrzKqHbq8DhCoSMukgg4CEQ32alQNr
VB2kU9NR/3m6GeviVDepRwh4VoY3OaF4WnBetLwCBnThGyOUsJ8N+luLZZpl8iXH
WeP2aJEZXTRopxtc4WsCY4oNmGsQo4miY59g09ErAP3x+w5YuvaAxikjkJ2CEzpY
diJb64MPCPOddjVto2Xjev7XIkMSnWB4kOzLor84du8/LOUE1cO8yff1Yb3nSEbD
Suta0ieCTdT3wvBgGv0ePuaXbhhKARht8Q6MwO5CdOIWETPujxMtQnS8Nsfyq7jn
YywhoT+knS4dgsUq2hivwniVEuqlCFuH9uBHwuzBff2PJKkxbygX9aMo5eMnD7D/
/1hciJjeNN+We9efKVSwPWodIwAKmv0Vzd2rlSOQUeu4Qx11ICdGdUeqUpj4A7b2
+GXLu4RL8NF3nmfkQijwSt0kYz8n6zmjzxStXmFYeJ7L/xc2CM/ypxBu5Jdchpus
N5hq4NfE8s27jIxvYc9N2aBAYSIU8em74xtEEg+FZr7FcxjmGDStekFgLqHU5xLX
YxfEnpKaBjxvva0BgteN5Up7Qjaa9qqucVj/xOsBTLgmIHxv9VHDW8w7OvQs5qBm
EmUqlCRREJXU4Ty1blZ8ltFDjtRq4jnv4q8gde1FgPcwE7XR07TQZbo3irue+BXp
M9LYm29tUj5UJFFvtzsD84R932nkBDcos+NefF3f5T8mnAg97YnNk4I8aXBt+jiJ
X0PS3G6YyH4YuEV42sAtR/fxZe+yQNBdb3viEVN2vT7pe9cUpt7PvrIubR5i8XpU
qpjLn62xiuiJTwpoo4XtVSehavh/mt6fVCzqk7/EtneBcox/HJZOhm+Wgc2s41Yr
COY86dw8Z96poIi8aBaxNb9CqW+OsirSToVDohJUTUv9rN2fcv2EzDftsNfJYjQS
KkgPhf22E8zsVURSfZYFqbucwJlScG8oMfTEURduUvxuODowwxZngoNEtBnCwvM2
LXNime2SqTYhl2Q/oNQxilbm0mBFJZCEzYIZoLrygVuyfasnxEPSjwDJk+OmqsJf
4xuOPCdoU19kk53U2jfxWykbWHWuOki5ufY+edL8EYiJkf4rl35e22Jflic/GJ9t
Xau1HbOhNuzH22WVctbfJ89NFkDhHU5Bl92NSKCQr58xCYCIOf+dNirN7Hvb0Ama
CIx4SMQg+aIx1q/tOsc0qZkcBGEvpRANCvvNoljlapXgShq78qcHwvQ84MrzaMH/
m6wocj0Aijqc9QKoY2XPL3FjKhyMXZwZ6E8nfE5CJgFdwgd3HaSboc2cvdtYr8QK
+VMC1d5zZLpRvowB14TCy0QgeMB/+llaKVZjrLUplYnjyHCuUnPNtmjabohr+vU+
yLfXR4EflhUZFZukA8/cyzp7m+lpJNtbTOupEDS/FrvXns/NPdQ7A/J98X+v8s51
Nt8hr9u9ujKclWIpkRc0wlwOhozz7fQOYNfDb/YgbNtrFYV+NJHZPBckTdXlXGbh
d7XV82IWjqmnZx+WUMY7Sqq+j0v6yMVSncOMiF4xiqJNgD1gVv8w0CDYi6iyNfu7
WFhYiiZiWGD/EWl5124Zywc7fuwyTeFM+glxGGnIxx+9MI9b5N3858ROeMSAPRp0
gufFjrTKSMdc6D0b2xr1f1e4un/4cbwDx5JENF7pYpbTkrKznIVt6Dlq0qYYEA1W
UYHa/l6ovjaf173W/mozkA3INoU9kcAMXfVmM4sxRiKwm4F9imptsEnBiStimha5
0yUB1yyqTU2muD/tZ+IakhRMMoWf1yplRGH87lD/S/y6dZCFqRgozex2/oIe6KDw
uNY38JcpEWDew5FF2Nx+t5+vA0D2LWXNUvmsC4i3MfXIqB7Tiqcp59T5hJM3TNyw
cF6nTxxTzadtT6Zs5u5quivLPkJQIff7EJtfgSP4JB+da1ZEZG4YpG0nRM2asCqB
eSYfNICSL8LRLTwenQ+XehewspsOqp2ydnb4PZx7NbAh4r053HjVG+UbXo9XsQsA
0jUVkIyVPPHurgs+icpVVaKHJtVUDzQMFDmss/RoCBLDLl267oTCSfGxw+K45DEv
1OU0Rqu0hCRwJ3m96cHsQGWUSHAH8DF4JnUhzAmBc/QbvzzTnEPBQmwnuaK0icY1
QNet0/7A6GlolEX7PeR0eoD9wvcSKJgUTaPYq6dZjL2DjTWQY69kz1HJi96gAVIQ
unFh2OFwceH0FbMQlKtK4rv+Ifx3bKaJw7GOytrkpfsaJxjRuotsRv3afA22Nk4c
qcyDk3GGih5KPxK+V8t/S+bld7uODylktJTDZznsSnq43tmIOKhxt+qop+GpgdyR
iMYGUnkmNgfn6BFO/7XCTtJSIxNqQJ8jx/wV3L6Jn2kq1fFPw0WDRYRoMwcpJoY/
qGUvI+bUkMatsz9OmkF7ov18xPtoYFbIzZF/QYT/s4FWMAhboCScA8ywicffkWm+
vIySoE3Ixfe4uhB8yyuFoqWKohY4RSQ5TZI+vWBH06R/v1eAUsOUglsEPTdF49xY
LjffeJcHx8JO/t76MZ7xGI866xG/OIemW3vQwqJsxig0G3NaVLK4untafi9QMYKg
bliqN2bsNdlhOGOLMuv74aoBSUCbdJIOsCaRseth9JSbS25QSDg2agh8eFrrGb5T
WcOQEC2fLScKFYDentd5oXXIp/IzF3avcTDb6YxQsIaBX9T+9SdZKI3Ipxzz9AOY
+ndH576wSZ1nV2e9kUZ5WP7A9PlqCddqBraqZNkZeluFxhAWS3GqAGGzUFgm34pn
NVCiZli56LruThz1rPNszBgCQkpn1aux8fUuBg2OEoIPUjT2loamcHZ7xy2QTE8a
SJ2VqFX33MEc03oQq8trhSit8hPEmqiA+ughDtNwK2UzDuMaFmzYCU74m8FSFLOm
AkCyc8S5AVS0MwSjtZZ9BK1uhziOXBeZIvINOw4zlK9h8yauMvOpyuoMmldbTd8v
qxjfBifdlw8pXQcpOYQFYrPuZ6cyt9UKz70ItdrtMHMNr36ZkhXuDbPt6fr+EHMD
J7vYpsER6PZIfIPpYBVA8WhfkTcx8HAGxz+86mREFYlueOn+LbM1aZWCgaAaiXqy
Se5sfiF9URljDMWhb7ULxOm44MFBvLSiQ4O7ibzY7Asgi89vx36LiTXtc7gyDlH9
jlkqhOuG3ExPZnwF0OepqRO8+9iR/y0pixOvOlcJLG6Gbb1bx8fEgntV5WTQGvam
Fz6Q+JEvZehOOcjoKPBd/qC2ghz4MGF2buY+oUGIEMAelpb60rmbMqPTj5ObvEkC
mWmDTR2hlNIB6Jc0+t96VEMP6l+QTmeH/AalW9dwkzQl/m23G3hVw2sNSKEauUts
3NxdgYDw4BkP8JuqtKT+/TEqDOyqdOkXPb2rUtIzHlafDxxuZilrltztGpLL3cXw
BieIu5jT/uwGiBmEjm+qoNC8n9lc7mF4NjVpyVoFsZN8kvkMcxQiDvg+cy8xB6bf
kglfBgwLF59w44yQ70JreSkHRfg+CAolevHyZmp5kCzAon4fSJnAIKv1jwmm+Rx9
xkBK5S5EcPiLZbD8x3SNvgfBh4EIczChZhR5SvgGjFRiOOcmDczPFBgoUoh+HKxG
T/4dUxGOLvxFUf5UxnewZoTVy1qfmQMw/YBWn89QB/kOBbQcC2qe7Ez59LY8+Def
rbsCUT5dpAUuDcvTZfDbYtO6QlWqMNFbFKJiLtpqqdMGOLoAoZZxY+dujCk0x3Ae
UNHLIVjrKWhOVGkJ37T2yHnjxeKmHhy6pINHSlxEqm4B3DLlzfW3qacunQDDw24M
IxNRJYchpoiPoCMBqVhcqkk2PKB9jNC60YGefkpkUb3zzOOpcLXKobTkfWJyfNlR
rWJNIyt41rU5GVO19VJAcrewqOk5KIiUCUgrJxFKZoF6Wuqie2HzCOIjA2JrkjEY
voFx915Qu3dMqK5ywE0AYcsEy4fyQ+Fulp7cDgYo9LYQqx18tYqqHrcMZhZwnFmE
+DfDRqtEcDwj39K6hbCoFBDrqa0OXLnPZNJxJiRt2WYrO5BvZ/0MnSoTq2tq6WKE
wpF8IC20D5KPAwlsXc0OeWuxkw4eqrAlzfjo/XcwLbm1pBpGzpPeBYasJWfuUFud
flZPXFKKXGbhvNL0jwUxiFvp8ckLJj7XFW2bsBhkgGRR2PIRgIkdfXVjs/4MPAw6
Tw7fBxiXCgWfE6K53OT7i466mYNrRWQ22jad4p+2ysR8Olj5lqfLT4CZA7pKD3sh
9SKDjzpGEh/l3LNjfdXuWWAR5klUt9AK5VchXRTBSzYQUzmJJPG1QRxM4MowRzbM
pQjVrWeWI3UPQidqMZtojL2c9RoDgMM3ongHerdLP10XpjQKfmDLv1brvcYC63Gk
lvQqv/MDdM7zTWNqAXyz7Z8JHj7936gKM1y4MqMdhXX5aM1hfVlv5cfwN9E49kWp
EZvioltIl6HASWcW+Cu3jiRG+GjROduhSXBkQ8R87zhas2memUukzftFGpacXdTS
c+RlCckiAwOhRkrU/YlixPqmocsDzd9JlYLTpeKXpP+Ik9YSaFXq3BvQ2uZHNrUb
0EI8MDV0ehBH1t5HYR5GAVhVuar10B42yeBLN5ptJaZXtvQVZJ9hP/UnEhY5G6F0
uO4bOAT7GvromLcXsH41q4agouo243y5hqjnxFxFSgJh3MB6NBh5+Tq7HriDH7u5
VqVic9wSyg+bWtohjfuxn/cZOLyLHjPpm54JaLQH2oOpZKLk5NJULkIT7wcT+KOz
gPeLsmJM0OLt71q1scZNQoqdUCTPooDkKZDH91IIdaRolzT67y6P3D7VkMdVOJY9
qFO8nTovbyZoi+diuztrNE1tGG64ziYjD6r5JGeJdQxdeRRE2D8quHozG5dzBF3x
VmR0JzXsPJV3jhtUzqC/W+LxbB1Y1SgY7J9zpurbZGfnxpRjlDd6NNfpbdjEUHq/
YzmrhtfaFmdh+AP6e2py8KJWz0ZiChP9/OgGOnsqwGJbx7+usINmfPZqPyGX+dvp
yBBYz4p+vGZeWtwP7j+CyBjgHpMMmSG1yWXBVHlWutiUQsK0ZveMEaQf9hu/Eax/
1po9Hkih8NMPt+QgSpY8NBX2Z9UlDjI5tb9p93vxfjBBuUYY2Aa25n1fLsBfVymg
j25o8rXKuQgHyHxGqKJm87TXsdeTKPWbVrgHjCm3Rmm4Zn9v4zBh60rfOpseT1L4
vgYA17tW8zYQrMXOhmxHgHPneG32I/h7XQPmjZ35+GHcsu2SdqGe0TClKIPkvZgn
Ro06qLqyQoJqHuiizUiwVyZXwioaFwPa8YtNMJPRjNVlJrrpqlDxhIG6kPiujGkO
5kDBVKElt2qxaBqmBpzQlWk+hP86gPB2JlyQolNLON7p2FEfSqmIS3JiqR017n49
gz9as0f00RqZZ02iXRb5RE/pR0dzsuAq3JIqcDUn+ga8ox8fIBrHlt+wWyJmtWU7
UI7QARd3M9SaS2OmqnuKxojSKuqOuFXDQmH6cFCW+7Pzn1VRvqYpBIB83Eqft30m
j41fLR7NAgUbQea1ldc6sPZwDbxj0uZa9KwlVh2jsWbPv+FtvO7H44427/ulZ0Ly
yf6kaC5UpsEP9iewYlCfGIPPOEBRD9HC5cuuBIlZzxw/teS4v9X7QAoODN1oIurP
sttLNHdLJPaxmvHqWZgfbad7zbLjysLlpexaIM5ojdnkjHhrp3and+mbOnbD7D4I
D7rSCaC458P9JnESHCX02lBA045/QvGfmcDpsiCgeNMT81LG6Gsg6reBRRkIPpMJ
H+osrEO4RhfrOFaYSq8BFPyiDKNWnXHgOmHTXtj5TaQN6TRX9DEga9/aUx5TGoxD
Ywk1io3aO9+nAnR18hZWAMDxLtW9QiyW/fsbSN0Sx9PtwnWzqjKlDVywH7/Sqkz7
6b1iUvcYV66GGeWF+9eMiXehStasX4a3TSmRq+8YNPfja6oqXTYJGJdzgzkByBFJ
f89+IyAFGAIgenu8H+PfMR2zWTmYBH1JES83o8lSBFpQklBbaevFf43aRKENT7p5
kOijnXO7G9wV4ehUZ8OOp0RLqcWmHVlOH+qi+QftsjgQqynP5kUsDjpSveaH+1J/
EEgHMH2RxxqSbPyJb8s6gVjlrrC4xdpsASYwl2bEFPno4F8PKFKykExz08oAEa5v
vwKYUdkpsNRMA4GRKElsKfraNT+wa8n09OS/ZXoK6BkLGXOoodqOVNj6VxdD1EEb
fSANyDUwWhulshG4ZAsTawA32U0kDXzYus/uOkeRU8G3yeCgArbc//j+W+TsaFUo
iAojU9H8UBu62nzLOynKexwT9CvIT5psWFVPy6QNQtQVB+aTRrkc15i53Ac2mAJj
hCjdehd2z69papE0L4ihAIE1ZawdaRxz7mKQAv0ZL2qoBp5Fz25YCXGf9fDZGLPY
PU2aGKoPertOtuxELq6hYX8NUDt4a6gIkrYN0Kviwl8Yblvt357/Z308sT5rko+X
Xu5wdMGtAixPLYy3ZtfFHMgV6Q39Wq4coQ63NpWDlnWJD5fydINf7ZDuDVXh6JwO
VU2Jw9GRf+qhQSzm22dFoPHp4mlg/7+NH+06oNrFHjJbJMYZeCRr7VROBJG8WOZ8
Toa+6YFTJKtrMpfjNCnfu5mX6l2BEmHotHKSZE8t/iv7Qmr9kWNSf7mqwq5kZ6US
ScG92UkZdw/fylQVprf3vlgri7zEZgxgmeL5h+m6D0K6cumNl1N1qd6BdD9YwQpn
XOtjY59WC1LJLVmPLvCFqat7o4Qu+kOKgIPBcFfh5CrzlPi0lvf/yEvWunO4Ijt3
7x4fKuFuOA2HWqjwKe8oJU9+WLWgWDr+Yeq/zovLh0KJPCwE3POXYXpMgUiaqSKI
XQKkdRFNK5l3OHhL/ZE9HR7ZdOt2WiIZfhAHCIzOeZyZ/WH3j6/5OYQ7Ow2/ufzW
keoY4XpeTboObkvi/WQUTwoWio+sJAvORo1X7875K6GI5cHw28K3E/VTWPwpmMGv
DtPap/W3Yvj/1Uw/vQTYmDBEhF269Es/E2TwPko4l/z5Y0nOgsbl/TXRjMJ8YpDN
FmOHlBCKKqolaWjNI+jzNQ/yhyaBADntqxeZLhGYPqmcMXg48mjYe1vvHfMBw5vZ
N4Yv/jmdqUhA1d+pENqBzYLyzSAn2gjbN/4DBXb3M5kFDzW0jLoyh82XdtzFHr7Y
jCTEpRByuc15376E4uOottxRMdkr9QRsCpzWndV4K9Lvx6nJWV7GCnjbSto+3EBQ
9f3MKtDqqgyzHEbsxry/fpu2fgbSmNiOtFmFLK8N3vpO5YlS4fZYHQO2qYGnsmwl
k2vTqwP0UR1PEyQ+LtPVya7ydnLSBpI1QyHDjU483xhDDV2yfgxsa5AclDsgUmis
WTp+giSyax4d52tbcEnoKabvX+cuT2VzFZjdiFfG2ixWtgH4RsHb4j/KTaJGPVsX
0Lco4dLftEacUQq6gM6amuNGVu8l4D1bgYLBblbEAX4LseNzYUfHNtyK3yw8jimY
72L6fORbq+CqudY3LftKDiU1Y7RTKpLQ0GzBddJpfHx7sJkpaNywCEjRMW8SK5BG
bWq5cNmQOygKWgOt8j9RiWWMzHRGt9vIFYR4r+Mee3ju0PRij5IWVb7u87h0tJf2
lQjpqt4vURheUhIHSLpI4xlGfXLZABJgBQir6GGwFi6b45MJ8mVTDsvhxxpaNCgJ
ti1CPJcXhuxky2/tq392CMQFKoQm3o9+MumRkURk9wR7GsZO8B5Z9DELD4riQtP3
LPhx239Fv0JeJyHeq9viCl42JBibKVYvIPKv8C9K4yFyqU9sbViWK2zGwofJ6pgO
YBLc4R3Nqzec88r0cuAKbVWdR/IR15p2S9a7Qqh4ffFxJAR1Kphv4mz5BG3/F9mq
hTSuQBVzA/mhRPNT4bmtTWgX9IOiZ6Q30AOumkCeKc95wn0E1jzWwvmxE2JaX2vd
ydBh/d1daDfFyt7zRY58AnhQu6e8E6ETe9yrxP3iQYRZ2mOtanXZlsf3t6bRT/YU
VaSOImL4uwdlAPAPPz1E+EfKO1rttR8Ai2XfXBGXtvdRRApiN9OznNPJxaY8fRgy
0xR/wKy9Z+J7RRNGlPS/39YQ5ky6Uf+myNrIxSxlIpq/3pMeev/E915iImDfbZWA
QOnh5UA02VX8UmjtbCa6+Xlj7TDNkvq//2gV/MmyU+lvULnfNO7caKiaKxzL2ys8
WZQeGpfsZnLw+0VtwA5MuRc/ED+AxD/SI4l2ix3VzyN4tb7Nm0a8G5EOljEfYuUW
4YZHYzEIomDxExt2N+aHmBQ9OP1RQkAzTNS2RR2DaY660AqGE95lZ4J0L9fOz2FK
s+fA2wrCU8DaS30rHZreqnZM3FVdIvZNfPPpla+oRhc8TxeskArFSZYAvwCScWTm
m6WJDJ5rjZWyG/XaJeuYlSvbKeRz0fJsCjBN43QdDnn3gpUR6MftFnE1YZPYayXe
vlyO9x6vx65CEPmTWDVRUGnzv3+osh24jcNKtDDffObwULXWKdG6ho0Sh7tCYlp5
0tvnvw/ox8oBoxIqAS7Tsq72RH93XmHstFv2d6pm80qKssUBoFNQX/6rUdTVSdJG
Urgo1XT/AwNqwHRC0zq7O3lIOqtM/4ay/Mfuh98+dn52K9POqMF8XXpE3gCAA0Ir
U04oHiWXm5o66Uwu649/ahFm2gtPg2ZtOaBe87DAGtsvvR7W+6Y8+pehq07LeZix
jr5CGU6HXymJ2/UCjt2RocuWw50sY/IemRBu4UwsRjgOgQ2Cc/n6KTLyrQmZgQFi
jpnu0WYsHQNViQ15M13nS+uNJTFK9QWCVk9odnMSQgGHuGOdKOjLWJhP58BCPdyy
ZFN4ChDw4R1bmjnsAeSQajhnHVl/v2YNHtxZEfwY0/RZs6Uo9UFILiTR+7GvFNxQ
xgF3ZHTQPCnLHkSsNwPkxYYPXhu8ael4I6PYVdESyrQKdjL35EJLH3IV6b7lOaC8
6qQLTiFYPFpJTtBng12Zz6AYupJimC3orIjnr3itC6KmUZyf+K2CdrPoYGwNJt9B
BYPVAcVkfhuprEZKRjXVyscIIUSg1Hyl2vWSqOVh+R4fZxSXxdq/cx7LFt1uW7RB
mV2iBK6JnZAGoP//aMPM/QTS+HfEhrFW6SA+8K/S/yWqhluDn8yvTHfLGtcQp37E
4WRLREQBRNuDydELxqC50p06I8fut9C0L0p0IWCjMpQ+Kpv8/vlhuAype5pUEryI
hOQwKzHGoX0eU36IHL7gROcOAUVlRxSGKK5WYPR/cEh/U3xKefrDpfxtcPIS2j7b
smHnho0Agg8G9SJjZEvhyI0ekWJS8l2GJOFSferI6ZIMxGXiSQl2K3jQU1V1GJic
1HOGUuBCGsJmgBztlPoR+cANZQHAejZ3yfjzhkimmsurULuOaqrYz5aEBhXzDTGW
Mpf/l7Kvs4q/F0K4mvQj2T0LJK9tnnNKqgVnNUy1sRVOVjqum6yS+eGNHTkO2a9E
+YPNKqOp5yRC+vbHxAYyfq2qcfi1/oP+1kfxmjVNCFW+QRyMlltawnNvWe29VvLo
8A97UzyQQMyCi9OY/6b8vQJA9psr/63oSr3C4qHTplxfv9QgHcutFE97TxsWGRgb
MXPxeHIoLnOEm4jH0JafB/Ik9YdDQYPTToAYdNtyZ/RzVQij+o2TroaU7pNjE+j4
5OFbxv3E5xDkS8Q9UFLhJKehKXnF8ARRhhZoZ2hIWXgJ8Iv2U9ef2P6cv5AfmuOX
puBoPhgdyN0f7VoQq5RsxXnpoiHaLoTIU5HtKoUbbY7J4i8o8oorkcppHAmKYCMh
dyg36xn5fezPoszxqK9ojGOYn9kgvtSShaSXlr3jbEuFclUtY5Sg/xINO4e7irr4
HMPW83SehD84c0N4ttY09hVxMxYLDGcRNnIZxsm5jKLv9jCEXWIZYCbiqk/GGDRV
zs5TNX4fN6qkidLNT4JyfmesGu9tVTfXSWoZR3L6p0B4771V8COOx+Mev/VwVEhk
RY7adzRc6WE6e1RkXR/v+6+6EYW4iqkXpoGtWeL9uXqa3DDAU72IWKrLHGHexKqX
0IXCvTcBl0zNDRyO8V5dtKVQhBJgDjFGLXcHxpn++G5k9nNRt/iSRNYQT/Bf12JT
edJaKxaNg2NDkYDJ6BJvSrJvKk9AN3RsiESdy5K6enx6OXgEkUopbKsunVEe6BIp
T3DGH1qLNGkyCEj/W6q9nF6QM+2HVgS9Oz9cYX+VmSZSFQaplCtHV9EqE68ROhbq
m7h99QTko61MH3uGZp9qUQY6aHu9UWsEDdkcYXcWuuZxBD53QcvabuCDyK/Gsbd0
AT/tkl3UmI1tbBRU7rsKogJr2iQN4XUVrbZhe6MKYU91BEL727cLCLC9U2g1KU/c
q2DOdeHzx0LzqsS+PqKgDVr46hjJjSWkR7CJSfwSHJOMH0gzdIyvDODFkyAn1GNC
eI+4Fbmge6iM4UXyYz/uTiY9SEaiXNwxLxRSVTJCETwhQBmHg7y6Ka5DLLqEryHU
POiMMlrLEnLA6G1Hq9BswXTEeTJZXxtuplhQH52yXTK5rC342S0RzM9t7xwLljWJ
Fb1FDSHWNhGveGyLPnM0/FZ9lEsfpi8fO4EtHLgVJJiVX7FVpo24dQZTSYYgQzPN
5PrfZVZvJisfENzADiFPBbZP7eKugv5U4EOCrYRKJODNPhEUdTg9OnwOnAqbGGj9
ZEPQaKNoLRn8yCD8lKlVRAMBAwC0O9ZeNT5DVmVOmF6jjO9vEyB0bSv/J6r5FoMt
slNvRY5M6pKs+XVO4KFpb9Ta7eZvTxdgI/Odwix7rrSiVbvHwUc48V8uVzrNDSS3
GB1WoE6N5V+AMYS1YOxj217UtEwhJeNG83Ag0Qr520vqNr1NzmQqEcE1XVgpFzPi
RIwsYjPYbHqh+M+shFjiM42+r4plza3D0H1YPI+JDKPS9GlRznxLsqtRSHHBUr5q
9h84//WuV5JrUZvcxOnbXM52Sad71QDIkNjqCuobOQnfrcg2qID0ljgHpMC4OssC
OGXngZrvI0MFYOyKvalVAfoHegwl2eTccjcy+MVbrq+osK8fOikziMxGVnlNoGQU
zC5HpkBD9EjMQa3Is09CPBg3F4xE3GDQS5NDCVd6V7H1VvgJA5kRljbGOCJUKAeL
0+GEp7hjvJR9MiSBUgte/JX/JZOAzwTK8V9pOqpY3+I02blSYivoNM2fQjUENptq
mMnXfKSMZbE8QLCwrhTujODLcWaWZGoG+c44POEAU99Xtxjnnxf4cgL4VKtpQUI4
rype36Xu78WtYxOJPwvIJ9lVUwebBMib6PXO0HVi0hWene4155ATJ14fMAT9tJzw
xRV0XNzhdgtuxi5SW0T2EOv9oyuf6VtGsp/saf+JUwfXM3nalOWVg2gus0Wipl6y
t1BKlZEN5L9ofZgLLXzqOLTtE1Y/KqicPMmQV8kN6Vf8rAe38oBu/WrouMbjwgz1
V/HfzprHg/E404gTbCfI9eD/0TcngpeaoUoaFiusIshFsmOtRxCm0oRjVZuCDOsZ
cEjASRsjikaIztl4hlqHs9BS6VoU5DAPcdctVry1c2kNfaySLdSz/YiQ61CNi+4X
xZ2oCgOL/Zmi676pner+o6+nW4Mxf/vkvF3y/RGE/+IS/gOpJZdLK91Wg1y9fE2K
Foeevx8mbzmGtUmgoh2i3OUzrS4x+L+dyxQxr8Zzx28wDULRNDlA9IuE2VilY5Dx
5xqzitM+P2fYzyv1v1zZL0+TNro08cQX04E3VgVvYFPeDjfCOVGbye8F/AcrbWnP
gNnHCPJAabWjOR38uvCxznnMLQym9rvFve9uqI/HMb6Wc+wkImjMn2GlIap46iU8
ScHSJzE6wgbHHdjc3PY7eU+/rGaYHJjEcqA9CwQjGKS72kpeqKLWtpIw6eym915M
J4e+94IsfQl0JBGhl6uR5RyiVJ1LaWvtLb6BurGkvP/BapHUC57AdTedHz81FfBl
avSoVBrxGUjuhBTo4A+i3k0XmsEKWfvqtpBg7Ut6UXff1rL6N3GCCxnrqiCOMfRl
ZmMn5+/HEM+zgUPw/Yoh9aWi3CZ0ngp1Ju9FO6pWNavZQ1ahOtO4bL5OAhyicPwY
U1k260pTxWUp0y95PKha1KHxHHZI9z0kfgOXbn9Ib7PG4B8eoIfR9hrGb0JyDHpM
vSjbiF0FAT8y004907vj0Jrai3XOluOQi7UaU/PHtlu8RM9jWqu4PAeVtbD46o6x
GU7+YXxtoN5DhXWgj19TNelD2/cGuSei1+JHZhZFXf6gsxlfD1tEXEO15N90PfYF
pHjXw8kzJaqG459sTAZuYglDRWgzjpsXs5XeJmbFM+9CpgAHfP0F/pSdD3HbAsja
7Zg20O9nDZ5Xjr/iPG4iBRq0mjZL9HtEvOPhJDItvWpmwiIbMlXw1aB/whH4exMw
z7tkkFI0iriwz9XSUUtuC/6RU2LUKNnDlb0NWcmbgiHsEmtdQlxQ94xWbwvaKRGU
kdTl4PJ5e304FJZ5Mwem9YnH/GCJkJNX/+n4JjoifKu1u8G3D8dTawL8j2sjGH4N
vG07NMZ4tqQtRfYNNWVt+8TCEktQAj9VvPQ0tsvzmR4MzSTeYUCvQ6Jc/VyGQPXu
dYZeAojHzVREEZxSxRMRWRPW40t0ts7RdGrEbV5JHZqSPqpyTfaPLmJS9QLmusbu
wGpIyDRrS1o5dFq7PEKUxsU7e4BEWwL2MxdslHqJUHTNvqoEdYxlhZc2yCWdplFx
jAsUZH8mqO3eG/L2ndJzGr7RQF1szDmrCMJXDcHNap5vU+/k2zg8FBu7fT3bQ/mv
9vBtYJC1l9tCd8DxPZ4zZBVQA/yfhogBY/448ADjPMP4xmkO5IiHUBXihoH+m5yh
ki3yLh7o9HSioPpmrH0CbFp8lWAUODFEVa5x2PRuuhPUJoCaN8FOe1JKMHYRFpqX
Qp0vgK7ReCgbTcdvibRKdlWfbigiNTcjLf+phqJukH9fPJgSJHJsN5uz9PpTAKo/
dI4B6z5Zo6SvRu3RF9OY/6FD6pg91Lwo/f9nEty90q+J8UhS6aNFwXuZ3tkaX9cQ
Afqr7J/aXp2ns/xf3pRxVxYoyOV2/w5WkEiqGr1plgP/W7c7CoNyUL7P5DvpCR53
GH7hn/0kYIJtGlyng40wZnZM1PPJoNMEfgeBAXZh8qCb6J2cbhaRH1M+mw3rkTEC
UMssboWN32gBEaxrrEQBrMCzOwWCjqPATVI99wNoxGz4ls3Fw68CDXxPVPhwEXTQ
6n/1MBB0S+l9SrGEWjYuxBtX3trS3SsLRkp3ECQ2A6gjDgF4Ai4eIS008R29b+mQ
EftTx2gZpXiqEcFdMbINwdbAwQ69glIeRrOcAImXrOWyLyTL+m9nci/6m0AMOUs+
kJD0oY2eEpA40puv8XlL0xkcbT8itZ3PIES0NBfUajGIjkNdmM+PemcRmLcJiZ8r
I7IABuQM3iM0/YXgnFPekPjdbJ2CT8SvI1HSaikw7+6/DKrx7Dz61HUGG9hkpPKu
oQkOHkkVxtPJpo7tw/di5+RTApfcnlX+30dAjV06BRO1WvqVs+HnWkiyP7NIdJuY
l8nrpzdBT8962md0YmJVADp+fD/NfbZFOOiK7BcYcQoRsCGuVq0Tdai8vYXr4o3W
9EiZgISM/iZEr2q332j2Fz3F4OwxcriJ+aj3EYlEtUiJoEhZc51ef8I7s+NG5R06
zW6rH9mVys7Xc8gY1BL7NwsQSuXH//ddmKyqCjcbAqiejZVqhaO19Rsp98l7AkYY
aFtR48qIPE2GVcB7ZEwoMkvzPPhYMBIEuU7SlbY2vyfvNRk3iYWDG2GTr+5nXHMF
y0bS96TdFagBlMaRWABCDCfxEi10USs6FN2dQDiDgX6Ek9Mc4R2ucJoE5ptwA0ni
IOG8PCvkg0SEnFuIA3DCS76pJ4ZHLVf+jErw5JfPgcQXkGYbaWAMWSx3EmCiqtYT
pJGo+9ZyJUW9B0i7zfe0GK9BX28xWB5p0/V8TueKPTZK4ycMXwS5r3DxEeE9BmVR
6B3AHZvUw5siJ5cfHpaX/SRma1PWwcPDCBCAyCgwPUeOIgsNSCNKacOSqtPdqyMC
2OvLR5sKt0CIS0npYGpb6NZe9mI4RboDBiJSfcNcGi0/oHW9L1m4kjaIpjxIThyB
beygCSIR3wB1NsSHmQdHlfGnZoXx65B9oqSwTp93/N1XWReViyFUGARNj0htr2DD
7xTcKPVzsGoiiWPYR76fm7EzklO7tg6UrEbnUed7WMEFTy6SuRxLHo7WtsR8SbPP
gBvnw8R4ZsUzbY2oBrJFP4m5Ie/DKFFazLHKixDnpGxbfpQ4gMLFvUngOISoDtIk
1/pa7Op76J7SuvWbxO3hMuA6pdbgH+V7qoLMWHWNb0TyigDIIjXFPRFOMMzj1zhX
6sQx4QjiFfcI0jsC3UVIiDY23UW9dQr8q1lqMVN7mTKWKN6zItbbaefPOlEHNsSG
fCbP5IqgfM2cRT/5rnKuzNct0brfRNPapr8/ocy8twuDnYbpQerwh5x8EjIHbour
0aBHaES0D0gw9UfbOEu9Akf2v5wf7StXRRSq0F3XDungJ8oR5xFovO4GLSMzr98N
kuF5mIFXenaM1TKAqTR0Sgz8Ug4/RP4DqaXawx2Nl3eYmxdPIoetaVZiYz8pScnx
vH2lB4JxbNWD/FKCdPE5nv/ZR8R50QnrGrt15Q+y5KIZ8KbuVBA376R+7RTdJ2mJ
gsH/O0nMOuN19s61Fdhu9kcL+DnYBinApgiq/IVOKrup5sW8nkybcmOqQqSJv19C
DV5jZG3P+6Z7ViHNXhHrqDd0L43xMtOszdPe9fEXYSFqTZS+BRxWiTAV7W+y4251
aWpJWpkxzAhee3MfbawVExyuGhJGlZgTqYmUbR7qrTr/1FrS/x4ET7RP/iZ1/lCb
O4W/d1XO0Z7Oo1hPZgh/YDRFiZuDekQ/DUWTrR4ZBF7qL4L3wYXPdFaVlbESldrn
76mIfriVmTh9fCURsAhzMH0nWSLwnAVKGcMirQkqr6tMm9NbXi8B4zn8F5Gwk/ke
t5gTkrbXjczc6W1nJp+4GvUotrBV0wHqUTuh6/3JesGq2wpoUHoTmIctHUaD7MKJ
vHr4tGgodXjjQOHavckbW9tYtfj11DPvljItHHlEh2J5FLLAghNTLoaio31j5RYP
hwojtZ3iALJxtz2t2Z8TVRW9axEU8+nQaNpkzmNbYXUQI8DxzIYxiimZVqW6xsjf
eiqO59szYNNDP0s4Laty2HNzR0NXgKcV2t4kvuNl/rJgE/gtawH2Z23Bl6chVUh6
h+NJ9mEGFdPzsOO9d7ot0UvSeSFlK3xfkcpleGKm68GrRDZc7k23H7IgABlQWvor
gwTNv24eshB8yr1LJffDpxuWyxCxuNsRoWA1D84AkFp9Q726Geu44228uC4lkpzZ
q3oPq/g4EPzklcQIxylYpJb8YBGDO6muBuVnDIvTE1X4PGXVL0xWMoqDCBgeTd2W
ajJmz8sxbulMAb7nX3+lNy9Lr/SnkU57ifUH8J/woLKR2LssvziJVjuy5UoGg2Ah
vCQvPj6l7Jg0XL5K3YLWlekfNhFdn7vRYcD8NZPzyMmPqIV+tWJQg0zSbGHmRlIM
7rUvpPpoy8Dd3f+/1gYCwKyxjBLgt5azH1WdImJjPVne5bwFGZBThFgtKFRUQkZs
selF4bNvhMKP/QVGUHkGX5/bIWAxAE4xlfZrT/p/cmhPvNY6AfeRjrE7V6M9axJ4
OjQsuTWcsR65dx1ubqj32xs6XkWordJlOZ8lzWjgh2u0ISjxD0GNOZjTwEb/nt2f
zEJv8WsmnlHjdgHMQ08HCFtTAxty3XPkmpmF2YV8etGLaauhZ0kH6AfkowAeBXeb
zS4Foidw4i3Bo/EGOwXNthgPx5Xes876y8/S4WaMzsZN8T6Zyo3wnttYeXaD972j
UzJjPQhhZizXPTGOwW/kdg9luIGTBdr+P+ySxpig/VNCqHhEYtPnWm0aLk/QbTAm
XTtIQM1TkAFgTeDHeT9OJuP0SD+WK7at1wsE7zD6uhOYP9gttICDSDAyJRi9lyeW
IE6eBg3jIxqfz85zdH35nA/tUiUYxAI/Ap38sPs9EiqerUJ/WWzxC4ycZmlE5vDc
Dxk4E4/1rETOrLnyfSi/fmc9ZAQwS+PnJqcfvcAzNoIHgpwO2tCzvVmdNtOOrSt6
BM4oBsDAd2uCULSYvTOXebdBVmxuroio0lPfDFZBuNN95SGMn+OUs9D1a5YkrkZS
zvwtdtvYWVAW6F4AaqjwbEFNWQaIWB+yfluPtjyIK3xvhoP9rP4UHCOWn3sVbT4H
tXq7XMOpCwrEfAZfYBbupJQojn7CPqVX0XSnpIKs+E7SGX1klHpB/91e9IQ8j05e
GrASJ49GR1hKAJLQAZxctmdt+aYMDeamwwzly1ifhNfCfk6vzpsF7QSnvbQI9pe6
pb83scyt6/lGxcGBMQL8tUiDfHhAGQ6z5OMNX5I96YY5tsyZVUmpZ/Z1LgRUYo2F
Kv6OtfPXHcDTzwLUfHk/9e/fOp4m4/bAWCwZWPey30XCzw3gDbG9z8AZ1oqAHfBu
4WFFRotDFR1RVZRACXNSfdV8dMUO0huAp3CevKPM4iuwtkGWZvpVRE1D1NvycOcY
3Jve0jhVZmP/eD9b27GjEZjayA45GaBDUAPUEortoUfYnrPlWez4IGW1QfiNWQ3J
iQmMSi1XTpw09+r5yEIZuriYKztsfgkJtlDhjMNJPFNlhjghoCKrCJj11QUAe5+/
2gO3X5M8igfCVvpel9aBhssWB+oGGdtash6wkH0G6BozpF3/3fo1h85d1taAbbwa
MF35Gpb5WGNDchHABrJy2ouQo5/QzmS59NCEhEPTSFvnJGo6CzitCDVLtMvh1xmO
D4jf7KjI6luNIyaccPZ6yAmMEuWlHZWmR3hEO+/O4k/tfZ365dsPvlA6MoUCzzDQ
3R8jiKVXDn2P0npHO7D8/QQYqs0DDZ8nFHrYwUt+tC7WZjeYajmYATwNGFY9JQuJ
RVOmaaRCqKyaBnT23FQpoYQ1gpEw1eamr4LzcfU0KPif0MAsEYBazG1wbi22N7UF
yVIbTzFzxNDDndZNLdB1WL/aLLNL6XlP9J6jZOKjqHDlLd1cVwlFu2A0wIzV/jAV
qBJDNAvLsarRHM1m6BhG82i+inhBdVv5gwKM3bq1Jp+5nDjPXEccRHeahmep3wJX
J7lPRMBjfZA/hqAFiM1mNq3JfGQZE8M/tK7eZrNbUFHVPE/fiAb3Fzr6tcwAFhgV
xz8keaFUjStGbBt3oiDUYe2nabTHHkctRzK56wKWSzPAHQHlDLRZtGdeHKLS7xla
5u68nwjZNel6/Z8FaE4PVH/O0veFCWX7OE8aS3zGO/NOrLhxXjzRdawZt5XkQaCh
Miojgx7kPA0Zm5k88tzhxOQIdlOqXzkVZ0DDLfp8oNSXxaY0xMzi1rx9XFwPL9Zu
Lr4wbVoLtlpSODV+se+F3d+d/mHL72qUCRYSky7mRxEjYCqkgkuFBONdUSn8VBat
rU43udMzoXy84PRMSuwH80ZPLay8XFGpvhN91l0sIuLCMCr7AI1nKJRg1ZqyS+n0
K08oAhUzIWabna+e4vxqYoAzyQfsi4lB7WS1naH4KVS7K5l6S6LniPgSVmQwK11P
zs9Giapr5ygBrzmqdzIe0x7snnkqDYIdQUyW3KA05sF6F9mzXnkLgugu2bQqz3GR
aF7r0Jinfdr4gZ7D8B0o6rrJGb3y1uJW7Nb+PMhEHYolepZHzcd8KGOm084G3w13
pKWAsWTj5KJc5+bnVA8VOH4t8F5VjHOhfMkQGBYp+IxuOWmGx8x2keARLrg4aGy5
SkYKa9Wx2uCRz758mOqCGgnPXKg3MYU+fYs4p+Lw1ROVCGNkZ/LcJK9OUf0cZlz0
0X0lQcS4qMEzWryzx7rY6EXoRpXk6ta55qeV/P/qgKjbkbK7iy5M7nvHlFMc3JiO
hfaEs8Mp0dRc/iJ6aqRt+NFisix0mrBxF8Yobbtul1OrJFwZhbB3M8+7V27AwEO0
YotqHbjpx4vfahWI3rn6en0eKZ2wlMxnCix5UE5toyeYHNy9plhg9VfUnNaRWoi2
2jq+IWLI2xXfdxXDzjBvsXzPr51c4CF14DFPyTuMO3OqhiXSCCAS1YCczmr8Huf8
Lvj+FQy11x4oDl1dvSHqQ6T32kehnGiMbGDcKjUOG4VyTYEhdM4sZVFrXMLLUX1Y
r8XEvsL9l2GQlFNgdYpKbSRkv+NTbUREmpRZZMJyMlL6wfE5A2ffGJMta/cTYMx9
aqZvsPabHDdSqkYjrupHbPQzFdy4uCEO4VSFIvXD33dH9zH6t0mrz0RlrJJLtZ2L
5jiQG3o21/iL40LjSlZqWzchDCfpmv46o3mBI987UJEVA/38GbeNc9x75nfHr7Is
XIRDZzzhHF330P8XfFWZ7dhaxoWHPl2NQJ3/DKH8YppORuSMgp7zIKvLd6+5L9VZ
zIrE7zep+UmzQ8sAXWYRjH2uIBGWH/r/x1+pcgWM/EqBjFJB5NE53kYNDkcrzx/R
i7EIAFRMhN+B5AQTXQ2GsL3V12D3dwYwAScQq8x62mK0bBpIL7XkoGMQvN2Ub2EV
6I95Ot0u//Qi1pwgVsXklgpoPUlrpYj0KjkNcmk/bEM8WwJ/pf8YAuodFyIfOrSh
lbihQCdqwEBPVvNSpdb/x5GxDyu4Zk94MvI7Y2DRjoLiik8zZTxjSzEq7zXb1+no
OW6qoZRFqV3CDvbmi6WrCTMl51z1Q27hHOOkQGVCla5LlL6Y65JW6xrJsQiE2NCo
xj1MrJjvPMq6yMMxIqPDsa4TjFlGkOpdvvNMTtR1WFa/txgQqU9GcE5y3pf+b4VC
ue/NvIlY0Rbe3nFlRwUSmc3Z7JGll0nDtKIMcoYwBd5VOV9/fi8wxyZ6agbJYmz9
sFsZEw+X88aLwes9MCHkbN9YK0JEi+m494iLAtDHrTolPqfzjg9KV7bToqRU4Q8G
7BFEkVCGNVWbxhvcmccd3w98ZuTG82TJyG28CivVACx/OEmZqEYeJ0sskhnT8DFg
LUDF4ZyeX9gvRAWclNHV+98tADHAwdtXnw5GIMwGfMhi2CSON0PC//KeSD3J3iv2
xFnU6ze/q3ggg1AOVt9QgS5/9X4qA3dsO3DLAyuoDCz7oJOyJGNN+fw7RvztHiTT
+GBT9xIevAEjVdqvm2nctPbh8tfvFzd3lchbxZJ3S2HvTlMWjVmfaS3AblOXOeij
L/L0tXj5jRjj9FF4huHgI3gWywkxATkOEodoY5xRNtTN6p78hga/YIO3Mk4Vecqb
NvFkp0pt19TN+6SneiBNFGqe5k+heU+HL08flyxbkszLmesmm41XyHe3tUExd1q9
pcOkQXelG2LA5F+VudABxgXOPbBMbCAbT1ivkZ7xofDT4pndRcsOg5ESmII5cYpu
7cL9lunhJ7vazaNYZ/gXqPlLG25ZB6S22WIPRIvRICIEd1A9b9v3Qez4wNSJ0k5b
wy5AvLetxNUCfP/OWAd4wDBAyhPXQmrvansy9RfrkU5omTIoqONPr73OPjnugxF6
zVihuGOxdglWqzQrodLIA64+rboIXtUW8t9XdAwDopzfYbfRLXm3R0MDK/RDHzHc
otAUeeuIPGCoRuUxfizkoejWt3a9papS7A7oiZObmeYIgQ5qL9XncHgrbmUTissJ
XO7zo0Lwlf02PJy/bWM9A3cSrdRh3uUJqQSdAsTps00CKae8ztsfeRRqAX2+2C6P
WtCAHtuYZXmDE/VXBBYKn7BPnBE0FJojCsuVdRifNqkQ3GM+kcb7NdKXOtrWiLNB
Xj/A7seQw0kUdjTj3ehg8rfOBx8nkoJu7E19O1Hq8gl9gR3pY+lh6x4WgBQuwa9a
YL8ylawBjfAJ8HEKEVgXSgf+8J63HSzwcaeI2Gfp941svC9HjIIhXtOmygWPSn2P
nIO9HOq3qwJtJFQhxxSCPMzhcqeu/UBAxQ58/8x2rZy8mqKmjuS5YmzMpKxPW9EN
k0l8JQ5Mk5Q2CTSdpEom35oIV9r7KbJDRyyHHeXSgl9Sd8C9r14rEwgpDABlSDeq
IVoVlhrshmSxDwcCcAytCfsJCBfGR74kTkQrtnoBnyRI3z3HBh0EdSsIt7Jy+WgR
Pt+NnCQJJ7ayIQthGwkydpHIDn4IRcPHigS/HfznRTXmCPpz7s0ce+zIaDKTDgrb
W+qDDxCGyZlX2cpzcIfHQjmxYdgrQpKufLIOmFkuYicksl3HKQ686DvwcO1h2cEn
GjzOS+xZAXo/dzyEiU4rp0UP2su3Kw8CWBj64dqpANq+sVzvr7RgPynxh2STBaBA
qP15sgmHCPdQkESuGTO7/3WX3quU2TzsFlrysdaLTgnE7pNaEZ4MoHvc3LVdV1kh
/oDlFn8ADdeO0q+JurVTcHirNZT6aGGPP3hAqFRlzcUcwNWakoG+nZj/pcO6hrWv
DO7t+URiwsOkO7iViMuTX0I0i0bCLRU0Y/hE0s3x0xr9hzsUNnbNP3ztRPqGFOui
n6m7OZzfinMYScMII36qLA5LGrAYpBhVEhzAtNVn/nnAfU9WPKE24fydbmAsVySl
DCH8RpVdBSk0Umw61pRsKRd+CHxc82r0Ym08xSPnCf4+i9Eq7wEh/erktVflL5nz
nZBqlxXxR1Stx7b2ssriSHdJqwrbX6TsnBb1HkhR74RNavHQT2jxd1EVd+yRiXgh
QnYySYoQD915akS/xqJUPm+clq+uJgoi+aoN+JVWXKf4idh+kJD3uLuT2nu6emXm
GQul6Igk+xj2srdj1af0KvPVihDDjxu9K+v9/sb25XMaLco1i75nZdisiPZOMmBr
7dhNtmlThuOyMB+K3vqfxtBq2cea/ZiYj7XhKQzpJ2cGZQGJ9gnTSj8jn6Vr5bpJ
k6ohoQBu+3J1I810+809mFHageU1KUY1FzWF45HU+d/fX6mctn9VcfiJULDuKQWq
AHsIxKPXCPJTThUIex503bW8CG3yYF7avWY8aOFaGtRqDBl28zgrshdetNVGUSpG
X/ST891W+7fFvMkBEqn34QfoAYlTqkZdgqD/1j1lAyT8g1Ewst1z+5LlStX/bxoc
ndq26a9iJTgVnms9HM9a/LYvL1rBuUUanbeBPX8Xqd4ft2tV9EAi4gelmNnJ+iJH
kr0Ju60LDNxbWUuomsXdSMC54uWsBGYhla6Cx1jfuKBT8o/3stAZuZYwpMepop03
Vdrpl75EddTWUv+hoWjZix96NFZHTwwGuEVeJ5kV7EwE6lfDVyN2tLqarlYkrddZ
LT8H9pZw926e83RrWcXzlr/t9Lqfg7T3y10vxvOoK6WVEedm+wjGE/PG1j59axS2
6fCgtNZOUp10B4oMAa7gDumCChtqLbkFylJzkP1vSNhie7LJ+dHvyxJN/AFpkKAT
hrtYIOsyJfaYaMg3YMh/mrE1eUvroY5ZOoXPY0n4ZrCDAZtTB2iLlLgfpEwMCTAq
buEkdgz+r1kmkGboUBEtmvATcQJLN+fc5+Ia3N9XA3D9nOUY9q43VQbPfns0mH3w
vHxM17c0i0m4H7hXIjsUJXSzIR5xX3ryPRFmLPU8nZtpnLiAUABfeyl2jXjcGDDb
IHQmUGDAbf33T8fSkIWBDNMhDUzVBxb36y8d35YD3fvu6iO4Smz3FBg1nI9qGT2d
QS/DcV8ZGXMV7Y7gK6qOZgDzg3EdepxqdQo8yE27rVsVPMERk5TUbDCy7ksGQ4Yb
lKOPclyAxH3R462VcZurdVIMqSiMc82TyxPS3EVNipjy28oFT3XZBK77W9d354SG
Emg6JnI1tmvrl/U/pokDEQorv3vPm9jNc8JHND+7J490PBhVwQ7sp0jWcqqu4teo
KwKoaj/Pyq+taG0hxI4/ibD2ucZKCAvA232YSHAqexCTBJEtCoUhG5HdFN/IS4Dk
1JRZAP1yReYymXJP7+4xXauHzLtBAkobnm86M2mPeocVR546Dkv7+0brxpahGCz2
WkZe9YL/jnl5FJSuVTODspiIN58A+KVbLoGiHaYDkENdmh0Pk6diukRC7iEm/veD
L5Sp7LeJKVsrcmshK/iQ7b0Y5uXcTuE5HIYx08PucAtwl4WKCWEv77qAq4Bzrj7K
wTB4Q6lElHenUyIlVOYvfyx6nWSPv7udsdvOI45cF/oRHrlAG7npk2uxSbqNr3DZ
llzswIzaBamNpp6B7FOBl5PBCVdgE0IwQGYcrtxhZRjeKsHDieXLR7MOj500h3gQ
omTuRYyqeXAN7645Sb0gjVF7Ni/lfsR2STkNvIUd+lftZ7B41NTLFw58hIeWBHFr
IL7ul2Bf4ax7OMrqiYvFnqtfAg3wVkUfxfllv+xYepbqcZfv+7CC2Ds6XTk8q3L6
AWsfZUe0AJN3wLLQqDcQTemBAqBImWa1urBWeDUur/hneOiW1NQls6PRR1GfK+p1
GIU1z3cD7J+V8mI+U09FB7K+TUssZBOmHjjn3QoAuCS7Ozwo/aA/kgn27FUFgjNO
3ujZAJKjmebzMrraQiU7M77gPkFYUVklNdlJYq9KG7/Bx4b9rGNI5XTvoqFglgBX
4Kq7E3Cs4WkDNObTC+7moPDpU/7MUTBkkJKkkyX3wyqpEqS4jDV8EpUo0CWvm/E/
HLyyFPTAH7JXW75S9+JHi2gDAP3B2tJFZVatTtSix4qlbDGkb4kbLRMV5OTy/ATH
LjIJkfqxbJ/7fJ2mOJqm7BS0wc9CsiU6Ue+pW4ikGA8lXNvln0nkL2UwgqEbxpLe
QFo2JFm/QpbAefodkwtnjCiyqOYZ6YAylkkOIACjLww1e3RDsHtZjMtfgnRJtewI
lU1n20WjwMLDMzJOktIgCaCQXJe6hh6Tr2wdE3ijKWbROmQJgelusu9Xc9eoqaUb
jWqPquNaHsKDnpgHqDazdOFw1KjbNoAZg3YZ0481G8KjlSkHGDbCxAKowVecMhGu
cG4aHgYB9nSWQ8Zr5IsIe0vpAdc8rum9j0p5JOLk5ZF12S6ZYeWcINABf4CXDQnc
Qp1ZMGxfTR4IsA3MphIDSDu0IH5cgFXZxrQfFr47udF6nu+IHi/BvPiWdNhal/VB
h5pXvWIOW1YI+YNYhPxRTI4G/NN89ehbfU9F14ATGYL/oBewMtCL2kJ66+t5RbbZ
UR3/JMnaTehkN95ESURQyJUo14648dV4e4fYo0T16fNC4nF/W3taQV6OxBoQw7xt
9VqvSLayZixfSmB/9mTeifV7ZEmiHO5Oz+aH5G8iynNdvZbTHZHRbgQypvw4+tyJ
iQKMBwu/KOifMkCnpFPYqCNvqOP5W/SwA3C+OzyXy/qG8NHjSx0yI292hS5Z32h3
kNVMrKi3XOfi3U76ht0jAtl6+5+SjTtKBME4wjoqGOU4gbsroP9eRM6FVSeB76h3
p3CybQfpWLMLpGSd8UTeS2r+FoI6iiGseK8DtmBXfiCzmykD3N6PensTts+oYlTC
0NlfDySGvqcnZzjFX942q+JBRSNEDSlnd6O6alj8n5w3548+utzQX+TsovkC39WR
BVfZECec9bAQ/r5iXORMd3zbeao0frRQpEoBkufa08FdK0TKIeLMLa0JZYMtvTd6
emoAuqkOyiqjJscTj5y1+d2QkhGoixZqixpbYbz5HLIqf6ZG4MkGTUh4GQU3H5Pn
O4gnFtiQ6rzC8BNMO8Zwl3q6zIVRHIWsfkDY2Wuxt0LvBMPoN3abJ7C3Z8//J7PY
p9nH7xdsy5QfldpFz2KPsG8lLy72lI9zFhL6NHkojvPWeUkONUTTRw2BkNzcyCw4
f6CrQEGvfXVcJoEZoiY1oD7LMpP+nYxloShV27Td5X+dgZFwjfCOKSuNMyhJ1Ae2
QTJkHlkZdQ1dezLBSpkEM1/WD9mrJzF8rCq/+TBPINe0Mzm7RsjWBMhIhrsVMlpU
Zcyy94yh+7/p8Pn3Y9QTKgUFqlgzTh6n4az+EOb5npcDvn7rUhtz4g3oumESpbGp
r3booXzs+EcNPH3QQ5XKii5EsVbIlLi8DlqF35mHWe3faIujtRaOKxA2DinrgHUX
Rn7XeRmGblOxlPHGm/nClDuQzA2bsK422JEu8UCSMzj+C2Q3kNIZXFotGHO0KT3C
lLlvpj6B/IyvgrV+V/9Bz8fyN5SPOCZCCElFr1EqWMVuGtFN4Ktag1MAtGM/AXTL
aGw3FOpSF18XSSXrXiembbFnH64ko5PkVQOpzU8VKlPsaHflFznTZVzr2XsexAPF
KEc8P3HZXOJFJRfwqJCLQ44bP5wuOES0dHVoLSynk9qFwwa2ms631LxxODAWo4oC
7vlaPJIQgdPtOGawGs0TCFDrFo7wZbIUDp8UPbxODFRNR/XUPxeBmRVOQtDs0Dfu
CQ/2hzGpShB1Z9ZsYGRsi9KLwYuiGPnQ8BOoAickzFkOrGF3V+R+IbsM767W/2t5
cJOgyYLfZn7TTNXSrU83do7D4165UFBF/FDd/oFcxxBEbny0w6FvR1Fqwc2dJaUV
A4BYTWRjVId8DBO9/lmnbuRSm+xm0rKHV/VTUDpnZBQNAVYl92fOmyDzY1S8Q6YU
QtgNaIMJ09UQxFdZzDu62eq1sdNBw3TuSiYXg+SEGtXZxPpQpPX05SPCjNHcSVWY
p3L5zreKhwpTRw+N4Z9a9GjDKjjectUb3F5DoJbaJlVA6nd3DHTx1v8NCbgQzpwS
vf1yj0ONzU4d2y+fs+KNVXlPjjgaiPe6i6AmXn3lj/Si4k7RBqXnJVlfFdBai3zC
XKc1LK+r3rvmR17gxCLkzTBdIlIHOIMPT8HNnEXaSqvXZEAXu2VtDcFefwz/r2Ys
EGl9B3wAr9bkByD9LSN1K1zVynZspgZ9onaPSaSymmRUgiekbCHVEpfnJgFVpz6I
83cYOJx3Rytp109aOdzV8h2rTdpcIbigEaAHmh+F/TJe4C87HKwbReabEHXulPyW
Pc+Dk07fvr3eCEpdCqWufAgyS0SVkI4WsAQEHUWytlMxffl0ITheW2RAmmFZupth
S0Qi0U7Hg6XPOAZKF1y/qcS0/tJfJhYvZd45UdA0VVwAglR9edRXS+GIDQibTZng
iV9In+1hIFx9rIr+90IfHt3ijRBM0E6ybk9LkK45J3MqOMQ/AewlnmT12DD2WDj/
9Ct0y7xM+B7fxjKZvTkLTZG+QStfmus1gasyXws5TxxFuB9exfMh3Lb+4xvW5LUf
UOc08BGGKDIKryGDRtZ7iUxRD61EH8qN0UCerHGSRZceaFmmCBvhoEUn0vhexj7J
pZCZmTdufn7BbJ7OlLUJPNobg2ROssWtcewI1zWaB6kByTA/zpX+3CVuxI2zPkfs
YsY0+oSVPhmZSW24fgXxaZDx3jh4fXEFo0Quoyc/Uq1oayTSJ6+oraEWjP9cWPXM
d8d2V0IIt6NDbW9xoSETaKYaCZFSNIyd7jFvg+r02QpWJB4sgIPM9mT+zWW9r+8x
QNVpg5unDeLr3FC3rVdREpCb77RKkMRahNiSjUUieF77K96gtfb8mFdmUNflpnm2
6STzrWjJGA8gO91B9OU/3ruk7QzIwYqUR9tTcbiwAWB63Z5XVgMqaA+g6ujshmAy
iaH8TMk+n1Oex5B9MBo7cg4mAwEZ9dv2RWWXnIKoFDDzbD1g8XaFfGPpZ2KQ5wwq
fj68n/12zaNJqcOU6NMBuhM7IKCjvqqKAxtKHdRcQBnkQfBmS/5FTvXnho4Qcg0i
tZly+41MUx8OEK5UeIGRyF8MULZMIQ7bBE0LSro6/vJUP78YP9+FT4djZ/DefRtp
ehX+pzvDAM1XMsQ92U3OfslNEmMsnVOvijlC41NRJDRiOmFeYFZsxIf3wAu8eGnt
1VYIO/Pq5OBnX5gzeGiMsmtk0l3bonSoMSOXF1qiRVV6OZKOUb7lrimEIa7wHCBK
kfpQeq0lh08byxc4XzjfjIO3jvo6/a3DsbUlOYrvdzWJfOLPpPO4C/cVLGTw1OIN
/6NkNE0ahCW7J4eMhavkmzsy16aoCnMPD4AGyd/1sFv1epplvfcXseYUp1ilDXA5
2kEIqrrO/+UdqwlsgIzoLs4A0YggdArJ39VKHkWxWCy1algUJN5Y8emjIbJqD94M
jRkGGIvHRVencRNfHaPBeSGD6RXWSbY9dn03QQIS0W2e6PCfAvaKw50ZeSYdlmEI
G7epBxnARLpov8EafpvKKksWme1ufu0RUB7javw4WXk4hZITsPAKLw6bGPlZsCyn
y/n6CrPrw8Uk1Mk5QS577PDVwUzyJ1hvTChuOp3hGswfjjOskYqFxCdUicTiNcXg
OfMePhbmnh2y/ZVazOBYjxwydmGV9cXP4YDacTmO+cAD5OfYTBZwDDEbxF5VNRYT
6udsVfnH9loePr1jKuPa8xFxa/9GdArK77f2cEqY3Lyfq0tV9mBM6hy7PBKO4jtt
yeJOOmJwYWEmYro1RjfXIVyvIJPJadqP7yFsUc43Mcq7yty3JeXCV85zY7qdwuXD
rR0kdW0T7QiXPWf+uidvGN4ozHkODJv6T7ao+Evi6Vl/ufZ+2PUl1WNC2q1PDhw9
nzH+k7AySzRs404AGCX3qEOx1mb/SdQzvvg5Hq2zeSB6XbDTRrUQoOzqyB1Gx1Z5
QxOkHJN9WruBYCNH8FZ1eGgKwBRMwi6BW1Il+s5OSZNdoHg4AbFNZCu/tNZ3t/yO
AYCnAGk3hANIzuGkngY5sTSrREM6D5WogCU0lXF/76r1DbayKQJ6VdhTWxfeHdcF
QP3qa1a8SYc9JzzeSNz9iSaG1UJw6i5ueT7rblHfkXn7ysdHhyulWFH0txW3mThy
kVsz1JvAlkKUIUS2pHMSKE9fbbGI5AlIVae5dFbyktG+X6G1wZHVSro39N6IgIzP
emMCDamaPUnE3m9gcilB6d75CrpF6xB81brcWdxgsigs9Dc1fyuIgLOfE1s2d5o7
d5vMIjs/ZvheYnH+yoKIBwPMJxyp5wO7d8O7zR7/25Fy/3u6NTCgccWTkv1nA7oC
8oIzXs2/WOaGW1UtXADhAWQQ/CDGwl0wIFQSsKLUSahXvE8UvklMcSpDQi9EguPG
vh53tvVF971mfqx0JH6RBhdmVhMt7lXbjhkRPYEXIvOFpvYN/u59P4+qn6v/kCye
oqN69FGmhIVEiEB57GYCK6SpVSktTjQlMGRr7Tbn0CpePGs3iGU3InxqRQVLf0ca
W+S1j65ShK3u0C4VI2pHjFaK0U74Cb9CgMeDfyukZu3q/3vlOkF81O8o3dxjGOFG
RqDOiRdHMKspIXda1dIxQsyDQTovWYuIJsFw55tV24cNBot4r3LT5WqJuQDCwzir
0H5gX9gS3DpN3uwx306D9a3Tye0xBk3VmZVx6tzO7yNroSdPaO5AREQESkJeQK2f
0wBL4cCMeylPtfXNcxj0QzI9YCm2IgtBeDPlNvFxhFR7gsfeIg7KMCYNxh86ngi/
+w9UBkD09T9bx/G5YPCwofBUxzePNqKrAkGS1gmORTtvBm88Gex96GW3HMxINmZP
UqYRkkN8kiaAYBCXGK0HWzikZtRjnOuzFVQKceS/86J4i58cKwxcO62l9ysdH6o2
zNiuGHUHO+1LzQDohaU5fSVplfeQxdto+E5+sIauxoruaysXV8xncCO1bbpo2u+s
Fi07Hih8k+YBcKR1mD7Z6dAPQFHRm3dHFdN/FmT4mVG+bRnNUlyQykyY89mR5UaW
ADbokFKRHbfjzXKv9mL1pcFs6gN363whMpXEbJvV4/GVNc0ill++X9VRlO2HCitz
lXsGbSoytkHoyHEZ2MkiPCbs6jyzey6ogV5wB3M9QMo2MEAJfpfZsxb6orBaMHQ9
31FXl2VIyeMfHzhLFvRFzrm9wrdjGepMb2tkWKxtNjPEh9VcKyLasqtfjDVipl0n
8RG5NP/gCTvK0aJruDHIGha8FedKltf5BSxj2SlMvwpklnawc8tg2CN5D5J6J42f
17J3OrKg+4OQ2IZsemcBmG6qJsndX9M5CDjofkAA7fBqthZY6OzytH8OSdW01gls
cuIKJ4n5a2w5VTZ2nmUMQv1595CWmzfMp5aGxjxrk66I0TVxPsWGu9mgK54A9Wxi
RVL843Ew1x/BLFd5rIEESZPov1UY0E1kqv2OL88oAJ7RJtgJF8rGXB0Rp6Hyaoln
K9PiadPDJs5JfjPewkEnMcPqmMvI9mrmhlAXoegl9+3bx3QpIuAq2ysXbEFmkr5d
8EK4SZWiv4xUEjXVQ9jhnRK3EWYMP8X/N29YVxg3vNdL37SI9BTO22Z5NcO9VAbe
AC0HooLVLitiTbx+3J0HUNBbGXq/jmd2Mjr0uMrFa6z6K6iy5zL4dc/Hl4Gos7WB
+PAUSXvZeY1FFh5H3bgf7qeeSryCfqMnEym/IwNq8z04a0r8c0GkSf+MQKWzOJn5
xOOUXIkQ1O1mvafk3Sx7gI+ouJ1GqafKUz5ikStxZzA6+3vKSRDoMfk8CrS2tmQH
cHaVeFbSWKNrG8jSO3cXgqa97W3i1TFzfLXv7w93fizZUPc+WqsfCofkGkgkcvIp
PEW0XUN0eDNiJRk3aco/lVmq0Fs6wstc+MbcXcQDNK/7WdQXcxsGFMJ9wYfsX79k
i/cHEIBIMBzHB1tAhQmaLyMFzRRw1lPl31QGlV9AjQWh+X3QA8qUinE+R6dk4WSl
xrzNymdckautUuvRDY7YQFPSkxz0DX7mxbg+hWq/rXAYv24RXgvFeZHnRueix56F
yX07MTAtIvRFL7KodMWGArIGUua1yz1kr68MsVcpasLBNK6KVhXPMlDfC1omjanb
F7TXAaOzmNg20TWKfIdK/VnsUOe6+ESfsWSUh6G1tAHde92Tfc2GCVs08i83fmQk
hAlBZ9bL+zUilVIpn8rVkAGjpc1y+hqa2utsVsV99un974d0/Zzjpm0XtGF/y5Xm
guqERdT00ibiYQZ7Gj6UNrx9weFpvi6/umRN/qG03TAEoc+iy1I0C+bkLkZQuN88
BRaAWDxshSmp1ZUtcwIvREour1mwysIZgKI426VBaLyXrVEqq7YO3SHCWc97whyc
sICpDJB9ejEVyxxKfFKaWNJaRy5/fmCQKgQBmwOuKj8QGItkEvLWbMY8kNR5927m
ZoWNEPLsbjmHlIV3ZRs87RRFwyKYlRoYv0tv9iRlWkK9ojMk7iVG3qHEmxWpnkxE
NW+baIvh6wFnTTyARr9BEudVi0jOOIlDUlJq4gvxAKosuRb3SIzClGTpu8/FI41Q
MzRrext7DSooBid8+YfSueIrGPfwg85nzzvcVsf6kJQgIbCQBpBZ0GB8K78GUlQa
vzWoj4/loP4+1Mg2yRWE8oi4rO4xz8ARSwMnwsCjJ1HqxOcsK2UOLeUwF8PPN+3b
TAnRPFB5BKBsFDa3xt9XKEgPzLAgCpR13vZRcyOr90k6aghJC0wm2mzOMhMdPLgq
BVA69lgUJmOZsdRI95G2LPiu3b4Y17SrGFpMzSczCkWK/g1ZkodmUxI0ACjbF2OA
rIobGJl+JvGl+dR9CVC1R3A0JL1RzAbIZcrBBWfxNysn1ifGkK2svZ4JOh0LAdtE
t2vNrko9nKwaIEZVszepnlRwEIjR/dJqS/HFfQMHkHHqD9NLJmBurt68N1+eO5US
IyqR7Y8ZnHbOL/bU+feghWX1g0ImejJ3z+6fmn8oN9UfPWlHZJym9qan3W5Bz+Ur
AlTFknfNLMdM8lVwTo90d8BGKMvFzK/5ViinYJt0ULUpF01b4ih7ubPIsvnQLJhl
t0ObR9ZABNNM0Tfe+7ZbFKHdxcVds541jn7qH79aM/f6edpDihmL/Fv0QjoDWuF0
1FtquBezrjgIsmc3Hp0Wc+08HDOMFqND/9N2QEkrwLGcMEG5O3wnWe8PD2Z+mmwn
IcUJ8E1RtSLVEYmVQdJrV8/o3sz1Zhd0Vv9z3zjXy/zGlNd5npkfSCnJX46I1FHQ
HrhJC6ppnTDernEpiLXfQWQimRfuP6kszkIiIQrv/9lBfQt7bp2UO4rsKytjWxRB
2cN1xi5zBkFU1Jc9sc7LkY34FNMnSnnDfsGyf4DYY3fAjhdyDATBAYQ4TDpfIAAU
tkTik+LwuS+F70Z+a7sde6+To6K03iJccemiHMsTVdQnLg5HteNbx7iKrRGvfnvy
CfxEcEfYQCiC91OGG5s6wT0HDLbOpG7XcqxOt/E4rI7A8iukUz9CZgnzvOvWvZe0
hdsHWOzBqXBaW7OKtOAWGmVSyy6kAZA8AgH79nFO34LVBkjoRStt5253E6FZWp2T
x4uDnGcDMRwRGR5j5YHWavbjzudLuqw9ubIOQtcFFFc5T77UcmHsWphJqK4Yt1Vq
0dYS0Yp2aXj1KFIJLfB2sOAsR+xKq15UCBN2WRHoRpROAcjR5uut6x7n3jf8NGiB
jX+2vjTEyGYCU7++tFezaRmQ/kv9rXXbEYTWAhudVzQ2/cRgr67JEY1eKA+2NDSB
gAMTlLZSbZLy3Kw+d190XWO7l9G0JhJ3jpxxPGqYjQT3otheZKX1RGn9CHgMQUJL
DA0+SgMSTFyHzz6bJV2adEfJAas2Nsn3uoAMw5Zn0AxSXE2rZ4IdJnwRGCCKAp1T
GoqSYWbXHiP5eQqY3/OVMSM6Y8FDOh6/rOX7Q8WnYvD6MoV23X9Qa/L51OmUTA1m
zuSgnfgNWY7Hn3XBiqyIsl7GZ/Mab4lr4YWByOf61axApmGnUGIZk/t1DqWlJPQq
CTyDmKUVByq5g65QgD1OOn1C8+eK5SUCamDoYjix1HyjcOH8LJEfhT4rz1D0d2RQ
NcgViPcCVa7LUrghAOXq43yFXx+4LFUytg5dWShltF3p6IpiCtvk+TG1bLAg+M7R
OrDGc2odLSUZk6nSq39FZ9+hziVwNtUXyuGY941uad+bRvdmJINsNAqueE8M+fRs
92O1xUZxVI+r1G9utwIvh3hRcjdMuLOq/3Cr0eCcO1QGCSpb01TG2zVCnrOvoqHd
ljt96Qp3RlajGd1EWfFZ0k6eeGj9/l+EdDt5D4XikwrqzYQWvCby5/lpqbS0LBJC
o+JbGsPNGDyW8QmNbTlufD5bMIRwmW5WM0EEZgmlXdPiAwSmsZOOWHp77k9251CX
zbtCb7Xg19bsnQXavJ+6GUQ3zpf9oSRmC2OU4wQQPd4elRGqnntNvyQzsNQmpruC
e4Q+oNoeM6p0jl+SpxkdWST2zzr3FnnpYy+DkNZqy1yQ0Lp7ERBHMI/Prnvn/Jft
f0CClZAidA5IVontF4wtfZz8lwSH+GeT37E0cACmAet+mwXeym29Ie+q3H+qEKaP
90WpshoB5o3Pv48KeQZ3mTFvi/8mYg7/lRRTeOUcefDNgwA4oUdDGo8Ws6Ydl71R
YMQBBoDkFEEHH/tseUJUWAzCHJMxlFY9/JXudKnXQTQDPF/rFRTYd2g7nPjs/d8e
/D5bKf7vUG5lbXjmYsIUSOd1FgqWFzEmRn52UbDEX4xVm5HxokohVyZjovd9z5zK
2utyOLptrD+JJWHaZfcWbbR/YuUt55fVCXWiivdEVx6/gCWIB2fRix1sjLTYVXYj
MajgRtf011H2srKdrxNPCx0ekMI31YnbZ7/8lrLOE6cHd6G29g6KEiM9e3UC/tPj
1+ItyqP9//tL9B1lfkxW9d522WForNfprevSGMgixM9B/GSfsCP2a8+/lmW/2aPy
gMhH8f/kj94wWmOOxXlABWpEb5PZ5FG8DudJIXUDx5JNkwOgvlD6EQnmxCJdF18/
B1jgYfGTZtlQTKahd0aaLIdnL+Rk+2iJk14xbpevj15I5YI+FDh0viikdivDRASB
7mcYGgFEZTSUEF+2h2XFI6zheM+/HtkeOlBbSun03UuKTgQF8obfVz/GMRdBqmki
kKE9g6c01ysbvtjzs2wbeMvmvR0mjh1le2r6caMgYz8QW7yKXz48gXUV/drgCUyA
y6cqYycCyk4KPFjlE3AnJ/vevlBDslLYT2/isAD6IRxHEZ+TIjuvqzCwImk/dZgG
jbVeRdykw1DLruR9jMfbw9CAVPSF4bDZbSZx2U6vEeeIAgjgC+KsZ2+9t0WHrPXd
CI8GTd7sJmCymT1lnQ6fQ8mD3xFbkVPn4svcB5FjDn9JyZFAn5tdrhugp/SFL+MA
ajNbMWOulyEF8tWmzcGBG12HH9yufg/KsEoXAPQtGF8zia0hi2GaShSxI9Cspnm/
T0YNrd4ywM9lyNq2L+lzjBZTCrgC1+1LkUqQL8z4V3OuY4SUq4LTM16xXCZFtJoE
eGlriNiJqzsXx5QSHK1+Zn8hPqRJ5vb6Ig7RDfg7sLnmogS+x8inWD5QT8lckS3y
02vmF6jateUVhquf99FwdunxN/pUA+jL+pli2d6DTS62J8PJPxVy14hypG26+5ag
DjVDDRfkpwLMYDqQLw2EwzfMqw7Psraq5qmtEX/gLgSvzCYVQmp5EExbl5iHAtL6
7D08Gv8UGvNt2d2tOmM2+s3+teDC7dlCbVKOuD4o2nWyt0vrP8llmS2y+pSLpq2t
UAm9zMe1R24c8hk53SRodPKWcuE1QIkCGVGp5FKi9fe4t/S2VEWJnHSWVG2CUrQK
bezO509TpLzMuedFrznxwGxzA1/D7L1eDkb+HfWnsoUicTuJsJuvQUN/FmyxJFdk
L0ccE9c1TH+7rpu4TLtPYHoyPKJSpKUX1tdfAWczZHveOWgdyFwzyA3p+6OPgf4a
MaFw3HXozPawNKPG/v5ZZ48fBvcTnKYOBbhXEHfUrppmE+2DMWPn/EJEuFV3t+la
vAWWlHkS/jThhCmluB1WX/LkqU/TCDZ8AlQhgOuR8NCinBBcxlOL7+ucgS5deX9U
u4zMLnIT1uw6PEYbN7VsJuhs5zBWhU7WA7YU2DH9lYtk1j9KO8rERfPIGZRyJd+X
HESit4lK0SO1oMHxWoYinR//wLbtrwUoJKRFL8ZRYzrKT+62U5cZDpxJiz5rM4wi
ktL5T5u+Ix8bxcjw7lKq8DZL4f+wdMYJHfkVnaIhoZSwDF8xsVbO2gW3ca931UG3
BPBZyZDvZJT6kbILdjYJopFu3/DArahlQAiMwXmfH+MRaGgNBI7BAHCYaweip0xO
FkCQKWclh1MJ5G1t28yau5Y0jhgNmAiTfalUVVTJf0MWNAWBva2+EEstIraKTxjv
eLKpCgBa3ixMNSorxKW7w3HRKQxopPBwYC7oU/Vx9I3ql0Zd5vAOF7GCHnQyV0fo
lXrohxsvBk3SLeTt5aGrjvSf/reuhO3509qULaPmn3oRTKTVtufeKqr4Xi5i3soM
LJUL+tEAJRn3G/5DiIjFYbOHElTjt+6tBK0oBcGmJ47VKWRLtJFRgWl/qyvBwITb
jPlFeOU2wumMgprBaGMFaoA7ieRdRraAoz+qIKpj+RX6dHTMc5X0B7QpQQnsLPVe
orHuUtr0tC8aiEMEosHK8TRm5pG2CJ9pp0gUUm+vyBh/9a0bf9GK+48nPpv5IZu1
lYHB+1J3U88rmF4oHQeZ6bzt4hl9FdmKcOz8tuijFRrzmCXjm057dB3iO7Qkp03e
sKht487tLSOUEEa9xMvEKbkrX8cyhJM5st+fxHEjvUALoK+lwdPzIMeh3ftFt4I4
iHL3//4gERxmRe9CW6mExKWFuTNQQSsIIOI2XfQ0d5IVQCYEYoP2xNvaE/uFzK6S
mlTJ6W3GnVN/p2t8XD7B4zt0dOQT3kj489D1WSGpFpK20rxuNlC5KHhEsdX4LVYE
mTOmtZ3UNmb9NahXxGLI+U3iEKBLCoM6fqJAnKB6HPGzOGSfJG2I/3XN4M1mAjVN
2LdcRk2s4nkcCNp5aif5aRLcXUIzyaYtkNFdQB6FRuTid9t1Ar6rmg+8DsZ6RZQ1
wMFNumoxp83tRAEm/3UQQqZq0zPtFM3LkYDfsmvSQVm3fo2wI73WfIm59JqF5I2U
Q83t/UpzrnJkMtXm/TnGLiVspRtK5hZIV5uxcaqfwMs2QGCTEeBNrjI0uM00mT3N
P9qBTSXEMN8hgL4/U+NSAuB/W6/8qkUK12IhIYK8VfqzqSXpzhBcJk7M7hakQsGO
m3+v78jL3Rd4rRG6ICwLvz12wl9Dny8Jz1kfnHPs8p0Vr5h3VVYC/GLqtQq2oY8R
kgJhflLCZ4iEQniMUTl9yPU7Mw5y93kTkWs3jvFpUhr9uOKFN+/v2Gvve2+DLDRz
fb2+zltaQjrTNDU8fJxTk+Xyl+bAUPmjiG4vSK8tAffu4critjUD42FxqmzKSRhB
nxelw5Y+rH4ABjmjkd4NXNlDgBkYKPNPsfdN19Z4WMQgaII2GHVQQ/g5/E/zRL/u
Ia6kXV4Bys8+6ZB/+fULisZwXkDkiE+2IM+arwvnrQpnWc0MElu/uP6Dv7SdgNiI
qVnQdQchTcemrMuJCjR0+AjQrGniLuFQAEB0+WxThZiFJTn88L9GqxomiAOgBMAW
PadA4U6EqUi9XHXSxZYFFcJUbchAeeqp4IbMBLpJ/4OSioNi57MxfHrgFksbieTZ
iqA8495T/r5OR1msDhIC42RlhvvmEmoXXNwq4yEpyQJcR5CPLcJRV7v2aA++e8hV
b3BhIfgPTNyEDFzWsUN9iD0a4Ro09+2R9B4b/wry6po8VTJt7CGMuPZ/LHchrAYP
1Xq2f4NQ1Rni7A7+PljtWhXz+6NRsUbhjC4mWsfTmrY7BO0+KSTTjMulSoSETTwb
NpSvYv0c0+dq6mXoSs8RzDTSwm9Uq2AnzjEFXHOKYBsRTweI7YB67KuM78ZiiOBX
xtQB66o+/8DfXVXCCAELdcFZleW3Oko+Ws+gqVBZ0S3KCUDL8lxsUT+MY/6vC9SR
gCCU10i7mvGSUQbhjNnBpmaLHVlPsPJgIDm0q7ntQKrZPCrr+EBqyJXNPuRzp00x
ObC9Kq0WWILgvIWg+kEPlbgMdPrSK7qnwU5jc0OovB18arszhsua4ovzxtRKr7Nx
/QuxHZFnKMVkwqlxOFipFec/l6Tsjw2CSI9XAbWU7nMkaJetTaRu3pkPDCaqxRGo
22cNVouiqE5Opoo1PaPYFLq3HriQ1Z9+SL4ljhWLwZLr+8FpxfA2Px56u2o8bDCA
Yb1sCn3w5GO4In/b0/gMXlZc1/rajMfImEsZOpmrB503vkX2Q8X+bIr9T6nYndgk
6oZu62OyZ32Iv/0wXHo38pNqqSwWhd93FMPB+fxjuR+f2o/QQ2joCIpc6cwBZF4F
x7o859O5MP4tFM/LF1fStx1VC6/X6DbmqK9I2+h6Bm7/D4vjJ5CSOfhn6rM2oV/j
YFUXalGwkfz3fbi+XP5jMUkIMH4oT+7/olO7m8JjPrkwzYZoTm23kv+xxNT0HsxX
yubSfS4ib8WOq60VNh/Eh+PXkUMQfZzWc9embvqj/n+YqnwGuzE0arpcueTfcb1J
EHCsiCOIb1RBBQs6My1L1tP0miYop2vPHsdHp0KAL9kSwYoT1K5HYYgT/SsYF9Et
iadjVmyNOOfHmwAcaGjU456cEvfC891AIvtO1a4EGqOYIDN0iKfBr5lZ28CAGzMh
Kx1GcYZXeMF+9SSuOMEWPSuViZSi0K1RyFEHZXqmlRVPynZCB3TdB3NT7Vl5KHC+
7bbQpU52M2dFght5+tD06I30si3iqJ8Fgsheypjf0w0LWHOEVOu5tW74nGEBUg0C
Ga7HThHnRESnPq412RnAm4jEIBv0KQf5pIuBmJFwnju6xqjaFWZwplOb1qR7Wb+J
uvC1pFf29aRd5u/nmjXnMT0SiiBxYWoWtEhxvyjhEMuumuyLsBqpdRYGR1r4tc/g
pB6v6scgn7ze1XBuez5Mw9uiEAgRCVn1ydFsei1sriZwZ9HYoimQcaOKLBg3AQjE
OF2WwhGKp2oUO0SMFEzCjivfqotKTGOxQ8+ZgNvD7TgYTGirIPJocpcEWrnUarNM
8V4HDl40HNToE6HWAoiZhkHLMa3AGz3zrpCJdFtbIclowmO+PxQ95n3CUBNwb6Lb
vhyXsaznSNq1ysJuEgbnuvJZppoMY/8rkddep+L7WU7WfYtMfzmAL4idxDlB3BXO
Pj5U5H8Lbl7MJ/oqqxNP8+zNSIgGzd6GOMayJwVNjIVEO4lt4/dS7H/0qGC/gv/o
/O1k2OScPcLcop05VVHV/Ea/C4BdU60mPmDXNrIhGlTP0xp7KpkwAK1O9GqTtDB8
Msv84lcAvkDsm9ye8hqL0frFMH4M8CJRde/w7BMeR6pgGSiVglcY++OKoU2UVGJ8
ra5j6SqdAIVKg2OBLcGSMTcsAqEVq4vIAX+fCa3MmI+d3Fde6nPZA9sxwJEZv2Pz
nD28ztVusl+jWvq3gnW7yex/MnOiUn8wzvByJ7dwP6xNBwKF4sgPkVZSVQFtuPFr
Y+cN+1e6O0/j+bxRt3puRCkQnjZ7A7v4pRICGfjflTO9udy3CP0+MsaZVuKVnwF4
qIhrm3o1qQuvAali2HJrJrfDKA86CB4NireZs+rku3AaQxAYaV5OWhvjxBo7zm8H
CdxlrG6ulH4RqOt3Nkqja+SuzHSjL4fRgi/mNb6BHMTxcYvSZHAhRqg5YwqBoD0i
iB+kEcu7xv8WT8I9PrvJgtEHBKir9DsKUOlQjgHSypDvTBt4J6bKHpsJ+inMxuFG
GIe+OgAM0sSq+k+ZvIUhG1wXBm4BRr+2hB9TphMdXv+7vjfEktaRzBGtwCBKX+mU
vvaZKtk7jIbtsxmeHGuxjjy/JPCO/iNemcpBnqFsxoPMqBAmXCop7ebTyjHy8fuQ
g7uA9+mVoK+XxhqVGlnUi3eMCL8wsHfx7QegwoKriQ/tZgWNAhfWjR40EsMDeAIV
cQ5hTchpui5G6O9D95S7bMAB+xvyOBfKo6eD14sBuRHTVZBoWw+MKlTYJsAB8ifc
iM1DZLKhqt5FiUR67hyILLVHKMErw8JaGdqa6D43wa8PgIdWc1aWa4HPIlA+7pA5
d9K42k+FErp4ZHJncZLF/HjLTYGzKQvvZMYK44YOCWqfs1PLaEZabHeOq+sqpuSm
Dt6nuG90OHe9QXh+oVLxx/2zMzzUWdABTXVvJ8FPK6RkQORtlu0u3Ak1DXg5efVG
JF9/l9pM0L+aoywuZ6JHXHBHzvlbVm4xFBGgR1O3nJCNrdmc22rWP/6DLC/Wwq1c
MdfVvO/eFxlxdkuxihfuIeAJd5amalFjqJvJgCgEh7x5uws4xbrQ+ZMBFiznfoKL
HCTfJCtXIwUSR08VJioNsHaN7cbWXCF+fODSTaEVcmK7Mh0OB0gCoUG+efG3uqRA
/69atezBbZwdQMedsFXPXj+d0cmVWysFeK/hfSVxZrI+0+KQOZQPWC4uA+QH6LKk
uwTiFaLiSwU4e3VgoWMkbc/16NlveFW3bwW0bjW1fBHtb5WQHAZVGN1Sgqq2aftN
a22YXFTTrVHqeh1OYmFHZmeZ86l0VAjrCBgRf5c/nAX4kcuQMIeNC7DpHV6IdGq/
u8T8OsV/9RIcXl1m/uOKKpGjikoXegXsL0t2HXjxX8TDS/xF9kyBYQdp/djYjcvH
1wXqzv7fg0XVfaTkBDVuCBxp7uMThSntOL8PG3Rv5CeOf2ixiBGw4F7i3KY8axAF
VJ+hm7OF+gJ1IgQG4EWRyiXhBiHBLhdPpr/Ydnn1VJZu5yA4w5Dxb/z1SdeUSw7Z
wWV3WPXvVcv2sPsy98HweaDVCkRnNUKFOFsT8mCOwIhvh34r7aGuebEZudXMErYz
1FxJRJf0dIZiAQ3xK5stQ34sKuvTRvolXtkRemSliCaNVM8cjijyz638VJvyuPBD
b5cwawJHFpGGKl0Weh4Mgh6bxvX/ZFjeYv+JzTZuW3VqeifCCEIW9QSGbB0EOJ7S
Uy4eMh4f05Lo/yIwXivuXs2TehpPkiARNM1qv0XQylWlx8O0qFPdk+JeTK+hhrRt
kD34XSnVDVDTqllZLPO7M1gDwAvW6+yORyQ5uzlT2l17RKwXqI3iTlvmSpu/PWAL
RmM/mGDRtYM8OAJ3pSpi+inJkURr7RQc4Pa/4SE5WG6iDaCf97oyzwn8nhBfEhKh
tWXXeBIAlX9/ZekuVOlpBs5AK3V6WfON+Eq0uTyQ2ULfPuB8ymuSjRlVHvmb4ArA
m0/2xHC5G2YgV0q8miKP3LecbMrB5c1LeVFThOYk3mqZ7qTpxL/uGYji7ijBpF7+
c/dD0JhciEHtl0sAGFqb/GbQfV8nbDP7zPlwv69QTni5PhFh4t9i28GFuYGQjkJ8
MdM7jAK9KBVFdAy+Ty1b6cZxjHCilSWtaIBs9Pc0CHjWVrEO/oGzXxzivZEgiVA6
9cMYrY2o3F811Vogbki0tCrEn9/9POYijemozyLoMRDzyy4yB00cnDUgjo9xYrvz
gGC6aokIJRZ5ScyHip6JjQ1Bfth+QwKMQo91OPXMC9k7kUhFGE0Y7o7Baf2JGQ53
l6DFakxAHycj6c4LM0oaHpZa7BfL8n7ZCoN2xvKtAXVN+r2qOjyW97TEshLXmYJN
dHQ0DjpNPNg7YTE1Z9kbM9s7pGuJswuaYqmPuvtE2RRh2JuLyjb0M3qmUl7cbA5S
vxV6MS/82/BLBoxGs7xnoHDiLKnqRzd18G4qdOwEyzW0NRbgCDVbc4aP3DZqPQsD
NPAqt7hoGFTWzYMY5UH843RuiFsT82NdS9GGU2xUPKoD7PRm60vMLrgaruBfg39H
5/QgLiMl3G7fq+xrdRXJdxBHMRqt2K+HU7wHwa3fOjD88ae/6R93HBP2I1Cr0/vH
TSBTdC3TDRzk9ft1bDKlcCBkxvmNc9HprD1PQyqmSWFXnv7oCPVVQSLHV2LRMs3Z
2lLOt+XHjx50mqTs4GMvqzrSsP69O/luepHKZX8Bw1bW12q2OX2QbO/BrDRhwrN9
4KTqUghUDS8/SctAONxNMec2EYcZcqng2XE5LOKd3Fqgmzr9o6ORsWHxYnRi+JZW
Xhk/Qpl7ivgfQy5vgTttXZtPILpacqW+LFFRY+wC45iqUngNZVboU5tW8c2ZDuKF
OSUs6W23Hs8FB/CAleaiWfO/Lzjw9EaT00XlgJP3lQoukC4Jmsq1kRwfWhqmfdhr
iGdk6xs0Rb4Xlz9JXWLNdXe1lVpC518FP6yd4mG97Jv8+ntj0EE8D7eNV/qN4/oG
fJLmOY70a0WurR6jHNnp8yf1DqxNl7ixHZH0+PYUQqFrQ/cvhqDRviTuY7XH/LHa
LwEml3/1LadJq3VcYgNsslBvtB2cn5SbnaGqz1cymDQjfN3hDeZFVdr0Y4gncOEB
5ii3sXcWlKSsUNbcG+/Hrnk0j/gEJGkn7GzYmPLhoqPE+H625EVvN9U+W//o2CO4
eqZfnbQGAApsfNV8SfTM5BSv19ZyjpIBYF2KudqVPm9Y9Wom0J3weCzWT0xKU9hL
glZBE6Bvt7cEZ+YFS6Vl3GtTLwPzDciNVJhYUe3oAnD9JCyuniMkedW4CPcQtF7W
XcfNFJqTkmKiYqp9kRD2Ojtd0wcnTf7Vjat4z33187gqRv7jV9dLHDRU5MpRlyVf
O1VqcV2jeGZq2tm5Db/QOR0Vdgo0N3RXIc9Sjs1fH8oJ3r7X4WhAidh/aYa8TbgA
X75iXhZ15lXn39wkY/9vSBqlV0VGUACkMHxmj//1ImmWNCUAp9OQplJNkgP2rAXF
l+bUcJbJe/cLRDIc2klHPtmvjnBoiz44ylC5Dzm12DpdpSw+VUpzHVd2LGRTkwFc
6sqxvLXkIRRq+TPU8k15ADewCz+lls8ORTOL0MM7QGsW+d1mKrZPGXppKJrNyieg
0cH6bsXM/F6r1pic5sE0DK3cMtA+P4eJFthk3CZ5pcW8seZYMLbE3cH4ZYZswXEb
3AYYb00i9mGetWgvu5ja0au2BJyiOGWB9vEJZTTFxz3nk8QGRRO2kn8Jai9VEKJO
FWuR2whI6rjols6frVLAn3QpA/oI8mlTrKjivd2VuLU/luUa7o0GeaLNqShrcuhY
Lp3Xw4RvoZQ8ZBtsJnZS4E0XCocAc+dEDgqWR6/WfzKprUpqONrchxsKlxyO+cJ+
9SbZsl5qTOoYSsXW4iT6ldeUxkI3l5WgcVM+sEZ0PUdffp4FrD9mHAEcYL+VkR77
BJcSf1Pc1WnGlQ379nAbddIJSL2PdCiPe1U4e+ny2piikX6M+yS97X9UUxkdYxTP
ROchi2lCBQ9yUNjq+NjWvTTDWrQdYfDQWz4RzIPAbdE+z2Jy1qTJ0dtU1fC54Zn3
z4KryMT/oW2GGGwg0/G8NJnArFu3iMxGyZc7bOnxY7/ORb00CoPI7+ltWxwepi33
ZQOhFuPayTZWcRT6xxzmc40bT5HtYQts3XYtCLjNJkGVWnz6ER0sdg2jExlxiJgj
Iu+BTZRSuoR0J2BjUbSGnUeVWhmgpBekdHO1Eed/p8Z3W2ZwATCE+hg2PxwD67nm
r7WtblhSj/XWz8BwDJNcxMcUY7HwzFaAki54SDx97vFG3SCO8sTY92TzS0Vt6M8z
HdrwejDwFCCFMsboi8Fp2i3LkGwMTgyVXRcxh4LUZcTStWvtFlYV9ZYzvUjaDvLD
FpIgY33NQJTpDA1CRHnTY8xzJ9FnB5pDNNu1Y+KAX9RZwsULChltOYlP6LKzt0qF
iUCPtgAQpgp0a1qxfHGPYBJa1likeISiPpfE5gpeU22B1iymctCzo50L33QJglPY
8glpcm87u/JiwxSJ0oFoSw7QF6elcNzx1X05xWtG38GchmZAXK9cKEclmRJTl8j1
5tcwNBAEs2+d7usFN8OzUzac6ztvW2gm+K3ZrG8fX+10kRLflkhbbZr0fH/j+ptK
3gV+24ShTXz9AxSE7JvWMbPYvGo1laQwSe0cIHD59GxwCX2TCi7q4VkY6nJJvONU
zHEp1KtrK3PJlP4QV8DovcAw3Jwq2S2DXVWJKWjj38YbCwJRPrOwz29nAPyszItO
qsK6073QYBRqpj5NVHnGoRL7HCWU3vAzrgEreUfOZOTLrs0oUVOlq0joT38TT0Jz
2lW6Cqm/SCpYFo0y0z/tc1W/x6UTZkl7bMPZu6jnjBmGBZYmAwINsRTaVcNCHyU2
KApNlkMp3rsZVNlHW+RmhixZ4mPrljcKyalMajiq1krBxzK8UnaC9FxoMyNeYelj
7dytpx4TDj+ZGOOYS3lWNoQopq5xT+mqglIa8Eg5B7Gd0XAZMa/YD4+jwH3VIgas
ouzW/6hEKs6lyvVw5d/+muSaXlV18YrqSP7z7vOPZIVr6d/GGXhsbPIwvpmf+ze5
hqbTUYj0pDnmZutubKlO/xg9bx7SI4XDy0JiTcdcaNrYE+XGgMPANR8c320BueVp
iwZUM62mQVSRlcyu3UmG43aSQGiveY2U1iyVmynxD7KjNme4lMZqdqTTzfp2b0Je
nCCkqBfkTsD1elL7J1xH4vvYYTlxYYK6wgfPxYDPHTZ4ZNq3ieIv/JeWfMtUxZ+E
vaeeJixnX1CqVyZ7gB/BRbXT2CtxRI85gV/VRH5Sg212B+I2PTWm69Mxkb7BqY3K
rU5dFnvimVJwF67JI73dnhhskVS3tvJqfmRdYwnVWnhUhPz9qoipCpgiVE5mIb6q
smvzo8vExHuP922muryLQST0ix08ZOvb4qi40/h1BaKQn3/yxb9GRD/YIBocoyKI
/jX9R0LRnQql6V0FGnrRRChGIdLAHErbOdoHKhm+2E4YLuTlo/Ukq9+GdcvMiVu5
wtEgH1OasSz4xNJjuxP/iMSNIE/L+RT0KAot8JYvlema3YnKh20CpXm6Qo9BuGuJ
SKH49jZ41ZaYUQyPMQfwzmZCqfEaXLIcELdpuhy8IQwkbN3Tuq59LuThfs/d7PA4
u3bxzLjR5hVLl0N+C7VRL6WDMarfOvw/wmZWMjFUVmmbZ/j7nRSdJEwpZ2Q2hwLJ
2rzC6lfjAQ8nKuInoZZHOGwT1Mm3cJdYpxr/rjDveKUlEVz4ZvoQVm42znZPnq+c
3vD5Xq/y0aVZ3S7vpAix3QFlxv+CD5LKAh2jx3cx6+kyO6WVowuqKsZxi4momJWX
VEKCTB5UM4/OeMO8DMf6tcX3RzNaathIuaRHGNyERv2mmkHp2EDZo2H53vJPcJsy
L5qfVh/NPFH1eq5FBWDeOONGNYcv9zVnCtBiNcCPzrgGX/SwjCTDO5L6jrKBXLoj
VObcTWVelvkc6Bdke5bIwVKGWEPtlc6WGrZX2QwuMg7pIWmcVwJurToUY9uJUFeJ
1YSwZgQl9N+CxQkPaPjwsau1lZ32r3RmmSIIHNOIpJED/F2YKJgezDGugIDRjGaf
R+VhKEMff9rhFcnykABF8M4Phr/n0og+obp7FkLAh8H+Z/lLGEdSpAh2QLRltCJY
l9Zoor4jaRknkQR3FKxOEMc3c4D2gu/kv+f5lbe+aBH4wruc8X+Sx0PTAoIu01s3
S+EuA2QBL5SYjI3layRIvONxNSQwOHFEsKacO8NhIUbmzCGibZHhxfA8QDG5Gryi
TSE+VUBS4h0NLc5+MdQEH+EG83UtQ/yLrTAU8ucO5r9Tm7GH1DqWEzp7kINy8AUx
HsvYwotI3ceNaVcUpWmOo8j+RTyVeZRcG849cU3M8kpZVAdvGSut5u/6sy4RCuUa
hEYmMm4v4aRsJKv/C4H2Ud9cwNGJ2hAxqwIq/ZQ13h5fEv5n+JZbtgCFhYDBgaW4
jv4r41s53RBDWjIr3DmFzFd7pjtVJXwsnPL8qoUkPdKA9FVK5fh6LCzYhoxIO77/
CUEijK5jsR6kHTnE8DRDnj4clJYKm8zrfoyDS7Y+5b5iRSvBDDZ0kOcSpwosIuTM
R7c6yx96+DgOsFjCYvUC1qZwtzokdv6bb++sJlcIeG0i5E64I+JwRkOX5d3FcQXi
PV0A3BM1rBL7SBKsaxOFxkLVR20RaMXPsH0I/BAY8g6Vc75BCsea7pbD40vxQaPG
XOjynW4UlJr3vfpPiQGuZhRfbhtHt/1nd2f6/fwqZMl4eJSHfS3BakKZiX9r5j6T
T+SzaXQZbFBH4iGWOmUs1nR3yej841+FttavGi5uwVg=
`pragma protect end_protected
