module calcRay(
	input clk,
	input reset,
	
	input [7:0] x,
	input [7:0] y,
	output [7:0] r
);

endmodule