`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
M+Nq2gz+i0JIspMQKZsr0dEqIWdHYv+Tsm1EHLuAMzCy72zc8yVL1AL9uyPREgTs
YPrnP5tfH79Ar5aojJDueDgINhm2WGz325XaPQLFqmbKHiaV2VMcMtFbkDdqmkaa
Mf6DCiKVCwLiyR5Ft6QbGhkza/A7sVm9l0lC3KtVnSc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
xnuOeIMYPIDBba2IHx4vikuUtAdXkxltYryI/e8yI86BebVU/qhOcCXwJ38tVMTC
c2L8ZUZEdbH/jiTnMnKUgIdnHcnzkQoXkOua3dGG0EFfmmJx7j1EeLUOj1KjPsTz
/Z+y2tbRWqLWcdHmEgZIAkdQfFIedKPZCEJ9dRlGGhcNttb9iExXd5THWGPGSl1b
gMBeUF9HQi0WlpsyJex+dB21/yF1fBBBK/e6OPqkWgx5zt0kDee31VZ3ZhdQv9IM
j+eIqruBlUvih6mzl0g78L2G7iG+fegBLWyll/5lboeQ/9A/8K9npgZuk9+ycrMT
H1Mr4ZPp0b7Mn8dJJRXCXdxPTleTV2xktWpujvCNGDRe8ia5NOkijA9Xq50CVI+D
AEWRoYsac29MslTTujU5LvxdVzg3CwqKj98rtsoM+qz2WpfG6S1GZ6Tpv+LOGbZ2
SXUp6cV6bQPy0mDEI6c8BH6pwXLU38SPSbihw07FsWn7zeb2Fr8bq4VbYi0/G5gs
mYZ5C2TGRlICPg2fj3qKjXeX2HS1yPw9UkzwU7rvaRL1HdzCh1DSREgM1173LGHH
EmGrPXFsQ6/YNTx5pHXmUXDEDKJSfBosSE5QW7Vm+WVXe7qHvgwOBi/gKChY1xPC
068Dlypx/WDno4DUDpRvraDw8ayXDyTpkhpClfNf9oSnsNyxThjuzm/UcBhInsxy
u4knpmcjToUPv2IF2dMix2aQe0XHB+9ulaEabN5ccLa3oC14Hu8aQKLMIf6kPkjk
6TEZjnz+hR+YVlYNLmo8X3VOm6p05TNu8vpT+YUYxRsowV7AwKokV6uvcQDkW7rl
HLzMZoYPKdY7w/OBDrjXv1PSo4OzP4uQgVeOiyUx8NT6YNw+YC2IcVbUtXXr7+CV
dNGhkh1nlHlu/LHILjdYLBhx4NrPS1ZABs9dz0Nw/0//SpygjxvKgGzn9MMxgzZG
1geuagWNgS2W+RXzarW3zdy0Np/9BFdpzN3eKRgwn5AbJng7MV+Keeq7GwAVQT6M
XjBvF43qIGNEXfqbfbUyWopLVTuzrE6L3gNXmRfMlhyLcSMrFyvI8CnJ+lNOnu69
vx93HeqNwbViniqAQff4fkXBD70swn0TloJSorntbXBDaDaRzE9tfaOg/J5mb0az
bwTNFaHc3QiSS7NbHgHPsG1DDBOU2A/E6rGidRgRdyKWiCMEVgt3R0tJfAQ6fhlK
sHC8Y36tplYmm4BMxWKmmJZoMHSIRDm2234L3Sy6ZANmIxHPdIquFqyIVz5dAKJu
wJqCQ+eHvdrgukeDQ4D5N1COJpLHNICArQr2s0qnk8z1UGE71mKC7fQ5+fHybW/I
K4FWX2B2OD4k0V8liM9htaPXj9cyPVMjh7Fi1YzB12O8nlCVZqlbkePdLTyiH5JW
JbnNrhcku8rYqqGyQ3sF/hc0q7eLhgWt9AkhiqDNaUFloy0egsYlpeXoY7EHfwgD
iK/+z5+3IMwMyiuP6xoLW6H42TLvv5P1OhEw0Svlrap7zsLGywabwMv/3LC0XeO5
Q6FQnc46rESf2aj10PHBdC3KOmXfqNdFlitrHGT8ok+1lhhcQBAmu0NSK0mAn7Da
nzL15Og2xdKbsEAWQTH0Nd1B/8fkUcuz8S5CgRLf9A7ZwhEKme8CAJtrO35vkXbB
UFpZMqz7jRm9vP9daWCZMgtBKKY9QI6rj7kpvtjMzvg938jQB55OipdzzNIqubN2
g+0b0F6LMztPn9I1k0vhdyCKh+rewmsD0H+Gcee63G0jkRa6hSKUTSrExre4Fsx6
RHNhgJLwkULMiBeAbGJecMDQMDPCjDgcqUtz0LIj88z/cOjmPUP9Hz+xnQw84plj
YhgxwaqBWHdvApgCXT/s4FTXFm1rZ3ZkTXHrHLdLKvLeY+W7cJ1/BoYTjXNsKoqa
3uj7jumptdPVcL7Ed764iEUco/SWMdDKMWrXJGGSb80yA8q7KE6matqZY4uXf6fw
zOEwEBnPvPWx0AKFmBFmt6YQ4R4V4W8TKSRQcDvW0i9wfpFFlRdwGrhgYdggADbk
iyFdfp+T/je4vVUvk4Lrev4d+xKqvLBVFjO3JZtXPsPdUqnu45IAhz6LLCQD4MDf
ceAuyr0vQBlXaf0ocSV9zFxvmjei4E3TLQvZAUkzv24eDVmEz+xJqC/TUw15CbeN
VtNJxZ7nmLhRpiMCDKn0J7AE2vMrXgyXpkRfnR5DFnSkgr+h0WT/FvMtf1DbH5l1
NaobJQVOYLFiyMVpMLnCmUBtVxxYV0WC+DEPNxSzaD4MkPnmd6ZrdSs4EZOjJUH0
fFVRu9geBmUxLxWoyebOdSUO4xnuN9Aivv8VV4mExDMqeyu9QVa0npcDG1noHHWS
8RC05lewq06yU3Trg7YB2HpzYHnlxh75kjPBgtq4/1cF9V8KNrR+FI3AMbLD2R9H
iVhfSKxxnZDRcayo6qWsIMqDt2jJsOYQ1ieoxqfsuzPktt9pgP4SC+aF7eTiyMu/
UkoMpNhXUpOEJui0LNNdxIKpInscxKTNWHxL/I+LxCATSfRC/ou43D8sPl8Kwv1l
BtJ0HE6EG0Nxdt3sY/x3n9VGpGploZ6a0mEBK/gScD14Tx99gQsC82LfdYH2paPD
pP4ald/dQ0J1Z2eAXv171CUJG8PWYR7wDgF9YVdFTE/aG8icdw0gstdYnPQAD4WC
ZJFd9cPfAtPmpiw+NXj0mIrflBE2xd2T1Dmp5dW8Yd2smE/fzh0BMNZ4Z8oF5KzZ
BF+tl4aZ7W21z4qpibBm161vh/gVYL2NF+UYwZLfI599UK/HddTDlpaVpnMzybIh
Wm1PaDLC5Fbu5jNNaAx3IisEjp/vkCipctqrOOH/VrVt+jEi29U7+LsysOnNHFh1
sbkt+BT7j4lP9/ZZ+T+IXJjp60iIcBbBpl/DsD5Q8RwfSFRh0Pd7zqBqtgYbXX6/
syP9PrW207l7rvmyiek+xS5Z/fcYrD2VMyxLKVzI/RGhpjVTHl8MxshqwXVTqybQ
Xvnny+l/YO4e74/IxwPBk3VvBMHlvlHPX4djIXrEG+4ml2MWEZxPwxpVdtVOp06V
p9dxGJkaEvETUwzSpYsLA80xWFBhGnzB5qF09FMKSixFkjPivilxyf4xAyewoqXD
ClE71AcjR0sTfhTX/E7qgjIJl9j5nQ4iIL1uoBJg+JJYTw91HTyZJ67JtcdeflGG
Fkp0IYSKrdLbeyKVYPVnhefutv/UIfzzMfDXFXaDUaq1/sNAWk3E8DRfIvb2vQeG
pPYCf0o89WHdQLiK5lNAoAW8fpSsoMs61heb+uADUpdLxcedt8rM2jyhh0y7VzYJ
FlO6y3SpIXX8KrmiYi+k23V8FvZWYqSPE7COALlx1h3f8E+iIg/Im7kyT3Q14Sd2
xmlaEEd13u1pXDhRh4W6dvpq46zTLYJpQy8FrtTAQ+/bxUCpdsCre5jnfbWTVGFm
Cz9q1uFtifp4HxxZCatNS2mzqHxEOepvTw7aTcRaEfP4Lcm/1IG84kGVsI80J7D8
ZHFRcOCNELlg4PBMb8vAtGzzeuufGLSWA6Ga8C5YpU5eNeNgFs2YI1Iip5VvVJvL
zubGuQTdp7a4kF2T9Pzn5sm8Rhks5vr10g99+/t2rNysN/gJtn5wuhUZ5v1lkj4V
1wQriBhHIpWmf2u1ooAFfCYynG4gc30NVxrNj6KanTPW6DbgQBCm00zrrpmVinJW
y4QGysVY+RWAwuv/pT7TcNful6VuZnZu2RTuGxBdcInBZjc+bn0dEv3ji8ZcY1O/
iCfD/yJ8cs6fUQx4NoUGLmSDR44vrHiePL/7FN1DqQfw61Htz3LwSX26S7PYEYh2
+2NkaKqX73cxhlMgbOQdFtKXJl5Lm/R8JaPfJAdmfWlLB1WSybmOH0JeKBJkvlQe
7Wg26ItnewCQxt/ih7byWDvosB6nkSpJkedo31qt2T48d9uejTX3y9jjigMJOP1L
4wRy9EvhDgmrJBMSEmcI02FD8tyH6GpP72A8SZGv79Biy6g29uxlg6RYN54uMGpi
NUpzQzkiQ+7Kv7N7tN6iN7wiZxVTZaiigXj6hHbftnzmYcpDmL3s8VSTYcqU9rXB
3cpApmpxdRmY3LZ7DtlDXqW9DC9IIm7HZDPeWCf7iE4IC3hC/v2clgkJsguxnjnL
spgOD/r5mY5TKmVA3z/7ifbnC1vQlWceFVQxzmW4Rk09pjYj9KoEB2gQ9ikXGpwg
NJBCO8p2SGw4k51Qub7kw4LFCHNghmq/7bdk7qyKK3hhnJOfyJFhq7AOJe5Ejp1S
/33j/BqGuqkIu+N0fbBChqxW97FtuENelb0+lKMZuMjX5WC+R3hX7XySpv2L5uID
jisGA0/cg5gBBxpzIrT1qlgQQORgKNe+781wFSzErj1dKdvGVQdr7+oNr0SWzgbx
iDQ3RVmafx66QMh8thqlew+YRBrTARpB7pQnDOBJw+WXuSmCybgwUKDwTnnG+Qw7
gy+irFu2UMRbcgpMqMe8uSvOs1cJclEVOSeXpE3y0XSqdbzJ02YbVq7mdxf0+iQ8
oAgNNQ/r2CWeRn9Qq25FPPugXImynb07tBfAc8YWZVSWhMv60PIVw3s7owAST+0L
XkDuzCaHEaEoFTOWzJULFPuVlvyQ7Nh7XdXeWJfAdp/YlJSm4/5ko7Ysx+m4kHlV
JCgFX1JROtgzMnG8yZk0AMeRMqlNAoL85UBenxoArY6K3CQq/noclOizY/2CYY25
mCaYjwqCG4kuCEV/xJncUtwiUcgyB3oSs1PPG4n3lasL3jx5IJOD5G5hDVSMQBor
Jy9eg71swSJSzq0ofDbCxu0XW9hpmJc67gj7o5rR2X0W4hluckltqmCYEBblyeFR
GHiTcxMS4llL1roKyc8GsdkCNzU+wuAtPunX9PD656ZSS4PS81FM1nKKLMBi/EeI
p4HlxxOCyjpd+5xcRmhMNbU+896SO+ZNMGtaV3jbl6h4BTi1LtBiURsAwcY5JW8A
pX46fe8bUAy0hHBd1siVgTvp5qinx+D8LAtezFoQho3Z8hrV8HHiIdwaEnrJq3wI
lgAJx6OaAVA2t+QF/aHHU1T6I5UyLnOX0mIlfDq787Fx38zAjGnVe0USdmLx7oQC
++7FQ0TFPmZ0QZVfpZvj/O0dk8h03rnY38QiY6DjfE3c4xbIuyYyDhy4h4Our2pP
FFCUgTvAIIAu0H5QI6tYJD77oLNmvQgpocxuLI9moyuDuQnjt5OXqZzB4LnwSK36
RAvGBjKdg3d8ebCfDDuhF51F5tmuc8r4ZWPG96I36pqKHmowjh3AzYPy6TzrDSa4
Ka+ObORHR9u6Z7wLBHxx/Uf7z0KrRDuI5VHKfBYPstBVNcfNy3YLDmH6D0QJsLiE
u+z+vX7V/VYKFtgjeTXb0X1+y+zEKquC0q7anEVIR/3RyDekKBXccuQ5rs/3OyCf
O74uOcR6c9/KD4K2P7SgGP1ONb+7L5y59njHI27+YsLVxgzUloM7Kzety77g0itE
cj3m4cdxubPFLymBQr1cAF+MkBe+HRTHofbaiPmP2RkioSjli2c/ab4LPDaYh9PF
O8oxkDQDM5vbSublnjtCcFzymCtFx+p6GNN1xYw8U5KTUQ7zxfilsmTbTJujcB+1
jnv02GAfLlahBevONII3nRxpiLStFkjUltrUHQxxdOxzkj/AvTe/ceIf2kFHmaoj
JODD0oRHfl5zKXV1MUTT2Wts18MSPkt4tsNuW26Khwdgb1GpLrXsoznJVCWJEeK4
zMvxztDwquSN+3Sn27IPMB/3n+dJrvnp/Wat33Nff6X5P1e+KqDY2M2SsCV0hAXd
ZytrpYevEG1Bad95MFvRhdsuz9JX4Dl712wwBZM821Nw6aw0b9DJ1NJtGoGnU4oQ
eRIJW/EHl6ARkn3B7R+IH5+YkaVx6kWxKt1VhhBCsxWpZc4hCxI1OAo06VmLxGMA
xvp/Jnx+3YWwCdFI8Rq0TttopYAuhOft1jwyTuXWvDAJjDvJ71HhFCf+xTiba5Fr
5ff52zs3M/UHl2pKqFXdZjK2gl0ZNlqXtTp9tOM4gK8HjmtAwr9EZn4Nuw3iUamW
np33nJcChKC7/NPdfQKXy3gN+dAalDysBaH9Iehe70jHDVdFn0DXl2KqAkpfoVgX
VR3iVJ6/YSa3CcujfPUrYKqz4q3NakqlfdMKslxRBHefJyLmuErxWmGdFIJSfXFL
BGHhkwGzgyfHIWv963G1ZWguh0GRlTssLsG1OaVum0AY8Qv9TPWuDT1nZrSl/oHl
K7+mhGoq+E34tGbkAnhikk/kzriGhZB5cL8HZxrG4S+lp1gsOeb8ls41QQSLoc0d
oz6zgjh8ici7pEcqkvcGucFpyUbutws54NLj8MQiIBMKSVpWC+M2nhI6nXQHmQc/
Wpql4Rl+dGKilgNFPs4qr7cnxmv3BcBCnElXjnNKy1GTmx9xt0fCu/Ihw97vWL7r
XgwV/3DK6yzGAcsSpl9LCiUpCyfdfXy6paaoz2e7m3lGOVlaxP4+hVZYcK3AAxM2
OVNyG+QDPYAbVe7vMdluWMPt++Ss2GDrAj1SLlnJ3LrQzEgI8mg0S6Od/RDzK9v/
q5CgtcSgU9XasuDZ7R2xdfJw8qwQPlUEI2zae/uqIQpwM87InRQ6HkuRt17qWGyV
656n2OvKII44/YIy5uY+WhcUmyxvkCvGJmWP6KQ/m+n17IlqA51mydSVcNWAK6WM
Vm8GMbTPkr6qwN6LHPLDlIwMRBR8iwB+GxNrWm27bZiNFlu30rP+vp1V76amCWcF
2HSgAE5V5aN5IPYBzaW/G22gMb+7iBK39X76KgLtvY2YK3TzEsF72j68bCBL0Q2b
RZrt75nkUY9U/cU286R31+S34Cv2xHFEXXYN8c/jJqhV0SiHVhRpssgA7gA4l7FA
irs8piBCuCGSp22mlJOvLQhRq2HkduqNulTOnGJwQh9cYooII7FM+bMMn17e7hkL
tVdoUZXtf7VOowm4riZamjMBOIDhsWmqIcz4TvSUhM6tQUOFonQo1ken2lfc2T2o
+kwiBTjPacBKuQg9PLYQ4pKyfvOOIEPgB09tWyXl8gXVRoWnxvShhgJAMys7Am77
PvEJIzk7Zho5I1EQMGyQcDmLIdp1iBS+YFZyGh5HOJ9nMVnGTpi9Bfr73FIPGTwL
Q9byhmTSfRAtbWVcdqf5+BwoUW5tWZTjE6tUSrGrEIxjtqVYuJmzhdwqJedhbGVQ
BpGE+vLuETMz/wMmPofveRhfoEk+AXm8cSxs7Aq+GtVBH1eKm2816t2xPcYtNoO0
zzfn0BYS13ZVgGweyHNIpn0WY3R2kub9m0MpLUHQBcsOXUnKUsA6At6uFzWi6XQ9
QR+e/1dpWIT2ZOWhX9d+zZtiEfQO3zrYn7JmqmPU8zduyMK0O7ptFR/hn3KArSFi
czVbswDMff4PE83xd2l1tCj1qTwGlgBcTzKBALKLXX3qjsPBrppsNkxiiherXaf6
mkLMSYqzkkp3oq4FsVhB+OxJZ9NfOSv3Tt6bDoxUyJtLrajG1k+KYtf3z9Gn1XxA
4AClGs8cYbLRhSo27eO4f/9ItPfgIP//AyoXFeydIsw7dVyeJcTh+x2iglI/+R96
/o+z/OsHCY3KM1ykX4LJmbCAhby8cOIeNIduSVaDqoG/2DQltcNZt2EfbZIiHnV2
zESBGijsO0TsKdWLdlpm6onQS4QGLUCKjLQHHu+eM3BbfZrXTNMgvnoFv5ghjEUe
29v2rkZWp1TRxi+Y6rlEhDle9SgEvK2WmcAa1DC/ww7VyooVvDgrrWAWojLGPQHz
LiePt5mOPB4jR+/bn0AmSvVcMmyg6QPuzbMdDqkLIS/lLUDK1opTRnZhfNkL1KDc
uaaDVaXWY5qGGbm6o00duBvnIVVOb6+MvlSQTKeaWTCppUWit3wybqpT6Xh1v7Pk
r/1vTB93onx8ez402K2e7KG7Ni/CX/V3Nk3LqqUgmi8oMQkGE4yUrcE5ZrjoQO1s
q1igl2sm7tUbGYbh7OJ7/GZl3xe6YDAmyyQTFFi43gSYnXQLm8FSvMi/MRWzCA/0
GWHUXijEqMJysIoQkpSwU+j/iYHTr6EV73nCGC0tWygXJ9KgBmDpu/8PhZHc/AXk
GXNQfBm2/xGq2WoyCz/f5F/a9/QqXQ6VwmPmPX5WlR4th4sdXODdkFTTd5XQsdx4
/5McXTsTRI4F7HXLgVH2rEkww+5qLeolu1Khs1pam2NyiA7CJZyziQ4Wdhytl5vl
x+94eA56nYOitd6FB0sH/LA1DLD+PubBlRy6gpZC+q1doWx4f56Rg2Y5xD0mQlJi
81irMleI98c7I5Hlu4X3G4DgByoXdTydYyXIirbteiRukv667/YpzDsHpWFeNIuP
bDm6sXR4rzL+A26PcYnPG+/w71D40hkBtK3Xta6FCiLD0pQsJMsrtEpOKoHr8iDe
PMC+DFl30SA8rhkhgC6zZCCX38znn7FYtpBKFAGCqTBxuvVX2ug69jNvr1+9i7db
aO0o+rssZSWPZQ70symFMbGW2IViHqgC/kUp197EZ6z9bm94jV4C11bqKKIYCFSo
ZkFnVytYlEQ/L4Gk+N1MlpKSmTUKBL5nBESluaLR/s29hcyLT21pB0nh0SHabxXM
9FL+a4/5huC1aVNrLwk9j6jX7SKaMd7p8ms9mcZKNeWpU2YCr4FOsZ2348uKIU5U
yQRxn6n4p/M/tHIbcehO2bVFzD3bgcLfuAL5AqsK0ikp1KMXJv4pEd1LifivuKSL
93MsT0efOvbhepGwCGujYtblu/YwVL2IQOlwDCnXB/YZJWqQOmG579YljNdkE89L
637K6IdMaeLx1C7oOtVZkp38PtLWodQ0Xnm4yqxR++Zw5Iwkje9odED3FMpppZKv
n02dYXOc8qDP4U0PDsJF/Kb+upyQcRcZHZxMPU79TTEFbaaoX5ZZQ1/NHCpkfYYQ
MkyAfME9ZSSJCOMlHEuWjGjBDhHfOSll9vaICZhxSKlUt3T0qvh4m/6kCUo0LpF8
Q9S3+4PgRQYjzgzk9K0YcNJyQxAD1HXfuCr5ivWcTqX/jWKwqi/+l90Ey4N/wUDB
k3NuQsR2MQKmCiRpO34FCKuDvJDZrFohZkhVX1qK/md2GPGazTuLNtgwi3KQ1rbg
lbigsAdwhnA6lRqqwIlIfFXXLVig5AyjVlrCF9lwOiu8sLY7pe3WwP4KBT3jVmIV
qU9XDo95aXyzHaC1wBbktJChuhOtE17NK9H4jc0Ovy/nhOFeuR+eDjOgZ+r3e2Wa
Dq423sLYG6a2ham3FGb56mYHyETcsvviZ3ac97fjAVpIndE8g/5imyw/P5oFf0mB
BpdwnjVpFSKbti0CtWUi2DDDtk3J3/86tWGQ9/uIRW1CUhJYfRtTwHeOl7leXHDn
ROUo6dFzmL9MBiZ1LcmgUOsm9hIw7FOvMuPpU6NxmA0XCcgMt+yBdd1CJAnDVwLq
VwJhiBUkmNC8BzkKX0rA8fm6UhJzQ4CcLB1siS9Od6ca5AOwea8cOdjzdkyWyBEL
6d90DWPuMlST8Vy2Kbhf7tOvxp9a8uyGPfGO/fc7SokdiuKTwCKWy/aRYIBQWyva
wcTC87Voz51GMt1e4dcb15B7Wh2dM6SMEwC1ddXkacpftTLfQ1Cyc6lpzxNY/XCS
XZxroa9BoXZJ5z5VhFl+OW4+3Cii3cj5pRwMyEFUcSuebKgIPvVEk16a59xVWM82
MjQxMpbByUMuKm1KIFBQywSbgzLcvo+6P7GJTIJFvL23/kiJ7+U5cP//1vYs/oeX
k06Y65YjwMnQvTlssqU59Ycjq618RKZkqKAJlFy3l8Ne5JDJmpP8/d7tXNRZzJeT
gK9XmBACgAoP4WQmU9NDKD1iCHAywUAwF0rQMsSZJ1aa0gc4E3Jf851HfNdihL9W
cJYXifkjAa0a1hHWl27EYt4SEuBjwwqb6b+KaeCsOIDVBoUB5jRhavyGuGszgoY1
5voERiouedoPQ0I2l8Etn0x5GJlW6edeTHQlvYpCED2pOK/9lqU8e3Jp19XCHKfQ
7SRj+jaoYCAyZM3TIdCs8NDExQ4F4c22B7nHtRo5zuOw999JVhavTZstjDZg7hlS
25T39DoNnvISLCB5+F94ZQE6QdJjwOrPzk3+uIuy80QwjjUKVx8Xn0qRrSqSVMuX
9Gd2+oGl8/eGokGDpQHSdFY/K9+ljovfZY8tAOy5YrTFqjK7vE9rbk16nzrlQ0IW
DhESVXwuoEKNeeNjPZGNTg2ByGN1rY2+c6pawOheZrAXYoxBK91zYq8aLkMacy++
u8HonYh+ndE28ycJDiYvNkHgaMg4zHBJEJ7RepIcXMaVnNkx2bzr9sCM0O7Cq3tm
h2IAvU97OyV3hyq2kerKFUa/vOKwYZMP2F3n3FE75dCNGucktMBc0D54XOt1s21f
qE3ig01M3ShMswt8jSGHNlX3lojyrU9OYq2SDHO06PjDDkCjNAHOfP5mGIR4uvVG
+Fi1nn3tOXX6GHByhsQVUnACgvS1wYqasG3q55932EmhgP5lkAApCTchbDZPDfnz
CFW5o5aJWTb86WT6umlEE1e7oGdSWha75w6VzCAPRcLgX5MwAPUJWPvzlYnTaANs
avJ12moyNT+1FfSKMnhHdtpe73icvDzcs9zUAiYnjOHMftBbdvAGclw8WRc4l1hA
nR3lMJ+9HmgCcxl4QrBnB1P7kmjC63GQeM4bh8ZrmxpIyKhLO3WDnsZ136egrHtQ
bzWHpGfiQVFV+GhmBRYT/TLQ2wpeE3YtMuiMtaVOmJW2/qJaWBD4sccd9t8xdMuF
4EgNvZKZQMW6Nb+uPwFt/C5lOXJ1/pFUdWyuf9B1uDebQi16s1jhCoeBHq8NWg/b
0q2Eq8tQi8TDTa/lFLn61CDvBv8RDOMCT5NTafJpZ6I55/oEJ03gWoBWRJi98S2T
PFblZEiiL+GpiA37cUZSpyjHXECirS/uryjEXmAjkxW068Sv8DmIFkEfINwyWLH8
WRq7DTUHnJpprChPVEsg2BXuKHzWmCBy3livdumv9Au//IBsDFWzgZDewYP92HxH
qgezpwjFdWTotuaA1YDY3qneGQVSxdScp6KZgDt+2LOh58Ea8VujB1NFDNCIwSy2
XAk44rFRWYf5cfP4jwuxnY89Y6Actm6R/cNAlb0pDb5SsNzPG+PNBzEdahzLT5xQ
87yTWBgIa6jRJ6kQH8Zakz4gjp6TVgy1NCGDF0GbCnjZAPBh8GBeVZcbUO7n9Eub
gYjW3wiFRVD79bz8pFnr8JJpQdGYTjTbfCkGDzxOwRHGxvBKFZ5pWMDKeJ3bLP/v
vYg6k7IjF+B2h+31yNl5W+IPJyXbqYc8bz+km5wuMY7P3asDOIlSpmJVLH71G0fa
hN61ycXdEfaa1YXVjUCyCFzwupeScW6/JakDjm+C+o+5ornZjEC1rn05KGWEzf9c
yEw39iRaE39x4Xf+Bebso8bMatBm4U5wuy9razJSjqOT5mWKSU63ejjaMLElq3Ik
Ugjq1XYfDb0vX6sjVnEo5S0NCeHqJNA+f7CdpOiTjnnnKXzMvIzP8KI/EY3YyLU8
kDakAnC4oO+646PWIFmPLJcWKgXN0gmbwRZyy2HLenrKb6nIRTdFMZ8NJDt4k1jA
ovId3sbwX8gBdl4nWDdusoh2RUjiaNiHx0bhvyKaT+Gn0g7HEUmfv9P7RvpjyfAW
BtmnAGWNRTiiPz19joasWCSvSICx7LFhJCWaoeonVEWn1JMiF40aXZZYUJp3EtYW
CiUVcj260m878NRPTWoPolVwGPwWpBtlJIoYBtPOLVTEIBa0N1U6/5zqcZGDxpRd
ZUod7+dlxdKukzasBRVlqayQR3ERL6KzVt1VkBQJ7/+6dzwQKS70/waIYK6ZtNMe
J6nuLp7z5BbZgjYHMIk6WRYNLqUpO3WsXOOlCrlpRLOfvpH/vYhAWe/SFoo+sRbB
66+e79FCgn0m+S0C6T+p/Su9AigXxmHh087C/7NEv2V6HT0uaOGLKKo1s5ZuRWZW
oGexi5O4+bNC7IOh8rdG22CL0WNU8i6dwbP3es3eCLPqlt8zKbQNdNN7b83Iv5FP
17S1cMw7nvxsWOToRXWw/xD1OUZq+FYDBe+CiuIfSALXK4o0T8fV1EFHXB1KITfh
uA0M2CSwzrvRHa2I65QonhlzSi3gQTZc+1CT+uNZQ/Wgo/egQEs6KLC+rL/V1h0h
uBlG1D9KOsU+2rJd7v4cj6vIBQr9usXfN1eljaGpSxjQVgWO+Jo+aR/UHlRXVwHC
43uNbBldw76Aab/bV2/zUzGNzOfCYjGdnerc0QUqA4bE2n0iQFYnP5FVrs+3xWW6
FPoU6kBNJwTqbxaTuZZEn/L/89Zn5RpAl0ffxLMDNsKsYh1fbePZG1xdkZdh/XBY
lS2J+VbHLoQuMhZjiY5JcaE01few5ECTJCuejrn0wgF3ZOjyt3Rh5UP9PEKtu9Il
INTxW2wBtPwD1YSzDdXHnFZDSp7SkDtygQoJ7fWcJSRvPgVleCiC+Unq2XtwJTWF
aaC29ecEIpqTI9qIvfSDna+Q2kcQdgA8D7qhlipJRMTbTLx16iJFlLyXsKKNsjVb
SEn3089GH2N5YE15AmPWFhybCcZHyArELp+xTiS/SqPfLqAG/LC1tl4zpWoByemm
DCYb3QWy1tIwJkdb7L010sjdgypT3a3TDOEt+FDir97tgCOfT69A5WjGErJicQbk
DSKRJX1dWCuRYXvtTfhj2EYLHpA6CJnQ2RqF3pKARuFh5IO6bcTBZm22BRBFFv6Y
Dr9+F4mBDFL5Ii4zAdXjqJ5Y4C/dHqwHj0FGvCFMOfi2iJ4j2VVgjA8QI4NCGv5N
l16W4qWeS6e8QnQgMgvYHc9bWx/J5D0l0zWs7XvcR71i3xis8EP8wQ+d84kq0hcg
VWnmVyn+sUuTYL/okOfNlE61JXN/+KRsEr1q593umKqs6wuZKH7umvxwSN4zZknN
TIsoyl2FCqmfAg96GRY073t9Tyxnm+sPcyhBs4RR+7zGD4uvzhcswarz9PnbIk3g
x9lVjO6UR5T7FV/XdJhP2CJKPinYWNd1sm/QNSmdvLghf4iGlSyiiq2W3peEth35
udO9dYYJZCj8eSlrUIw651SOJpcgQk3HmGcG9DmFG//Tw1dfYQ8Szpk/FizPbGYP
Jgu0J4SMgJTMAiuK3uqNQPFHVRkS+pWjBMpnqa1E7rFV4yKK/2DUK/1x58goYMKw
tADSszEqrASE3SgHmQjo3+TdCM2L9tFmm8nGSgBaCI9JCqMeVYDxggSURyubqdIz
JsktcCWo80dYj6gd0EASaf/uwqXhqdZij84PoQuE8Ggcxckg8B274Yuwz1BWP3te
hnnXkAsQRT1KZUHdjVOINUbVHDF7MEL6glnsOnPftUr4b8f3FTDEfUgqtYxuMGpO
/vgjymv+4k2YZTHmbcWbZJaA5bQ7O26p1DoXTFnbkx+VPMaTXUeODuBoHy4i6ro4
oz+5rgJClsmFuMR7XAAFNCoKPqHHmPe0Wo1V3tc047hxuPBQd8daE43hhHkAxpSq
yPaXp1jPCNNg0VPWpoIvask46XsQxImJ3iQX2LCdn+o3io7aHnHCvcshPIPT90AW
WZE2dGAmVpZpMF7+/25KmnTuqIQ/xYb6KPYoUtSBrNKp1o0vHZk2M/tqBA+Fejxb
9/Ha6DxdvU1WRHUE6Nk3xrkI7k9Q9wg2OGmOC+p7I66wKC31kt1Y60mRjF+Wt9mu
ce4XAjZ/2Qb5u5ZXDn1WhjjJEME8IJlvg/f1y4udE1Z+l5tV5hk4pTUaRiFDZVUd
Egjyym0RTafl2ejqgJ5Uld1WZ5NMUY1CJslO3agqfeHXavPsNYMC2HVbipaYmwhY
V++BvQ18gg8kHJ4LdTf+unkALrJ0Tcf/x2EPG4QRnOTutrKrZFwWFve8kLMCjdpQ
80ZZP3LzqdCfQK69JduK3T+pauCm9xPerfoXt/4I89GD1nSlgecbVc2WG4rllrh6
Gx4SvkQw93P/8z+Mt43aSQ97hXpfccUsZ3Y+NVX7lKCXjAznI0T5qU2hYrocrYBx
WW97j4yHFcHNmN0Vt47Hs7aW4aCJUtdVeVLwIJt8VdxICxVPcSGr/l7Vqx7n+STY
v+QERHtLzHpR7lc5d5xE89TZdnVRiRnAcxaiofPAp5y6Dbb5m4S/CvQ9Jz6M0JDd
sE2GZjAoI8xG54ycUOkh50+PwrtYdHkWrxJQW5GPs3lmEm4n0ymDnaWUA45wNgEa
111pehnjo6ftKjSrVDB6Z6HD9qBc4osg2vw6OoKUvyDnKrQMzyeGxGJeGUdbQwaZ
boZA7JnocUINGBZNY17wZ3vjBP4WO7f5ekkBPBpSlcrpomo97kwr8AYbpo6lillA
Nehz8tYBxx9cHGwGtvsIKQFxWWPWm8Zo7WyLCFU1t5m/ZUsdqURwLIVHjB0Pfmi2
vERNEBEbHQggSAPmPRSxUEC5ApWHhME8mvPO8yl6/b8pW4JY/awWjrcicslO36E5
8AL1DDwakmQE5hCz4swkoPc2BPgXQB3S4Xxf4fcIKvY6Usuu/+FPaDFbPrp8KJws
MF+KWHJ9lEbqjN+a00J7GL9Nx9uYmcsH1v6Jdfux50i5Fb8daWBGA75qlsi6rVgo
ttN+fhcwYalnfqCPZ0RUDgpQ56qmxrbYnPMynNB6tPTGl903vfFgpwL4jqXpjSnL
pysOt6nW9Ey4oAglAfiYFWBMrCjFzCP4ET6fEnzFe070RGkPzmaUGxUNrr+41puC
rCE9/E41JIsbKbya1sSSSxQWtwprEmSkVh0Ve4IsB9A0z2DlXwSh6bA2ehQZnyQq
iCM3cxtIRSNoV5VACWJPP9fB5igcL4uZqguXL/zAUr/7MfR2ylAg5H2jGy2EI7Ha
5oOh2pYmO5fCtb1G+0LSiuyhtp0qhU+LhscgYSSKHqhduA5QjjUw1GzLu3jEMvod
27wTFcGqO5WJwqFsgypDX5I/2p4xC6+1aO1DjUy44GlQsC8gElp6nL6E3kaRAxgQ
sNQ4KYwuO1fxjeYCuVJ2HDMVgz4VrS5SzREYYmiaBuRHwHRerW1OUTx/ahbeUOOD
zFdQ/2anNjEDgzuNFmU3ekJTRPok0Q3aOiyVebnZEHJZnSvwpeLUpIYPDUyFO5OX
qdX7VZu65WwyaKnPpK+6qqQ2+QFwSfS1FE2Mt7hXI96oNTt+t8SFpRTV36gX1QTO
xtf4dXkeKYV6Kepw6ua5c1HiOWV5ebj+e3BqjlwAy8fNVdIbFU8K5KMV8n1Y30ff
O78Qf1GxkJhUayfAZ7Hshaxk3T4AFa+CknF/B72Szt9lvsQzbKfN8b/fvlWEK7zP
EGYta13FTaQIdrPbalbnBVjiOvmzlKOCc8dYmkyQB6ZGP5hFk2ySE4rIrNVUnwa8
BOoOPChf+J3//IfnZe7WAnEAiPfR8UfSLY5Kgxp0e5FekWvlNuea4kZBJ21iLLrs
DD92UyWCX86bMAGwDlJK0DMemP5CuITNAllzRqWOx639lgeMuXt19e3I4jqu1oJD
3hNDJTqQUz2JHNzSWhmKaoezYMVRAuLuyHYQBBs5S9iQgusyqA9tEwwIaDqPeAXr
lJcS53PVUVSGAkj/Jf3gclc45g3U75OBzOop0KizHsHtZfmQTBSUVUSP1Q6YVIbN
P84R5NdcrQrKd0EueDpboPKEKjvhO4YXKVtJKnwE0q3M2BivhoLmUy4s+tO2SpOE
NVyRKELK1C/JX1/QaimjV3beOYk1iWz17XeCPmQFHt1DkFPbP6R2T3Eqo1x8j9iH
g4W+fmOfXx/ubsdhUX448EP5Ux5y0rCaTddG0D2JT/69I4QcZBrD3+G53Pq7vbcA
t3L+IFPIszUpgfyo8TtbniyIIMJ3cgPXsQbb/ljRZt8lNVx+Tuo0lSDmS+yyCTdG
lGvolJuztedR9+BrYld1vwHSkBtKDRjv96w3Txf/j8/TuMP6kveY7vqs8phSiPwu
t7fSkbmc7pBzJquBXEt6uAEqyUXZ2HH1sHsASpBAIORvj/agRJ6c6vxuIu12wTRI
7mB9BV0Q5MDtvgf8OFPpSvWnC8fk3ZC+5g4lAetiQP6udrhWpghq1xAC+uE2uN3k
Qxchgf/kzxI/NooyssmjvgL8iiKro1ARz3teKzPGe5OWZpogQ8x1oV0lmo1SRKb9
QCTfF8TrB2Bb1/sQp8tSpqsA/Cgfp4Pqf5qfZ7xipQc1sznQjUpu+WoSqjMWDACp
RX5eJXMsRYukOXDUVxbzQmR5P/yhQIum0Pej44oLk68daTkyhM98i/F6S1lCm8O6
r2trrCVg5eQNVFnCGsYbdbksCsYDDewLC7X+g/gUdgRhke4VY5j0lwsCOjmnL5f3
dGgQRtYaAiY68C2bNCUlk5w74Aavepkrlje8F3TXOyYvUu5ivHQx1anUPhQ/IGmz
IlZGGzM5AJsv4sFVbJCpbq4WytZc5lK43+I3YxXIRhNYk6BmUmIKbL7/69PV65Jc
OZI+W60QW7eYpu71dHEqJqbGsbXCHFz0+MS/JeM4yJuuhxnQQnLl/rVIEdBeSLqT
abaP06mlCW3nNz5Fb+hkN8nTPKtzbp0GkaOaUtAzoTx4i8XNI30gRPM3NXM1C1rh
/7zOx2PO+yO9tL28gNG11KjnRzy6ni+a/w55ARa6B/RGlgAdPam/q0jRZA7ZJ5b0
eJDCYB7PtOyyFqw3dwL0LZmrz/niDbYcom6gL/11yHME+Hae9mnw9A+p2sNml2gq
7lcKHIUoXXDoq0WbSmkfbN3Q42W5FkhMEof4ZwHRB/pm5l8cK3Rs6d1scsXYSldq
W9dYA5iERASpHiPjbXBXmFK2KAD1hZF22vfKHZt9p4NmQv7bqDPjKjF+F1d3r5HW
Rjsn/BWPV7B/43gZU2Ue923SfDO+a+ifMXHuX7eGLTPNjm+nVjHZATLP8s9OyshH
6AzYEM63STxLAPELxO3dIERfYIcZR0keHcQQ9Y5dyuHaLqjJ2Gl6o8MqcCWFozjI
lCme7jeL0tvvIVkvw35hZrGOnoWb1fXHeUc/FGfVtwjovVV+IMcxUp9WD2KTkAJa
uQ8aPJMaMa+HZvPzc8hcKG+yy30EKRXNhqN1jSHohISZPVhrlAf5yrljyJyb8qSZ
l6pPPjwbuP+jJ67JBMowzl2XQjBGRNeb0xXY8dX9WtN/F5hW836/mMhGlb0T3U2r
/Darnp03+itLPUDImCh7LTnpUwYHNVDO2hKEoD2wMx9f2izYKCpOwkrb1QqA+QXv
WkDEbPMgbopOcys+xI1glpagd7s5s328r/E2NQ92fiVBmAXI4AuLQDyUUw7dZl4K
lXl6uowH6ZHAoSua/m+npqj6tcxHLH8mHvk1U7FfJuBHxrNSiz0LZnepINCG81Vo
rwRJwL9FwWKq1+PadU0q7AF/3Dk+8zLdy9bX3Sh36Gpludlzu5xLiTCMak6Wwcuk
mQdV15rY+GLlpIaWuljXtKqfyxEiwv45klOfVpng2YcUIV1ybl6d8nhA/VyzTQqc
yyWbylCRQb2+3LUdTQHjhG78VL2Mw4tLv3AX1pVUiv6jyQjRMU/wUUO2QF4ZTj7N
X8DDjvxovGmLxYRuT4HBPOVoAc/ZtLspNQI5OElzcjC6NyeRKFPTuT8sU+Cf+N6p
2S09WQ/SNmN6tcJqGqjUXABU26DnuVIJguOPber0D6lBgvXdRAOOWUi7UP0/DgEF
fFAYXXwR/rrFqA258E4X9jkyRUmIQ0Yormz3UnegDGgthQH/hSfnAz/GkSeOxbMR
`pragma protect end_protected
