`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bcYjhV304TXE3sEeyfiz3MT1dAWkxTOPsaASNrqfnRn5/XosL25z/0v/BiWbg8yA
snrzMW7zvOYBtF7hYPwENfcGlEnw5fiUI8j/G9di+J5crYKPoSt/P6EsKQNIhBpF
Av2657h7LC3pzeMMGYvUB/xBT+FsWf4mPSdiKw83FUM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
9CMjXa4OT8+zpDXLANhnJX3scIJ4rH/e4/xwWYfrnhKWxS/vFsvWL5wnvuciFUSO
uBwYVfMYpjNkrHg1rvwf9wskGaylyLc63fC7SuX1Z8Wa1DHY5BovuHG9rb+K7kSD
kuIBqbw9TMVsekpnIKl0g11/KzEtCm2yFhQUzR2ksvUrxvIBDgjh1nAxN97JZObx
0Pp9O82IkTwXGEcZ91OeQJ3FoLwW0jO0LER49CNn8ATMLWyd8v6rZj3iiE5qHIS+
mfRmI9ai754uVbUERJOdRypHqwGlTPk4yLQ4JucKWDWTutzXM9Zm2lZ55R+ilv8/
w9vzbwZ8P+XWCHfbavUef/ranIE5Ti5NqTFmLYRa5CwU0xQYvnK1JG40sktL12UQ
qCr/cJHoUy2IdksuM4MrusuKyeeirzuzIB4MzDmBK3ss5+jzwb0u2TsfuJCXKhRw
U7/gIVo+aUYzSc6U8NzZ8CI44a8yiB148bXUSicRwLv0o+mFv2wDZ3oQsTe5f5rB
V4m86Znz2m2nfnMcvu41PtpMGpZvkeKsPKgJNVjubArs7IcejDXjzpPdaTrcLQJQ
kvx4ZvINfkkevEEOvwhRQm5XYaIeovfuvlmGnQO8uyIhBTxSM6oR1sFvDgqzjBnk
CT7+87aB4+dTbsku5F7RNFxdXaQw7RU8Oi1u5kT0xFMzppQMIEzi+KKjKMWq3j6a
0kgNLeKUh1Dwkq6Ts1mkm/GcN0eWNtffJzQ9ENbg7V8mfXKpSe5QXzG8bwlkolHQ
QOx8hVAj1WZS7oPhfo53xeerY6O5hLsV2lORaJ4T6ezfRNqQcr99AhfrZF0nnbti
jDOk2UJdlJCwOQgOo96qCy8dTErRHrQleWQDA0mzR/6WHt3by8Wm8PvlBFExaSD7
oT3ky5oONr3Tj8Us3bdQaRlco9phAUv1RRhW20Jx6mbx5nPdWFo6p3NH/FAIeuIp
7eKmZEUnlkRZRqbr6ArcX2HHEGvWGx6GySnNJTlVAZIcKnBLW3pBDH3/5ShXY1ZL
ndkR3yrUXUVXsqGzA7Fj88zxSKeYkwf7E4I3q9mQ4v4qptceyGb+qka4ttCVblAt
fcnqkQGQhNtaFL9dZ8T17pxW8NgyZqSQIqYPR5f/3sc69m71LJn2Yi1up3xCchEO
Q/zN5q1U1PUXGxjqxdooie8XQiOWBX1226bg8PIWzI3GF/xzCBsfO3WD7Z3sc7VZ
knJHuWp2+kwz/OXoAoJNLIzK6R5S20IOyHCxxQ5C9mcoiTQnYdpm/GhnWWaK/ANO
y1jO/OqBM/79yVMPN3wiUV1dgGY8irHR2UxRdj8nU1i7y4v26CPdkayYwpj8k1v0
OPMY9qmPSK4zi6rzo9mQWn5gukzsRKH+mx7Is96pOunzlbMUlGyfezfiCJ0+3oD5
d2C3rLavQGf9wSWPjr2gJ105ZJlpIm92U6YD7cV9lvPmzm7FcwNvQDIX1hXTgguz
XdXa9Da5UbXrdLIQBVAUSi4FpjuLHqTW1YRXL+dCLIu8Xt6+hIMk9CiTH+3vWcT/
p4LQexMlGOy0IAaYnnJItOOVBKHGH6o/L5Tm2IQzRaERPvCZ2M0IARwNftj0YX8L
/xj9ew3bLkksR7eGwhTB+oZeRfdNk+yQHaiOYye1mapm2BMfyi4Be2QV4/dpXer8
kjFS2k2cyNNVkUFDHWoNXiy+LYA2K+66c9uve+/t118uzTI6Naa6uD4BiZQlJHfe
obKSHz6X9P2xZD+thAIrVw0h1Hk08KZ9sLFs7h5MndFm7T08x0DE0X5VOtTCk1hc
nKRS2zxYHmlPzuAJ6DKaLlKIKKgSYL6a7WXZA4qT1nnCfzzAV+mHJEHP+gJB3yYd
rtFpf4xxKYXu9Uo8qpxdsv4F+9dI6v0s7iHikSOCYFSnTuZGNhwRVWZsLFkDO2kA
kMgQfGRWhvFZwJoxlW7bNk7b93n7DUB/vcfJTesgpPEOqHmnXSO/snSLUfbAYQhQ
UgvEy+fHZ61kyuVM53vS3cvRQjD8mWHHWrvPvgASrjwxd//NTf5VuFFWxtgeBtHm
1DfzLlGiFh5VntBi47WnAShOXqJs79UVJDi+BN0NkV0if/6omA2xOYWp4Vjyxlua
pIXiU9TuSo25luMn7E+G2wrQkXbxPT55EA76TuZuf1u/SvhYfTPcwgPhlNsz0qrf
k7Xko4ysPrUNNOttj8T6jskgqVBe2DOD8HRbmQhevlBCkgcNkOKtekIwn12haKfk
Snwg9hiYRspGT1XQEF1wvubzCFgBroMNsKoYy6uMQij+pKMhqESCLRnp5Abn20oD
8DOLdaNFzR1hwYuveHVr52ZM1o5hTrVS1XJCC6jrh2YntdBnMk1tPAeczt8FjC0Q
4LY1nDRtbKNR98A7wrIiPWHSHY1/VSCWam7WP+YgPEh7V6qsoFw3il+fJ5PNiwyO
NbR6mRQFszkAnsq26ObbfUJ4Y7NkHPI1H3hZs/e+1QTilzV7hNe75zF+isP/iqPx
Yol1gxxA7QIkTtM+O3Suc8lRfDV6IHT3q5SG/iZ1P+v+aymI6SpGxsaBEQiQE+Qw
aKD1NKfpIKUwp3eC+1boZx3JV4dnR8s78wvbevcwshsahB2WkrAYouwyscgRBX9z
fre0T67D15h334CuKOk3xI29QYrZdWZXVX32AEE3IV62yaygmtnDG7FflufIYGdy
5dZHG5Uw0Tr4PU4CyhhuFcyrohf4KQmretvrVUv5a4VB0jaH08I1VXerZy7k7K/x
lN1cpx8Lktha4iVIn+xeJHJHMHY+ZOVk8cuu8NtYA4B502UqBxxrPbV6Y7wHEAgo
BPHZo2mnAfon/fDDGCzhm/TdLQUg1a9AnTY4CPAsNU9uy0QcYDA3uWu+8sXQgmzp
Z4M0X3dvaeLWGVVV71/fDFDlzcpaypFHvWWcNClbANrVascQzwx2lrQHOZ4ip9se
X5QBkIB02IcjLM9hadh3RJLF/d1D5oFuwpGwPJkF0oBq1GHxpCFVJtr0iSTTSPl4
qwHOJE0cFgCM/5PK3qlXUqk8Abfep4U4Luo0+6FBjs3ZYeLlxfYxWnClhTfubcw7
+WQk3Xkn+n19uggfzMuFu/x6fF3lL5n3NfubiaP2lwxM+7pv0VZoj3vqKQkbwvI6
lRZUxlsIF9kU+lnndZJy3X2XjcPCF4/y26KBorLYoJv0MMKJBYxlE8135yzkzXbX
MnmFcKZe6YQFKuPNMl2ZepwMjx4aiXu3v7qLxSClq1EzkXu/VmuF7zGTYaVCxeQb
tpKPdIud6tZtYdcYno1BUS1c6yF9CE6H+HAz7hsxyD2H9p8zrlesh2EHUfOIDsm7
7sYsn3bzGSJxuxF8OSc1u0CK2Ti5vhBjA6K0rXY7XFUh2B3kXGZGCERwbKno556I
oOo3gn1mIlGy+aOJ/mpSqj+phzSGkpdSWjf14HS69iNA842qSqliKefosuCYAmLu
jj+TW9XA4ofQu1JKXBjJDVBOfVWIbGBloL/0Patp4HeoJpcxYlVqOS6OV8u0HOUK
1plj/YaCkZE6vunEtzzPvqy4rfIZsyCSvI3wdbTxGuyvqHooYSncyrioZecLstpv
DV2oZXpR0NQSq4I6dOnpN3DCYuiW52ywX556d8YpeQU8IwCWVzi7qFXMBVQjb0Nd
jJhrpG7wgXjBBMucEKBQcY+IWoQ9wA/NxdS38hPYxtdzpiSyFtyV9yB3bdaIAjta
afeP119daORwMMb1U8Eucd+zewMJTZSH/ehScN0gtWXOp20GVd2CY7cuJEOqCrnM
ZqZVVZjUK6XwgllbeEg7P1m86LWiW7kzByWIwe7cG4gQzUiSsV8OWLP1qT1ISaRl
HnqRgHOCl08sKp+Kp/Uxdjk07pOeXwQRbq9i5xfOBtfw78R0OnPdU1RQa/kZPqRn
pwIEU47aoZIKd3QntMOVqkHRd4aS5M2RGcW2JeKLZkdJ3KuBTgyADleeC+P0Rw05
OhcNWseTVCX9sR6mbpvTlUkECWMFFiUM6Qj4tTI4yiVA0SgS8eiXeZWQgVRQmE5r
JTwJ4nNvlmtI4Lfz2LKwlWsUny7uCOFkKjRZn+0LX1QhtrQUWmJESNYjHTeVFitK
4T+0WrNab9aF0cYpIllv/ZMPW+BCkUn66n5nckfzP089H2Vsfao89qZIsbGELZvn
EuilZF+eSmTz08+0Yc4SYrWA9iY3i3rykhIJFEWw+gmfRH0CbdPGr6bw6UJCsK3Z
VtqDb/nRZjJ9FJXSrpFJdG5AETvqepaMGOIhh0DIzq1Ar8POJ54IDnzsibeSzUCu
6a7LAbAgVOO0WzxdSDyUvjJMGdFXajnQRIQYpIX7EZR+4FrmBv7zc94oNQyR3HLJ
BOfv/srbS48xqCJ6yTDfmfvAybrTgfF03Auwt8E1yCu9uaFAM/zmY3ahN9GUkQe5
2dwj2aAZTx19SeZtUXMBkZ/3X9yZfLwXqwMyxhBrfgCIoUpfKKV0g7gJ/60HaZFl
QfICQKt6VkRjKererc9fRg3bVurqpV7CJRO/oK1QZe2ITS5a3W44Psmo39VPmCrm
9/JUIFHK/3scKKoBgQok3CdSE51K2MeMywXJn7lz8cCewi2rdTV56iNAZACvi9y7
AOauowKBisFJ3PLEDDyxeMkiH3iLe3MNzt0ArCNG0feh8EKytAqDY88ERh/Zc24P
zCLR7vLi1teG3jooDMbxUdOwLuGMwS8nzBNLyJgfBkVcclFUK/4kv5mIP4We1Siw
z/TPQtiof8DgwEkUJTnrwT0tWFK3cDDnCtnFZ9NOoeFWgOgTL0B6AFR8wCn/bpt1
GE8f3RIXBJa+NUUa+rdkccyhMhLqE9oyersKO067kXsdrVqw3chpiVIdmmlM5Yxe
2r129+3rF288uCwKDPaDEXV7FVmFpN6KFHlRcJsepax+cylcg1UYhTFAI/5ILhQV
7+ip4aEi7GcyehElnnHQp+jYGriuPvVlV4qS9oe1qlML+sfMV+NOIqUhziiYXhn0
vY5wUVqenASr7D0MXclxdD//qgd5FUtFeYwhEw9GKZn+z/M0rq7BKf5PqsfYkVeV
E9xFjD164dPjVaMJzaYTB/6pQs59i0m5ZBakr7XYJfoV8/mDXMGSxJo4pK4YMPby
VVnv8y1wjbSkCpNsOav6NIgCjhxhPIjeGpokptnxgHmFqfITzjffe77eDR7h0h3u
zmO0BQXmS/uCYIjmFfkmEi6vz7awhwdtWvGZHebMb/LrmbY3bzbDiYHI7JnoRFAs
IqWyHg3ufkahIp23kTzwHaeJowRf41BNehHMz79wJpwE+qbLW6Nerodqq+7y+r2O
FHSm3adgJ359pItKfViLDWlueaoMr+5DyQi1v6QT/HvTOzTdbGte4t5scKRyD6y7
hEmMfF3rkzILDFl+5f7nG7x8MI+Ifb3iNpMLlybslmqgFtRwWMEGag8+a1Mi9A7u
9l/BHa/jVNRGgaPskHOmy6bMAOz+qYxUlxskoSjaHN9ulEEbky0IsnTgWVrdV8rx
B4ZXcMT0h2TS8nnwwjQUjZJjfGU9xFBuJ4ZXau+7jn1qs/devPl0AVksaDyMZy8N
T10GDWjZQR5dLDXFHUUB6G+YgPY78Y1HM1YXGrFH6Z45n5sjN55/+Zr8JDPB/exH
xd35/KSp6ISuPMuC+TryZ8s6H6ienXEVQG7sI+VhotxmN8HGR2YG0EdW9TAa7xq7
+WQxjC0uoTcLE5szEqHIUDB+U/QBhhwgiuynBl4YmXW8W4wlQrc/pBgYENJlQ4vJ
dkLhKto5SICw+2q5PLaMVWMD9y+mW9vWFqWKXnGSiyF6MUX9vejnwoF6M6BeXhMJ
TETVucakW7LgRsC02rxagraRXnpDX40mdDHRUTCyZ6jUVONSv6bXq36mLftf4e5C
FBJh0+6JQ6wwMTpwCHDnK3+6kX6sDMaORpFjTy2GWNp48zRHt1NedNS84Qevv/gv
8ZarnpB4ksUgvRXSp4x/ypWKpkkUp8I9wvYoqtydxY2dtmgNQI/Wea/QDzedA6b8
gf40a3LMLwGE3RodZ3MNRx0jf07BHRGv0ZCNUGFN3Qutq16b4gXU50+4XwFSaFCI
x/I+V9uUiQGbu+xgrxG8SNhLPZrVwWVD7dfdiooRYjnWSKYxZFtAWN8kSZRh/IbT
BUuGcuklBUzd7FL9L7sfXVHSqYggT7psT17FLsz3TTMhJqL1S8G9Tixry/rQgg6A
Tq0GCWRbtou1ZRbQRqhpxMoHRnpsjgu7HAq7Goo5HADMnBRgKBS0O0HDVnUqJSU3
EcJZFXNJT4dA5a08eimhhk8AR1yZD/BJ/0vlkXWC4EptBDEww8zfpkW9se1oFJM9
TsiaoYtmS9p4xFvyUXG0s+/ZPhDR/5o13tfmWH9uLlsIEyvOlLB6aN9f7CUBSeFl
dewQlaRgox/4DqAh+lHFjZednv5fZ3iULE731wjRGLudKnVnAXNIyR8ol2xDEHgk
oXWkY6xyjAKjPStPWZyiHjxr4CqRL6inv41BEJ9YUBY/QYF0NAsYkDfHF2Z6ob+T
Ke0xf5cVHY9PBXq3tUgLomXCUQkxef25yBwvsxe3jFrre7vKQvfgFHJNKVoJ5h5b
4wwQan1ENMWXxXe0bIQ2FBGf9vPCtFDMl23Ac0TZvxOTzZuaM9xHKf09oVlZvgiL
zqARe8XvOLQMoOMJSeQ2EjwJ2uth1LNReOya6PA06VvXYIMWHrvcfNVFWHvM1vI6
rZFEIdzpiRakZumtd1CseFKASEfUFwYrWxkR89Ms+oMVc7DgCBbFUf/D/0cDvnp7
ZKyJwG4t23VKsSltEv6MtrHYchBNvcLT/VJ0iqpywMLQ+QOY6ucOMRkKBb0nb7y2
Y1WMkJyQvL23ipLOt9F+jlT/dD2bWaMrGlcEIRf8Sz7XL/fRY2E9vCEMouJKYpum
E5PeCXDF9heKMgZ+Lxz3QqX/e5DKXzZnprz+Ux86SZxwbyOyD3o9oYlo9w8E+SVB
69XvpORU7AI1mzPmgqRhfhm843H1O5IP2u889i9fHU8w8UGWJFpTYxTJLPOpdIHX
SbpoeUXdJ5byKPFAtUbdaMw6cHzqmDNwnmaG0o315lUm/m11UiRCxz73oMRdoZk6
SZb0VvFFYChamQQe/1/yNWPRYOHxMhL3IKSEdIL9EnPdtfog1nWzzslD+YUaeQPu
2s59nExFJ3d+ryNmTBSTfXU15jbPzGrFOWm+ZXG/NsuIClgAPM1kdTf+ZCOo4dIT
tTdXmDVbtsQp1nEc94tF1+1F6UDS+M5T0HM5K0YNZLq0dnV4N72y521WmOiv4SLF
eV1whTwykZ0inTpMpWJWVZlHFiTTY1M7ZfgJmmIDqN1nMrR5IcyZ3oWa6gQ3jH6e
RecdsgItYlqPlqMwfOnuvFibjnGbNm1SuvEHljPUCY5bfWeWmCcWhQ70moBggZHT
Jxf1lz/lB0ycd0FMto19p16d+jSt6KdxT1Z7pxee9dvFfMjHUwvNIBIkp4L69eR1
RVGHSRTgYg+00xJtA86KMGKNrwuWur+27w6hU8wi0Lv0m4ggzHbhOqDsnGnMw8bG
P0Fo4QRmPPYBfABnk1NL74nETWdbuNlnG2lzQf7kfODwBCobQwmitiZNpAQpcVH2
8XEJbxSoda1W4ixHp1yEM+uHA546VnT08AWcFY2KcNULH+JQBEt0Pzh1fobMT+EG
20bl7Z1aylikRtZ5SYsuQaUuqGandUDLCLNvK5mThbMySdS9choiTD7lSuoefYN4
v463RG0WeuNwORtPBuFZFIMatw27+68dBEAYAfqac17W4XpkKyDS5qsyrslDkANO
lUI9sSUYbiQAEfhybEilJt/jcrGcQte1OSbE1NxG/idUtZA5KKajQEt2+8DlBt1Q
Vf8JNYt68A/8fJXRmV4ATKCS5r5HY43OHSes5CkChBVmNXqZkp07TInqJY5tixf6
B7wwj2BPHZ1NqQ1nbuzsNDq+VjWsVtPHy4uIiQdKHixSibTKckg26DXJ+FluzowC
04t06rIyOlP9Kkib9ym/laewVbgV0EnoHPCkvRJ8q9c74TxDg+VMJm0hqGKU1Wfr
xQo4eiv04yaGds7JYVxFcjXfPJE4ZHo8CJ7qGTTxZg7+uikKtxRusYlPJsubNgvF
L1NNY1lC51uF/wxhk9TIqykf3D/SdNTGg04HxXwDDb9Pvk5idmN1IDDy762e4EYL
I3ExcT88PEnAlIdJZHKS1xFkljvuAW2FFyFrBBHD1w7G8MzkHecTGg6oiyXNYyTg
AFQVi67b5HGHtz46wUsDVu9ggS5RckD0oloc8sFpGjBvOjqhMRl1halLt7HzqPoq
viW3UCrUWiN3imH8nRfTins7ezBmYlqvMZLVaQW89viBvKBWDDhqLAGKwq+BGtdb
cMSweVpoEfNLQ7olBiFyNknbfzHejHc1sYcP9cTg9KxJ1MJTAYgoHML9h9aoaqGv
69QfC9Y3dKafRsSKoL8+UGqpPA2H3orKXs5QaiBNbM2ne7asVNutnIRZNCTVEAOk
Xv8JYDR5Mj2zJApHc1kgpA==
`pragma protect end_protected
