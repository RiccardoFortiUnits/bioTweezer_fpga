-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
m/vdu22YmQVTFIwNndMtPGuUjwMZhcDjDnBPPOJMFu3E6sPQqUnMk5SZNi46WetpakMTFj1ZV0zh
vpoyPrios18Z36/TFSakVO/XOy3yqr3zUFj4nAz6ZY6VKs0NAqcJSagMdeylTFmApLyltIQ6GH/h
+fVkrAR1WontpxVaY4i5QFFlDJeH3RhBxY767O0mdIN1ecipwk67S3Gr1KQxuFYxcHs4EtJf5SUV
DEfCaMhTvUBKB2+GzfHp5YUdb1jlRtv0ClPGArExSk4+LvqB+32m7wimpPGAJ3ks7Xcvq9sFFgQo
RsnBS5/2fpii3QULrSHWfzecb6wsEacvpjqW8g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6224)
`protect data_block
gNnBoXsvM+lOPpkxM80CIuLIX3SrtucwtuZ1AdkOI/kwvMVr/We7nbAtI84//kSfnfdgusx9MPmI
U69jd1FhP1NMzl4K8xXhgbgLS13aYQaE2r3uxmbl9S8AOoZ8vJ95kR48Ox/9uc06drkrNLIunpXI
g+18Mr2kF6Rc5w/8RKsj33yKKKxY/X5ZEghK8IfmlNd684atOSJS/07AUJnL27whQJbIBd/A+pD0
F+ANzGDJ71jwJfuuYrPVF7+ieRsnIv5CiDQg9C6ZTE3ej4d/eXdmKzBHrvfOGa++XlfkwIS4mmjA
+wbsqKtiEDCzngZ0Hu+hz2lKTLChhcIxmLy0N/Y9WUlPmdRUQ9hTCCidsZ5Oo6T+7XodD989KSvi
yeagXC/3KdvRkGkucxkKMRv1gXqRvCMH1GTRXzED2Mh7P05F9oHGe9B28dTE/Qd7AfssDuBoOfcF
mbW55kB3CiGRdg4QMrT35cNgF5nntSI/uvFQ0lANWbhASXv+sIFqlnOF02TkBUFtgkI7nX5j2o9d
mpb9Ry39Lzc2mvK8Ewh6VPk4+GVlR5NfIH4yuQCv8IHehDE+g68xT3TQFKTNQxhisUPEXPdNl8VT
ZZNO2jvX7ORasnN6fmGQeG2Vpx7kxCxqT7culdzsYPC/Gihn3LEJf6chBZGj/WOANchi9NJkSAM2
TR5usdNuZHCbOC5pFIm1yWW8WMIlC/xESI1oiRrIUZKsDjY8ege+Zgya18cA2iZEA5qht9B5rV6s
rNQvMsU2GLA+a2hzVbhU5IeKifBnHrAFo05U0g1iEa+QCnn3rx/lGxlj95bKMBX+1ow6ih3OPbAt
P4c/9Of46o+A/agIubfa1Zt0wx7Ew1A0DjPk/DCJEjYd0QnRR7Kc/O4z5tKBUwsiq1z5AJBL5T9G
gGRFt4Hgan53LCpE3aBs8B9z6OsmQQttGZxtqvoR+kLUgDMQ7+WxqvZwZTEqu4EV6zFhIju/d0jr
tKsqSarViDWwPVNIu1Q25akGjDF4F7t2O06Irz4M4tlsOqjwBmri8xgMBmnJbXYL2mlqzxFl4UD1
47ofLEsqKgTYSYWQHvahYAw93YLGjVIyUKt8TsuUbkQ4YijrhbC/dpuy6HKmRPxqLrPXr5jDEJZ6
ZMVjwvPoOOgMy/cmeIBwZrCKH8Kklo2+8LcKnDyLHx9GDXKLVGXSd+xfqA4uvqdAJuUlCarDtKJR
A811HkmeU8MpYebX6VD/otN3fWAz83N9m8XHx5I5+0nxVgc283jsstKlV/gSQ9TynVND/ynIGxaz
D5F3i9Zxs9R+i8RZvNiPVLCtErsJy2PcpfMeTvgBdd3zUXY2oyFrYk0Es9a0jwDWlrU8sAkMLVm0
EfkJv9bd9WTofBEZZQfYD4C5q5qguioJ1lmTY0nfwHcmWVsfkiKo2TjnHe3CZMj8cFTiZJAHvVkV
m3MEHEXOuV04mrxNqsyWKrHmTgeHMn8rrFyo/p3w6Nt8Ym/ttCnM5OOSGbrA0ccS+rqHyOHUQf2b
k08ZnbdjCCp//mjyP8r/8AXWL0Knavx/LLRLQL75k+/HzQSF7Fj453JwXXG6m2/ZpPPBam5SaX/S
0UDIGbJ8yxpdoOGqGeDvWvHXChbo5Jlom/mq+XKLSxmNMEamXcS7ac63tZec85mgf1ea8bgIqzqb
RUBHbBFM1QY/XbNx6uIzvnOI8AMje6+LQqGj8XcyPbzThafQ+H39fsBERzryNpU5AT2i5mSB+M3d
+GSN5HxrLu6TfZARDlyNnJpAwUk1apCMczgx1iede/jfMa81qhIMQcGVkjanakIAizisqXbWHW7x
I5NE+Q+sWQQmdYL2T/ib2h00sARNCA8SFZBdDtXDW7Gzk8V5KtE1K4EpOcxpl5Bi5dO3x8gytYOr
Aw6eRQqEnjK2AhuPsVBJrzpE1SQEddWxLM1+tq/OYoKLvhqNvKLlJnkWsv8tbhfjLbZKCr6uREOf
T564DczI6jvQj7Hp0xu5LEeweBUVjfr4GPNQnytfqYeP42fJxYuokwNfc+ztvoaMT1C+A5LtskYB
UozseZRBh0sNXFJHJn6u7ZdQP761isKdYFeS2e1clhfHo05z7IH8BMuhmdiHKORijnRqapmmvQH6
WVabxsiC1QpA2xKHlZgNwk6X1B1J0B8Gn9Ml0MdUu/o5IHwJtk+viEW43mVZvO5mlDXNDruthzGP
qZ/V0SS5r8k79P8tj5i1oyqTNfzl666uaxPPr8NWgE67cmpm8WwCkVBUdhq+gOcRF6ytRPizX3AR
olZfcbA+ZULdpkL5KSz9nowg25AHdYnaLwkMQXhJHjGb30yCYjnfY8U4OIyY8f/6OVPHw/cn2WV+
Dp1EIrpCtbCUWKNy08rJYZ8L74QLEvfwMfsR0ag9eQtYZLQwR7x2sBI5j1xlN5b9dQ0Sjxtwoh1T
Q1SnlV5HW7+6gybH1yR1txXgWAFVgQjyxgQYL1drsEwXvmHs1JgmqtWi16jG5rcA7whSbpYea3SZ
h+t4NDHO38AY0dqnZ1gXAA8uOSQogeh8BZv0LpXGcONSYlWfDPXge63L7yBToU0ppRPVYpKdjMvU
sSj0uLvEAjOtTPWHVhPz/JsTN47uJAdU4BCzj2MloEepIL+v0xSeQgR0oVPlfPN4DNSALjyljTHc
vkYeAEtRLB5vI5V8aY4cudIhLU3/4yppEabyLfUfWpvsYha3e0gKSEeOOWZ+B6wcmf9rxoHYM8cU
NKC76OJ4gVfkaLdKhNTGTj+5jWabXxzJOswCCjr4dApmfiyjTAidhCD0WsaWCBXVRJmeiB4FnAbi
flG9FirTiG+CAEDMb8uuGnqd1lzoA0DiNTkaomH14hpW7iQGVr13RtXg2T9ZsBazYQVqrVu6lPsm
tAb+fo80y57Os9Yn6RcRj37TjedV1I23nK/Lh+uok0SG0br0O8/nVIfbEmmvnp9KAPzzjx51ICWe
Yk+O0LlyN8tHz02jy9cLHOjKL8ghSuRWLtHpijLKxZpjHee8tlsD3ZNsbnhb0CChEsIKK/vIg6l0
YHSgOx3qXeOe/AxNSoQVnGCd50LngkrrYidF8VHNDoE7IrrobB5cPToxMUCfx9HL8gkpw2wMMN/1
BFX1ZXt/yG5e1VA8WD3J7S/0VU+JOF51z7sfnKGid3ipx1aS5L6J5vaA4KhHZBFTRa9TTizUyynS
nXtFv1/fYxv1ULN3NmoyjUvfzMIAwpSNqqiS1hntpQCpv18PAx1uuyVs1vt9HxTH/kCpOn1kKalW
ly2pW+OT2wJLKrYnTMLBH1AxgkyONWsUXWbD36rd7mJH59he2lDWhJ3kUuyevGXWvgyOpfL5EmWw
rfg4TXo22X7XFr5BZHR1dQnUMqZO1OoKX8FtR1U2gSqjdfBKN+NPWApp1mOuywtXCFKeMk4IrJCD
YTWk7rCLBSahzHfszJ8YOaIA84SwFtDMEEFXHcI6qvFh1ogOIdB+kxz/B5PuYNifsnLJao0SuvrV
xeQaKSxo1UBIFe0D11Be0BHqAWzAIClh1Y2aAKywvIRfTnb5KL4U3LWAgg7iPmn965wLk2iyliI9
sGClHUzQJHi2eR7tlonvHzO8VMF57+xcAVconh5gYvXZQCWorecoZ8Z4j6MoaTo42gkTOk0ZcNLW
OYoTSCn2d/XGFGuKXDxKvJ6bh82h201VgSRtPqoNsmJtM7wE6gwixsIKyYWsxtWOdyoJzNZQkTIx
7ZjSIBG4wnICqaOjc0uomB8mw6V2q2h8x+FDiIjN2nyJSOyBhWt8ogz44NsmHzeGFhstfdoq7g3q
szusRDsdzgf3g7SZph91L8Jxd+QVZVvekP+0/jMuWo/B0H2EH1SQzds/OViRl8oT1XOUb9PPzFeB
FjmYRd8sWfAdA1/purwDgkeivE/jB9fu0k6j2WsPgxkRhtgRWO3tjkIhX19aQ5H3opKkV8LNva4m
gBJSkDRo3ByjyM0dj6p/u1av6A2wwt2YHEL13mBCbpmRI4uYf0IzSNDWqvZ0byJbm3dFw9pYdnh4
KKS2C+2zsUEaPAkwYJYzhg5XOG+C0HiWRe1s9VMF+4eRebH4hCr+Xt2BzNl08qKaIrcRLaEAwYK+
uomxzAF+JoG8hnexzqat0pT/io0OyyvrFk3TrTFdbRz5XYXOhiktpBeYMXR+kJUN/2n9E+KionYR
qDfn/gW1pBqMbIfqF6TYq9PAptWxzHiWwSuJ10T0pOI6gHZBES28zdUfbmR5pPkU/G0l4HDpCfMb
gDd/rhbnr5kN4j/6Y/8ZP0ySoFi2r6qq7oH913vw0xIWnnf1S0ixxbU42PvHqU88QtM6hP/vAoNt
XJr2hM4InsdSvxqbR80bYSN3xODsdj1Sanp9z7mpxpzlBHt4lHnNoPwksE2gUl9gxSucOlbNNOP6
QqlELxU1xsN3LYovwW7t4cCGatagKziTbrCWPBs0/QYawWXjy2e4plIxkQMBRwCq3/GS6HLQ43Vu
DJirsPqiaigkqlkArN+nC9QCA99PUWY9qtzSJcTeasvpSKF3ynBXRDieBcUSUZvieAHppRIz87xB
mcTBCHLgIzScOAC7A8iLa1k2h/LLckbyXyustB3UqHwwUs3Gmil9cz1n4jdJufItiMmlIUSWaFhA
hY+OAzojGKn099pSIW1AlXUP88Bio5adyHbAEjx5Yqx/4/pMzMc3xqoUzy0HYumR5Z2GsEDGD5ee
nyAekjNxnkYyvXb056MgQcTIjI0Ywxv564JmVHOTgFqZmJdC64bJn2UC3oMfGQVLDS2TgpEyFfnR
e31iGuV8lh5LxZpRg7dEn+6wC2vZ4m+FMfXNsc6M87lCSmdPXlbuX1xHryCHcQ6IkRvJQIxV9vj5
6QTorYMEJMpVtM7T7EJiVVFwL4BGIx2DRP5yIbLox4x6LrQuFPkO74tVG4j+aAFrGt4it0Q6NuzB
iY3aDWa8OcCuY+WBYO7opJB2oYT9K9iB4QB4rnAIioFtpDTV7Z5/qrJZsJ7vdW33zpctbXZvRH3S
B5Fi9aPt0ujwICRx9qVBNIW9uv1bmsO6bLKa1GxybL51wzb8yoq0MN1/R1k2fx/POhgh5JSpGVwO
fwlBMZsyGsynNn2J6ZMaB2JC9+DlbkAmDV4pxfQQBP66/sOiNsAOdIvRTNvGDZB4qEefiJzfhrxD
r1kxLR+5QjfuFQCfigHyGsjv9tCsGBYFU7Hp/zW+PQOSg9jLgZnhN1HZNdrz1DwEcxRZrtxhlL9j
+o/4xNpR6y3F0/aUZTpD30FN6QIAOHIuViI4MmII0vqFuDPIQyaIdU0haZchDl1hWykjfJQvYAUg
J+4UnwE7KDH4FCIARc01f42xJRcTc6q1paYLyXpo5eUaNmrFKeazijT7m6puQc9ZZOnQ2nEuR3IR
BN8ryKfIj6MWv/QAUE7P5Cq9NAHZinfZFsHFVCRy28rWvEhMANmn42Zl8ZauIsMnbgjCsPAsfviP
r817Z7kTNjL0K84LovxLqByh7INNoIxGnj0HgQkNQRmNEl5hEBopqQZBhgS6TnYEh04UMn1/ns2y
vUhooZk3pm8w7jUBXtK3zxC3eZ5cDPXT7Rxxmz0yGc+t4/7/rXLiDK5F7vIQOTaIT84y8TtxdSGF
evOnEzUFVs3IYBLrn4QrDkN/StJ9p5m+LJWuHtIyMnTFIJiv+PwFLJ6aT1XuvWpI4wgQrb2HeBuK
XiTk+O58Fecuv5CLADb9bodVYiROUgLVZvywWuc7hi4gS4umnJMe46Ax6pB87uJhq5FjyNRMD+Fr
onrFQrc5lWAZ+QdqrY+a0u6XEOAWBvCTZlfJJgp72j0vLSpPamJmiSGFgn5s0q24Dn4f5lD+gTkl
X3raQzv5UyDh5hDlMQxwFXwMLPbPDJOodb9ro6Pc+WbmNjnUfR15cy4UhrUzcDlQJsH0ZGSC8lGT
qkguUb3vtxbd4ebYq/rPG6nhwlbYJOzQyzRGk5SmjOeFzyjxChwmL5LPe9mqOSoTz+Ocy+G4lYrd
qr98i5AsFRhlATtoUMFDXK1dHn4VNKoClgyrQbFx4rdRO6udAiq1usIdjecFEjvDeau10zE0xacz
O/mejcaHjQBmMlZn6zE+83QqYGDcKF2hbWnOC6Ug076GNOjXG+Bmuldka269ZCKf1M2+o6Y529F3
nh4c9lOs6j7MGxUQ0lZ0U8SSB9YhZCwG6V0YMzP3/W27Jp8Wqpf9/aTtKEWuIjlOmkrGgQ/4Eja+
Ob9FHKbZLP88Mrgcgqnld7tvFlsWipHnXigPe5a4pAMBTefeQ2FhbxADb454OnbVe44BPDceGcQm
2XJZ1y1wa/nTrKhzPTU6/WEM1tFWLvf3kjS2CC+D0jJyjHhrWjMvDywpWu3M/KctIUfUo9Bjrn5w
RCLe1592BdtItuunFdt54kZo82yHNChu+gO8OdKML3s1shZoBJMjqByEiVM5rbBoPPTyDTfKqtnL
a6X/A+uF4kMtftXrZ1gOjJGbcxs4xVsbhy0HNwSdgQq8G6BAY93WaoyyTme0VJviGfPAaSTDj1UN
bbFhgEQwLjIsD6mvYY+REGIJ63LVdx2xlgZ9IqbZPSB68UdKtdvLAlmgkhWDmuPRfHYavKH48tU8
zRHCPc9gsvyGuOHv9hYpiXKmY5E12/dWNhTeGI3wLPKOos9XOh2g5Y3Kronw9LYPwsxf20wxNmy7
KiAed/iCPplSvo6eDL8jZj38WPBuYNWw1uzFt7RE69PRXF2x7pcY99PzFqJ9m6vQ/IN9eM4Vcf6j
u6dAGBs5cph033FX7gwR+PCtfL+ngDrfuwitkgaFQ/KDLW6e+8o96Oj6/zTtYx8iU5FiyfwxBiti
ssTbNiVdyEM/gDMPyYuTJ1g85lQEu8F2ljdk7z9Y84Y/TXoGVhO9DhPY1pjGbYUGS71lls1+cN/N
BYZ/4dwbsWiaZm81bqkiehqwb6BaSrs3vNKAvxd/G/I+FxbBamkm+/MxtMPMnUy3BfmL+Quly95b
Xh0wZlK7KTeOJdlXJpvo+lD39JdHfMeHUYfj9mytCiUv+kAZgEmTVPQt2eMQ2VYIgaF2AA/rCoPN
btHWhA0Z+sj1vJ4CHu47S+W4YVAZah05Dn+mPZI7IZ57K+naI8aFNqfBE6zg8V9HpfQ2Rl9w1K8W
KKepUh9osR5v3aexQ869p9wWCrhojp5lodfb2GtYf0xRn7dePJWM/CdRn5cY3NdHUc/HRcntWynn
Sd13OhOkLcuS21WdmDm8/mO9iNXP+J1wjWFPRMFHsn9nIqN7yX3h0Luu5kbuk6j7CVcTz3Equo0y
JZBxs/p59BpSzjWgJCZe3VMWhS1cw5jSEf7WuNdwYBe6BLQyJTeQiCZOFj6q5YpAILMmonIUavJa
UGytZOqqHxE4C9CfFL20Iuk6HyvSrCQ9k//3OqWCQ1193TuUcw1IJf5IKv+q/8QCIw1FAf5mr5HR
2qcJjHnRoDau1cpms+tSGWC+vnBwIiuAn8Gk8cdZITn0s1IOYH1pfWjNh3xhddyOXDUQCHj0ubj4
UkllP1cRnVMvvVP7He5mV5t6DqpKqiS+PAQN/IT5pQ/CB8ABEUgj1wewbtwveFizjoRNXHRAB+IK
mHl8MoCPOEszME80ZQPNZJUaf9J5E8IbnP4mFUYB6/Jiks/l7xWH7PphfE78D7V/zlTMEjoPhogk
bSY7JbR2fPvJlNggcE694zehkPCEo7j7+IMtuBY/Y+utY21gtpLXSkBkxxVsYZxRC3CgBdU7GXDZ
uwYn0b15+7zCM7JO4Lt/vE5ZlA1+iDx1U+hvogUkdt3gxS6jPAs1W9jnk43WRF+ma20V1IpzAg2o
z5lB2xQlW1eMYwpGmY83c0fXvDCbZ8d3/X7SbQSNH+/ueiAEzujnUTyVzHjhDSGMNlz/Uc+1bo1A
bU1Gxi8pF6XSLCGjE0zKjlK3y5CvJZpem+2U9DjetGPABAdypQx4lns7AOyOMMK+VYcFVTuqmthN
lOUyxdyQZRlXTlx8m2yQqZiGndNqgLrVAUNbR5BP7ucJpJYB73+v2ySEnWs9JYsoMAVR6mpc+Bi9
cEH2npDbB/7e3U+5u9iqNLSh2U+FgPxX22iGZPwy/XLWCetEkH8xS4lKDXM/iWbHYBdjMuEwoOPz
wKAktUfZ+uovBp0po3S/EtIwHVl/6tjAjnxpOjuMr9W+hVhxW+jjkX2k/yLC2NiOzwYC6L/eIDLC
vDWi1Hdr2eeYBFJlzNIzkVicHNjJjuQ8BIS6V2YhvK+a7Yux3WgAOeGWiVlMQ3hgDeIylexkmMNR
vBW9g/j2koXxWxM=
`protect end_protected
