`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YyFUlbu/gRFirCzLixeirCnLM46e8kdIXjYk5ZiPfEbwrqSLPaYL0VFN7qceYXE/
WOQAxh4dh/3J5zhrqH9fWUO90r5UyHB0lwY5WwOnhKJHLragv4YcUxMG/rUx42wi
WDfx6YXXrHRp+XGizxmZAUI1tzQdCgmuy2UBlppORoQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 104688)
Ap7bXH92wr+0tL4vUQWeb6v/tgJEETYsmbQwPkm2LtgKO0zG8EZsaDJiXHeWmWUq
ALCHybPMqG5j3ijvRQS7XekumgAQK2kFtCv0A8PRV8UgmaT4P9tQ5tKuNm+f9Pjo
1jPSYMsjkK8cQqZGtuoFcYRZsEGI1kgQN4mVxeizWOjcQxa36E7Dopa40KKd/KZ2
rCYYg67GBNRwVvem47zBAU+De8uu05REYaas8g0JqqWoCGsdjoOn4TwqLshIJa1C
hPU+NR8CnGaGBPtMBgHD99OuX3R0iMy91ExUmM3TgwPhs1maqep9olqWbtDRi3MQ
ojR0tctHJ3Ux2ma7vSOmHc7obkal2t8/nqLSBKi34a/KA/AWorrxqpd77TS3p6Oz
4EFtm5nSUgCwhtFcg9+vih49IRjtVo4BgfFfBB+6KygFi9XMiLG94IzkvpZsUHbk
ciLkq//Jm+nF1M57aLak4iWj8o2zPLVm156KyHTFyrfv6gsiwdYUlWgqVGlP5A/y
cQfY8tedpwLT1tVTadDaMsDi0Nr/HzIuknR7ZJXswX+K+GpNwZCgDETob9nk5RpH
E5lTwxp2Ujip51hflafdNCUk0BsE1Wka7GV0PZnwwaX+ZV1E4wuOKtaG3R6TtTvw
UuTSobJrkU1kJUVupzv8BK43uhgGzqsihJ6n6N6nCEFjFOIrkJrzXUxBmjyjQ6Nc
Ei8lHDz03XG+l8vSvKwrpZzUHhPVDZbrRWOzafxAvMn0kPB17KEDobqwabpjAJca
BlZWJzDuYSK1plTCGrfdNmu+JthAWkg5csAVl5zzxF2udDoG/nKeqKsONftMoDkB
rjSTu+gR/ah/jKvEav/1TVmnw5UJURjWf7+7LKnmkyHJ6/4SxNU7UPIwDrcxlv+n
AWGQCGorQXXMPN+0lSxmlhUUiJk/GCO3app+UlddxeCLkBRovThMzTSzblISQmFc
cfkaUZkr+5IaTljZTy9MMTS0aUx+VC1ycqilBUu4gt4YE9yy8l9/K7/t4Rj5ku2q
kdQsG+iHmAOnC/uXl7dGSPy9YgQjMRH62h98acytvLnYGqEDFWb9ssLSMivBd7Ut
LaepsvVPfQvimJumFdlAXkX77ZgKvBtfkZILuxMFjs8FB9I6zzryyzXbY2AVA1Ea
1iWto9Rjmiz6ergf3J5RLekmsJ41iPK4QyCm2nCl8dTnrQHYcWWvsh9djthPGEYG
IxJWaK0WYP4uYQCRgLVm3aP2d22GjgVPKnXC9ap7PPPnTuWtxqg5LuYXYK2Klp3v
JDD0KtmWLcCANaNDQ+g6Q+EAC40LIvkGFKjGGCLXf+RzNbGbHVdxxq49inenuxOu
B3UcURIHRNl8TZIH4jC8PHUgzQE3AaP+y43ZwTcjrfNMq5x63ZzoKlhrHbBiPkIk
QkRxorc/fHhMlk53V5OD+FcgNwYvIlvfBc8tpKREs+GWGqiN1paVxzciB/GaDhHZ
uIADIXMaIUIxwoRAEg/N2WNEoGAUjoKKtLZ8q/rS6Rx//9ZYSQZJhSmY3xIULaUx
F6501AhkXVHiJigkV/Rey3RPRUPIOlypNDexN28v1LimFRi0yce1oXYYudu96UAs
1DzIwJZP7Ue7oV7sej3FOUXY/3Vz7Wfd+MJa+pamOlAL/HaKmBgLITpmxg4GxaTF
hQagsOAcxtUQxrvEokHB63+mWZkCaLu+fo0nDvNBezoJrlPSs4eM7vLQnKOoUR4a
XJ0Cm7uKXFehbZ6PjNa1FQpLAPF2OerwQq1UN9Y2xBJC9Rw4fr5gCiu6DIYfKVyJ
yf29IynF692WunafZporZudelh94iYUCexPXGxnpfeIAPrtfsb+xNeg08MriUEDm
0zdLVJAID11R2o19EYL5IKH5d1tPHe8uJgo2o5Y8E7nzyED3b0LA+56tJ/qfyqRU
zlvpWVXSDHBSbyNFN5KIIkVFXfur5cW4AkiOyacNOdxqDBaak9GMF0zYlt1q781S
wwUelivlKD5em5O+R053chiqeMh0Qs0S2iYentBMq8L4Q8m19FGM35c2PTef2AxY
pPE1eL51kIkC0yYy6i6PXgj0/70X0LKnRc/fJuDrkgkGu6sGjGzmFwvrfKvylgXn
/1lVZslOGlqT8oG1pcqrNk1tvFXHmIKYJbKOl2cuOtokELTgePxuFCNnTPZKfmei
48qxDHtbhoCn7gAWAxi1YhDvlxN8E/4GmPEAVqXfdOknH0tXGSi1WbljowY4Tvg6
dd2ZA6HcAn4zIBmRvLMLRLhENpTB7yvwShDVaUfwQf3GXvgQas9+6f5t+sSFvFVg
0dwNy9gkmFN3HuS53RoX7nR+isXRWrZKYGBHpcxWYVPU6zZuZJv/nj0+wBbEaBct
a44Qa/4c3GGMYbxlWvH22r65IzBDoMMogQHgHndw5m3mVzIL4BdJI8mWO2dQEBTp
YBotS4W0gJgZeNG3GjetrbxcZgfOaEvYtkKFrGyZEQlCTCltFXvQUqoNo1kjbWbX
NbNdqa6y5yVscIaN4kyy8G3cnrBJb5cPSVBb06KNXOFu4EZSDsJrFAcAUrVM2xDW
vjFRwKw93bwoj9V3RyOSTRZM5s/sD3vt73RcFXcjqLH4a4YmdBiBbx1Cxdd3jy9n
j1kHaINJ8L3XTYpZaYbWlEMORSeheTwl5S09jQBCg5KXmdTkjixP0dqpAgIgXhht
AGwnmKI9wezJqX/nXhTjfV2kPmFSTIvcR73Wn6UpkHd+SEj64AGMz72m3hAJjOKZ
qshFOZjp/5p3NzU9z5OH8jAjGTqpLs1Sqz4dV52vDWegHzq4+RR/3GGV2EXnoyls
CkEOq2xT01XCNLCFzwj+p3I7Ra62CSjcvKIlW6E/Dlo0OnmeR4ElzJpgWguOkcQ3
fRzyfwiuzscJI2fj2B6/AkW8ISX1zrCnS5VB593kMOQ4twbBQVFgnrbGkxQIXbwI
5cOmDkmyIDUa31v2YuFuCWJgwVP/RnmOzfSJNqkaWQ2qUZYUG+umxxwcHqrzWasU
HoNrbT93I5RYiqpsjSwX+qmiDUIm0QSay0Y37eHWjBcCSbV+rOnCHPBtwUAGSHAi
8dx4she8UphWGzLcnmFyvF+OoXNZ74I24QX2mnBy3k0R5fQ1WwVvVWTldwzav5ay
WEAnPTJvxamCh5rRiqlvK8YQoWdbVWTR/doRmGwZfb3XyvBxdqeVmKlh5sy3JfYW
rIRrSoMbZ6kgqKz0sHYFdOl5iWbzQzScS7hN3GT/bSzjrCDuHIKDFZavx0amlA0A
er5U3oQluIKsZu07qumR/0bku31ILt7vFoieRZdLuxOAOwN2pW8v7H8fgb9GmmdW
htUJESUMM/Gi4gJ+sFpn9HOatqUM5uJOFgvFPeeHxxUxgCgNhlKTn5W3LaB7LG7D
x139ARZF8Lfr7YjonfTDtuIhPAuQSv5N2hQSZ9pbrYSYe16LDHdLI91UyCc7BghK
xkm7eM3h9wN4CpmRSZ2s00sKlR7067drcrKnmiCmUtbf9VTfUnRMp1vUiB0svKt+
lac6fuEKJParY5kU1xCUA2ZWkkJ1soyh7XcpSjGQGs5gmLVVjUoW4bcedXqd/vvG
INGegardtsDsyzowO/Fh2RF5Zztf4Y1Piib7R+P8/ZdzyJNh2Lbp+pR+cs7b3tON
/BW9F2kzshEPx1bzYt+DJ9TLcBg7lKt5zKppfy7OUFZ+XuurJjLPDwFCK8dgB4n6
fDwgWQayVfOgwm9mKFAvk2Oz7Gzpc5YYkN/p1Wpw+WFu7xjmSQgxJ4oVRN7JAKfB
19H5DHh8upVkyaEjoQRE5bRbVQlXi4uwtyyO6ZJjHxpSViq4YP8VbZcDV+R4m9Pm
ggC9mq4vWVGGJC7dNFjFi6+t2Kt6Sb8uXIcjT9ZgM5IGKhu7yyLvuh6cDklrQ5zl
jDFCthlA7x0MAOaMdAYqrInchoBjAUREpr8I7A2yw3U1zQ5hDTiCJB3p78VG+pCM
lYJOg0uFqbvcPtbZrhrOtTnwKh65FEKlUoL6GZiYCLxOCIR3GpsKL9UQuXX8o5Gl
gTVlRSEE8qMdOjFHAe1Dt7sHnoogjxlZqeOzwfxNvbCvGzkhVP0JkjVGP3OFvT1j
jou1jdQhpyZTPF/lwWKKknS7vx3sJF44m+zo+4vsazxiAITSRaTQEThD+HrbhIVb
bdzE4ng5RZje8khck8B+trz+rXxQTBtZpxPP1nuOegvlzxIsHuNNbvR6gzQFsBam
6eONkSapQUJH9+3YRDrW5VkzdAT/Nr8SLQvZkdZfgnmnQE49pchKQfpf4LdNV2RK
lchHLwMBc0W7fnpcHpFe65Vaq6Em2rkNjIvlbn4F66jRD44urMWdsEXxyGPjIe9d
kc7Vu8/k87lvbSvPHBxw8AI7kR+BRbqjJ3+jfTy69dfBUxWwdiy9tZ15FhrXDyQt
TPT67HQc5prJ5vigCikEuzTVfQUSdCb+NfnGGSycRHmg74LKt/4M5uJ59EfR6nUI
Uk40SjXfNx7HSGI4U4qxmUDdRsUXj1XBFqrV4w05gYY39YpyhovY9N0GW7WgOw9g
TGMShFJIh+JlSGRKkdsYgJy2adjphbUNesBnyomCk6XvjjyaBUACkejYwqSuMMII
9DPajYbI6g0KbtPHZqNH2mUk7ag0FZqaLykVnhVdJrgSRz9sRByRA2hEGeaHxQJv
4qDC8mTUKYqKVKpCAmO7f3m63Gz/DQuxU+WQEyt/OI/X1ex/7mICMIiFnQN/1AYB
p5G5W06OvJEf61+2yhs7mw5d+sYLNVH67XWBb4kTB0FPKRgzXyGKVkpq+1NmKDsY
BMqR86femQvxfo304+N4fXqoEm43ysZxSbFwgCy3EFDUrtKScsZT6k1+xCJCsw6E
TecHJHJwOVovoMapvBS9w6JEBiBM3W30rdf89lCiIN18wG8kU2VhvlZyYCqZQZTO
S2xMAm242PUpzJMrNv2eTJhCUHC9Nc0APcrWmE+L8t0hNLzPIN7GLTrzXlh2s4R2
KG6LPi5oSiNvI97LUK9wLCqEi93ZRQ+W0b3xv4pYadkMr3qZBSK61E+wABpdcpYy
UTqFFA4czjFV5V0RS6fEyfwh5TvLcESnTzyva14o9NIqTw+iT0WUoDm0+K3jVF9j
bS6ofE4gg9X3DP/CASVe08xw8OKRWlyoadiBuJ0tza8+pevgMF8YzwTUrMyNMkgq
vZhNGCF2QKTVr6IY1p4EXrID1sIOOrv9M/6niwqzxAjwMfUfzmHNBQPiAm7XKeld
dKL4/hn0vTmGDsxVoeod3gv/vlgrqhKBxBPKnHfOr8OSM05DcHP+889OJ07WF+Jq
l9CfjTKeyK2cN7Qf+/BVR4qNVExLUnu3khRAZARFIdH/sbmVcJ7G+xw/2It+Mnbr
qd01y1jVtlizZ9wBE+mcryB8scveF9hOTaixeJhIH6vl+fPqgrUvtXhGqt/5uPTv
2lQ/JardTEuAsoydsIwhEYL+TyP5bGNDkxNS0a888+XxflL+L6o5pUHNevi6o0oy
FTeEUgn2wKb+nNGLm11wzqqpif1mPWi84V+Pz/V/r8jIjuRTDy3JLaSZ8deTtV5L
nZqHMGyGgDxi12okfsrVaZ3IATG8cvWiE4/btCfAyElR+6sdNwoLFwYEm12OZjOu
CPZ5kUnDHbOI6BRz+K0NEXOJwhhp66/oYw3dlatYyQOHyFDzOc5up4wHpVE/b8t5
HFLZ0dRmMGoaeArS9bkMNbdp1nDLkRsiAUdQyrWUXRsAQBsdJiaGz1RqV9En9Wml
s4R0ri1vCVeOikmhJ0yXO9+DTwLWQWw29Sa0/sYMzQNrsWAeRnjwGLNacSVOdZqc
H7tkpgy3+Chp2GLyEecEGS39TSGxZykhsmBlABBlJijanME33Zhv4mM6Xod0qaem
xKHPcIsgAFWNBTyFqtnjG6imirS2OpYafOn1URby+k6pv1NImUkOUuFthQHf6/NK
0gTU9c6ShCzZzwjQwP0DT3jGu+zeIitbyuRCakMPz1QRitqkAC0dGIuyOPVfMve1
1A0nF1bUKR8ikJH76JEjbuYTzq+kPGNd0fvHLjhPpIMUrTFR924R8B6xiHMaKiyP
TNfOcXA+cx2fXC0bTpKgakPvZYpIU/czUmbXWWF649W4M+cNbVy8VAsvmikNomd7
IVT0vbtjcjRsjfSkgome0+kykkF5pQfGfNRHs8SyQQF2yrPFiZAsIU6YgED3wvH5
XToNSi3V0sUH9glEzK11mvlPp557u7/HF3GBTfcNGBsErBUVhTX2ziknFcQlw2Ck
UyJZdzLacwfsA+mleLW+S0dIYylLZu3lya7UzbhurCxfmj9V1/jjvLtCZ9RCHULI
A0OgU6ooDrQ0SzncT69C/x+p29CG/6B68OfPZ6cFsZsx+xFcrH/ButFwSqiYk5x1
aAmVH4kz+Ync/17EkMc6dL7LfMUe/OvIM0pxKzKs/ox8pXLcckdmyjTCd2SXdSsX
sfOOXEWY85pJ3tDk3oYaT35jvczjg/sG8J7O1/IzhgYP0QRl1N5ujxM4p6Xi/pCB
pF2Hqia+3K9aSFbCy6iPFeVm2TvNCAiOarjvLwxbiNFw6VeLHfZ0NfABPQc8hRSL
fzU2Yw0ILT1vy1630EWmdBVkQZH62Q2tpHykRhRc81QFSBwaoAccWBgJi0hEjA4K
8zOdEeeZU8P5YZhKFzCr2eIs+V6Fa7SuTFJ4xcRx5YAQsnKtWHdRzJhWzjAcIu92
YiqoX2n9r8BYeG8UEU8+CnYvWS++3A2qhLSUSOoApPAPJKUNM5VuZYXaMZJ/oh7k
d6NJ6v3hpK7SaOm0Kz52fukBWiVeaaz3zzN7UO7gaGC0MeTxaWdpMRO/G7P1Wdfb
RmynzWnabn209XDpgvKZEX7zBD0BXUDBUxlsaJF1vXJaEER6UVPQumTTbYIWF5sZ
O8icZVvYLydEWtaMa1Pm9VYOixqG23Caf88uEHT8YRelYA7P8jCfTdasbbORnSTK
q43lV9sl7azObKwA8p/yZ04BRfKuWJTUQwNNo7oSbRVSeX15kp1xKDtiwhKBL+fd
EtARqVKdLwJrfmzA+gBq2x2Cy4eufCLot6XXGInUxrsX9dbYwubURoblDr7UeTlK
gO4rFbI28EerQWRPZDwD7mX6cY1Fc7VyTV3lxif7X7LhilZ5fwX8iKUUKSn76nPw
hp423WhB/JGzyI/pFQZgM6BiSLtvTu/Gjy2+ZjU44Ti1rQPtFOQPMRsGis/U9YgN
NyRBvgqsn7a854HeRDmfh04bdyXZPa+Ax0YKKLrcAlajSUrbT3IzwqcESMA+nqGu
UViLhjXncJu24OeFYJqGq7Y4AX+kW8vQsr7ctMIyJoNKel3LGI1UNsR/EBgTOwdY
ztitrTKP+I7Mrc0NoGLe9UbAf/r4LxsnrTV0+CbfmcQau795C3sMVsjrnyTZWqtW
NdC5nk6Ivt2CEAU+BvCgZBQ7Cl1zXrvt0q3Y/ps78RQy7yreYD0jm6vlr6iChyDZ
HOWjb9yVtqtyWbo+aE3P6GE+My72k6BMa+AYNkHLwM01w/VRRjd3izi2CuAhHaeH
R38tk1qC51pRw44HLeIs5hIVYXTE2bXwqw6Zl67bqgucVhE5D4/jpVfYgsd52uD4
vLpffwhXyhxbFUd7ArZeLOw7j7+7JzgBh/ZDdLJD30Cvdl3pyqUcnMBjJHPheQ85
hqPSdFcWf+LCRRGsGPoh6rM3HiJA1UBvNlTRh36kxD+fj+PhOgtXPHX9M7BAdDpS
6qu9cRCojltSJaZreae+d2rm8yGybE+DTHvC8yi3RxZhzQUj5AnGA87sL0urVCP6
AHvab0qYgA32IIO2ggQZxSitEjQmWtPdickF//nnP9l5/6wW1m4+ZpIiZ49lWKIB
7Nf6pYyL7OG/3eBNKoUH9n0/ga0NCF8OfyFGoTn66i2oprAKr2W1C99aFzC+0dCk
S/fTnDn5Jbhc3XiGjkLgGOLQNA9bmLzdTrK0mwqmydUyeeKF7DCVEkAGKLGvdKK0
XJCSmLyikVAiVvYWTCEQau9WTCvNKsMeE28522JMFcPHnXXvcLcqNhsCJR7zXq72
RIyuzCa25xcha9aT5dKjcXZ3cW6AFTOoWTKIb3tpedETZwMl2o6NGKJF4QRS2lBV
OpfuquSbHXQQX3CmpGaA42TL5Tip0icWExv404eI8WxKJJ7trxq83sNdKmeoQ4yd
ZZQ1Kk97lWH9emjU8YMw1Ws/+NDed72g8NMzh8l11K75lqgiUrV2kyYOUl6IVGwh
+x7pvKj8d0TNqNaw4jTtDQeeQGuLPsHiprmL0hxZVa7TEIrdPgFkdoxNjcRrf7Yg
IpL1ufSie/jD8CFrBWwsqJyRYi6tjdC+1LJvkuSkFHm0VhinjOow2eXeOtOJ/zuS
xsOBGX7VlDDfMWezoVCnXJSpcMQK12yqeMqxGQCZ3hRk4s/BDxnEmzp8iV/8IFmC
deamsSjPyjRZuJYJEoSFfRbcJdofxAlOK62B3BXWSperYr3ocs6Zp4Hy3Fa7OMyZ
zgEV0ObUWi9CUA8+IX++Hzism4cpRfwSvPRFX9H+3e8TMa/qwTNMn4wQDByfnwWl
TCMxtbj5dVs6JiqGZcW7vXbw1riqTpwbxRPOTsofTgEZdjVZyz9Bz/izSI8O+9WJ
uEGcda1rXhj95JJdV4ziBfunfXt3IHTa75uOsVR/1jl20betfXeCqrY++eDSxO41
P5vdxy7h57AJ5X0UCW1YEFpuQViOO47qKhbR1k1nNyos3qD04zGUHHmz5+sg/yKW
ylnlaTp0x9blqtMB/rykmWOLKKkLLMljP1mTSeynCSR6FpzOKMz33I0uK2Dk+Bvq
RGn12oqMtJ14sMgUkVWHvEL6uYTikOlXu4VTiSROJKAmqXsHXa3uOfro2Z713HRB
wQblTY9hSwypybmREqI8zdJsfqQ8Afg8SA1kLy47g/Vg1rAjqIEW6Kx+FYJc75f3
gZ2xp1W87CC6QwKZg94t82KFgvaxjw9wFUvenf2qqILJg/G58kaht5xTixwx0FnX
BS457W1JdmwUSAnZMrRNrqpiyNKI3sEVQC0VLxdgcoqF/3jOIvVUrXdO8lSctruY
1Qj4ugqCkonSoBYywEc70iQodIT/a+3WGAR/oopnUaxMMU40qjfBjbbrNFsICN1k
8ok/Tvfp4djRm3CxyCkig5iK+1jhvww36wvq6JKcP4LTSUIg7Kkw3qUTFpoqsrSS
6j2/w5ZM4tewNAi9oH6JevtyZMOZX3dLNUZyXoKb8QE+bkXPi0qpqRThPhZN5QLh
PKFKInHPFRmL/umG4xPU2bPkKkf21ki/sHpGgcuHQOSViP5cIoeWZ7COBJ9Z66Eb
Q/9exrLy+q3F6BqtfYo2mTnesjrKxAdw7BJkA77KBrCJhFFBp15VeaZUVgFw9b1K
lrhQHuafYLuplArOmqrrnY+Ct4IcjHMc8kT5u/Z/2wa01YX32Jr7XinKNrcvGcQK
OOp3TVd7VnNUmki4DddXmdl3mmsqJV1L7KYIFivy4wSFa5fXG9ITDnTcRPzKT/7p
vcrqav9rT0HWT3j1Lf0eyUoAKuCUMdUIUwA1XBGW9sxY5u0WOg/Om4IcBHkGpuGb
91LNWRf07cOLZvQJ7FbiDMvMT3KqICEjRt7raLpQc2KZkm5OaN36vNzN5OpfzMBm
J0v5ebkjIDpXFuUPsDFIK8qsHdg4JjrEOMtfghFUDSAolJ/p28qX+l8B3McgOgYr
2mcVRh0LZXMgGQ0X6gm4o6tktISnVhsRJjltuUbi1rLQt+BLLoJ0DM5dkOM6E6BD
gcOJqCJMS7OsUTW4dMpeNVtuieJsxsGYFGOjRvhy1TLrSnRILyWP59Osha1xTQut
vHPrSmoz2eWpg2BxlYGQBqDCy1hk/Hle8+nxSyG/PvfsJCU7DU/NKxyGKmsc345x
Bhh5M/nCxLSx96PuwGELmgT4YCud1/c42o5/ecMRRxFrPMuJSqP6qO/Ph0qoVi3k
R1Ca9/4Su7aiYP8ZFApY8A12GzD2DhQKg0ZDdXnbX8NiyoQAJnmwmDC9/fARcMzH
Ys5sKj5pcCcRIe2W8PmHbqWEgOGxY6pk2LXn37DSH6DeZg24LwqTW6upadJBoCuO
q7hUVyrk6m4DKmclhbHWyLoaz3EPJ5SulQevP/6qZJ3oB4hH9GjiF2BprZnd+jmI
JmzBlA/ojWT/5EjmCN8N0ns37dPXQOetM4e4wGQK3EH6nVa3rXxGYNLW8SUehAe0
wuG887YcxPBM2DPEiW7X/QBnO52rahbWKv/MiKZ3e9HE8RlqjNzyFx3zMjQ42/rm
glRVsMsUHmrMBWh4S9muku9/f5YgUjh7qKom+o2sJg9nabsuoX/vCZGzDpeo39r2
4f4/SHTrntOs+PaF5OlRioGpizam2ynX/yv2xdF6cWa20CAlFWmmZJcph1BYoe2O
mQvEGbApXsYptcCJlIgRq5OI7odO6BISvxCM8X/8jLgez0U8a/3Y1RsGqlNQ3/GA
IAFHhf7yt4uM6YKAoXYMYTEjasU92/1/GtU0JWu5EaZfm3dKtn5slpfKUF0Q/8jB
uqWutWSMDP9HfXzmlY4GIb79Je8kHkec4IUQjFQXmo02zJhNuQXPGKv8fNI6KBN2
BmSxiUDXVu5tc75QcCrCuJrR4p+cc6K1KxYrLSrIMXxOiKy7k6slHEJIpsJ2Hmgz
keUjyFEwb4yKVybmpvGgXv23SNsmY8Cm+BWp171Q/e6bhixxNZ4Dal+fRoH+Dgm9
sDgoDBvj/aabzD6Pn4FbEesSryz6Xrl8gZ+0K4NAbRFXwYP1se42f+z1dl+QCgMF
9RPoChS4qRUMhABAZivXAhdHTW38ZDItFp7KJUyTm2oMhUYrW0V3CsxnBumWZhF/
EJnMkzCDdUDvu6jyrb0C6FImrP2lCb+Lq9Ua9UfTU+Y7M0CeRSNuPEwmAJ22WADO
xc6bCkWGFO+e2cSKAzUtZxhmF8JQRm8sshb5G/ZSd/8Gdq/uKIgN2qfDrStX96SG
5aofRMCkSX3iBx5HKW3On4OAsGoEhUz23AxvDxEjNZNnGWR11O4j6xXohxy9XtPp
2gCXksD9XMANuHG3+GUGMryVLGHCiAvvf5fOMH6TSxr2+HVhevmVODmG3K4+UMkP
khUR/DUzZ73gt/Nc9a9xlq83WtHamRAtK6y/34WZOBvnckKujBcaekYb7hsiblKQ
W9rBmwCILPDtgfj8iO/3lDoA+3W7jV1YXfBm+UNa+If6gyqWQ/CP3SDkRe6Goaed
6MWdze/VmMoYGNvFjGZziSAWpMfZsq9WleidOZpGj65XQhNyF87UcxZ9CiRMhuNz
zMpsS3TnAjhXpA5tXNzRGVV641xGyt4JZ4c/KeK4He8Dm0n5rGYIatEkwW2xQp4q
DtRXeN9KlLA8Il+GGm8TMi3kuT8DEqEXoiXtOQNexlK801N2t64TfoUpiRlNeG27
S8an/FRJa7pS6WEFUJpa1D9WoW/DI6p7ZmNnshJpq0U1VDgHCyuyK5srGeUbivkQ
/sanPOPb/RFjpofL/9dJN9n8l6MKUA98ODF1iscl/e5LXxw1YiFTEPV/fT9T8zHv
lhmoiAQhXwOFZSxj34QZCsDBDAxRrPfUpb55dv6hZlqNSKEVXC47fZbHFaWMxifk
q+ftW0VOzXk4XES9v1V/bJrAJ8q3XJQISu+IMLd8c7+QO7LNYRX5Dz46tHM+6MhE
rQOjTyyBS8QxAqVkbXpR6/EULhB0cVjZ8FXWiN89OasRR1kfjOs1H9lsnmHWVK2p
nAmEpx3NYn3rEStDFjYxGV9qg2ArmMSjV/4HkysmF8xMMqmxuiuMiT7vpVt26K7x
CMUnsRgg82esmJ+rD/iof3qLON9lc1UR/3OSBUhbIB86gqlyMn0Prv69gyrA+SZ9
lt0AKKof2eMAN1YnrivFnMWnDtiNKBkhSG0aLsuG7Rh6e0XaKtdDouHltCpkBjYR
j4AElB4sMhxzqNc/jmyWpdlc5gCh3P9HFV+AgioDx0TSAn7yn58XjfUTKt2ulol6
PWkaziEUYXsCO8oj9Srcly6ya3yPeFx+dH3e0DYn3Jmb2lgVCxc8Rb32wIMNsBwC
U8aqT9JhFvKeUHscT04M1hr5nTCrO1zt0L7B/OEHAaDCVNtMpUsEDqV3TvlVOTGL
t9yv3MM8fR9ELDXmW6Qwf0g3j2BooP9QFUQ7b3p+XPajQGQscsJ30F5LDVDLO9bT
yRT45dkLTfAG6Sprv//VaEMfjFi5OBVHAYrmU5oRy2QZMxQs9G0rZuPE8NXYiL/C
ePSTCg/12bOb/pPOvOfKGxu/nKI6g4nHTra5MdXDvC0dxGAYzzF1aFMU1+KnriL3
BW2akiWdlmOlI0tl0tj3YWYOCZu4U03K3cgLTZNHhfRKUNH2d/TWd867CzzWEgW2
pI031QqpbtlDROShaCgzZDAcY32ILuI/yUsfe6+0WigHHEHgvX9xpal9me74SzJJ
e7nDnWN+OLqhntKRCbgu79/LKRKhdY8ANjgToe9rTAj0fyUo72fh+EweF4DX72pG
W8l+9QHtF+pLxta/UZ/r/kcJHUCbWTHmuWynI3UjowqICeQCP/RJFGB5YdFnH72l
6t8RYBqpc5mBE9yNGnIYJ0O6i2A0RfSerxcOw7FIVSAc9OjY9OZ+32P6raMZ4qKg
UGrDSWiTBVfubFKCyiRMtFqQts0KPqwWYny6ugrmcmgnmuGmzqGzYx/vH+ChwRXZ
5btKzXr/uNz8fgtXv4NBlFPm09gdZdEFXsOfQCkvVGrwiZdkeYjNJD4NNKkhvb1M
4jHf0y3pBz1pVBiHfZzzvI59rYcVJE9vCblL+ZG03U+7Iwl/qUqNhe15tcaj0IK/
KdjdWP74rdgIeDYPhU0lkTc0omhoBoVxbM+exAIJ2Tf25ehChWAniGCiR0pzvoZy
EPsPffIfieNogOK5077G+cd2xUpJbbjmq8LBFGPLyQ6TvBe99z+19DL7jX/A1Cm+
INQugCIcydIlZfOvPAm0oxvB1jD91SXJN8kreGOCWAtGZQrTVqhfWEl1vsZEzOxB
pA44fBafvDbcyLI/yB7uFc+nT0AHrs+DoK8KRxyTZhm+nEMJIjcsPimwGvMQctu4
iwqcRWfNyQalijgJRwvbceAtijS/9LVWmshG4RDIfg3qkm2rTH1HNa0WuVJdX0LG
mpplIfKhLSwJCJD5BmSejURTIvroh/ymUJKOa5oU+mL1mrHtHHJpD8SUYwvfB4qr
0GNaVXJ/Sw8sA8NAHtp3XVQ5/mkw7rwuFcqQ/OoT0jGXIaEDmOqqs/xjb+Vu+4CH
upXEnPS6dvtF/2gN7X2Ec+0tRrL5XTuobJwe2FM06LQ+1SJiC3TmiD7ZLQzwW0I7
XryUxNNs82csAKCcZqBVZagHloFiw1rDcScfx70EXfKRvJFi63bSOBjabZUIXph1
nWa2M50v7woeQLYNbSkp6BmoQxbwQ4s/H6/knkIfdXU0K0NVN4cNdP0sm//3ug+v
w6LY0tLjyWHMkKSe1+x4EqKrTrGrn4zDU0fBGqd/BEGAYNq1al+TPY+yOJPAum9a
IvUNJtbV2EzGmieYJduvc4m2ZUIj1kuldKaN/YfoULIuXLFAE8pzxtV3ZqIyEm/h
7DbAsMhFqhhgPJ0ZZei/KJraXCd61+dADKbsdAN0IyRX6B0BcB/yqhNcD/oVdKdt
FqFWtyxGRgLL5l26uFzLsZjj0hfDAe8j5YutqjG04ZXcYxGp0CodXrtlyZzXKWmW
8Uvj1waz+pEK8jixVBYet1YqedyXEIlefb5oiHFWqac5xJpt+mFBCOMNp16idXDX
eYBivDhVCk6s8eKzIlv60qXV8yYunq4g06jsqjjufN/MI5FRyY8LDiBCBTiNnGHw
U6a0iuA56EEuk+/BtG+4G3UyC8FC25cDEZXUseezVjDQSkHUfh+18TzZqbx4MkQ/
T/OR94g40B0oLWwb285t9e4zWFLQys9hN3AkXtRaAwj8nil71CEeJ+ZpJgIdtO1p
9oyF2b1XyPYJ/Uvsu1qntHrZ7nTkE9fYBsALPXjlXPJ1CCuYDHDtEAfnNSxmaoDZ
mik4z56qEC4l7/1PFpM9Bfaw6YYWqejDLcGxy3VhDn5JCz0qc8N4Pb37nx7mTcbo
ivli0hLiBsZB0ZdJwakGb9xOhhs0oHssF8ApXnEGW2SneWVuTSlBYf1nFXBeJfuy
xnmANLw2pKc9vsqMilNXnTwHMsah0rHWRzYbXbfdsuxK8QkCYbp7YOACAwq2MeRl
MRK7mqeyw2qmPW5vtkyCpjCqFWmxxLT8UIaGVZl515iLSSJaWlj8irW7w32ghRGe
RvKhxbWBlGC78KkLms/5ulToZDazQP9PxXF2rdcb+yUqF759YA1j+j9E6IEWGfRK
PndNxVN0Y/T0KCHXbFDnjRzbTrHJHjKZugD2uXEl+1OSmP9pzxWq1c+hncbtlPdv
egGOzx88RJ8au5FdzwAX2NVQSzeloQ5KeO1rtvSjvfFb4L4IWp21H/XKciGLe/AV
gqy3uMi1UZmXpmx2ll0pvJPRIv7c4lT5liz1Yxl5ziXFgqOAthTX2BzFFKD7e85E
YSnAN+gnm8ck3UfCIPA5jbzhPYonnKoNTNj9Ir3Yu7xKSwGRct/dsbIfqCV5PtJv
sETwwMmBY6IlAqwberDiBtbiWwwxH4eICD4IcN8clJ7ghlbAFr/5RUHoPVEt/WEI
OiRtFznrj6rYSx7+Eqy3jb6D5hZ3fZ1XV15LVFTIErAtOly/2iXr+kiy8fhzW8ld
Kr76isvgTEyMcGJxlPvDmX9Izrlahjz3qx1JEGbTU5YQSLNeFRsCmIUMrYICDne2
BkmveFgNgbm9b6UPnuo/H9PdG/r+LT5QMdFT+GS+7sAA4OjCTuw4+s5NrRJcukrF
EQ0oxMEWnKtFqnjkiI9d8mQRJ21h10qDQAe7nn+Hf507UXaKwwJ5xPHNsueRXeCc
STX1Kk+91CFbdanRWYpghjLT3E4dOgOqM5qde70k+4k2bSJFzJFVWIBP6wKDz4YE
xGaMt0TM5WBDi6/UBTps1lWEQFYeGO5XHHuyVANxJvDFz/GleJPOJv04IkJVsZZm
CXv/Tpz6ZurpW9xNQa6Ti6tEF6XPJdjC9y0aXwUc7m81it3JOIFa1UgWiQKmC1+O
oM9Wa5P+RMTGK/xO2xijP2+HFxky1zoQcxvY/9g5w2Ola5Ru+Nycape8xvwib5U4
cB7piuLW7wE2WEL5LK/RnlBEuKQX/wmBBqBfgsTlZe0NqSDyKs4p4zfwUh6ZYBV9
yfFP3/Mk5I4qhqtA9EAiZ6S8wq60FNqCZVaSoLd/Akn6MDcISP0yjQb2qENnWqea
9XiYCDt9gkg58bmleEzQxQ1P9D4bk4G8UwbIoLwcUlIKvSbGwAYUt84S3xzuuN1W
gCj6Le1oWlfn6jSNoF6cS1ZlAGSs03iLv2VYeX9ScNjZMXEmaIraIR3bB9gyKWgE
jqqKkzmqC8/nS+3IQ0dHMtKnMBYMeuRHEwPrUT0+NZ7IDF0k1+Uje5ChLtQioCz/
OEdz4UHShWkLTOTV+eqpTiMY4F53euRmIabqN0LpnH5sdu76GDmXWKIC1rn4YnUK
PfX6grIG5DfXqcT4n+Qw4eLUfmbo5G8OtWWmIKwVJ7mE9JRR7n40kEbemVWwGG0t
lzfKpYkfoWCVM/S3mBNcXt4ajjWhFtvTHaEWIb0fOOmHiUA3IcrbyGKPBUE5/RdU
Qx506kh6U41qCemy0AZKAPPH2bEoA5A9C/J+uo21OhzyubKZRzRZKIzc9vu4QwRr
dFdkkrOGcBf5FInm1dCbsWYqwC9oGk3y/U9NQMuiatYyV80zT5WlZ6xO6tEAXqyF
oCEuW0KfFKLPuFSr+/83nD+fPPJAT+EYZKV/4p1yPx/XAVRYxz2c3zP7l690vdDC
F4B3QGInqJkoAdeUzjN9m3w3SMn8qDDjOSdyAfEGFCmu2vQFJYx27jYIxioYp6mj
ZtEgbd+/HOfB+PxeBB7Enzrb/Wjpgj2+m0SLCHZZwSzxiwt+Xnx52OL+/K/LWcIh
rEMFqV5HlXCAnZT5uRLihDwaaJHo9h3opKzK5tXAcOvypIQBUJtspBq0ElPLP4wa
vcADLWb7dVEfFzULAoG6f8qejt3ioqxTksvp+xnMKPwob+aLNAtMts/NQ3dtI+Mx
CXaajPIoK3lQQC8nFQ1mu69dzpBocZFHevvqu/XIi5LYtSE9V4JztVWy6sw4r1GP
It+z7e4KCq3KjjMPVlViCy/mTl1nzQump5Z0B/VR0OSwGrLnkrjBFMeXaeCNCv6O
V0aMs2zOczvcJ1hglG+7Wly2dAkb87m1wLhqjJqqvdGuybdzIdH1TXc0ru1hhgzK
NwLoPAw4ugkBrc3r5D96ZWQPNVZmJfG1N3GXbWvl9icodHyocLy5YtT92A0v50jO
ETUV6kV8KJPbzIDr9jwiQf5VpYObQW6F1c3ba3HnAvw9Lys/kZz38H4IS2C4K2yn
9GmPGzHRCnQeStDoNNYnpdtTlt+JFXhjTEhQVZRKT0wlDwYQ65J19cSu91hnTFrh
GlLy2etM97yD29uZ/CzZCl/sq14kXlcMf40kHiVLtKSokDnU4BUEk7jmkuOLX188
NfBaplpctsVXBeTF9NZ6ltWXbywXukg0cmyid0s2nuB9Q9rrhnJtsnlAipOkWzsE
hec0QgzRF4HEtK33dLBuenKLU/WP6fhAMMwe/+TiQnKqoOQqKS2pQ0mltlt5wdCS
Jr63kyJVxSAEE0GDGiSEuJp0eAbkIPKJ2VE3droOZcB5ZlJtSL50CZM02HgpEtFY
OnO8kNHYcdn6I/EjqmC3dMzdpvcHEjfVDJonQQMdaHmj6zMfxD8na/jp1Y4BTaAN
KiSCD2A2he7hTPhHDm629//OTiBiVYcif8wbR2ufMZ4xsKIcYCYJWh+0YGvX9n3m
KartFPFyiBrcR1F8WGzLU0vkgrQIdemDns/SHuB+7NDki8ccnPJWqXhHAJne/ZGl
aPgyMt0CRUn7HY7lnTbTp1NTF+nlYFEaux4R1DDip0j7xCwWh3rpzyrV2eM1UYBP
fdBoJ7mTf7xRrfM7R4GovvhYL44LYSzleA4wgljOCeBxHFBC2cn7QItNOS+XEMJG
19Eyw4jDGNZAdQDoWKaLSKo91XrFG5UHSDGzfhpPIphZs1v9MUzD/uOBH2t3zva2
9S+OuZe0gN/zRnp7uf+cIQTFKf7A+6yLEN96IR0MxmR8cvgCX6HwQxSOzMnXRmlt
ZWlyR2G0t6aDkk29QuUlH4/4WtGplq+RDTrfFwradF9SkYfCSgvv6bgnJ6mQCTSC
QaXMnTau5SuyDmFvG19g/RfrgT/zN+8pzwqRV8DF7NjL5lQ3M5KbscmbouTrCeFt
2Ej/1KoJc19zSm5KjC8VpVuf7jhnAXDFdCXNMpAEcB++/+KX4Cqc3eoPXkvkaDiH
EvJZH7GiltMrjEjFgHdLsT5XeO+AM9Zn5B0gHXqMZdGc33FyJqLviZLrAfVCGFAR
qX7V2wEuSt5o3vB1K9Ah1gr6O5cLBXuwxtfsxazU/UKWlZiaSqA0ZB4zEWKuWNqD
K3486l9mG1Vj4MPwoqF/2fSb8/In8XQBTSO48mBaJLQR7NTBm1c1aaCOsk3turvO
TETuZux7vgokpeXpRSie3FrNaFc/Uuujb4FkAjCgXbaZ9P0kNupXbXzBSTMDRO0m
T59P8Xpqpnk2oQcJBThjt5yPpTnnlovsOl3ymoCkbW/eejrt9hvdER9f6LUkcoL7
31hBYbn+0PZdzj/7pxejlBmluX2cKyAkm9kpa1/6B9exxNefoI5W1/lAd74Ro2+k
LPvSCjxZj+zzrMThyniuuetfLHukEs7sMmJ8I3cqBtgH5Hgq1o1+3LMORTtizBha
4sAMCfDSx8SJ8Zfkeqq8WCkNEw4frA3YGCZgEKLkWZxCoc2Bj7PId/funwigjeRM
BdDm+fT7reQWu6qbl99EiPE1bbXjwOw232TWrLbhFWItiKCtYNnNEhrD4RcrKKYG
TuIDvIUDjgQQyO8LDlaXlnnD5hjRaKxBlD1jF5uQ+Fokuk3svls4lGz31v5MRcIx
nhEmJN8itXUb/Y3OXdVQOb8BMvsBZo4vGMdUjn+PDwtYKqBTeElQWzpnohICrl2V
TL996+Bq17SzIqWjKhHFfNylUGVBo41Vzrvtb7f22qHIxu08QNxhLVhICK7A4plz
A9zS2lGJT9IOxkIJxprU3GbgY4rZwtM/axJ4uS0q2/kGCjwRvr4UxClAEW8135xn
d6CCbbEL9Ir/fhVVlMUcCsCaJknyNnaG9vbyGOXBi47DgMyh9fc9vGCN0ZlKPyJZ
Om/+wsIvCwc4Gy/HWvgm7VJRTUbntKpcXhktruGPaVHZJDdZQnuhnlVApS6QpBRh
IvVKwX1n51gexuZbHyHTJ3MM7UcMrIK6WJ0UZBFstyKtvrYW1uUxM9HncpqiFCLP
IDeBezLKZG2eHP2kl7orEyZnHoC4S2jgIQ2+U04KcUSO5Ewd4gDlwPB8wHaunVbk
d6lz7w+Yo1Wpc/nwLkV55/1JoPDABulwwucgUrL6veEQ6DsRuS5l4cjy1sT7zTZ7
xNsKQSjF5zASX+9BND3QA+g1GTiaGK6FwkzewTlETjbg+D/uhg99I+XvROhpW/KX
InMvZ58cuPzhtUGalpK3R0he56Lt0xbzQdU/uLDsSt6RlsLjGU/RXyzrGpuKBPES
CvjWLeqw7a15jE2QNuV4K5juC78OsvdXxAzGKLsTptotJoepnJwWh0JBQA4Cwe9B
BKyFJlzxwRA7WeLYxCOhg0FxIi5oqOgKjl1mGIRhdEJQi99GbtxRCIAj1IBmeFV1
0G3mO04pIF4hOu5tmHCNzkleLNYkDatypks5HxH5JyKnmkVOtoJHfAG/ugsjHjYn
pLHd4fHsf1K1jqQ0T5YBdjZA1RKDwi4Xe2U3uamQRP7phTVKeh46YJm2ZanIhY7J
bxSk+aFTz2UJMAHQLyIWlNhLuE6FY+8R/0pQzbxQONfvhIYyMqjR1gyvv+zoGguj
FxhTYoNJ/oPohR35oVxm2YzhfFecervCZBTLjXyvpRH3gNmy5EDQljuEObId+Z23
3iGddMQvIzjl4690wx0KtQKzNfiW+A5cM6LhLJ+F/4XbWF8aTilD8MQG1ftFpAG8
a8HjsKisvdL1ShPdb98GJSb2wt+rft+9UU+v7g3EI6NuWUsL4Q6SzKoSlcoJPwY+
P+BLOo2KIPpANynaqiWgomyoTxvKn/Q++eqaJEWF/6J1VOArWNI2zSf+zyHt6+sl
JZwLVNoiH5CuE2pCGgaBhJAOFjV2mSi7PN1a+UfSRGZIzrVnqPJuq2X3Ryh2FLFd
HOZC2/kVeSS7OOAoOIfjg5OyCmjBi9YAOhR6kyEGossardQCMF0j55wZzmUqi9A0
bnd/deuLUTWf2BsFebedxci6O/VsYorSBEGMXFcgCi0Y0dETefNRG5+06iTvgWKh
+sLILPbcvBI2xTlkVG2DE9Hyolg6WXkQQsDiyBrRcbWvNEk01Ky7vzwGmjGbQ5DL
xgNK9kW8pVn0xvS8sgtaiyqa96B0GU9Ycevty66d507wPCaGhG5QxNRlkw420TMO
6vkvBnIs1Hf7iOFaWyBh6Q5fMCrVEkwmZZlJguk3HN1P3sWaGFE+S8R9VVmvPREk
qEwzlXh+fRy8/WSypf8A8sEWNk156PybEy6m8GPWmnPAQi/XF3zbkBl/8wWNKKV6
zuJiB7FGggBncZHqERaLCZ0oabOoW7jX0+7iqiQ37iaNA/iZthBSu2kuT4uAm7YZ
FHKHnSTPwvqyjo/ma0pZCu3VlVNMnSvmFHfmH7QvRySO58V5tC4CRbq7u82vx80x
5u8XdaMBIafI2QjGY+oNft8UtLJ4+6VpyOY0oXF61Ih36dtYYvyV34WYBzsRE+aS
LbnhP1OndHlNp5vQkN8nIso4ej822/CAO+boSHjhLnkcK6Xqx0qEFg7E8BnPgxxN
P+xK27l5VZpx+bj9Lt7M2K0MqnRlg7+5tPXQJDeu/BgpT3XcvzyWtu/I5thvHtMw
SJ+2XKu/O+Ni/3jzjug0PPMtG+uvDPf1y2sWU0eK/Os8h+VGqwNx+XBM5kJAodwo
yClKhd8JTkX8xZD8Ka0Q5vd3n1jmVuHaChSGmBKTL2taHg8QnRoqzY8HUaoXNJSD
uIwb+Arb4pb4Uy7Uz4oE86fRNDXmbr7FrzDXxnwgKTJyUEVER8RIG8AeOmW+T3IP
ZpUahjxYSPUwsyhPVBGPEy91rnKTM5Oxh/AwKJn+pScasXY9+ATzF7U4wMwcexYB
64G8fKq5HQxqZxed28BxiamJX2wLrECyqbUtLdYwAtEFVRQiYE8GMX4xoKRtI11R
KZ8KRDZx+a2E7cHLfqyx4+2GdCe4VLZwDkQG4frTohEtKSJA/G/FX2+YXICnsH7r
tV9PJQtESn4fnkAmyYZ3o4NErZ0H1pGBs0k2BsLMdDMj34x6ZpjeKR4TZSVt8SrS
TfvLsjEb48IGysTAIhxuWHDgZk5jd1lJtEcwoTjLetnnlXTcWH54ORUG5wWpgmtD
8YdrcYa3yymo8C54Np7IV2pvLcy++6+gh5RSKYgp/K09WjukUMtZK9d898ndc8Mn
NNJ9V1EEyOdfnvaDib7v0IR+DpL1j7b3pOMSvIecerso8U8mwgumlH4k05w8YQ0L
hsTSJ9SoBjEQtNiEfITCnmxAsIgrQ/5MqwZwKDV0KD9Uie4AxOKCQ3DmwDXLJuhF
4KBfiOCpppl+Oa9Rh63G2NBvNtOmE+UF7gPGIbr3I0Z8lORrPWcLs1egozDp5M30
3zw9cHitpWkt+gxUp2FKyCjY3LhLAhNkxyFKW3+VNOaDlrxh4JBwmOlzPMlnvNvd
brnSHEtAcLeFJgYobHitwXeMbtZgF91/XA9o+5TyueVazbOhUCcby6zL9M5q4/bW
th1hH4gIs2q4SxR3Ry1bysJxC1qNuAl7/jzOoG4D3EmwmFL7XwR975tVo/xTzUUd
Mbnsc+0z9QJuvZUmIe9t3xKTPi26vXBUQer7/RXNJziGJwMwpjdP7/9aQZoMNdpY
RvH6lXQbPIZ/+RIpIgJL3MAZZxhEsyHtttqYvV8WdP4w8d1TZ7lY5Msof8VcTmEg
5dFcMdloNfsCh3RPdTxLwnzN0qGyiYzRNfdpmJsbxoNOyaQ4ezetmXcobG3BQvRV
L3zz+O+pttnzhT43LSJBMyWLBsQCo3my+1bqoxW/W132+R8Iq68SiyI58tJZXrQN
3G0O+5U9Eei+NZEC1o3cSeItlIVAO0fQUOQF45P/7fVxbARq1R5DnrMuA2xMdRmn
eFb4UszmEJlVRbpMdJsfgiwoZD+9sUMozrA1uNIS536A/uzOJdZw/xbuPyhDAcbc
8GFFqHZaGpt6+ehC+5F+9pqM3Fk+DQ+/pkO5uUJt65LOyhNuJ+U6SwiAVWtSZG66
+oseXixby+nHhnH6RFSkWhhyit+Wq80jV2bKAjaXeGuGNtaC0Wpg+BwjGJGEDe0D
c8gfJeiFaoU6BNuLDM+efxJVpHpGdwn3+skklNet/rGjV+1Zi1NNRMXO/4dlvwgX
vDOEBeFNox7QEtwBoIU1swAJ4Pi/kqGlx6po5zBFr1o1+LgAb2IukonGl7mjXZbZ
aWybuYhZFccO/GWp7iYCb3iqmPxAZ+Pw0qnX24gkC8C5iNQDpNYKoHMsxAhdO3xS
NRunLjTJEHxelhmVgVSGRoaVtpvhhczv23goyxBXJQITdp5pkOpt+dOdhApFj1DL
CsYpo13F+MHoD5PBSrj7XnqMelew8tCdrJeeqbSfuNPxPBeY9qnp9ozjoGj+JKd8
B0u5MyxAsueAfBhewJiXuIFUYZAsPy/ALViyEILDisIa5/cwitaUsPf8QHa3HB5M
gWbU50Kc6aHsZin9oRorkaW+K06udeQVoAo+Q+EgZv4PpJ9dvfyluKYyIPQfc5tM
4BpbvIMmzM32J1rTxTepyhKGvogd6pwiSu80augKqLgb6rJeFuk+KlllgXLV8t8B
sKxDU6ERptwsnDpCH2DncAZnSEySfTlB3UXll/4GiacPBYySozpX8D6JgluptxpI
U3FT4GzpDP4ETm8fbfvtNdi+O+8fXuzBLGR2S3JNJGB1B2txH/Ss3AhbmSVRj8d1
IzYbxR3t/sgU7y2JSm4m6tE+QnJxrPWTCEchLLqXpvDRlRv0cyjv4RmXrWaotfw2
XgIlvs6ULBWc6R9OJYvxB5Mi3DKPiXYTV6vQAmFPGMQyZavZLVtoKquVOICcfHJ4
Lvi4kOHyO7xjgsvy/7uiONkr7kZiq9RO4AClw6aBqe94PzCEKv8wKiPhmqKzUFSV
7fsp7lHaQWt33OikRo4SEmro2fmM077Wd2BFz22iuABw0fg7hPpUBOAjzISMaAFR
+9dg9d+qXKQCv18NsvpShPNGEInWIzNsohPHk3ErARlH7Xez48rN6FEM5IKBmBdu
XMxzCjOQonPDeYFB8wkTDz/h/k+hA1R7X3R1h6ruc409SCi9StefsWRBaxk8H6aV
WAL7AdWlaWC5HmTBgWzFRhuwUl7yUppYvO7Iadp2aMV47/CoF/NQQ2Dnbjxwz21R
5uUq2zdWDLxQHe8hET1+/oCm1lEgXXoBwPTP5O87lC0YDL54zOHOTAtUqOaurhMw
nRenpXeFa9F0+ZhxFBlZoDNsPbiUefN9dIA5iCK05NVnWsmQxKpfi22v7TQQx7Fo
gDZ5NvFud4uM6IJuOZYYDMu8v4r/xmWBkcx4rn3o/94Atr0erHsUktGHNgLU+MDn
XuK3OyYJKYAMOVwUdrh2FfE99qiVdLqqYbQ42/EfQ1DvIHQ1fzr2rUtqYgtJ1IdC
VeR5uBZS44bxprXHv3M0LHtkl8S7sLwmwedCldtO6RRgFyDL8UgRlLioyDknycqU
YQeBs9uDGyA2sSi2eb4cwZhZSah4Gdc+y/ka1rC0CE0+bN5y/bUTIW9MSFfE/haP
RoXsp+cIupP8dTIRwnL9lxVJXuANLsYLlvhBPw6eKcLY/DtsXeqYbMOcAYwcAEuV
L+FTKFkMceA9I5jxpeqpkhc4gNxA2OiQtfzVBU6lSrID6IRYxM/AMTyFcwsBiKs4
ILa1ut0FJgHn6J5BbW42U7syTXSuI4Vo6iUtmyL8XRbLV24LyXmy/4MCYqwTixxc
h1hBWCCbDgBwdCgugmJZM+fJa74gfAF9e6eQDv03+neZjQrV9cjyy0mLl4v2oHBc
XePeRo/MCNvY5p+a+tXYFXPZoFc7BVr3kvf7NSNTfjpB/q2iCom0dlr3PAdpHbrC
fRM/AbCkRrgKVtw0q+BVHnc6kxjxuhXDQeKd18k77UtoBYVxOsMlKxGS7buCvsoj
6+koY5uY44rX9OMXXfHHQEhWDX/sUp0zTmsZTwzu8kS6eIggA76NNW0T703K3hPz
ApRYZK6Emjms44KE7K7sGIQ49rb4FTeNqdr8im8ysfJClETxCtIWh003zctBbXWY
EbB5MKqc/WL04434HuPc6WFESl3JMo+QHMhr9MGlsB7e3/gfAv3t2swpT5KbKBV4
tW7/yCVhZTic3TYNhHL+XZuWl2btd/mh2/R4Oy8zk+aJYrPysA90B9sfV2Q+h/r5
qjvXP8724A6BrABXi0RtPlBjtFa0I4xTX7HbfVUVnfGrtF0g1Mkq9uCsd/l3tiKt
qtaFvfq8OtSJktbKF6Tg67Di3VD2gkR5OWuz443IhiCkBb27M06sLUoq7MpX22R5
quYFAH8ATPWpdM3ZtKECAUYpIjz49dDMkBeqtBaeIr0HF4fyStJgp6ZCnJKrYwDI
4PRu/7MYR9DPws+TukfwMBdiytJVbrwg5osfFYOwp9v1zLokl14UuUklqOFqrHhF
SnCQPYZivq/O6JizbY7ccTH1VJovTrF8J5fJhwM4pJ8BUxMbLYBc0lbUJF58dYr8
obfnCqS+qI0TnflhuPwOEtfZRQlgAhgqjNWBnosfRK752SGO0GRIU6I4Op/uUvFX
rFUNL6aSnrN0WCEYLCkB4cgW9JFkjZSWhIZqhJ8R5sEe0KFeCpJ+pwUP1Cv7ir50
C2/NPupiVxL5skqGKnZOiHeD7JRRBJQzzEBYtkdZfzpjNTLH5UfIzh4Q+LY+EHM3
kr8GFphNwruglInB6h2iwV+DduAOq3dz2BwpnS+n59+lXuf6y220INvi0F34Syuw
r36fedwj2rzWL190IWXZigUJaxl2BBxyUKFa1W7jZGA+u+um354KhzCAka7Uoxg4
BbdLTHotxtxcYNpjv0HVfo8hF4YyvgPBSYSGHusHKQK6qtrA6wNizmwtqCZllYnu
igJwUKPEnaAx4VepVi10P+oMDJwx39gtTmWRtD+7NWCg9jPhLnlbvSqZQKmDRedP
JlMxxOPncLlCzTDzswfhP7TWM7/SdvT8qN5Enb23k3JK9CtQuG8hJoLYYCjigJjA
WyYy8LF4oYrg/Lc0IF9RTnosdvzRoN54ZOMM5Okc1PqvX21CZuQvTAGMfa/5Yv06
lSbCa/SCTIiyETc3d9eGBHVdt4O26VVCHZShKyRCLtHrQ7+hY5Bjy1u21ga3jSh+
d3H2LFdGikltsnOv7Dp/zNV6pQtV1ETd4kWx1mjNnfTBVFRAvF2MZerOd8iIkERJ
bYd4ifsZ3KpEs0GeAGUNWN/QnHG5mUAdTkZV7PgqM4Umf0WHS9qFxcbyDwyTZz4G
AZ3OJkRUgCPMhqxGqhBWB3IA9+miOew+Cu0mw1K/WG4iOw0OU1YwCkI/zDUjO/8j
8otY5ZNVhFGaxkLT2CXc4FBdkEVxpgDjDh24rEcxpSt0Aexw6wcGU5xbNY7V8pFk
2X8SeB/WU92wEi7+bLRgjpEFa3X0PTU3+4NNB3dBYSsmkIt6RWlumz4Wi4EjgYBv
vYhMbtgjHtj/eNpJ9tRgcRnCa7BkIQ+Mq2VHR8MnP1x5Yq6HXbIDjINWzduAUs+e
aol14ZeaEqF8S4JfLNWjnyi8N5OAVLe8mqitCRV8SVJnktHCSu59eR9301ebLj8X
wC3Yc971VfdVervMRwcq2qXiVKwTlcfXT9BqArUUHggBf8a7bXNPZ3K/8jYo7nq0
WpxEYCEA7BCzGYCAwHP3ojtPW0O+9umuepSo8wYRfnfjUb5BvNb2tDOvXU81N/hA
R8BwT8laDDeccL1Wv5QuYTxkvj4cDWNOan79cG7GAUjg6ugfnNejYwckUVLPDa0S
+iNFPfiSVPF6m322rSycApT6uK9r6INriu1mYj8d767QM9hbRmB/NsqOvLwkyljO
3DaKy3/axpuXaZAOnbVTJZOPBD+pKEUt08LGqHnPlcyf/2idNBAwS2eKl1fesIaF
JXhmAizXm9W/ZWo2UsnIYyCFq5Yh27jqKMbp6zGWhPbLYBoll01okSyzY2P05cJk
c64x/QzMXPbKM7xpz7ZFy8VnDetf5kFIQaL7Fgbl79A8QZAA9EcAxPSuSvjITm8A
7GgGjj8+85etgpZflw8ZLFqwAfNv97Ajoy1EX8HFOrT5BOX9IWQqMgt+TAsCYw1w
NR+TjyFn5HTWKj3Td02VcJZr4YminBXdnJX9amcAmlu+VQitf5tJ6SvNSCkQKl/x
c8lcVMJZ1ssb4JrqdiCzxan/28LmjWOxKcYEC6t1svP+HHsleZhyK4O6/ch7PPbS
HZRbpmbtDmy01oIWp44c+92QOJIf0nzsnk0v6J5LYzQeEw+fuob/xODRbMFviX/l
djM7W8Iz06h3g6/8Z4/aw6ShGp5lrGJhsRNr45y8SUFqSybnAAQ5XgfC8DDmQyzA
THEv6ubo54YOQ/0ol8G8SbC6fLmIuT6kJ7MXHPV4jLwX8ECkNLkFTfcqJYrE8z78
NCmuvJG3awcmzCpgmwjpc7LBS+KvC315L1SI6NEsZR0Wwa8D0lf05cDOKhQxnzLY
dHCUQbltnBbhx8ikUL/+QJlGI6JvdTeUObpg+mRWOmUW3XBTcWbJVgPNz3D7qORD
7likemLyHHTw/WaFFRZJ8MxYdq6EfrJFkdUSRMqhs8QWG9/eLWNZNFA4EBIOwOqO
pkXucsV5VvnIk9V9bNX0J2J2GTOxj36JiQVI4MxwVRmM2YDFuAdx8NnT5ZO1YDjo
d5WzwbhJbidsldX7OJzzY4rO5aIS486JcT0CARXM3uC65TdCTBhyyUrXoNg7l8Kl
tpFMP/3bmv3UkKcdrWaetJfbtR3Sd09RMbr6em/G3FdoHbzVUZEv2f5NgYIYqQAn
QADfDzfqnpAIVb2Z7cCe3gkh/cYP8VHJTugs5NrQSokJJAebJvvFKqh080wha+BE
7vzSY1+HMqfy9SIQrb+XZ2cmIo8c6Q4ivR7Valg1Pr+Vd91hPeD3fP18wnIA9Dc1
lhaAzraTm9Irim66TC+ofs/WoJoctZgUveqteliDrlGbOChUvgIk56qFxK/c7cod
UibexHVSqzbIlJNwHnYGNcJUjjdyM3+9PALKH4D10EzcCYQKTPdYMCEJfygNZiMu
IfqJgdhNmz44cYdznN1G9tHfYMih+gX5KhbdBYYfp0y43hL4GSWWnBSoYdqLoizM
eWneTIX1VWcMMdLzCDDtaQF9daSzPj/OmggN0vKUGPWxv+nrVBWm4RpVeXwRbyVF
+qJAxLgSY2zsImLa+QZSYdyKmCe8K6xVnMVZwkcItL4gdv2ghhyPfr1+pla+wwlW
VHQTaTzbiOCohNafVj3IqbJ24u6g8iswSDRNV7dv72dle/Kg0DAfAOW2ZsCY3eK5
c8JRwgMSMsWMNbyTDGpiRshfS+/2B5tzhP9OWpf1tTnXoTz8dGye2kiaV9If763A
aChJxcngcaE/zb/nk0C21VyzZCzzs6g0wUiOHF8pjwAWiQW8qeMGSkdiv/9ljV5j
i2NwIkNBz+QTyOkO9CBURiOfdcFsflT9sbyAcggXUEFzte0cszazC2lrEP3eixks
qM9JKM2Zi1WTtxQl6ZKWQzmMonRl8HjbYRbWl8wMNSTkNIwSdUezDiPVR1si/Ctq
uTSRP7GxRBWTqwfGIiieJuzG95Jq6kjyQ3sRO9eIUmZxbgWuRVcikZjC/sEoAieD
U4MawjAWObMLVMaIgsqnU1cHXdc+16RKPcz4+HE0Kdk4NrigW65rVsHPQM0l1vTf
4iZylVGtI+8NB98+U1JMVQ2HdGTEIk4kRuNdtnYWLq83buEjo5HLqvF472A720Zi
8wZlC5Egwuzj9JeZZegzH1Z2Gz7xsmhDIpnEUH6S1dPQdld1lwyyIc6r7lI5mrl+
jl2LTpWsLwLze4KHT2c0ArklHFoxqJ7M+jX3ogYYcPMK7TmbjfV0Pizs/0JE5rCQ
CPilfD3JUo8csFmmN3IJ83C0agxwf9IYwgJXa0JFtdq+EUJEXVwn6xxAeu0zTT7g
S39gaTprIxRWXyeUAVKlJz+NYbIYc2i2kpm8x4QDNda372kBoZvNdq0G7F1ylJY4
EAFedelcbiWtHcwR7aDlEPoUW8kZGiwSUKin4K286ArGBVJNa33VDIgZQJyLIXru
xO79OGcVC4R8dpemn6O0QgMMLD4vyV3LM/R5q75ugw9G2vOXcd8pWCuJp0ctjwu7
hDx3l4Lh6PUWszSnIP3rTZhlNekIYI+rjHlE1ONJKYAeLUI2ZmjrstbvCdprTi5e
K+5jRAEjPtbi1ND7LENMeuq0+m2mxedhWZg7US9qlxrROEVcPsnF4R+Xfj72xr0P
J/CODesZ2tivGDruFXz7x/h2LDrPfj9owwxfmf0VyOorwvoE3v0gT72aFcIQ3Y1D
tRLL/Ejbwhu4dz6ks31G/H10t6oT/M/nO/3aWdqbOLRkWN+G0ZC86B+UIeNLkuYj
5NOvOK6mw2YDAW9JKF3DA42j76kmAnPvy38t4xLfIqiXSVaEJgWJ2vYc2L1UoT9Z
yHaVNq/ihQmQjKYkUII9EFN9WymOPV3gv0lSU43wt7AXbKf56naREuZumtW3kPpz
BjXxWCWEr3ZzpCxE+IIPUz4zhnA0QmjDjpm2/SJ31DnWKXohyzEN3vvh3jXFNQcT
wCS1Ok+rf2MJrz99tbvsCjNs0OJiiBnS/mRxMFU9NgrWXwHfMfbVlSgHmeOCCNfr
9lZhO+cZwVHH82aqxYqJ6kq+55fJLKgik3vI6SgfPSgP64UlnSy+V47bIhsC9FUs
zhOs03f2qvTQThtRFizWmNP/rn3C8rKcAwMYg+hhJK4K8kio+hN3cYgXXbSC5JLW
DfOZ7nY8jRX6esMl8XzZ+KN5/ybfuxyzojIYhzKBt6V0e1WqvOFPYNubuoptSlm7
SJrpQe+GCdA15sP9iWD6wF5oohL9hFjP0i/+yQ50Kq1kjLry86dvW/dj6c54N4Y1
zTvDldEyMAyNavE/ihokz9r4lnMMwC6BNWFADwOfMDnzFH6wSP0qIdQvqjKF1D0p
qYw8nzbm3qpsCs4sryJhxmN0y0s454Qe2KCWRf7puMBCZzvsMfoPUw+01dl8b5+d
J1jyeDrzCoIiSU8VeVmM/KmRzJmCYjmUd8R0Ww0MjAQshn4fQCHoH6/kkLAyrxIR
MVqCZ9URePJOr9Yr9l9bTwiLm8cphRkCr7kt3KBBYaMqR9OjrwbsUdMzt+PqA1zC
omfpeuC7DeTRUX57r7oYP0FcE6rRLfkHuRTZ9/4B8SJNpZT1Uh6/lLACs5YqHzEw
uKt4s0HHFchEEFd1O91aq1aIMeP7PkfkLmAGiPh1MZ2g13qn0xTgmA8N/lLt3Fem
89XUU8KoFZjboxKvorhFpae2MFdhWNBikdKSZhu+MmxlwxWmmdn7BZTFRLUMkzLC
CLJCkLdXisCRzg+0ziAEsjXQ0Nn62orko0YwlwSaxU7TpDt3APLNAtPdALM1KAh/
8WYtf+tdIwgGq0rs1AG4pv4IH7DHySIywPYW1OK0VQCC7gV0XjC6+MP6Zp2yP259
s0XQJlilLAIsn9oza3krykHwptWLCO7AzkWIek+JetswGDou8dF2PBTCKew0rTjd
Xcrsd/ZEng3kllyekwLSDRm7yGB3io5qJ3Phrf9YQA/WxV4WPhRFdlc1RFwV3p0x
66t8lF+SL+KqAVoiJm0rBcyf6/F0UGa67kcTucKEn0DGsZTBICsGyrDRrZHuGuHW
N/QqpV7o6zBxwdP1hEmYaSwGooNqSgdSzhqFT4gipCxtQxTy9Hv2c7oiLTQD/boY
2U6EteyL2XotF/g7wQB/rIFgLkvS0QVSJ5N2runa/DtlykrbxrUjgelGwMg4vf+Z
FCYV1VEdzwePxnWZZTWtNIR4VTleKCHozSy++kjF1sXMFLc2ey0pq89J0Q0ngVt8
ldM0gXKJdHeQFj1OqixoDURv457L2pMfd3QpkCsFH7X7GJOJUMGVGR9YENJAZcEb
/gh5GXSl9FVn4kHj1JXLQQlcNDVh81urL1h65sGTCnmm87wFrzPtiSmfwKghdnxy
67lUBsIHJcZs+9X/2ClltZOqwJei+0/+AqA2Lv6iktT47hQnpRmVsznkMHjarGVD
zrzICU6jGNbho4jPblWDbOy8dwNahJ8VhLJPoLyU8bVdszFd7vhlUM80YVg2SBNp
uai6uwGzcHUxBgXVebMRrEUEUxpKs1f8guZSrEw/+645uaDtAQ6gvSeDgy5AjJzh
RHpuz0XYzHLyZCmlCnsEcs/zcnVFYEl4XR8OVAafcI/P7kRQ7Z8yVrgcaPZUyMAm
vujW0bhZXh5T4aF+Y5JI0B8X+rFbXSly+DJJbmgHx1S7BY93K9vB99TMdQ5moCQV
hNmOkFu6wz7wXwYrzyqvfu/Knkt0b85Y92rRupHN6Jgi7qNo2cm7U7putu/xWZTa
JTCILJzewmEpTrIYfkbH4EFJ5UfVP+4M24VpSeACxCgrV7LEREubUrSG9EO87hm4
ueqq1Jy3SOHcyKOdxcqXf5Mj+WE/q+BV1k+Muhw3EogMIYjRuzklU1Jn9dEBpCE9
q/z549/rZ54VrFGSmrptEItnvgTS4yWN71cuAyiNN+wZuvDn0uk7pR8+KglDGzMC
9h+lTqkMSpWW1AFXMNC//R+I1tnLmEifShmJe9+s10vU+ZTE46jlLJm4q9UY6VCq
vrIp6WZZPBZR7wqitXNlGw3W94+5/7qsGR4g2bwjy2CffdlsIE6gDBH6OW/WwCH/
lez8N/tsI+w+fDF+e59yxfdGGqJec+z+I/QCCEG6NajDOPbnhvfswoLA5SN5LebF
2D9ZaJf8Tr6qJ9pSIwcKvPmFPeMb1V/dYku0bXIzWe/YLDZFDMM1/oEFV0ZGXMdS
eBvrr/LXIs8PuCLKEA8f6FHvkGOQCYMjm3DNGpCE0dQGeolM2QMXQQ+5zJuOA88y
/RkG3Yd5gAPgmmpULpJGioT6miZNUhuIGORr/l/NQsEhfYZcDrXKOqLXt9C0OcP+
pGehal7ZwfkrFQUSKMnG7k0xilBFSlvUd6Cj0JZVYEHnTq9k6AHzXAxrb1aIO7Md
kmhxX3K3NDqEmXbv6I2rJuJGKU+lTuvtueiK5cETIJtXB0dXOqbPfJtpDpTOjfZQ
A3zyWD4q04R8xsmMlHAkj1nxvKm+YdPTrvUERibf4ypG+YVM2SS2U2Xy0B3g2bAd
N4jR/9T5aMGUkU9hgbVdAlTuCGZoXa+349ZpaS4K0RlukUbvhmcYTzBeNQo3hEJK
JcD4V14HHaphGwMpFURQS+aB3vwbZm1IOFfd3XXS8iRD8fX7nVTP9osakdid3Y/s
XrNH5aCyRLY968wSvvOM7DUin0f4Wlvn3nBRUiBeNLFN8Rc6lxlXzJaF4zeHd7v9
myPpSnqqV3kb4pbq7aXDiGpUA4dAzsPMrz5iQZpUY5AFLALSQzqdFJL50uK2wzrP
7+yjP2S8t8b1rkAa2i7zGQ1xhzm3Hb9YLs3Nd902VcPQKWjGCpR3EBuwvTKwT8KU
s7YsK8awCcGa2gtLBJMlp3lwg3qMKI/Qsuro9E3MJnvY3YOy6JvozKY3OL6Mjv3x
xrjxsMWjlRKKmXWHBcH99ykuX1qeQPwrzbhVS6DDLXWQX3CJzS0AlVpfkKJOV8k8
tppy+0uYB5TDQaVXgWt3DKQedFEU385qnwDGIXVxDNCaS596VVVVXeSSUbXIZzaN
n4yUys+dzFFlzkQWCFqiJ71t+WRXsGrkqboo9ZCJ7itny0XXSWlrPaI/4JYKd8U2
kmjtDReeyYG0693jd2aQ7n2IPyhsC0AtkdHoabTZL7QwfW0s0E+Py9IbAubqRmvt
sQlw22+8gpyS4uQcVgTAW0sfR5R0Z9wTxFfec8qBsJM1Oyfk3qZptpbkncjorgda
J6p4kEIT1ebi5KOb6wTztpYIjeVRA1BgBauu00wk1IvN2BueHeT2GyjLzUweTd2Q
AOFLz2eizL4AFPZ6e/oD8QyoFse8WHVdlZnO95faCKSHP+5oWL8HkUPyGodtA+Z8
COBqsuN5YcNjFN+gbIv5gxUMG5gnR60gJygUtXigVlaUOqc+f8UmPR6YpbZNhhFv
WoyWRS8/j4XjYnLvi2tjU4OHfxXO6acezoa0vrDDSTEfgZnf59Rc+36tswzjBma3
9d6RdLevHubwIdySmJG3oyHRFlMDXPp9CZdh7G1KowJptnUBrAsMTRIxQGiXiAkl
6lqhPDacyy+SGMOO7CO0D61D3Tzq0oaGkjCq7kLOQ/8IY4AC3EblP7ikf5+8GHYD
yg6vMjzrU/FWH7iWMP4xhr8QlF4g4JzkZIjjRqAFs+WhlHvJsHXTFzi/CoywMyXH
/pYeJ6qhOYicGqCy8y1cdzCOLLlpWJfBuwjYRkNpfYaICHc/5bIaL+5Up1aeV//Z
jLEr40DNFOJDblYtnHdgX+8gS914aWHsFqhp1Qo9UAmebhZgFPdFq6YLpgd9zLpn
cV6l73aSm1nazY3EQIL9r14KdfAett9z8T2cxKSAyEpLuQgjOmS161NWN0xMIgY+
X+jEK78n5DSprcV6RNae9g2DnhibTk4rcCwCZyyv7MKeYYxjBo1R9koyDIljS3WR
bI9/Y3TOgqx/BSmn52ouPFiAmiQg6ANnO3ewBTftXiNrv+tr1fvrE0nzQdjuwvnB
/kU7+FBha0ZQjJlZHkoJKfbuGQNatN2mRAdTgoLYzDPOAuFX5bNI5CtNEqeOC7GF
klC33sP0LeHxqSAMv32fD/H0T2y0f2sDyu6NIcsE+spxpRb82bE/1jQhIOinFOrc
U/Aae6vjwJi4azoN178u1B6bJp/TomUtxRGsh6LwEneWOwyhoaLux4Kw2bbyqeFO
aEEstI3oLMpf5ltwHp2AGCqkqJUT3I5MUMNjW7b5OCE8aP/jP8fzTdKSIPPiMult
Q2HOlxHZmnprGZ0ZATiQ1sh2TxYu5MsfoIoFQLr7T4j9lHk9MS6d4bgCt2Bm6pIt
ZgXOGBOs9/KjIGLZtMcAukbMEGUvkK/7FDu2t9YWEC+26SRTAmzu8aKPB6uHwmHa
jTbzjSRQGihAr2TOWZJ96y9HzIQDVh4adHVkqTuvQEbcinbXBz3meYgMeswB2/yX
mPAVDh2Rtl/T3y8vZvuL2F8T1BgeJVWkg2cel8G7fx7ZLacx2WID29EUs7hsNdjM
dlTDBAakImvhKG0g7lPrjZ2BgJnpBt3jKFZACgum5PxFl1XpVG0A7q9BtnI+Twua
a2EUfzjOCPWtRmCoIrELrhgEKJFicZAWhhjvLIzhgAvI6NoDdOG0lrL+53c9F7i5
glcELJxKfr6qIlHMMQLAfaLLcToVw1BlEKNJM8qlPst81zA+qbCGL7zN8K9XMKrQ
prFPeNeDMa+zHnQkU8gewmbxCPG/Qo6weEcjT+GpKvRIOsLUGO0lEqOCEl9rgBt+
HxaJlHTBsrl2gTJ+v/AU0azMaxv9VyLX53zqScX4TJGSMuHn8wRFYA90iP+J286B
8dOb++lwCbBDnQHU6KX2778vbppU/D8JintyX4fceC5qAGRRgg/3WZaCXUr8JYw3
YhtTtG08MdHB7LZzmt86JS3/i8Uv9u8jv5btGvKV3oFoMdZAZR/I53AQer02XuJM
bWrxYpEUdyy7+nZevx+GRKNbvOrEkvvyV9HxKgINNt8nrBYAX/eeLQLc3yHDM/8J
5Kj5qhLTPr6D1mstJxjFaE0a7zhUF3xpnuTENeNEqArI9TFGq5nUh9I9mL8DiFnc
CUNMU4hfs3OIsAYqifaFBbc4ixRMR8W7yx5niMUPm5SZG61qAGiWtzYriFzOh8Gp
u4hgYXpNOSrqD2CrhhaZXveHm9b5d0cEQ/mCdgnDV6QjiRR7ezQ21q1vI2qbYwwb
wN0AIw91ushBiTeOEudsj6rr2OD/WODnP84vHXdsfmHkXbdi8tDoJiACRTCG/nP9
7HTfgWBbpbMiC1s8KG2gbYC2lqMX0x8YySKaIjs770bGidNn0dMInkcNo+3wSZDG
yIa05x5KK2OeTxBURpyJQ+XH/OQzZi6VJqfzwbRGCyU10GnRvObJletg0iR0UQ8Q
dsSaIDYS//pS7x4+c05YZ3pODeYWKiAzcx09nvjTuUXcsideYgl91QC2KwJrGE8t
8mInf+mKgx5JMV+vIkBPsRwFfkhL5TayzFF6hJzGjVIGMEsrJg8YAzE5XQXozASO
bKxK/GKHyzAeaqmIgx1verCo7FzsHAV5frm9onIxbI4nv/AUPipVLzUgoHhO1/Lr
YQfD0SVGlwOnY6hgLMMe3jM81b2uNRaIDWSmBs4GIDeRFaUa2Iqzv3aXWunrccCG
BvkFs/J91K/gb70BRLmTbbev+ZZjBggTIu6LuQpLkKZxkbJjxCSBVvSQM8cMyXVf
0psqThmxjJdYlfP7FZCcZTrZH7LnhWg9DjWTnEASM6aPpgF76AN4Hro3P00m9Q67
LuLKxrEY71xG8dkiki8VrXn5hT7UnH+bBjDRAExAMyL55jRqhC8VI/v5sjawnaHM
LXP8QviDOiRy+YFQwtlOP3lwEaslIEgHBpyRn/SbN6/FmB0zk2s/8Fk4PkJjIjc8
DU1F0R1Dnop8Sfl5TEfvytNe9QqFTl3LMWHuAYIvlse1WQvA+OyBdLYeYWDDnnkb
XVAs+9EnL+lpvzWqEWMfaq8FGJkesIo9+/24G7Q1I4tIILzwWXjpinFkNUNyKHSK
nzh32iz93Gxji1IIH+M9FRz/93eXvQ+1Vt6aukPUKWSKPHoupB2EVePXEevhAna8
jDs0FU7aAz3FYt7+4JHOVYwnUh4uNi+Qo6f26KW7kE+9l1qV0r87a6f6y1SINu16
p7aJWHtKYCd9TMvl2q8oA3WJTJm40NhVsyPG3EXyzqMuYNgaQGRwmQkOIkyvl34u
kjyrZX3g5xfzPmK6Bc93GHZN9tLNr+QacteNLok09t//enMzIVMgFbmwVMBVLtRG
+yuRpm+r3m1KCphKLDiddPQNP5xRt1KLZS9LdimcxdFDMOiMkIxKbQ7gNYAXPTNh
lOJ6uwZf05RqNC801BjW8tzdcTFVedDD5qRf8u/noZZQqxrnPjBUTdKEE09L8gnT
hl+uHxu0J0bm4P8+vO2MVKTzq9FBmL8l2iJ9TWwhE8zfJI+kOmBygkDqHPiFLs3k
Pk4s+pTbFEdkahLtR4viBmtVlKOAawtX0cumYm9HNe5ghKX+sKa2/WbeCQnt/1Gz
sfHvZ/oqxKnhQAd154WwCwbB4tpvhEaqDVpk4IXx+XjiZTwSRMiZhiB44+mFvAjY
Jp9n0BtL9d5E3+NiFFae3CQfWmP242PYk1BQdY0QLyzsB+1wvKKsK3HdMYcEap0G
LjpgmC0FoDgokMO4/NOBlaOikSEgGtl9H2/w9wMPg2nhhzfZcOj1f4C+Njdam8GA
pIme9ficWUodW7PjV66Xeh5RlAf0JyO02K1b1iD4kJIsq0/c1TgU5BnH+AgqSa3N
6/r7iCOHkKGFCu23/mPmVtPrN6BkVj9pcKy+U4aXavCRzqLrqgKjbIC76Ap856js
NY/9RuYW51tVvJgIR9qf9uh7jJIuARa3aHt4OT1+QGk1MvK7GXORpkMNj2kl07Um
X718vCX4pJyanHVQCIJfg/TwsX8BhB1gvXLkm9Tf4ObSE3Tx1OyrPlBrXIVY4JZr
DZaaaEb9RIDknWc1kzC1QytrpjDGDgJ6miNAg+KVh6CzkJYw99r97eSngIgUfraF
i5Aix+JQz6OyIzB0RNkjcLlE5KGyQ0FrxW9sD7xWaxUGn2XpAOfAkG6g6RrQoBls
tqzXAd/LvHkbyrpmXno6xwDIKQAIBlPLSEwZtLeclrUuKrsCZbxncmwSnnAK0sWJ
1UEpipUlt7OhPhppbcHkF64gdXlsjG3/SCzHbuHbzROUdCkdmmacGVDaFdMixAO2
sMtMB2NE6ALM1V51Czc/ob6jF/fqSuRzcCFCmIkOTvOt7KF/bE5yIRwKDdfKZ++E
H5ev5lfRolW3KO2Nx4Oi47/r8zDfFfg3E1a3BQZ/lsp1C3O0x89DCNn/GfgvdVkf
kB+VlNIIQfvBiCA5zcJ9422Fg694EwCQ9oPNACHZZXTU7LLf3cPqSoQzFXSlTtLV
A6pScoHAlI2jPk+i6Av/w2wBTZhxDLFr1CIaHij6jc9cOu07TDsxby6kUEE8Burd
N9Nfr2kBFmuh+xkLsTLxYXLRG04uQ7QxgGclI+BMQaCWTIxTl5dThi5jJmaUFGc+
lT1RITOAL7/bfJs6scXsYu81iviDJP5YsqDeL7onfGMk2WvdQlbCZXjHmBPpWU83
fj8uO9iyazrgWDmUbvKcd77DhQOfQHN31WHZOfvygf56HlRoIg8S9z89idOJX03i
SCEmu1NBoyP0nFNVbi62a5ufFGx8YzlErXv+rP226XJcIFeCP6foumnA8vLftrBD
IVWBzjXJYTm5GEdrcgwYdCeWngrXrWKQ1sbPZiTuBQCGmNnuVC8XeJcdHFWHAnRQ
dN9EyAp7tp6lbbrVBfN333z+oaDBS04LyR8S1GYts2+P56PVjr386Iutb8RAqanW
HTD9BT+ysOvwVEQwRUhb2v0bdjxD2CBzpIWDiuhmZs5NF17kbuQsIE9e+iW8y9Nb
vyCcut6BwnkEaHXtmpi9qL4+9LBSzkkz9C71GYvqGD+ataCCdxRkFs7Rjf6MWFrh
QAwAsZ4gRr7Z6shDJ0dOrouG/IXU7iU2Hgwq+pH3fctzI4isizU3xfap1cPuYxD8
/bc1caJBbp94Yd2h6JWtMj2IiU18WTTgAfCtyo8Sw8EDQD2iixTH/8mGHyF7VQET
AIs6O3y7yxG8HVNIoFe0bFCr3hwBjuUNurJSIuYj+C5uv9tGszjf3rF7HReaY3O4
UUVOXMMafmTg8z7IkgCBAI9GmVpYTVbYnw34rSlDD9gDOVpFNuNTIk2gYsFQ73g6
118aZiyIqyursAZLiRdbNMjHSwQBJzLkA0Oump6EUYo1yM8XQdQNhwIQnmH6r86W
W+28d0ulTgqexgjLmK3pDwAVLvezTh4tsLoMpiPgvum5wb4KRi+13v3gi7D5vM1C
QyW4CcZm8MaIcAp7AETsiHJorEtjP5y4BlLQOS7uNO1k/gkmxFTiJ47iByNBX+Cr
ZLxOH/KSFzheQsR0Szj1UtQTDRFCvDh/5bDrpADsGcw4OM7o5xE6OQzbWbqXaoPc
NWcHy7fya0H1gX3QuGE+yGfPEweqXtQjB7fL8dTm78ZRq9S7jHCCXsk2++jefDul
sy1y92IlOaebeHpao70kC3BjCleEqt+Aok/MmzYBdN3wu8FrzDc/GqA3YxPKDh9C
S1o/NkY1f0IrYJVXv86g6okvxeTb8Mrgap/uaycpSseIhiXl+4RzyoNFEIT28v2n
sNTBk7QNiJLpV6rYpWfPt408QohJbWKQoAIeulrJdkR5VtY3lXiL3tuYAOItcKCD
FxjeZm3O4gqp9sMLwOWiuk/OHrzxqm7bmM44NPhV205nQTIMSUCQXmX7QTtYMnXd
2t0GfpCSY5sCYgBJ8eyxyUeojloRi8h70rIqT593AfRMQRSIex9ED3QfiJ/gUiKO
XukyeLKsbzgX6sevTA/ufzHhpSeSAAh7IY1rrASFbMdzL6pRXe7TGiOZGd9OZ85o
9dAPkE/i86L7nFxVB55j9ZrrAyZg8BWqxynvQ/rpWtHBVC1ojnVWuwJr/GkemMRH
H3e25MQ4Z8rTcjvaYdbbCCe5G7ObTMCJRCYHbaGgQxv2fTNVkcftC0SVrzN1+wQS
hUZVvmBhsTGbgG9ikagHpS/W9SedTL8iLWCpsEg/smDW0wockm6LjdHeqkgcRPb4
43vlOnRTKNze/HTjtgrXn7kuRPxQTHwYgTLOEEfmuDriSssbu2f8uJWRarn5eJyP
KsTXZY/OE7twMZOs4jDaOcOEEIfiZvLntkiGWcuG/YXjFQDeWdr6+jMNyexwW1Yz
Hsx6U45kiYoajka45bKdbzRE+/JC+YzL7f4nj8oYkzvNfAI0WUzWgLkGx4SUDGIA
9IOE8f9yRIEfD8vg7lwW4f58DWthbM2sgKGeOj4ShrvulcC11ertnPQFeUnGEUV0
uQwMWBy6e0lxDTCZdJDZw/9hpfU2Cz15Z3gP7A4H0hiadbw3tjXLjSPSiouQJESA
gYKBb/KR/Funuvp+4/n8oYCuAX2lLQBvsy6Qvnu/n+KbS/ZUzva0LL0Ss63Xb+Aw
4DJlC1oqu0NnytaOmyukH92qRnJK6v7ligCn24AO10nddw8PGJKv8QKkNbyt/pLI
myb+bTCuulphb/u4nnl3fwvZaH0/7wBTJMWFmQosXy3NZ8hZhikC+TvEmNlZdfxl
ATE8J4LhNDUVdbPHN6HujmIzMkqfCIv/k9Ydc6DuxP32Rd9jxC+NWVrDP7cWjVwL
4oLVamA+UC2InQ79Q6DVE29a5SFnE82Col96R/lt9p468WdVMSW5+2iDnddcMFf3
DoR6HrlJ042VKifOrI16Rv/7eWwsdwjAW8Vkf3l8UuvEyxkA0bmIrxJBoVbLKGsi
7xV906NuXHqbkW7exWE+0C++u49wlybxJJ2uP1zzDoHGIJOZ0CZdXyMJZutPFcnZ
qGcpZSfGw0ogV0sj7WdFEkt8QtLrm5hbc9dmlLOyeqpKx1nX75iyZxlDwDefWp6W
rTdS1dy8hROTAkPW2ivSXVnY5vZJBS3vCnc8J8sRNI64ausP6OFG6JsuaU78ho0m
OMNj4fdZHj11M4agoDxL0LB7rYo+xsxmmcyVxHcGhS5NOjNwJcZlzTqw8QyJnKVU
CnUfzK6XOAwJ8auvKwFDGEGdO22qgDBzvys4dmv6YuaOI53jW+AqTxjAV95UoecX
O88mnqHr/28Jk8Nz4clDLeYxMTjzBEUUB0RI1QwiSbBZiKg+XjIMzvWCfBkYZbI6
GT8W0IbKfQZJVWyTA8Z7h142yMmFDh7F4aEvXEXnYVASgtKhyGuXFZC3W2zm5SZT
EJ+xNTVwYN6B/x/Lmk6DGLTfYzG1axcsz/pN4TU2jYolq38EjJMo+YT4UvW+BNNf
QTmZzjwGV+JWi0QCGn06fZ7HSAYTwgM9BpUdL8st8ntpPsAg9S5OiKWbRBheGdkT
MmKRiqWoQnIDsSlHty2IfbDSYOsoFyU6CwN24qeVzvjxif+IjHsmBkuqmNJUhlBT
oxjq2ugXLRbIFN7G7LyQmzlo6NYJe/dP3nohFvvTGeB6ipSpNlVecmzP3NtMAATR
L8iCN0OLuEbGyYfHwgW5yYa/0QmISCyq2/ntXPQNcwBZkDyNDd7uVdVLyQUPNTVn
fPvqHyIfs0ZAu4gxD8yQIoJ2ERn++kYUWAey26MCAT/ad6adQyBKPUDpiXf20lPM
/boACm/IUMXNxXwMDdFcpaws7gWchzc1qWO05MXLVt+5iggeoYGfDijxGUqqSTfR
yyDhOee6rOKUDFIfvrvQyl7+LvVGwvtLU3qKMc0gEWklaQbVaupZxEqEPl21btEf
tq7DZ/tlTRq+1olU05ov7g62hnAvYVd7g/dA3WVFLUpRP/F/XAvPjoUEgHTCDfdU
FWt1nZ4GcwiR7QGvM4jR/AOpsvfUuFiu6AP8M30Bk952vHZ/ZPcbwyn1SQ5OlB8Q
VwJWqok9iQrxTZk5HUGibFKCKkkiFv5AaMn6JvNY9WJyb0J/PAUx85JPqCcnw3o5
kp/GctDE0Sylx4LHZLCha6d5AzkB5xqku8gGG0ZB9Ufvp74y6k5Nqb8tL/vRF/fS
u3EmWn0kF+jc/5rKyGrMLgqPIOcWnN6bPM4SU/HMI/nNxiEymY3HuYXxb71ddbgo
zX7GVdxixF0/xISMTSMTCmNC5r1RM8gA3gOv8YplA36M+Ujbk648LvjzNy1fSjYp
T1seX8oF1yA+QYs3s6rDeWk4AQMkuixiUUvGupCRNI/YJ5z6vJWzTGvHC057g3uw
nnUUQ60VvMY2VVQ2SqV+o+JPFUTO++3WjOrs3oiCycWVna0iV0QNpsCdrA3ZUVjz
UXVQPDOkGb8PvUF3zlhKshyat4Pqo+axvIezRwU7zM8NwhnwKJEAtnwUByiuklxj
swQ4e7BXSkJUQBmnalrhV8gsBW5b+Mkpr+oS+RReId/LJeMOCKDHEywt9hVK3+Cd
uymz71WJNCs60JbutGKhLTZ0/Z3cG5uu/8M5e2hWFFj1qQCjb6s/gCwSwdyFs3jL
I/udRAo1e6o+K16GSP8DTqJxEjZy3DLAE1721f0DJIZckXnJGKNsGi0WB6gDwKeS
ub02vlplbmzOUC6c74nN/6L0U1KbFifPPxbimn0wpmLvD+mkEorjuOLBJsYZx7tj
5AHF1E/zYv05JTt3EFkN50kZdrX6+ZdBhSLKaiU7qwQiAYKdKaFGAOfFzhENKq/g
KsOJmuYO+Tz2ChpjjecAxngJ/o5Gwwg8Of5FLzV9l+AoSezwkJmefwdroosUvl9p
U53tvoxYKuqr7KCjflbrlQfMxmjWHvWw48Tkpt6KYPZVNnZGM/EMzoj1N8rcIfdu
02nF4gSZwgaNQMXro/VVQ2MxKQ6UFAtXArMCcdcrCuUl1/jATJM624saFfl6Agc8
o35u3KJdLVqhXuma7WMFyR6vOsQC5pwp4J7Ez2hgmxZ4kIWsKz3X5yIienkPjoEl
oQSAdHZp/IZ+q0jPVR5FvOM75+yFbMvTboGjyNJyx7d5VtmV4rHzanqSNh1hsEsP
rWK+qEWewNC7mqVPQ30J2BzaQXm2T9FGWdd33ib2BNhRnZEMhjoXsJpwsx7Bt8zx
1zFxs4tk3KyWq/eC3mSqB/sR8tmsH/9gF0ARB5G49e9+AoHUEBTTyYxyK+n2LGHl
g5I962aUvKbHk8WwEeX1RfztDwArDRzUOm0qPskzXsfLUQqAsu5L0cF2leDwbyk8
Pq1r9fAJRV69bUS6NRefnsGtCIdKDVYybsWiRvwr/0U+0ktxA9/Dc0ygIZjMn8uQ
AxCHeesMstf1xO/xawcLBW8JOlu7nrmZlZXPGs/LYvhsV3FGZ20iEuN76ets/NPy
nHEkamC8iv8MK72MZDFfomGz2fHkqAcPXfjMgAGLnxAPzf3fMIaikO9nFthbAN2o
HzzZAeWdMXkT3uumWnjwUIapNitZJ/WfjxDDcVT4AUL2p8jhu0KFeQfxE0GL9LLK
vyYUgC0faaI5IgR5O7t94Uq12XaCGwft8T9AE/1W/l8+RFc3Np3b9NZ0BstjwQr4
jOn9BCAoYvT9P6Uop1/1xQL6kvM3eduJhClazbx1gr7bKAZ6FeRjinBIRJ55xATs
MUqnB0XQZsdJ8Hk3FFnCjCA5xzU1/elxjAMWq6n26b/VpfV9jV29cwHBcTFIEGM/
dc2HVk8y3kJht8ZBFU0bsZiAblXGxuoOO3RT157Bx86islqBaPSh9fR918nI+moN
5MGAD3idzUiyd5F9eHn1De2ZRS/zihRBZbhrdSPao9h26OJRDgFnX2vxTMz0hV2k
oVIww3behRJF3gHRGHh79lKYIyfrcXwCkgzsf26H8Ili7ODuTZTK41exT4XmjOtT
j/+L/OyTcq1pOGhGUXHciTRF5oP+w73dLV84AO7XwZsAEYiT6MfPZtZIN11OF0GE
t9Sx9AVj18fU7WsBK9Bagn09riOU40Q+Q5xY7HotXlQaYNxl1kI0dcIW+wggUynV
uAQVc4UE1deNFy3L5nYDPFQndrsQXvpaBOr8ZIJCttjQ3U0i3PhtABTlg1U1f8tL
DlTaFwYJVNmWrW1q9cil3RnCTVRaXuaOxJpmMs0jKPILA8+FW1u+eMNbOxxqTAcO
iMXCDxT+DbyVcFjnQSoZluuKm194FWnp7o2d9oSEsI33pR9FIdbErAeIMTbjBqQs
zrhvSuiC4QOA6J0tNzf42rZv3bEcpYfP0wr1zH8gA2TesorGsL27zc1+pFp6odO/
UXo9K5hrknBHKYpmEznkFNoCa7Z8EVyyJz0FbuRGuPjlZvMIe+G0ZH3y2tatmL/F
Xk5lH0spffh481qilLXxG3WndR64hxMg838aUp2VEcr2TOwtVd/F0ttH6o5uVReH
xEnq8sQ29th3wmqiz9aOD1iPt76T43WfgBaMm2wNmX2T3hLoOd86udAnz0JHXU0f
CBWpRBE+x/IQdjibzcLY5oBZ5wfR7zi/5eAIBmufgH95kNToXE9vh/utlUlQKy/K
X28liIfZ8qFVNp0+WG0bq8u+mdtAh52neatogb7AxzpuEO/NZQbFdXa2MiEEBD5D
dOqvEZfqo454bquocTrWihZQwn8HPLaJw4gKG4i8ez9IYnezsQKN8J7QLGF+JI6Y
8YT+z99YMkK7YwYVV0A7Wpaf6/BB7zzYK8LTTCTh/G2Oe9lmYqhDBmHhVuDfxJoU
9ErtX/5wIPSPxP0jD5Rd/hRiTll/YIZU3uLYbt61kZxxsGsuzK35q8mZDRrz2GAl
5FSgcvB/wKY7KUxy5sj5uJMZA5Q4mvxKCau42AgKmeHoT/aDPVlJdzwmJ3BoSttN
kVIw99fbJcQrZTZ28HHNXmhg6G2BvrORWIZLY/xFRPsK/xq8wE2yO1nOtwD2F3ET
fWvAbFkyQfq1ams76onMpaXOZSMVGpyo7eAMMTYOVkDIHZH0ty3Mrqvdm1AYFI5Y
vclrk/TXZUt5bpFBM7RLyGJSr2hrIGg8eO9oGvMq3KaeE4jixXF9Q3eQVMKTstID
jTXkJ+8A+zB1cG17eaHHjkfw/LRkqKaCL8wEBH1HyR3iV3c91lQv5mx03XCYGj1F
8qRG0egBexkP0xBCqA613OD0g15C4Xq+CCFuuZL++zbIZQHKj2zW+E/4A1Nzx9yv
0Lfi+f6y+f93f5zFWjdrozxwTKMEgtFIdAbQPxKZRFHd+beOJz9vvVxvSb6du4SG
ISVTLrO37QktNb+atvSui89HK+OWbIOhkp2v7kDB9fbQTqLe6Vkt45lFTj61hZ5L
XhC1zlTt3pM0l8dB4GpgHxzxiZP09WUhZatcHE6QAbzlfDNiQBykMOJwhLIW8JkU
/9D3ugkpQD6bONRgkmZA65x4VZg2N2DqHH3zh13xgFdSAJ+HbTKivMwL5OHUG0iy
5qSlze+OHPcznhmU1lnEVq4dv77jg5rOG3tvT6s2E+/81TEpDksQBhhEGbEEMXTT
gXASqj3QC9NqfzTbKhZaFvlf4s/WzHKLmhBemDvmLtlijwPVjGI5sPy8lNYU72nB
KEAxXbga9a4hQ6VHrFti63LYjf/sarb27JccmzhkjyaY2RYy+EAZLXurYEVtdVIP
mEo7UBi3hHpIIScaU5UWisfA4dgE0leP0zI7kJiG2UzepM/ZYgINKPQt0EIQR2/t
EaAqTYO2C1swvmHqt2hFlpH5gRXWyy46/Mh9bpRePJRpMYpDuoUHNeRn7Y9cYzGD
CAuM0HbokPT5trYN0+fP/H8ClTWmc77ZjvsReELYTej12OqLeRfXG0NpStj5iqb5
k1x909yjppKN69gyEvGfgezzwSW66Gkn0W2ahw/8ZrCHOZJjbmZmEWxEO54D5/ij
g4+w6dDyyv4pP5PWQQJiTgWL4tfizt2CGDHGrmjo9ffNZGXdtoa45qzOt3Amf1J/
pCnhYM1As0yNlvYw/ppbOppaHcjLagFVyUkAJLpaVq5FYaKbTEX9hduAwHTc8DPH
AZYxvHnYsiIGZkdXu9oqhVmAwCDizWj8+ntkUrQdBPFfj5GaKNW/4D0fv3maVCI/
KMyAwdRLOimJRv7CAvMqFpdax2M+J6P7xSXhWstBFDpKYPWiM4i7TV+Nn9vDKHkQ
sTYyTqM2fGk9qYczyU+cf5cPqEufV9lpP+f+Ssc8KJ6/3ZwIw12SLF7CKm3q3flr
mu34Gv3q0YwovAbJRz324o+V8caUyC16662lijZ5PCiFEXn5S67/G9zklaUR++L5
JGvPOPrzj2DwpP0CsNdokMn79SKEfhIIsK6cc+ZDPQbT13t1L5TkddemsdVef+S+
HorXEK19kvEcmDM8pd6hk402XTV4Go0P0m4aOF+Ye/hdGu97Pr5SqSJDIoWXaw7B
CNOh7kbRbhGvgpUUjrXyxhDf8GbC9kQ0Wh5yr7yYdmU0kbs+BOM7htrOnWQfXekl
cnUzCoUo5WrD/7OPFq3NCj8esfud10fVwcvdrMSLPF47lLrJJmZ+Tj1ftVTmZJuw
QXdiwTeKzVhGCavKjqWO3j45xaWzNA1KNmSZBWOcy4FopblE2blyEAJRhwhVcd0V
RNvqNHiG2+7qURcVegaHnqG8ZFIkCT+6Y+J+XTor/Z1uNLr3e6ddcFSOwY9fB95k
4UXoUjIHGlzyKOPedu44Y1iWRi4hIFaCT8gveF4wuJpydybZ5c9w73tD1UsAUnaH
PAl+D/Qiqw1P3PEf4Xs+gYLIgE0Dgy3mB4lGvYoFVVgK20w8ONCQITlM+4h5gYej
o1kIpLmFCqzPUnYwbHevqmPNUiivGG5w2AhfsgHZvibNQWurlThZKhIcRkr8XAFo
znBOj5F2WvLuoZB1TkD8beyNFLZyJ9NEXbpSY1VqhM1l1CDRqZuhaq2C2ZfEosAK
m/hlo+1Yp2MuV0NFQTo9Ap7569yavIfm93OLXt/MeNy8b1c5w/17qq6jLeAPpDCt
DVaS6KxAJY7bNyr8ECf32GB7tuMd1SEpaU/eiqd93a5iDXoim6/h9RH4vh59gW+u
s//bpwA8wHHxcuRyYbuNtNAQPmiwD7GIwgOqammLfD6sRh4QVIfDYzfZCRJuEIi1
/HApF8/ZBHIfOSaWDvAg4zhGb7HdAjvPTDtw1qt47JVNKwMlj/lDgSL4TeIpzyl2
FepbeZErYMPJUqZOZMD1Iy4EAZG7INPryeM+4tiUZgOlGXQqEMtexEFEldMRVvrA
rzgw/Kqw16uMiTL3Ucq7IQXlGNPr1TOZdP5fFmMh/tUmrrDmv5my/Aai5lPSx9G+
yyO5wW6JQh5XmpBoWV1HDglV4p4lWEmCdrqMUuRI4MfPnifVuKmnhs64y1SbPzv8
3FAVGIiBAIoHLRrvUSYWw1EuP69JeLecgLXBSNWgZt5eIsPw/c6HyVDC2v0+sZfZ
M8zIiSNQH8q0v/Tw+WHrmgBeITmChzAeRLS73iX9e8vFHqF2wANXa0N3JStWw64E
7maqx9vOboORth8co9hdWc2pCZESVqmVFJoyplifHXAcRNB5G6IrOC92Urd4Qz9K
C1OwN8C4L/PbOj+/23mEvEzGGYok5b50UN8XQYBERvyEap25hfAAt2g8A0EzK0p7
XOQ/b79JzfHSXrU5xewB3aU1urL2JJHeROy9SQORD5O7lJ75fXwxUXR6nW6gbx8p
13WCZbor87KdTdvMI3DZ/3cSRqSgnw9nJVRdMVhmJv9Jmv5m8Wq1tyrAEoAnAEWh
PkA9WkY7/HG/QOhyhBaMVc9hxA15HdGBymMfac487d4LGhEuGFDUprKliF6Q/dhd
xIR43zXf5C9mNbwjHaVtCOdijVzYk61F50EZdLm5R/RixiWdrpo1pBIVc3tfuoC2
crohNtKvtw6oMatoGgk77gBCLDjjS+TPfZGvvFxBpxNKOWNKxlHCwEBG+J493Kg+
nZb5FsTSALqIno7Uk9/6WqPP7HiCYczbcj6mWlHG5elp7Oez456rKjBPyAaosJWl
OAdau1ixH9AcB8E7ylSTOfIFAq7cGCbLF4Bu+ksqSH+lcQrHJJh0TwgFWHXPI55K
9Xvp+apBzebUEF0GkQVFEuAdadk5H3qYr2IfJmosrzVJpnUsX728xi/qbuDFsBuk
5bIdW1pGDgmlLBK/icoClS4eQGzolI2GMC+t2eryMXjIl5AWVEpRc+41qvsTBoN2
5Bxosc7ZGS3aFLVtvOaKmNCCj/1DamI+9wF+U4DGsM2V7zMZcgJBCa7mkqqfgVYM
z0Z/4VQuzsbt+/puTsR6TBI+Q3S/go/au6UBNOwObPYe8v5hQBQcVUxruIwBoztI
L5ye66Qy30IzIVE6qPTwp6hWiBag+UgvTrQE5bQW8/oTjmYU/Gwss7Oygb+40T/M
5PPu5k7o8k4jtftVbBQwi2K8MrNK+DAbo4dmkdbfnfqOWV5N1S00D+JzdFtIlHtX
XsvQFLjGBAi2ilWQwP2lFRljBaBriM3x+ZIwauMDPQfx9PMY5zBjz20MZ0/oRDbl
7vl7EVJy8gEFRaInbafEfzLBh1LZTRjQs/dGB3wfJIOy/wFbU4se0/tGyrZ86SxP
Wm3JJrwxOWs46N3mQG8tmw/rYl4cbxYIYY64/Kva2FPYXC75XDWTTo97kCMyZTA6
BLNEGg62PRJu/4UxpjWm6fEhKyr3ygQI4+27+mQz0VBYClCGEKsYCaRkGZcYTf4i
oUA7L9YUoW+WNg3N8pdVnED0DLokH9gRSRLUX9yAWwBc2idmliL02vjLYINISPV8
/CazyfSRmM+bG+zyqubrvMDKKZylkAqFjJhSVws3SqAxpjAu++wF6oKM+UGmOjWq
uCebP8gfTfiKp05V+E2TlFmvcxEi8pgRwlbCu3yh1oB3OKNAIFpalVsvb8n/BLNr
E3fR+337IcVHV533DSQ9J4/T5b6nrRygi62+Sl3AjN67qJFcGjG0/jIABFih0JhV
3iC1Mi2iP6OeF8SlEwRhjcSVT4bF2+eQEq0T1cw2H93v7BzX6NaKrM6IVf+GBiot
31dYZVE0X4hfeUJPBF8fxuKYCLESyNSYh/uOP8VJ+vDfNNfSM6NR5Cbt2ZX/a2cO
LfTVobl5twzqpfA7usJI8u+TFNFekNzkHjjHPHlrOpcUCZPFZSe0OvmTMYBP9oPx
flNKbM1DxrfKWeFAa0MyYz5Eyd1rvjVcGU0TCZc+K0az27UibQDT2MbVveLPFq58
m2mxI8sv85syOToP0mMZwnk2th8fhtva9UTtaI7FmeoRnDUW8rPWLrApwnbi64X9
L39lF1jyiQcrO875IMTt+Wo4zMkvX0J+OKrkOtO53EYsC3p7SqU2PhnZYJOsnLxq
RU0v7KqI4LXOeGjMJlzerfPPWYejk2gXQ3nYTcilb0hMIgp1SY8v9AOvksQ+Bi22
BXAyODjrk+ItK3C9MVk0iP1zlI8ZhBYHA+2bV9cAOPfH+AogXAy+6V+UAmstorIN
hD9NEcuun34JabI11q1KTkmD/Rl6g4r6Mr3UsQH5M4DWtyXBdFlgwqvVw9yA8hGi
iWQiQMK3hW6+YELGPN4R4GhquWAV2NQfAQ2bNoR/zmcpTalELIlBF4r8Axrkxgae
7vrkQGEXAGMvmpHWAyskGVbXzA7GFYOoKRl29sC7JJjNaEhNN8xVO4P7GNDXGO4u
b6BRl01uA6P3JT8OBSl2lA48J1xnjEJhvbaJBkXmkHYEeDbqsMVHjq+VxO3w+qgR
Ocg2X4u51WSzlOyU4HMt6akTc9PgJv5GEAvwTX1PNsTbtdwXBz3XAkC67kQKUqOg
VhU0ROanuUvWzMqw5/2DKOez/sX5lm7Mn1kpkNHnUW4L3ByKeJS4JEgOl3XXJgEM
hndLQU+jYHdNUILIBp+LnCF2oAJBFITorJUi4QzGPRqr1fa3diOHoHNOMEFFzcnX
vkP+HIOW3Viu/2vDyHxDRcs1UZ5OQ5ev8Rzt48VMYhffHaWlCqnFBto6UUjnlp2n
pEShq4+OAWeYNeMP1pwjA62BSqNvAujLEBsQCk9xImG6Jo9FrGM7jjMUoN/9vNwB
KPLLV/R0KI7+2wFn8QIZK73uN8w8nr8a3i7S1n4xt+17bqVBgnf8E+F4iXDPBxEg
GCbJkcF1QlkmkBEjZJwjAr3zbPwfYUdn0SP8lYch/QroJtj3EZSYfOzqTnrZZSRb
mMW69Eq260h/RepYGfchhcci3t/8SVDVt5e8qZF51NQwJGbusVwh/9ZMFUHwSJru
ZBWYJrzs3a6EDNdsdJCk8jgdcGDnZil+MLGFGSVp8wSO9qHcj+coSqWtRM93r7/T
hCLRo/DXL3/AQaeomOrxGRYp3KFSH6JkmlytjgyNhpFKD978CqgPlxnI3ZSyavA7
TEq8kEsZoCPq/3y9/QOcrBEsmzovkmKGCHJNIn3+V0bZ8AvM+aHOG7XS4LB7W6Cy
gZxicbDAREjrCD798688IapPIKugfufWdlmXqrICvem/L8t3SmqGqBKYXNyt6FNh
w7JRdjhn6IlEQSMiDnHRQ54NxP+J0KZP3D98caTKZSTPdykLJ/oJHcAx3U8j+ayX
8+iBxs5alYXpVxI3Mv/sy7vuGpqhaiqDSj9IWSlSAkYkK+PmsiMU9qA7jYUPzwXh
h4PL0euxOIDnQfbYcceC/5txYrz/Lfi1ELVdQ4cIjiUgYPJ89pYGqFvTJpWrqP+L
kIw6n1dceUMsz7Xgobe4EfhhYl7PAoRSzyOvhRMUomEF2AzJF3U2/JuID7N86zVP
LqXgdSaVZgUWjZECbHjXX4UDeUOOnGDwemf5gYQow8OmUWVDCg6Oht7QD6t+/77X
m/TypmY8kBJ4fZn4DOPB6QLi1DmtOQ2CSePxzr1eNI6RXJo6HSOovI4MOMT9gIhU
+eGUWHmV7iIxstNS5Czry98mw2M1GDl/3Loqoa2zwYCNsCSbplqpkQPpcK66Iw4C
pbzhSQ/VQ0EY9dWNb1Myam+zyqgHK7Y/B/j+lpixdihtDc0iNnBJg5y06xRIwd1P
bP9C4Uo6NYXpFeaoadfwpnVILf7d8zfZnrv54SqMXeMmzGvnTpZZgPvku1naraVw
G5F9coEMty8eEtrW5vJ2gxfrfjimQrhvmotsAG13gEFRjC66kIwalgn/0BoxJ3H+
NcdtslIJdaIrUkeqB4AO7eQhx2gp29kXQbIbgKnioyDcMsERw/+szNHygKEnssUw
XAV4W0VHDWtiDVjlUVk5zYv+54sdGi7tj/VqVkK7K2s3ueBZrlw+A3RT44idAQA5
5mEImUR2Wq+Xu0NnrK9cZDu43OLlHYwPrdgMgDRFGzssT29SysVGXNjYILVtbxbf
fClPM5H6pe/bYlCyiPQw2jaRs0etV//uZOCTcBli9USdqt1SX7xo+Q5jEihFQYTh
9ysRq6Q3rFfKqgOlFC+AnhtduVgcSsrjtrKcjLqgJgFZIKdXMzPG1iBcEZVTSyqt
6fnUx2R1RdGsV2v1UcXJeWbfkLmpQ/cYVQVT3K9PZO9G/PyQhVQEQjDhN0HgXqb8
R4ekgmizd6MnmAY9vjgf7glPmc8aZ40VtxtGm2BBZqn0z/VNcFxCGBz4qyjjXlfZ
prcgNxzlL+2B4Esrsu+z5SR6hO+qigE/+UZ85EvL6De5VyD2fFPCiSGwSUnLyJeV
0QAaphmXWBYuyDNnkUeIkTdcEt0k3s5nVEWFz5WkCRgwIh0L6XGgm3v8PGYUYUMe
LmhG+0uCtvgp/S9b9n/xK+PxkjSyLg+hIY8owEgbI/HrhnFT37G3XPbbHMd1k8AM
SbsaCt95TQOebMC6PjUCJmMXLZ38GudLRUm6jffAYLdrrEaHAFYwZbGN0eXDBM9q
LqSPOKLKMrAkaBvSpg2+SGYlQmq7aplYS7pfadNzpX0U3u89NsZULVmYQ1PpQRg7
E1CIJqSPHvZI8PHyXbGXf6PVxNhWCPb+9zpllgqGLbSYWdUdz6XUXmh8Etu6nZYx
xrYzmCu0GcnwECrBhkxD1GBrZSpbC8uCesc2Yl6Mi1vbMouFZmd1BW9SJWvsTPlG
7+EdYVM2wySLw3qQ/YM+9owfUTP+J4ZWU3+Bz/vxoCkX6xBuXAiDVEJKyPOoH7qz
SbgCkRodbfQAIP4Pk0dqDuYfRLejxo+OhjpDTP3C3zgE/a6FXbyGWYhXj49GYCYI
lzPCW1oEZSt8QC9cKAAPj44mzD8Pox3gjXCnXKOP5i5+o+KY3fMCDl8DqeyGG5p+
IvQNhqjodF3ehKRmt5334FdQtJNIPl63d4iJa+1Gdm5+m+XasHazutKFGaR9DXpR
tVCy4rjPXJHm5fAk7S1z209zjNSULkhSbix7QdZ563aMKd3obXGSrO86NVXbacDN
IxpJOAcQB+2PrpFwcJgY8yfEnlfO2kXzpKIlNjWLXbw/Rmja6YYQkCJHuXpINAvJ
Heqn9WLNX7F0LhcUsu4xX1kWyWDe7GbRdcjg477OeGrG9Ou9EKbublbCgto3z1XU
fx/si5p+EUPKUlRcA8W2oh/oHA5VYq2LZahA7QvDeiRsy1Qx8TDTKPlwBioVYmsN
DByqJTObHNEp7L9QlR2oA7J5xWxfrLGwytWRsS+KErlZsbSX2ENT97YxgfreZk2N
jKLobIDenPQ6u5CU+3a37a6ORTmgBO13AAugOGMtiaOIHwsOhJOed+y8fQxCs30P
TUU0Y1BuUTHuhAqOX9t7UvJ8mvni4FOBil76xDUyquJPEOpka1tU22Nc84OOfSJ9
mL7mUDcCcWyebYkZtBUwXjDOspaVMYBKUDCuaItDTo/7QonL1AZzHULhIif7i4ym
48Uy44GlksMldHPZ9I4FOT81psHcR/drOK9gNxHnAI9nJzhom9ivni/gdqTt+Vbd
7hU+uVWqlZoanjyt2MuRBPZzSKPGqfKXsEZX+ztHzqcFo+scbM9vWdj0Jy7xbO/X
dCe0emC9i66dNThNPGLTFdbezQjTnOWNdwRkopbVCreFe+of70ihjJBAgiZLJjPp
5ccjGsPu6OyCdemIFpmK7DgXqpvPXG909jB3MUPIQk2f68XiWzkPPFRms71niAY0
5GdwcxW52bX3X134mpi/V4RL+kjQbXCHroEi5dDBfP/hAAivZlBjCLeWh4lUBZd2
7VVEBpUSc22YF7fyWdYdpREf+djb6R35a1PrrhMnJ5bGIMgaG+YdlusJFcXpx2D/
pNuHst4avurlhwccUPqNM9RkAxIHyrIMhLR2cYcg+ESqRIgKe27087BTWaupmFmm
hKmiXYUD4GPHCHde5PHFuJ8DDqH4hTyhUum2R79agr46dPeWVnJWYRnbZPvX8Ekc
GgbAeRHIDHecA1qUGEbSQ90IU89BOyYl8UXneXzf+whV2TvxzwOuCPZ+GrQflYzj
JwknXIRIAtz4JuYHiGQ5Lz3PhnIYkEMfWBOLPZQpktvTR4gYX5ogT0k3cR+3Wqt+
73My2mYiFwl/CsTfYS29u5FUH8FLdOyO+QHJQiRh6zIv6Yjalt887yJ7c+2S9Mvh
1em8CCDfqQG/Eh37uGWlHQ0wLXERBc74kYuXcBeilxBkEK4eWy7CtpdSQUF4lyPh
0x1QZ8+qdUNoUMsQyd8dRxo3p+i6obVUh9CYuwmC1uNt33LR2iU39335cVDB1Fj5
LvTMS43+Em/sO5fQD2dArFg8iPDW0gpmT6nxsStw0dXZLFXJrszJWe6YZAXu3XhB
E47gyGfsPH0EaDVBBVElryBFaCYQd3kuOvPVo+PtAQJL0g7xETsQiQL8M+woICxy
LgqYwaOdUSx1QAVA20g5P1R+TVCdssya9+MgU7iu/Q5Yy49X90JwzyRIru2elBcj
8aczTvXv8koxABtpWs6N/cGnEAShIBt3qbWhvi3NFP0GB4DuIK2uEfaC3ZxWkbF9
t48USxHbwL+LQUbv/Dg7mFVikSxqhTPnFAjCWYIgdwwMExGF66eMs/RmSlLENPv/
AbhNGzaoEopVS0CXbjw+0WD9HlnmiYZR1xK5Avq8tn7yoBioewhLvDl6DbeEMudE
dF9lKEyOGUawKcXCL35ZMKOjF90EzwB/Fv5IqfpCPhS4d/D8qKSicKx/oF/SucEL
YzJBCPIo6WeQc4ljs8X3oyRvpiOM9iH0envmTmfy3JoC88TII+61k9vqzhurhvbC
yEiusuXqJyUexzESlpzVyYooBY6tP4LGUAZ34G+8CHvAvyMkWbql1WpeEOYSeZow
vrCV2uTqCbj/gFP6Ga/VV6Qz9wKnUbD5gqc0mv5VRFjtQvPBBqkF9FLxtcK3+KNt
Ipmq7TLqHnfbJNrRlqDDplaw0byMb5CR9ywpprR2WkvzXHqhkV+7uPKrzqRln3ru
hXq4qKPMgAzROOGlo+vETKICVhB2h2t25ib13Z8kV6Pdcp8Hs0wRtRf4K55UipLr
k3lFdeSc7WBE66ZzGepO3X1UbSETWWZN739wXupDgsw6t0IAPFuNxvFo5yT8nOtC
1Naf07AJo7hkUBmCfPdXeR2QOTjqjuRfGgCM/zOYB/ETx8kizCLh6S8tfZJHFaOm
aGYQ/ejwKUUqF2yXODHwz5nHbSjloL83iOBsnttoDSkopWx8cygAk7QCMkats51i
OkmBevvmjqpSY0Mu0XHa13sA380ZHJdw21dqpGolrS4baQYHelb4Eq1oZ8X0yrzt
QmyqaBo138ZYnzg84uC1DFt7cb+LA2V01HdSQaMFmwrqNxcAApK21L1it6MbOuz+
F+iGz9EC/oX+TcvqH3OAH2B6vbX1JhTgkidOFBD+Luq32p46oavG9bKgk5CV1vLH
BZAARNOppzNutdVAozsbyFTOAL0ZYWxiyqg68wobAuX0WG2M0v6R4Punj3Uz6ayq
YtYIAHpTf4WViO1zGHAOj70gjF+HCASApu5g4cRcR1UabKCmbR5ipQE43SJUzMYq
06awmsBd1DpNYGjVO+ntoIF8WVn6sruJ24687lvzFLWsRiOmX+F4NNy+85fNjT4u
pXp8jufU274ljCEcBErI8xYt9/ebDpmrB13spjeZUVYPNCHyNhuocv3Jy0LNdIVp
9EjUcJjXb9CxpKorpTCaNNyYSh8BaQXGPWdvoTw9cy/OLfkoKD3TVrSZuQm4dF5k
8QVDyGAtD+tR8AX/fuL+V1ZLe6om83ydjKjYTivv1VdQU5KkcPwbmJG4mdtEPUcR
gXBR6jaF9QsdCyc0MIys6fovbVgc2w8GD46eP6dXRw9sLqhpKqgXPi3SPuZ4Jmq4
39QzwoDj1Q2YeH0CaBW+6emawzi51CoaJSknoHDm8+svxgCmWn1BTgh3eZHTHTfv
X8ECFvax/y/Bot47ibpjfNSdLSO6IyqtbkT0YIaqEoFvFNR3MXBwqSJZC0oIGI94
plRWhUXU5Hf8rvv1olabBRnrFKl2UBivX5JgXCtCwDFMedxEV1ECnpdBNN8kghUp
4nik5u8WOpDXifXrJUI2J92QvrPa2FXZxDBhh0jrzne+U0Vj7xEVosKdNEjc1eT0
QOwmGtIJ63ai/LSYNYairr2CQlOVO8CWdDzCNXxtqet+SJHTYt7PAxRYwIiVhXsP
9a1SfO+mLnnIq3O1n8C45yxCYv8eNWL9akleHi5MT7WW+EUFYgBSlRj2LxC+liPW
4XDGhTZ5EcP87aeW9FPOMbifjhYiACY4Nba0KerohBycaOjAN7D4MHlvccW0xwQV
Rqwvu2XIBPVVQKt/WCgSLMtlA3xvtBeuOH1XWKF54FxZYfKqYXwOiVAG1eukES2H
grNFu3K4G3CFRMNkLpKuk6lX3jsdPyAzjc2sLSbdnwFAmlJm2aRiJb9IfNY0glfO
SJ790JNMhSrJBzfqgc2+76braYed0Awu+HJ3XfgmN5dq4N3nvEgNeVEqtyFwdlUD
pr5pPp8KCs6d+i4hmj0w/vpjlHTyxIz8p6WdGDQ02JBduc9KxvTkDTRJo4afuLX9
okdLoISounNLKexO5K7ou6YqmgxZCXeXB1vS4wxo3/4xYJuDG7JaY+YlwQPH3Lr5
VmLwwdeY16wLOwfWUGg6qT1K007wj5FEHIhovLd7lsZPqDXpEI2gc/z1gXe5s/i8
Ja0M90FdZQDoimtUttNWoequVymTanoy+hYAMrzjm2HeqZOT6eXsk5dK4EtM3Ajg
VlUt8UfPWWRubDJEpJ9LaM26KSZ+DV9trwyw70duv+aB6gQtZFNey+u054qhrKvQ
anbD7u0A7HG9JnwecTLIxYQFkNQ1upXBl4dWlOI0/KwVztLOFgiOJ6w+ahK+lkwc
Z1a4AKgb8yGV85eX0STpSLQ/hF30jzOsjC3KoD/emrZXTJMZj5t7HJ5opm76G5RU
vTcaoOqiSgj/gjRuzV2B7DoRfkWfj4HXEKHtQOCBfY8V0/OE5f4bSZwuurhLygCz
DXFIzgbzn7P0mckeiNfO3f47TUpaDEL9hTl/2fCIVkOkNdT4MfwE49XnQHwym0E8
YPdLt5qws6hyJ2yTNyrefRfAEzAV2aNtR0AKO/D6Sf8I0tv72dMDpJuUbvJST4Bt
MZaim0Ufwuf+roIXiFDnhGAkucXHyUiOH7BQggFf5yLpMWeafKwRIwQh83eMfQUC
9uOKvdlg5MiezX2AF2pQH8qaA8nzMUY0V6SWLXq3z7QZhNNA2fafJ8DlDuZ/N5N2
S9jM0w1PXz5PmzAJovUoztzdzdk2ZmSpoYap8blrPw04rAUOnhqNJPzciVDUe5DW
cQ80rYtiqugRNatQLC3yhkkDbSHdmxaFJ2h281Hum04qRwtrTbBDwYFZgzzQ29bR
8xc0Mv53q4U27AxYqMGE0oOMI+0gtNLbHefNoH6xVfOJM4AVbQRIrTujamH9VB9m
Fg/9iXcEWYNFlc3Ogo3qHvA50GuF01CmHFmLWd1MWwTGBkGPjlYsTm+Vly4NfFiD
8jeYHM+yIArufUl60eYDCFi9dHXZ6zSjvVMCyntfTAMDfn/KZFI/sPFa7KGPdAxh
IOcII2MPPryOIw5wDjartbZC743pRX7NSXz6Lp0b4wL7SvUKc1s+yv7EGrQFJzAI
/BKNS24sHzG0b6k5O9mSun1GGeLewZRSqKD3DJZc8SH2PQ5/c5COzqtlNuckGace
i65EnKnq2pFnh1n7Qnxsp1zlBklnpajoovLm0+v5LGkNzIyMvpe5XRsS4T5MDIJL
+2Ib1Hz4JlduAxLIEY9CtZfb/57lRi7KXcwajPpG9J3MjtsftOTwUg7YkLYbi6BT
S2WL0/uDSj+8xKGsr2PJMX1ASLB4g0TMfUBYx6YfL1grSAkTxN5vq2rs6e3ZaUoo
uK216dhsBwe3uYKp/6J4keETIyWYPZ6I7Ci06XpK7N+7K56tw5lGoglrjRXR9wTu
q2WDviNVp2OQWuU9+A99BzzQOu951HFB/iTZw91zvUZefBdHaKBFUOPE/+o12key
ms+msrwyl2cs7UJ0Oi0wdK/MiK//sHPUwjOrF9n/UXaj9eEkbFKekDJG3w4YPxNv
Bkj8inMvnafiqIaucYT7fB/s7ff0B6WggCriCB+5N4fLn/kUWbfd5KwzAQFl0bbv
wuHmaLfoUhnKWgq5KGttsVmrG7C2JgpKlohm/gkzS7u70N+Pl78mwfG9RXh/Zz4T
g3lG+5prpvzKqJ6sn1+HEZ06yKULh7QlLJ9y/WoaYq/ZPE3J4hOpafoiV/E0KsUu
hgWyjjDqGFssSxwD+HtPlHYIsCot2ShFrjFGT+eqZG66SGfLH30WlgiEPW212iN8
8SxsLosqfwQ+EIuM/SQwH1/UT7k1LeQ7sLP8SFFz7BrUZ+zZ86Mz+DQ9r8dfyApU
uNhOlx9aJVhMfhRnvn9/MpYMO3bGhVS1g7rp5IxRFa3YCN9fKlGkSHn87oV6ktS4
G6JTRyNUMmiqrHfq6InWbXoz3OQVu6knDkPfydz4VUtkGWyn7pTka/VXMekf+jQj
4rp9b4x7tro+7idb2H1EvnP2ZuyVkdYDS4luBgwPAZf2+7C8tshJQ1ApQBt/a0jI
2vUclI6pu7NhWWU1/vKKISr7GM8KQBGNbFQyA88Hn4ikUcUpkgFgTJbaiLZ6wvYb
RgrWRM9sKRuVGkaoIOQZWQPjpcAaUtXAucA31De6O2Cv2FxnWQZHiZFoHgHL5m8L
4nJIMY9P93tVTpd9mozBz3aup4KrmWRNHkT+YiyMiiZaufR5UW66sVfs5gFRCfz5
zTM5JlLmWZU0ycTlmWX+3IbNmdVPNAMXbEpoOQzoMK1qYTtj2C5TXY3lHjYgfwm7
MMHgjGPpLy5dxAEkI1DosfG4k6fgh8SoqOReUYly6TK0aQ9kZd4yto16sXmx405R
n38efQGHGllJnxYl6SXygfZtBdFLlJm/zNYNPNbyCCpzVy5XCBK/7Sd68hlIqTs+
D58jN/gkyP8bhLq0MgJW4qSJiq//csRUhTiywdSsuSkgxv51eywi6cQjnnSdYyxZ
vyyLFqGCz6Rq8TeJCoTf9xL7UhFJVyT48jckTpiVon4P+iMijCwL1MAjiMEg+hhR
mrbcRFM8yedPBkjYxqtjrSEWZ/OPmIMathNQCwIn54Uz87IGh/+5YwhcW3dTDVpg
ZHygxqi/LLlXjJzEyAB6Hwres4hAbC/Kr0WYuGPvg2WAx05iJcL2LHO1cYrdswXk
VnQ+7lgwLQNDphgCsXKZUcjXCijxWrW9MKUx1wIO4DFD4mTkZODDnpC4tLiCR64c
ORPt4vbyQcGK98/eqIkaHDCxYf/1AvWwaC7a4lBEYTjRprx3HXsTRWHAtDdDU6dF
wYUkzWZMfttqQLUNLmdFTWIpYGkF080qZGhkt88d4pK02NOQwAbMIEh9TJwgBG5G
e1ZT4Z132pldVO2pIselk3nvnBUJZjZViFl97He61ZQoNfhQ++x/yEWaG6lLY8m2
zFj7D9bD26Yq+uwTtbnbxI4JPR8N5Hj9SW52l73lH3buTrI4tsQouyuB1sBALukv
VjqVQvpq5r6fIOJ7ouBUBXnmAb8R7fgY/5dSKuLP933yn8sPiA7AmmKXhg+1gC5R
DGxBmwenvdOTNjVU+TeeMSo7okIb9wOeTJPZx3r0lRC97baJD1teUAZ11PZ9YXL2
HpI+x0mP154A33pgFYDZKBtuGrmOlDjK78svNfOnUcgdTTjYzDWLRkI08XZgIqsd
5NuYuiFFWebM/LUCTCyhnPnKqCVlD0kfo0NL8YSP+6nlGZfok9+S2GTmzJLOZ22W
GjKRaAvh7K2gORnNVdVQGCEcSroPr6LRGuoMifJ51EtYG/3Lga85XlYKVwF55nja
ndjYhyT713ic4jUp59kdSAZMTHCnNlI9FJ4gPjWrU5pQZCf0stYh3aFVJ+8eNngx
hZueYP4vfEs58YVW7VedOOPk2NafOUgoP0aX0NtyAGDBF2xpnfGxhQtUGGH9g0XL
DBcUzRWewQjtAB7LjNjW+8gFCuBtt9f2V4fEOCLi3eDdLLeuWoaD/6Z0xpYC0nmu
/yYxxLw+ms8FVkKP5ipxijHs9nOhWsnXESJ+PBBJ+8FiMRCepIQXr8chGhDip0if
gSA/UFSztcC+nQ0Y75tF1LBvH2G+TtHZMYqrU7wtaT97Xib2U3pY4cswsj/SGnyP
EtTgo97WtgUWYJkLILr8qR6QwZhPxcSPOxEd+Cqo7E+HJaYO9ndae3PiB0KmHLuO
jDIXSMBlmbwGjXIbNDja0yVoUzcpclp+3fHIWPwXzAkieEWcXBRZXjvIqBLoXZL2
irY3XmhhZnVXXK7XeQQ6xviRfO0OQZU9ZWOQ7vFga51yjpGV+9QDZcChbmTTmk+Z
jD9QnxX96hAEDzUvFyZ5kOoLFVnslS9FOAYyy3KjkNWaCMiokMC9hvuxdm86pMHC
Asp1A+PtEWDfXQPOZVdi7jHopA4GIamHqhvLnP+gm4bVIsJpXWFMG1RZKixzhNQd
FJvW6yFahb0QRORX107LrW+FBzscKYwnxpkTq+FSUDw6Ol+Evr7z2tNRbcoZP0js
zJpmlR52kaStvbi8WeNtnbHSnRWxS7lLsQVawYAj4hLHG/ep6eb5f3MtvyeWfC8v
YpF8gw7UkbtSsbdnOlZjqWXLO5g3X5pbGZYSEy2H5wNuBBTDo1aHyixsjSU1Q4qx
23p/vujauN3aoPR/Btinb0XhyPyLgVq0IeltFSGwDN5vhT3/LO8vGIGFO97EZq0/
OG2ldu0et4s1Cd2AybVi8xDXoJ1uhoEnX3h+VTYM7y3lO5b7Glwu19PSy+0+wS31
0r1OmG3SmvwpjCKrHoudFqYScJIvtMBH51cuWcHOA0ika2dACY34xHnj8Zy5YHC1
7bzm9FhhTtjTDjIgUqQEYqv6JcpZYgym+ZtmwXthHkcE+3TeXzzq3xV4rnb7cZK6
ltBZtckUerYZBbGtcSYDjpXOv1n7+vHiQy3kbriNgoKrVYvZbep5mX59DGZ3aOLX
jIFHsg97ptH+ymTWoodPTypUHkqLQ+gKAq+NMrivhuAQRAzuXl+XFsSF0VA/QlLk
fVUkZHxy9A0VmooXNLqlYb5eGREgATFtN2RgECeFtPxbO1snbcQQHbA9yIJVZEAK
P7bijurPMa6RNMrR5D4MrjEj9jIg0Zz01kl3d0JAWqKdvZoHF5dNYoF6a56glyic
/Do5k8nZ41KYOgjJk+DYH5JDy6LZdnhhKPHTChSMQVGR25pwrdHi0y4CY6Bkrkas
CwYxOag0xtqu9sGsh20oxw3XRwwolj1ioajT53M1g/ly1VDw+suS3AY4Cz/RZt47
7xMkD773oBWBfG0h3g3oI9KzPiTs00O4laP0nbBO0d+k59vwK+2P+itshcyqX8DB
zr+JZ57E6y8M9doOqPAx8fjrSAsmLKr8xRnz9RthRUkQgQjaG701RgXEXTIh+x59
Z0LRBsJsQvpLkOS4XEYrVorDH4uWOZV28/QUL2twb0Ji7VN6A5QoBRXmLDAoTClI
WQPEW7tgrDMCmnGbJB5sLoYoVaOzqW452fy8LTZ9vNA9NMk/O9m2polG6jKs4wPY
e8h38O5arJZrqLsgpqdC5kvEMgEaCuuZBbp5yqFCs/uh+hu6dKtEwbJ+32x3/Nqw
VOWNrhG6W+YAKi2DcpvTE+uqMVW6Xd4li1KZNfcpDlgLn39g+sPa6LQ2Nlyd+nBZ
KL7HIlf/7zCYeZDYZHvlOLr8XnV5GRdZYNnOkFx8Y1DO7g1rIMYcbtwxm4CqCzwk
zGS51HmfbkMhFN3usqVGRQcXKx1nPwhcQxV0uChyWgSZB0KePS66U5fHfvmMvi6r
qy47eKM2vXrXo8bs0nRvAEkWL7rlezD+y55gXfBOgbXIPW+Q2S7mr5xa6IiImqbe
3iMjv0NUyaGNHgl7w/suyJ8TQYXyqA56bty7CqHZfA/kuypBNvRtjimw5aop0oiv
gUGCpYp+HgMqg3aXI+pDgHpOJRBwNfb0JTrdb4mffbUFP2GZC3e+01xsq+hPo8sa
q81Uin+lS017MPmDwE22cfYurCDsyCCHq+s337I1zkn1rV7Jv+vEpyCB9W7pUidO
bkoxTsJflyIs5cYyjkbROwM6dcyQturiS/FOfyEz5iAppmUkBip/Dz4joVUQQh7k
w5G7PPDR1pjClAznp1e+F3tmrM0dSDccd4Pub1lwXMNqdzq6gXisjxMOkHOEgI5y
gxEHwVwguzLIieRNaAkcV72wbfNxl+BN+V4/P/NoGUSaxETA5PZ/aOEs3S0GIeAX
42PQJ5UMH6doOqr5Hn5KkAQlo9Bf/hD/rXcHA8eShrMStNiWDBd+CAYdmgZzB4O6
yRuFYJfwiSISzR0BVJVemCwsh/o36RLtaTV6T5cmSdZYsALH/We1f2+2DA+7j7CS
96KMPfIt2p4zUXtkbulNPXYsCIbELg02ZKc4WiupYBdQibzG9ZlqoHRA253q8qrJ
1rT8sSjkS15ukFwga6aaci1jMWTytuslyYu8SKjdsgtG2aY9sOkyGaSeHNp/VBM9
3UIb3ViuTGjVALZ5zGp2nUhOSnmFHFQA3aD6yqZXM3r5BlrOIGJYVX+yk+Qh6d1Y
m+O8dYPE/J7znqKnxIculicpkE5lUyR/tyNBu4yXoEW0ak9zf4XYK7ckF07blISx
lrDD0pFAM1t8BGGoZBklte0iqxTF0pz+awa3OGOz/SmjHFrrnGtFIyiBIcURpWE2
SopLOmiraoamNgxibLF30CxXg9JhZV2e0lZbE44iYSBjRCz4Qhj+xe38xDFvm2yI
LuP4jZXCTOKK6G1f9+YR5qCGWUkP5ux/yo/hn9MHTlASPkRkYUCTRdDUWuTUiJl9
v/rl/4hcvVRkTlJXq9NXoEY2nCWrRGSkxzsb4/Bf6pGTtbibKE/ajgWhQX43wjdY
P9tLd8wl1CmURGUvt8qvu/+grYY37iPWpFuuxYb3Utg3EMQbqsQp35pghpRfigdE
i3Ho1BC5CMouPS/Z0u7ytoYq8QiWAbeIkpk7eZLpDyNC0pPDyKQJJ/SmDznSo4Tn
6ZblzgWUj67gjymlr+sajsl4a1KD2B9tLN6rjsGToCVmQAcAPIuTA2C5gnjEPYi7
zhqO1n+BlZ/5Ogvn8+oVMp3SUWrxQyxez1GqYilgMlrVKM1mJjK9M+3jfXbqPshl
Jn//HS0oDyCCPgw9fjRsglmXFEN3LiwAmeQNIk01nl4ul+l8wu3nLrC/Qa8k3C1D
Xwels2LmFlqtxWJL1zuO6iESGPTBNCy5e9z4sv5Bb2qHSDyiKQtKr+8LJys/1Opc
/hA8eokmtTJXpS4+Aomj8TVMjQAeoiZmuHNZvdraHn7ns/S5YDRlHzhTmCG1krB/
1Xw0+Yh0kAC4L5+nsVpN8kpvJ23brlhrOusYAD8M1TAhzyNFBC9zcXs+jWfloZ35
hH23q8YK0XRCQKIuulLpSxrS2ea4UABibaJfKlprnFq3wRey4cMbddML1Wa2RJtF
J86+PhZgdUA1Yu0xwy+Hbh14jEMU/cHpIsGQqipi5Vg/81ohiXpUQD8zssD+aDkP
m5ATNqy/w5+5mT4R9EuNUGfnrtc7RWSXNL4cCyAUsG4MPprWc2GL+NAhIH+qZJa7
i6qcG6UFVHQXjur3lDJ5Md6KAp3tlGk2y0ZtYIeSPxXiK/h9vYCaKmZvPo29RLx4
ejVcruU8k8RlCtES5h8WdeXK0b+arKrZ3+MxCITtmq3N9XrdCS4z/EvbDYFxKCx9
y9vM+/q9pmFmtqoGcD0KhcEdtK8xQ/hnfNdrQUBWf25uUMFJP8isCVSPPuJDLTTq
Yy5piQIqe80ao21g+5NZ6qpDRXcYJ0SAhY9ELQwBWZm+uSoTzLk5bwk6L8rnE6Lv
wj7KvZms6YLl11OudYpMBJiMlFTq2aoccK1RUoReFm/DTYhpEH0ge9RDcGbGAEqh
6agWINIUgNHSUhTWVM98CE6JLfM/esSv5AV2OYJCBgVbjEyqHMhjcA1mFQEjYmfu
UFXXrkKSxKN7UZJd9ssYnvYgMHOFihIlfYMPAz2rhMfmOCcEZzNa6IqmCUScdiwY
jBMLhBN2hPX4bXoglLyZ86wB/p0xDK+GR25x9ul3O1jOfn6mpEQmY5L713FE8bws
EvFAqSfKtL5RRnKrYARQulEJh+tiCS2kc8I2AalGpF9Ys2eCx2X0QC1okv6fmAKm
F3RoUbudF1qXregIqEL2AfJhVJ/NMTXq0/E/qMg2UcA3lMX30yK5CG3Gqe4fte4j
zItiSSQ+lPV30owoMJ5B1xIGi4Jsi0uldrwQJ4CAhof/bgey+28qlNxmVb7wgFEq
Up4uBvId56M/vnNBwpGEWUypDaG17I/IvbK7MLZ36MGaZgf6o8CmMxuYAN5QShr6
9iVtqHC+Zo8aoLFRNkSIW47XoI6G0oO7N3jPAbXNPEBML3OCcIEJnGVEuwnR5I79
CQ63z54mXbdpsNtM0yg6I2KpuZnBlFjLmuZlyVJqDdQcw2VqbcwptHKCt4q+FekF
bAoxbxlLXYKNVUr3Mzi9+Tc8jJLYybZsNZ52InOGdD1vxVl3G574HRrcCHKbLfJv
EA+X+YUn0qvYFPpOhKiZ2UeEpF3p8GFmFLKy0xkzap9jrUQuV4Y37sO9WtWx682t
NinB+EpGGTRtbc7e3S8jX9loOhtCWvdpniScAPaL1r+5S+Sy3GrCQopFGcxs9GHn
GYwNIadbG0n0eeBPV5TcqmaSD0dJbdFjLp7pTP6AUnoZ5NE5SZsV96SOkliJ5Gz4
RRSFOq3pORrNiVRkgSHr1mS5Xs3nYZZkSPiRiR23Nw+NspjiL0Y53k5ugjIXtP6O
KY22EMppHCySZak4AshsTxsK/5Bo1VaAhh+XDsPrhJ94dDDXTtFAt7A33M+K6oL2
W2y/dE8nqxxu7MzCBe8Y5muM/oiuKeSfZ/lApmSy6AbqFQJjfcSg+U3HkvsoN9Vl
xFm5Dty27ZrKc1ZEKxpMMqP64S6ANeAAHCHUSWaBo+1huS94uT80/vZDhCXiLZVh
NdYpwUFrCQLuxHOzE2vzQclA8p/6wUQWiHpAeJqJgGepBkrM4zMn0STF6KWcAFd/
yqlsIHse7tJcdimbTRC0Bqwqr9+inreJHhLrTcYDjqGADw7kVMloLn7Q0P4YG55J
gZJBJBXfFju70iFnHqyT6Xp3phJGprAG/withiWvtV/oKOZwR53YkixZ/iWNBbNA
oJvzp5sYkapgQuzX0boIE8VKnvz6Zslr/J8zaLDcLMdDdcdlFfa3R+8TBiRfc+4U
tU3lj+L/rQXhctrCC1uidzr6jsyVx+wMCSIEBDHSRGJGB4qUN773aSGi0WwHXtrw
Z88+WTXO/ZoQn/6ndDtpJx8eiADGYg3uWCNFrCS8VZ5F+SnpbGCf/WBow4auI5x/
H7N6T8WXaqS6p1MOClz2ausSfwpO2Qj1FRNaIgJFSdFN/c8l0x9pLzdFdI8Xc+IM
mE10HNE+M7EeqTQNBpzsnp/JW53aSwoFGSG8a+WP1reul32MtXLNIQIJJDwAR+vT
wjJXf59ayx2442FWNsikveMoo8kBdOwUe1ldkDnXizXTtkQjoVQJq+3FtmkPt1G6
P5wwWBxnCIY2tUIOW7/ZHyCDe9qZd9ilPjEtw5y3ASwz3XajTJUTXYE2w6Eb8HjT
CqQ/5acA/B8xb3UO61/8SxYv/7Te8K1ni16ogEzerJoC76b6WvOnyF93nTii+wsa
eXFhTU8sPT5aLI5y27qjx8rocWBQbySPZAcKxShB6TyGwUbQdxvC0SvCX/hcK2S2
TPfsYgYBxXrlnlLc2wqZ3pV46ctC15pNd0fuKWgQDTri2uD848rR4CHb+G5Kd8vQ
V7lpExI1MHzZr6936ankJNLK4O27F0msY2001c0YxG2VAmV49MfxmuGphjYaB0hI
PUu43Gv17Kqa/Ci/3QQ3Cc1ZH73KddOQLz4cp3aFsDJrv0D2Z92CTUZdgwzzXIp+
pawxsAEjFNeHZLBY67xJvgkUkAhdyNbau2SbVFAKDjex8tpdgXzDHHN9hcxtPzXi
qM3/sfyTEQPWFxn2TlcZV7PvrdvDiWaWiCaBn76sWCmh5/BNF/i/VV+ZoxmbLL/V
N2/AHXiRwwJMGzrr/jeUTcj+rCZ6Hw/zJ5a1T625Dw38WAN6QrhGq44mAYPuv2ZI
RbS/F3pZ2AlXduKK8iynA7IQjbn+duynTmKVrHcgBkztcL0T9I3wrJ2kFp0XyO9b
2K8j7K897kF9S99diSr6F+yJ/RtzgKKAqIoiuslgjzzr/BztzGgOEO2VyfR6TDKX
jq6T5zr17Xi6Bp+oNJyKgFDqhzJF8BBstRjMqN85whjWYo162egKM+chI5mRnFW6
6fy9i+CrNLFif5rPWNOzN1zvSxXiIkq7VAkZNgUKESiZuTAt31su1H4nbqhQUvs2
Jul3FdjEgBq0latjMI2kM+nj2yHmOIvqTdowSiS+ktQ2pkcKvcgg0DdUvcSEYHCw
5VN+mlN0+TK7Cji8iK70ufu7xXPWFJRfpeDIGC4yaljE0RdWEKAYknbiVFyO/tJr
xKbvLIJS0a4CCECOs7w0nmViSe7SYep3+Bfl68hy1KE7UrejERV6H8bycbPNHTYi
UCE5O8lX931C5JJV8E5GUpl+rliDAxryPRanqdqFj6hbk/h/IDw0b4FycappCwUH
9sOXR5DzD51c8xmzriPjmcUJD0uV/jTCrblkbKVbBpl8dP8elWZKpCEsNW9yQjH3
qA9nL1sIVBlP2N8BHoTnkXQbPtM1OkgVEfRAMaX5KW9v7iciPEBBxhGyBwMm7BdW
MVwhe/ADDhiqQRYUt0STdl/zExnjiqPRiDY7FAsMLmIB7XHpomwHT1NDthugIsi7
33JvbGn0/CMpeOSB8SNHmG86lSHHjkcyEzn2J4jqx0lWEHpFL2BSR7VnSl3uOjIk
g5/ncgO4Q9FsIFw/5smEFcBJHFLL+ZtZavgY8yxP7+x37kBlc8NB7UyiPdbtjtvn
gu9nROoWWYIPq7tK5rgk51nCbZvuDPQHPA8zBXOSCb+kl7oaIvDA+ODXUAvqEBjF
kSIj8eeVJ7IeIvScQSRwGenVm8eQSy08xlNlYbSRaJCFmDWsCZ2JBqf3/+KUKAf+
rCnqcfwkqWL7B6IV8hhOnMHBaNHheKgvmxBJB58HFPDjYj+iwo54BdsBGhMWMQxk
cUwoPCrTgvuyTsEhKjMQNoIBA7sOXblo4QwhggOY3u8ccCwAlImVXL2vGLVKyxIM
mUkCPb61KVHkH1GPkya8h9OMJbeLAEjeTYt8V14P9ABCIx5eRXOoLbANF2sPoJvZ
BI9bpBbU4BnPv/zLSXoDBnm/1A37dYSWLlLnAxWnuxfS/hwhbTjrOJQjwzHYmDwW
ziHjhelV3v6KcEXFnEY7OAxeshBY5FsgAVBJ8ANFJ7f7/N/e1gjHKSDzU5E4uJIY
zS6dhYVmB83NT+CDP3bmG457IbP7INh4oNsQEXGPRy1XJEZDo5ZhnYWOCqVKs2JF
ydLRMYMvt6L6pbugwGO/i2B+DmGmMZh1P+nabJKjhjHdR+P+7Orps//IsGG4e3Yx
U/B9E1EToyvPvmV4O580ygkaexqKSrb3GCNK7ozP37iP1eO9q6hgSHYoPtZo8Jez
TTAeljtJ+E26NheaXXHCl95oXvkfLyEdHsyXG8GcZaMZIfTrYQJT1sh/h4fKv4Xb
QRFQ8T/v6cWQEOThHoWOLU+S5WnJAF68Y1ywp+8P3K209dK3UFWmF0nND/mJTEWT
s7uQD57ConVW4u8empnbJzj0mWWo4YOR6Xm56Q2PfJhzysHyvDBHY4b7oma3XYzp
eQVgSwvJAgQ4GamV59ToKH734udu4KDi6LsKJNtDUl0Byd9/KH+v7+BowoG6PogU
vtTofcimIoteWPeDpv4I7zSA1G3pYAtwXPssQ/xzbsy3kug+tIhvjEd0GM51eU9i
gmVDEjVqZRN5v+qvQsCgBTaz8EpWKdo1xWZw6+3OAR0oxaRDG4gqEmZ3ZZwD/9fh
orf5ba3O7JzIV5LcpGUnh40diLT4Cxn9L4eYavd3tJhVCkhvWVuRqch1a3poKfJQ
ooNaQqYC6ZnSwfJQOVk1rNH0NC9YL9LU640PvSQfa/EskwerLUmY5TZIqeYZiD+k
yaDme5Ud48TB0mlnsSq+PYcWi+uF1TRiWSDPVGOFB2jFP3Qoa1xeMV9SaXmoXoI+
cYJ167DMSYSPzDycGWvml1HVFTljIwrBJToBtI08TSswF+Q22f9EAM8wBeOqXHKy
3ye63NQs/2iTatmrGrbPdh0Osx3bYWUpz2vMz1PTXigpVfKhHoiwMroPqw2Lixle
h0DI87wfvy4YNM9mBaUl156CgjxlUAv5Ig+834XAo+U3nGJO1cQQz4BC0Dlrtdbp
O/ydVN9CQmD4uxoWH6hXemzFFtC/MRxUvDBNVREXovod/ucwowHJz1xQHMNHgkIQ
uPgwc0RmTFKN6cS7fF4L3zELaDwHwCs/cu5hGAawN0q252k9DT4RJS6QY2TGG8l8
SMTM5hn+sin4Ucbgk/PqWg1PGdeNMYJ7h3HEGpuBVvOTvbyewWiY8hke8zG+fZZ5
xKuNGAs1O5y1GkEU4pCqbOpZQ/ZOjG5oFH4Wy+1KfejWXl0Zqiut7TgEFwVzbLHo
r8Ydm0N90A2gh+KIQKSXKeejan5l/J3w765a30DRuFuqjF92beQjvijJ5uARMn0I
mlbtb9ZgCxaN0wVKpwdhePn7d2Ae2LIGpqsoz0N0Yba/uwV973p/OkQ+imeqELdL
19TlQPqtkH+Hf0zE1/HWBxCMF5616kuBWdD+vmGvsBX4hJ0kQvL3YNnpkUCK2qsG
iortoBlCGqEX3BVi2ZVVTvmUhObSTs1WQySC842pWbgzwkDJ4c1fZ4loXaYIT7Kl
6g8aB4IQyEqTxLdTR3Yn8NMorrp3XOVE2MAp9tc7TP2F7skVV5l7roUb3t4fM1z+
sF5jU9mpB2IIQW6kWPktf1j+OZYaB//+DBfLpwAlxcWsfBTkrWioYDzk4ZlTDsTp
C6aQN1UdCXoHzQDuezVnHaCgyog+qWD0wlyLBRWgGAoVtoqlq499t4IbnWFsXnKv
D7AeynlAg6XH3M4i2Vd7zJZtR46k1KCL4dk4UTSPoHcfb/4LeZfwyHqIFnJlINY+
j1c0zDAjbjy7js8MjwoGDY5B2EAIXtPFqp81hxK9xjG9gPNdpr5Bz4jI8nsH/dO3
WY9npXRFeONJ5gE2WVr7oYubUreFljsdTpaH7kjnBNCWS4PZgClBMaOJVfyXTlq7
rc3I+yLmxAxuaSXaw86tP969kta1WmWyPI1CYoaCtPrJu0NUQ1m3xFRnouapEnhi
Sn0OzI8P9Bej1YKhViOUp0jWAbOWZ0WVbBDRMhXCkSPd4zpJBmD10OJ1BD2jzuwU
N5EKt4bF0s8C2r+BwDp3u+zZ7RAM0uW+l+GsylG/pvn3ulbS4499jpOoot6aw0vw
nTPZNCXBdupzY7n7aDyek5fOR/VoJcZHjJt8G0lZpY9a4qaIH6gM++elf0gzBfcl
9hv+c2a+nam4rVMiB6UuQSYcddhdFsiATMdV2J9jTpt/xdStluXbjSQVm9LxuACm
Q2Xa9ZW6zAQLm6hZtDVfssAA5IwrUftma5seZK+FJJIG+IL29+qtRpZdNV441IgX
A7jFdtK+B5Wb0PUEkmgvr2U22uauqPV76WhkEH9QaqEdyL+aYqmBVSyPpoqMD422
qp8cp0Uu5zX9SSgBARSeDv9pjAdSa8OokTe1yJMDCibHdMbe+wv+i5XMwJjk2c1T
PDRQWncy4X5ID/PTMJGU+3+LT2n48evDbT3ziUnOVr1w//b8xKYlnTC6AMuAXS5K
oUUIKkKlyDARgECl+SNxnwu8tfK5rEGj+nkZX+0WpQkNH5cbQjDiIB+4Cz6Afdm5
2LMNCgzBOp/62BwH1oBvQQQKdt98o1CR7LhOBw2WMLO2DH6pluks00rMzO2l7Bu2
c7pFgoLyUrEM9W+owoMIAE5SKyhzrDKOu7ZhGvsimJGzVF5TWeK6uZBHVWD2CAZj
RnQGPGrrNiboOR62zx5yaYdsWhvWJBMWgQPwkDKcrpNghdKRytlHSK1l+SapO+KE
RMUEyvDqTjBPem9iceUxm1hKv+ivWee2pTNmDllCVj3ZGKjfn3mOATbF7CBNWOVk
EXDjwvEhgMLaIwA2djMcwv/NcGby3bLjo8myl7xKC6vFj08zqZ3XrH0rSSMTKLxw
HQW1rT0tw8Xi5Lm6MP0HGilwCUwXF9k5HojcqjKZhFqFopvhIToY7/Dxp1ODzuO+
HBHWgKe951JZgNQ9v1s5A5dKIZm9REISLjcRlOkTj3K9oSlYGAIJLoufmbOrXTRs
bZM9oQnvnXiWDSBjeHCT6pRImPLcwObdXDEHM6m3G5It5pFDn9h8cE0dfv0MoDgi
yVwQVKliOHKt1L+F76i0rPYVZOAysmYLyz0YWPIaV7hsJgiVw4zvgg//ApaIn8n/
OfhMsi6frW2XLR5A0xE3eF8S6N3bDFj3cYSjpnLfWvAUztHFfvA728NlmW/lXLLA
7PBuw2z/Gp9DQfTLZWE8sTOwfcH3elTRjGCS+r9ZtiGZsh5XuJoQqer2hkHwnJX5
SpR18erVGBhw3bnFIp68+rIMUXBAvhwy4QZKWPf0DmZiEjEkNRn1b9yiFKwYwJTb
BSGJjp/VCep7PSDDJdE0HyaDnQgbeKVEKNm3lL7uYu/Rzv6WnFwxTwu6FlTKN91x
wunko/XIyY/ouPP6rHrZCF/YWWsKz7GltyLY2+XabziNIWBxpn7kzsvFnhu7EuoS
eQu2++R+X9tzKf9eYDmv48O/xhRiid/bM1YJ9tFmBaSy5vO+Ug/+iHCsRrUzmbxa
xlrTVcjoPc7++NJGmRfHqb0+huZOFGjzDRI3IIt4na8qHvXTZtc4SAY5bJFJ2AO+
2dfYsWshvH/tI52KhsIbIEGU36Sb+fBdcOhp8y9MohsHYkqDcmirJ2B4hONZ9yWf
xFSLRbA+xtkNbP4C2jY5iynJNDevi/8i47KnDFowQXEHoNDpSU1sk3rWjMl6+rws
Xytw0LyB6Mq29X9lYTxSRLdCry2oFfBBlvVZwxnrVbtVlX5X4skA8arzqmXGbFFE
lzVuWXz7/ja8/jfWKJgG7ncuIqsUfwcFbl8vqp/v4V60xvDgVJZpfXwtQ/myKwfl
h9yGuj2siJWQPnh13/enwTtxQSa63X8Rl5OpdnCV/SlBIsZBEPPqgPcq9ltbnec/
6CxsZPXtVMhqD8tlZltb7RQwVIEhv2lUHHON+KZ/KhB9EE2ABoWSwYcHyzR2qxsV
bpGq1NKAXguS65SygEso58Zzl2+ZbgDWUHyJOkW8hrJB+vo8ZsmbRz60TiiFi3NS
kHA1WhXXcyETX/F7U/2LMwIS7rvugSNVhlE5P9pzbSNyTSJYZFVy/TPYWP5k/990
X6q1ua3OFeUWuDfd2ZPmSTGtQ90k0pN1lRq+7G7okc2vnLGNmwOhdNsRSnJ0OFUn
G3RXsL26tPOfNfZDIz82rW5fZa1vzLvQRFhSJR4dLN0xhLJHq7aC3t7T0C82lPiq
BM7l6ZP9RGFGCP0B5ENN/7C0JPAEiLGcXWe6li5IEKc4w+LFRLwbbj/DGFdq6OYO
rNPIPmE+WF6sJxaXrcwi2aiaKBWuYgRuudRxYrTuPYCMhLabDue0SPPQUAz5N+yO
jaMjU3WZQ2rFNsZHa0E3jOH2xSG3gSiyIJyecplv0DvOkZWiroe60tQTiYJSznoH
LXJq2LKlH5Ybpg227lrAetyvVtgEtFumx4CdJvQo68sqlrHqXuXQCyg92XfzSqeU
6oxYRejxAdRqjUfCVDTe+icH+GLchkuZXOMjMaLlbP1Zk8ucsu16wA6PoFhn7kuk
Fge5ulb4zromNLlJke0eLqBwgVVFWxOBOeQXfSMAYBTRMrdWu9Z2ZDrmoz9Co+xw
AZddxZsPcgX2Z6Qv9EVj9VUEKLEi4gS9Lv9B4kqWuG9VLFJ5CGAnb/qHEcrP6MJe
YrGBg8EnWVDrL92CQjuIK2NDsOt6Hq2fMNZyyJ4TbRaBsM83eDD3YyjscPNUWUxy
dt7X7j+sQrJua5095Di0h2XXxBPgb4sHM1ALbbT52CcF094l+K9WezXMZ2HB+Q4v
ndZIT1HIZhTcDotN3QaSOi88jvxy3lanuWpFWIgEveAre5znvXEwT3FFbU3nJ4k1
eIUL1ub3ka8DmzHtpy8ImKO87E4T7Or54sBtG1LvQGbCXVaXKp7zK6FXYpdsPkvw
9kYe1i+ENHfNshO6ikd+xWZvwNMHA27eRzoQNpJiVdGpmEftU385AJKaZS2SSTAz
mjmENHYlIEQBrWUM+wSgfQHOTmUZQfcKWTqV1wSbO7k1LJ+ZVrT9ASPgXYOa/YzL
fWZWJW0cJgrDT11SuAxk2jBXj4mo/hUMyAdAobHUp2EMbCQ9qelZ7jNimF86F/Lx
rvAvaotpotjqPGUtqFl/6dBkyDfe/qjM2a0U6TuYIxwvbAU5H26tsZjF8SmQ0uVw
t25sFO/2xoqQoJ5ffza5eG+V8gU+Bp7z5ReiKJ2HSMivSi1MUQG5p4ycDTIsFEYR
BfG85Zzeau0rAJoy3DzGIEWu9NQC/fM6NAnVWEcE9oclqDhNMi+nsjY4NivHE9Wh
/r8CKpTCsEQ6nu05ciAsBQM1EtIeFTHmKUH5zGEu+5BwvStzn+42y1HC2cfiXiHy
7xl6Zj3KtmwfDvpq29FjJkBqInDOq4KOrvUhyiPFKD89Vblb/bAo0WSwxQ7g8mOC
X4K/M7vinnjpW4MWKz44GGmqjDH/3zzOKg7rWK9ji+N7+FEL8sxmeXvYovZLEGYM
pf9jZuJR5aJBLax6B/tEcB9AIvZlECHIgXmzJ7REWbgsyk19CthuGZU56iajijxn
SY4Uc+c3nyTSs2vfPsay6gBi0eVQkeQiwjuvTx4hjggGhbXprXL8jEnlB2Tya/Du
4HJCK4ldL6oRWECJ7MEfkIiW7nIMomRF+VqysRy+i/ZdnjbMusA2TnVib+KlR8Nx
orcT2W4XmIfjvQhx0M29jYFsA5Sb5nVY+cC/0nieiq76pbr+1fJfRBgu/ilWBKSm
8HeG7Tx/n3L1TV8ykk+fk0H7A3RBfz1OjhTv/ry7oInqJ8u7MRV13fzBlftFWjwb
gbCtAAF5SSukZ/mV9FXYL926w8hglg90mY2Duhhun1T9Kl+U2ZBMG7H+fVg65oP/
qO028kFAN2xS0kfBhsyoM87buUAz1xZY3a+KyAF2fZOmVKZN6O52XmtBJZ/CUVc7
fp7ZFj70nZsmk2Hq9LOcJGVD2+rybAhVVgCQamtC6sm4P7nEVXy0Q6uX/FVF1+cE
tLc73TyBp3u1J3nZIYPrlBd33G04S+LrivAml9rke3BeqWtUkEFuEd8riHXbYazk
3NLcmwZXkJrhfiYUz8IzoYWDcBQ4e3l5TOkDJeZ7xZr+JDgzWI2asESZ5nnkHA7d
MO3B6JfTOxs8tbWPL1CGDEOuPrpNzMkn0bcF469ew57ChpwGzVFsi8fVeWvxC9mZ
shsbJuxKmAHFpACVDGoXMJMI8/VtLf4UmVPAjdytg7lRfrLMNUBbs3vouHfqkWCI
n7Lj5eGT8jQxx2Sz0LSHV5tDM5H4bDExjLzSykPRsxrvPpxw3JAxLaE8l+2JbA0A
I/yy0DtdkL0NuNCBJ1Xss5t1GT4QomxIWxUmSBQdEg7K5UB27d8egIKAYisvswTZ
TtSy0WBG+fUa5FjeN/mTk+CsGqMP6UFbW3IKd+gVr/sqGlEEv6cor6E1RZfzryBo
bYQMq7W6liDN1E5NZ6HYXcbpgwoAI8M2eQUumu4qycgsTEVmIPvgx85QpCqlzNqw
l8fl24JzpIK1EbSD5ITx50FuYkQc0JMg+8OHAT2n+vvAGBqWQWDpz6rTGTNtgPDs
/bcPljpNIigIv6K1LmpnG5xpjEiHNpE6tmaitrDwGC6hvDxwWmHsYykFricMb8OU
4bSvtREiPz7birmjkuiRDk3TNwxe+NdJDmG3ss4g5NNyV+XfhurjsAoXy79YFSXs
+UO47BM6aW0dlJrKHajSQE8NWoCLzIFmg9VsDTj7KGoOaNzY4DlewZ7++uVgCZ5m
T+sgEoiAfItwdroB83I5lSRM3+kUVT9aM24rsC6UgmeuT328TQkYL8uvxDXceYkV
yPPvhWg9OKQdyoaDKjCWVYWANpLKiC1x1JCmqS8S8xdGOh525bkpkaaVoN1cLh3N
tFIxkR/Kp7Z/IRmCGr9ywfusiI/X2UklQNqHoPIcIfS8cxaYgTlvmfUSqiJaCyHR
98kmH9gy6SOk/+xJ5Q8deAtLMLp5wdv05Us5IqXjSr3PiQlnmCt3mpsx2H47yqf/
S6jQmWPgvNPm1zCa7zUQpqtmKkISnXpZZSiS6togUm2PJPtDf8DHwOO0V/gAs7pU
Jjo1W+mihtDH6skYJ5TVmXY97VfYrrNw3dXkG578v7Dvilq6i0z3hFxT5Dq5n1gR
fpjjNbwb31PpkdH8xi3BjShfU+TlxjCMhW/Z7jWtYXcTFPHB+npKQbJbuH/2GqAo
DtVPYsf8EisDsCn/5ZFgAjnXM2BVPZmb4d4ZfPmnfGyBBs5ZfB+1Sxflt40bNEks
RnWAHKZosEERgN412bLwI/rq9C5/ItDllcMqI3qWoHIEF+3TUy0hFafGCfk++J1E
QYaFgLtVl5kc+taf8NsoD6rrTNPGpji2fYcYZoZCWhoGmjG3J7DCh9197+7WCWu2
aknP2lIIPGabsrKEGVnGqzWfXcrk+J8Ki0+OLtait1xK//2QEhaARR5bbjiYWRZY
qdE3Vv3fnKnbdwOrVg2s7QghSLVlxmb8dzxVavHk6xcOVsoD0YxWRWXIwTJtOqEb
boVc3PSWS6pCYkqfk/fdNCevN6MtMK/uJ8+bMtCSmKJxbcRwRSp3STCr0IF5VruH
DxqA5rpl2uqc8cdfesuC6OL4pL0+fLqGzOgTitJpLm8N+AWDBIgFhtBxlfWk0vbj
rmlx3RuswizUSRNJR62OnDXuu9mVszoVszFtkTjmJPRQxux0UQxOniJVzh92zkfe
aRxo8XCVLrFNzKyHYurhNq9o0kDQPlmEpunTMC/racSFeOmylXJy0rheVcNZyvRG
PCtcumLnZP1NHcOQ3uE6pCP25reeF3SmdiqrmS2qXvCcMGNSSTt5TZuaIJ74PHJs
2mceKu72m7Aof0gZv+jaiR/zI9DRMeNdQhbRL8B952rhVRdyLI7mbXOI0gTWQ9w0
lvCXJ7Cn+ssYWr4ezH7BuHb8wKOWM26qXhwL+pWTnPr9T9hLwy/BpCxoQxDqwQiJ
VQdDFjTE8nfKEh++rziRK9/mIZt3mFHYOOLCSE7MNYVti9V+1SpTSMt44m154TDE
GT5339kXJ+lEnm7fCPAkMotJxZSsdenXkQRt22Y2z1HkNsiA2kxUNzaDQ4U3M25m
h0j4nhV2QF3K7CUXejQOrFS7AwgIdagiUqhOPblh4roA23Kmk21Q0wZ3ZAqiaHps
bFv8ZaO+/Y7LjKZSrZbJgiKBv1s1UliVAgqJJnK63dMYVgPRmECctktiDtOWScuo
6s+/SaEP3LT6isB+hGMid3GnxZE2lu3GrmYkC6SLrsOQxlWyQej6waWFPi/NfG6N
yzuwdgPN80Zk3XTmR6I330BQTBqjk9DnRB/17Xm/Ho/RkmPYi88efs/vec09n0h9
SKzDhpseuTqh4EJb3W3Ed2Bi+KUr/ItIAQ+mjEnuxSzIXA1ihdBNEvroA0SW5x8v
Y1KVzrj3xMzxaLxRXHIrPNDb2N2kaEM+VvBEEUkqRtLE30LgA2DB9ZCc+bmjbqRo
XESIyp4n35ibNxn4PQp3gGd7FTgjsSZj0ArWz88QF3eYduJBKs5VZNuciqnJRoD3
L6UM4kHY6Hz1IYhkvpsttKElEzDDqClynte3t+kLJXLLU+pUHZiRkBetjzUrRs1D
z+pHrO/LvGxJBfmISKYTZ5LPYKTuLp4CIAGC5+XVLCLStrbUpMcoUYy21xnxRHWM
NSOCvrlFDfUll0NZso55ZCeBt78V3jLW+1Ghk+zO/Bztv4Yiq/2MbkeC5VBlDhlZ
+pE4YZ2WiDxfNoVRGUSlh6C0zF+pbK8YqBDjq30TAGEnUJYGlqMLiqfeGMKQq8aK
quRThjBDYgg89HatR9neUSd1urrM8U5WuYK+z5Np+R/kfEMvzy74mZhUzbNcwOmY
dPlwUPDf21H4cbjyi8dqFK9A/bJntHsiKwIT4EjE2fwnhhheHr6hdIqJVQ4EzWat
KOWfzr83BMHMvOEJ2E9ydfWI9t9L4Is3iH5V9Illr5PnG8erLbfurL2G3qMISW4j
LWNOzHKOXmASBeYDmiWDJRyFKwHylRhErtyOJob+hW6WsQnZwFZuarTdXjLDKPSM
Y2Y3vSEYDt5CaNspGqsbVaPVm688PF2JmnLnWx6RAW1NobfWwACG+Bn7HRFtehi9
LPgYuqsaBEnvnMSvdMEBolcO3cRaYkWl3F703alQ3yhwptj3sCMRVgQP2W9MTM7B
dwqyxm0l49JGyGeUweXEcUXUrPNOPR0XPCevLQqeOBhYjYxDDMLp2rEoC+gk9mMt
7DmY12cKzZbUwwg6YTnu5Pem5VsVis1NLqxbZvCrkdPHDhBFjJxybSbIr7e5lPzd
nGCavwzyaI6JeEBynAdRkMQwmqghKqCyLI4j46Ud+g+bmXjVrUJuQHmEkOcR/BIk
v6emFT0eTFqJYX9XpTAe/POnhkCpMtkKpdC/xNUW9AMOLVos/OJ2qXVvOBBs0qTn
PBynHZF8d77JkzR9KAcFAomrf/EHAhecKRsbael3GLGGgC48JJS5ULXRB/iEcLuL
jnFW/+FQk3UWQmzz1uzhMwQj/B3Krge3TOkhlBjtlcVTjoHydEEKfOheZbrb47eh
HLT95AIEL7Yiat3se7ExC7gvMc/j16KiPsp16aXpxDr1JUlhEUiAwfPp61JOhVvV
3uI7PrNJhmS26y8lyEzEHIykaPDekZS9HWeDvBejd3Qg5vWrhRFRjWhwwKHji9/C
wnEE5JlDO74ZTrbM6zl1INnliqcFaucRYWgwRVpnNvuupLZB+vabcT6MujOQynvj
XhF5Lfw3RWtSlh8/e8qZPy4VH/8n/QUmJ+OLfAqfmb6te5NwlUxcvJOO5cJmXuLy
JBdNi4uuyMC7TWlxFMkg53HAVdAPZU3Z2B8PYNtHAnkLULIsax6qal56aqndJdbX
tb5+Lk6Zhca0DAedKtYQ+v45WLddHvzgTPfjJ6HII6SKV25GAuT1puCwvpIhTZf1
TtQuWubLJlZ157mvKGjpFWusMg6+xxnq9ZpcfL/u9P0VgGRRKI4dTC0nPAcYL5lj
E4aVyyCS0LiVAX/4pf/aiZB9YNmaPBpa3YcvckXLeBFIE8YI4q2TB01/3Dd6yXUY
7IOmeL6siYnS++kdHV8eQu8efTAdt0wG85NL/H+szp8bIWAXY6m2wT8hcC4TYUnA
5tM26zmogtPygLtutv7E5xS0Yn0ppyZkxt4oG9ta41sdTqkXMkF9gzm4fN5D1Azq
aJoouU4+CsxtECeohCJTaC3TOg29iRIy1N6i1gELiJEf3wgnMBPWQ1HUJlAeC0Bs
UJYjkxi6d6GhQlnYQkwC2PfrizUvfFs8QC/X8cPoPcLiHLBVGg5oZsbfTwh4TKgL
ckpBR5HXul5EvINNaSj4ktkIAJHXwBiKhZ8ShFua3JDHkbQ8qwtGXj+eBsk72PM2
sPfP5Bafm1xhBKLCCSz/qRzaON6jfhzJ0pip+aREWVugH3zCSVjV9yO2i9+l90Ue
ZSiqPyq5LOgnYi+ZB5MJ7Balfk96+EDGqEEETn5Eet7oZltu/VRT2Fcx5Y9pdEuu
FMEmjzs6EkK9TNF1zMQ68+NOwlBsudBJppKoBgrBsGAomXqf7EJY6Mpw/UC+lfrq
7O4BDZIE6ZJtLtFIXtKCUuDRY9GLAC92+7XWvywGN0rYa3/VtLfS2sVZZX5Lu+jj
QYvoYf0hxRQc6vE9QuC3hK6ym//06Ohm7//UFpS2mVZrt2Sw//cZR7D9ziaWcU+o
Qf67Kh6/ayUmJEO76qMknkvWjRJliAJ5QPp6ViPCZ7Q2OCu3ebQoOo0gVHuZycDc
vnspo1FALMeprO2TLm1saEDkfRv9q0lsfUUnGL2qtCvw7qteSuQUyH1x3LNsO4sf
TbHKNvlRIOxDATWllsni8Az374xcPX2llk04ID/2kFfDzJ8OW574giTeo3bCkwyB
YT3TJBhOq1UsBQylYYCDT3c3AJz0QDi2FPB/XAnfj3iiM8yX4NLTRqrOAFCg2XBk
YuViQ4jsDg07ccQk2TssIuDWDTOsDy1kschxuYr2zwKOBpW8Zt/bhZ8lGb9RO2nY
QgSAMKGZoOLqG2/bqnABgwUIM3ZMF9FfFRxtY0+SMfWZKN6PxvyiOZ6TCPBIr6vM
xb5DMWVpeOD0/9VA01JToFBoO8QJ1T+S59bRBdPXHi5vKgGxBNibvxJxYe14SaAg
ZtOntOp2/+o0BVzDw9XaXQKPSV4Uept8EbHkReSroFei5CRAy0ouAOhYIsESZM+U
g4AqgQs7OzA7rw8Kxd6isJVKthCFNWjftOjhgZYsVq5dqTIi05pA7NDI1/uS5xGQ
LSWqwEIX3LgrbvuQ4RFdHT8vgLWL4sqtI/c+0BTbJaqb8njjJeeZdBsUQ2cxqAGw
aDm/2L4F1QF20F+YqXeCnA7yDB2Qs+4BHIdJmce0HwxhpeL7batc13ZT7YyOy1bW
HTgOcQQ62LuzldYySbUu7G3ofNU55+r2vPkpLkJQancREIZn9m1zmy/eqs0nkrzn
O5S7qsQsL+rxrQh7lFCVKWAThCVE2u0GisBA6qCKYpsoF6P4CNoBWtiiP0jUwvcO
3Q1hstZniI2jb49ShJJYzw4QBzduUVVFdyv+wMwWRmmwbICBaMv9hmcRP1Rtw5eV
WTrai/GbjH4Yl308jHUOkM4EAipuWDKZui8dn6gXNaCsEnwpernyQ8IkQ4hywcr/
Ec32FUb7jz6uSjBDlmdsMCr2d9s2fKVVAwB2NR1l2i7S/n0ekcCybXvPR7Fl/8Jj
Api+IbuzWUM2elE077sCo36bKJxiMCIPD/mYnKwFrWaEqeeXD15dyaRzOX4OXFWG
7ditkATFhKcORFSTofOrseWwX0aIafoQ6Dr2APd8cMrMoS3Zy8GlCU8CQem7kIBc
oQ9VkKfwfLytcmEfAMuMTkSgeaB43/mlBEJO4dowkxOiPaYRgqp2gb0YU2FU/TLS
Q1hzLPkP1R5TSBmYUKbuaWEzw8U6T2sTH3LhrJG8QIV9z7DIQsmshLIN4zygKtEv
zLITJlXo9Q4iaOOts1Wx5bywmideUI0671jUlCuudv0r4gBlY7zFvQW1bj9fJqGg
RTxBACiBywCkmV/BH9GKIHlAW82BxmE0k+wrYFLyMQptzVPODJqi1a0tp3HM4+DV
psxFnPQzoXQH9MtI++WvPigsl+Lu4ebKfQz5yVA6Il4B+AC/iQ824OIKaUUZ/RAV
ZzXvJ4M735A8dYmTsV5e+Xfj4K4WFFh3HRzC/il/kB9sct/5b+dFNEFGenD6u997
QJm6pDTflrU/Ru2OSEOU5CRtrtHffOCJVTXoXPYiGw1qKcisBJNviRpnliPfHaZh
pH98TsBlNt3wyaB19rM2HSk8ZZr/eWBGbBzUL7kSD3JZubVRk16rtRPqEodXSWz+
Rufy4qzklWhtKJkik5O9obHgroRCGZOt/EHnrvXOzCYXYMivmcIp5SEeSqBMLfcb
rhuaqPlC4ZNl1gU7xmskHqk4c8hAR3PFam80FlOq4V5WX0+oh4qLkfnCOW0I2Fgm
SnBuDWGQcldZWAy6AmR/ccwyYgUSvc25U68kg8oASSxNLDFJJSEFYPVCq7mSBMKJ
yWrEn+Ff+5EbXpyNWV/VoAtKi244Wj7R/HQ32do4ulKt6x1Uy9CucqTIDZQmJphq
ph8snoAjeboqKkpyGnqhmSGM2V5gUP0VjGmKM+KC/PRIAopdUv91Dv/SGI/EO4xb
cCw9nS2pPaCMENL7wu4gbfaAIoAmTfJXnbL8mobRuG4NZUq3JELRO45fIYGFSiuX
/NSr5ImVMsuEFUSEzZJzgZmPgAv8VnsZXezIl9tnDGasNUEPNhI9eL070TZsH25I
VYPxnK0lPceNJMM0MDLzsCwjpFFhkd3YtUYYrR9lt6nMXhD2jguZSj4ZC5dT57l3
diSYtQ9slfuXtbWkR88xaJjnlYjzk4261+KtnVba4mOv52vsrDirBre+E/kZ/KB9
Wc8DJwJWIEGmIPfMlcwk99CE7oCxNLgXsW+7SMgKgHZ7y8fC1sZUCJmnq91y4Q9m
/tOmczYby8NbA8IAHPKfbZHRpWzKKuni0UWD0MhZyuJC2YEH7qcZx6ElCjpxwCht
fqC4lV7ehCC4ow0AFgOZ6GtJQt/Gn6OhKnPW8cDMWGBW+vIQ5WpAiRdTehTKte+o
cZwk6AnRMt/IgesG8cXrVBU/Zg24msJfC32EVaC/Qb1xUXdUTOPVSHyZLEFk5xbR
7SvQ9swK2C7b9QqFNlj673p+54nKhQFmJYsti+C8+IbqI+vVnH6prY8+Uog8aJ+n
b5jw3dBGWjt9OrfbT7gUpqw+W8QYomAiaBjJDYZnKmVzIWagjh2FqmIYDgBMKcIG
YdZL/a7YxM6hXEm2aXIeB0/+OxChHoD5kqWnsi2kc5sneL4jSRTs4IhD2GOLtOYL
pEj9+6sbzL8mCTMO8LpDY0htfNQIVxr/iyYMDtgSbUe8iEAGCtHcQJxgTL4EtVZr
6yOrXY7qRot7IuEFEGUzcoq0KE4nkAUtacXlmT8t+aySnPNPxwdD5SiOq5kQL67/
92nW+l/T2ga605l+k4dhGDauP/fbX4KP2Go3iKtNVWyInukDkczixSZCAVF/mDfu
EemXcn/MfresTAQ0DfcM3GqXJhI6v/Cz1aawW1ffTSW+zjb3BOt0egSjJs/E7rDM
ED/bstTpM2wIRjLnpUrhNKnMxa5OLa4uOGBSfP8Rc+H9A0Mbs7rX/8atU9YirJvl
IMNAKQiMknsUeAN/uTYBYq8hCovVUWyHXzWdsvxiF15gMe+Y/wlkyEQYVl+lpXCq
uEZD1e9aUvolYSvITkxFE1Y2ZtyuxRb+5J/6riBx2j35x/ijF9hI7CWdrZwIAxMD
DTwa6UfhwcuzzFizrHfyIhvRSRRsNGH0jpz+bHTWeZG6D5SIbmJAIkFhf7shhlwH
X2S6YKkr8T9Y9+jdKu+1nWV5S6iKu/MHyLrZhHRIPwyzq37Nvd/2EMSeNPn435wP
ib/8hJWxQu8gs7HriSOJiIxIa1EVRcQaJAuH0rEUOW2TCCQxZCyVJ5DrnX4AgBUn
8WrI9fKWgo4pJ66ghsQkIGAVTQv19brfHHLYb9jW2qxKDysXetqeZW79hCCuSYyP
1N5wqO4UhXsxH+Qm2g5O7MEhklfOVrdpX1NPdZQ224cUA4Yf6xM8+DBRWRVnzNRi
vteN37JyaXzEHTQhPj8OW+QPuE1nDjARHMUCENJ23Gje4G4UXoWnKQuF7TDT4Uu8
/Xtcw9cPrYENEgJDkb7XUpBUiy/PmIUZJlxBgbCKzi1nBYPDONE/seT5nkpuIpTL
rfRmosr5OQI6qP/+i6YwRTGQmqN4LaOcagRxMh/mPtNNp6okbwzQCBNh4kx70hKJ
ZHWtKuWZ4vWRLh+EaFxm4ZBrrj1p6pxMhFZyQVgMROY7IOzzYAF1O+NdI+2c0JMg
gBov2C2/iBr8ASqelAGh56CGN1meazNdr7LD7bHzo4r07UDor4D0MEv+jJh+KwsX
g2xe1p/eJfz+YesqvLveiimB7LmPAosbb+QMR3Xx8ymHiv6wmEEwcD7cp9uT/hqI
UXQy25DecZSIX9sVTarOMrOT6CHr5OEWyd/mBC0p3Yg4tTokI2e7RjlbzCv3oPvo
H01+7fX9OrLYQDzoDrTAMuFcN1S0hWVeOV2NfOrj7CrPu5GksG887mNqVyfUDi2j
6+JGFFsOFwv6WnIJm0+UTTY8yrCGZ/Dx/URlviNVWOWDfGAMr2TCtooRBySBz4eA
gIDiZcn+Yp2CsbOAk6sz2xd7468uF7sLx2maGnZy/+BTSSYucs8mhyfNjI65XNXr
kZR1LII3acDqiirWuHxj6Yz6LgvAolRNeooXft1W/KFdXohcDFVVxuQOKukcVMSZ
8IcFxt9TO7LnKRkwvRTkMovP3tb0VDAF6qtqsvA7zE1oJNvDTp78QRxOUZ6Psf5K
C8rtyROrodoRgqmSpEwD1cBkk+x/fGH9RLwELaxf+cw1erKELwmY0/cUs5HG0mB8
nqg+ncTlzcpkpyXRRjcGxBFKirIj+KEdRcB1joJpqg9HO7gBvRWNAMbWwz55fuOT
Gv6b9PpbBi+7qk2qkBJ6J7i6NiGkBq0IiogqOTAP6Ck9hPnHN3Bpr1h7y6FgAvjk
FZar5YdnfIbTg5sQLOxujXbmVNwnaLcKisOa6gV7llq1CJDugPtkiCglFMa3I4sm
ts7wRhHqN3vwcWSrk1A6LLJXDKGGUsDucToZs+S4FJCfdP59R1avfNGdKTcU3WS6
MHR/FvIhCumD7PWhe+ETVmul5/U07PODOpQkclooGozc4mAYgpDHu1Cv6LGgke77
U0aDY/oRhCeVILXpBhj9oJ7LKPA8kV3N3zDKdLY2PWru4mrb15C/HDnmJpXPN6QH
1rnyjWDdzG9vKa3obPImjsoEi9n8KBxD7P36X7mWl9UROn1rjQGXo2rfn5rkeN84
sMJnceV/pgN5inbXJMq/PmJ0rkognKuXEoH+4caZEcg5ujYKEIAfnhOoIa8Bmqek
Fqgeu2ls6onLIQpXwt9ef2pZaFTyFEvXRLoVvTcq3Ta5jl2ut8UbXQ+k7NvzbqQ1
N2xPWdbayP1lRRTtpiRmwbXI/osSw+9ZbTSuLtJmokEASpsFBTTFYWbr4vqMXwxv
UsiqAdlHPsSnOlUVyds1Su25+fjbSmsV4AI2Ync9Z3N2heNUXi+1CYrLQSk1dRKp
S/6BOxRXvFi9D+GUx9q5RoNfSNE1anwhdeHf6yipCKjdgxk00VlAI/nc4zPPYOuZ
ODTxQ3ayjhS8+UkGXgmorGTpq/fNBswKupqXX0LS4oDlCD0h6NtRcv/LaKkP6UBr
OUgPRTOFua/Uz+Mx1UKr6YuGoYulFm3GjnqvCkrXRsV7Tkqr+MiL6pIdqzJXmHhd
Rw2H6ZySnQ/y/DkIWSQs2qiIJ4+GJcF97HtkVxKfLgaA42ss79wZV+kmhr5Sem/H
sDX5TTv+9r47Nke65f5W+JYfRRyCtYrC+Bw19A4VstpO2+MiDZag23+DQhZ6tgPf
0KpXGwK8CeIB8tlTPwXT9jWb+RsJimVUvP4crJGpjFLDKzPQGWSngGYmkRR97DHc
V++UMzRXqZuavj9fCDofDGswuZsZHzk9WyGiH00ZdJ1cvLhdUFIa5iTR7J+Ajs7t
GeuGUMFIh9UDuJ3LFGpQlARAEs6yuPpQKDJOnUfTE2eKEz8JwSVkPpvlWt3XXGyV
LmmDqIiu6/D9VN2nvEZa91CpNgw9LCGzhdROl5WnKWnZu14eMT5rrOYM/Y7XUqVH
u8RcRuf8jO3FGjZdFHw4yHYEudFGCQBr5AB7nheihcZRC7DWd+LMUl824yCdpYtW
B9nkWa7KS2wkL+HgOjdt80u8aIgY+J2t/8SpIG3apTKwD9RvynKvGcFa1mpUvb5Z
aZoD6WsaUCOvvLPOJq5rrLfVMdeivdLDIsZsckQF7+gq9hWZr1cXH/7X40pGN9AW
JTdG4ZRyGCMLYPudtU77iMvh6QeHTsZu8bs4ex5fPIq4dN0sRhlxneYPsw7zUGrs
j7VdY8XykCbekVZXC/Dh7I48sPXOjtxrjKP3h7/ibDgH+dfv5KkhInlict07SOau
Tbnb7RXqoO2yYuSrO4Hg6EHWNLjZkwRLSpBw6/pYXEEm0RnbuDFZ2GRWbVOTAp6H
akCxBNRtQplK/skGMXPrvjRoAGvvcK58woCuYeon6NMNhndOVnl1uzx/WSV494WU
7KRsL2KzxDKh6qS5Vz7PPdIMCRXnqwmZHAo+TLiab+MPpT8sebqcLcWe78lm4e/D
xHVRg7bYnnN8MEcf8vY5LOFFGwcJnE0MqdUKTV0AlJhum6X4mRqp6bCZw+bbXgfP
j4WrT7Sf54aWTIWKNhKellnkcn3sqbGzseUhXM3Bhn2lNYKncXORErbp9e5soBO9
uojGHBRxu63fhUp1kT2hvVh+w5cTDl11zugpY1RSs8nQab/LBOG7y75jqGuZrshc
sAuEJ1mvGDmL6CUluXEAsPjw4r5Dn/RBcQ4NdEZXhbEahJJOC8MypdIGU0yXpIuA
OQE6D7TjJ6GYsSEHpWcAVU1lGUROBB9pc6jNnbQRCZ+S+e27E4DK5DJVMEyARpMk
nofDkWUW4McZv9TjetmKQmHbOpcdTfrVAcX+CtrEjQ166K3wEJdjQbyW9SQ1PSzg
hGibsbW2XT7QYx1xyqBNQOBlALw9quSJREFvGOzM0JjCBjpR0vDNUJzdY56geHnE
WFf/0tYamxXO2qzRXO5tUOWmRPWDoA9liREE2EQM7UC0R+mS/PStWAat4jhnD/RZ
YvOYb3xbh7Ly3+Qj7bcgNV+Js+PBl2f4yTxW4fxAkh10aU5r6JmsLzTtYPGAt0QY
Pz/7W6FiAyT43FsIe2hP0nNIZmro+Hew88K4mvNNYdhvfJ5QvZiOV3sAVwPJHeUH
zh5lRt+4vD4Qtd2dHK14g/L/gVbwXnTseWHrRPx5GK52n2wi7bz19OEj6H+bbcpz
WmdojPhDZ4ThS5/114QHICHmhuFwYu1uhHmu8JwYMr790l7znqNyzoI4xFOqyrm6
/71bLKO7LaonASii3OK/CPZanwSRUi1fygBX2MdaD9aD1ROg67zd61U8tFC55AqT
h32hGhJAsGAMx4dB8oBaxbrkjylid80F04oOTd6jQGcrwJfmQMimQ/QK4qkDAM7z
twIQmro/54XEWcO0zZQqv4jKDovs8OVmIA9zefg3JlP93kKwwA1n/PjtIDNamFbM
p0NdEofMFHel6iy9+aaxTLMx450mARGB8zvyD6RbDaIuONbIQIioBRQ/mJ+c865e
vdAs+zqjyRvPrJe7Q7D97kqzsQsn15ZX/qmxTliiSQbqaCpdFDkvcf+nFVXUpQ2X
PKamRIkM9Sw9Qjw05OypMZOfEeVsO1u6k+EyM0R0+QrLOPagGTs/qeyX/gTPAX66
mNlvk0RoPjSxlr1jPsCufziEx1gMnJJ2r/NjwmI+TEIs3/LYOj82dggtHCdIx+Ku
l/OUpOVDQMzuGIFFW6jjeNUOtCh7vwehIIjUXC21kwjZFoLKeNtGRSR/lKXudr+j
hGlN24xPZS+EOQSmJ7L/61IhhjFv+GFBN44vdY0DK1prXl3iqeD6K4Zo4DaIDCev
Z28WcK3swBVumneMxQCrOyANC+ezb8JSyvjDNGZeT02Jd3TWsF1eGVW3oqPaLX5V
eX5edwos9aFTLAOpP36P8pUsMMoOAv3BKXqmSaDH0TKkBFfzwVeQ1Lt9kFZrcJQW
JfLIgiVDpxuzaZw11V2GZDzLVwmPWpJ630WinrTMefnhTj+bP/AzgxN0FTwtFol1
iKJ86VJ8dc3ugLCVoVLVvL0YAOKEvSI9//siZkhTs/WdoGFZY8dYDUVGH1MzdxCh
OqxhKVyK+FWEXLFCArn5eL5FHeOSzFYdNpi+AbyNFEH+RTbBVio1TYtrZWxbsMdG
k4FB81V1GNzi+87WGKNHMZsdCwPcAgvAjmuxHOLbaFFQxmyGnnvhP3eOy2e+T+s/
p3qM0Phhfax4QpxX+yr1j1D2p4EgEVBYdfVWTe2FRzSW1hdojhQE6wQjxoEeZx8G
cetFZQ5fwtHt0/0VOWVT8PBgUd0VTYVIaCzv2XTrC2z6XhAsPKGeKA8n9M6V8rZo
/frAN2WtAmurs1FgZeVP3AEuVHzGpaINDi9MLfTwyd3CQ65WNDGiL9a008Zs+F01
1DaqEmVpp39vgEsv6bRCSruJia6GvG2GoMKlYyxakyxYIldpbxjTx4s2W4MSUYPv
SfBgVMrSV3ZYeIY8lRGReFlseDKLcHvnLk4kiDHSerXnjE4J1LMj+RxwifNihENK
m4PqoM2eHrhgd+tOz+3UbImR8W/PgallBCdKGd0GB5ViNkhoZts3L/9iBTqMe8Fc
9pnCSb82ouGvwVhjiNOOX9J0undmQLAcYFm0d62YvJk0lMJ34N0i/h3DCBIrFHAq
qqNkkD6vnjM4RgA6frTQkdoF8mZ9PC00oYr3zdtXrmkvIWtbc555U3ATACDvdYsa
bamJ+ly2+rUylyR8ZyMJ7W+VfzRBoEyqWW0WUi6J51A2vfpK9DIb7MJfB0AitAJg
g6bOsgGOnhG8klYFnOcds3l0NEbCKxcTH66ZBzSMMn2pvlTeKtsvBV49AgPwB8Ny
cgUvYtsIzBybT2cAzQu3uhzfeY8/7tAY1JLL7ZvnWiLEADscz6w67Ic001y/glXD
SRYTYVpuWFmnrBI16PeM6FbTo5MTyga70gd6fsPBt5nFu08fDQIIhFuVwBhmsH6t
PCFN0s4FTyILZxZ3a/Llp34uAtC8Tnc9V97are9EsblNnkDaRMhuMAKWTUs7CvOf
5Iceyn+BPyiM3c+GO5jYUeTZNQahl/dkPC8hk7RRx/cnA/B7890kf66ugGMe4Cpc
g24dcZ7L6XDuEyCUoWB4eYaAucUM6iAwwdaM41LnVQGKE1NliLgdtWCca7astKdL
C6j3hP+ZerkEaQNKkCKhUzVdnvt9RGQ//l3+CKz/8sTVW6NvUoXCbOhcpM5rD64L
sGF97vJJCcqGmAqZdRBpltBdVnDG3h4xvNhvZv+y8Sv2ERxG/25x4dkAiDgRhxJP
jBWKd0rT/BwV9mPEslnxILMIm1i0xDxsAMYiYSEuRn0aWrL3J/5EQheGU8zSVDiX
0gZXgnYiSk5oMF/69dFX7sHdzbMlO1HZtW4Se1C7Tgfxrd37a+L4V7sd7Uor3TAB
Y5AR3aMRBRDlx/1I2Vkw4+mgusgADNGBl38WPp39eBBmgysqAltUlh0agFLNO5RO
ZdPgEcIucgUDT1UE0XiH1B2W0G9UaDYHxVGwFp0wyYOamuJCr7YLgl0QxfPdIR0f
DIolL5TpqQnqmijF3GOSCXrv3iLIOGbu962PIlNhrsu4A19SD5NH64kw0tG2E3hM
uiisDK5s5WL0QKGqQZecr8cNVEh/rKbHmwdF+jcA1h+ef/Qj5Ts6LPj4bFnlEA8V
gNswXz2zsWikm8vVr3Zfso0HsrzHQYP229r75aeYf+uuziKQs8v1KFoJaBzXsXZu
x0V4s3c2pdIx4N3sLLKYQQzvTuf4/gNDECGasMoJSmhTSi3+ql4jM8BXPPhjlotN
qt/e/ayaQOwBDiFahHQRp3DxSjceBcnLkpafWeUYx0Dn5iPFdd+ZwrHV7x2gawOx
/LhdRFNkFqarWaRhmyBtSK6AtK0ddkUI0Urqsn2cmJcTObjC8vB7E4occ0PZR2yz
/NMYflgY69qmgnFgHXmhcXjar7GoSM2g3uNjerxXO7rUpjuFylo0C/m8f9gnatXD
RoMfASLMVlucDWNLnl0pVb5t5njr1gY5YxEu+RjhCtaYY/1pvyoEFYNfcFH9Z24e
jaQNrezVRvRY03V4Dyseqr+7tkj0fMUdQHBy9VkQjMe5R0CFAG3giTdVuEfVDD/z
DA92qUt34PQ54hSY+iwKrAoQTzcUwNB/aBK4fsT2pnIGzrwXMJ49u7NyI8voGYBK
e+KTOl9xx5d6SLjpLtvziwiuPAFXhKDL02GHoBPyjujrTu5zI/xi0xQX0gTZUBJj
kjD6NT2Dz6rABF41OLHL2DmhkoaOHjLk1W+Lnn6VcSqeOm7UKPIsr8WFFLEJM3bq
iKfsJw4r96Ndn55Z4ld1HEdvOqk09puIm+wuTkxLD6xTz+ElL8js6FOZjo/5WaYe
ZZ+a8dbXrru1etZKrQRLN2DM0Vg7aGm2iPBpZzRCLw9NBF1Uqn94uxkP7PGhl5nu
UIG1VrwYAxiKhxugwvFAsOs+XtStpKHKWBCapsq2YyrAV2FcHIh/AY2nIxpkVJHT
lVEbuu8FoOvC20WUobS0rgUmQXhxJu0+l3dG9/aaM5Z40uYJVNdfQ5i89DRDqXbf
KA97F9zZWLb7qwvwdNg4aluzuURN/rXYXNpkHFditPyWHughT8cHb1rUX75WdiLn
XXdFvXvwCp48wrpjKViNlU8TPtgwFQ5xJAMtul+378aulOG7OKpka2vsi0UFlYa/
AX7eIj6hu1ktsNAhMXhjanjuFIAXVyQGLhL3YKdXpXxPcMWZdur7qVbZl0xbei6F
PMOzHXnxMYXcJ7VCOKZ45KDWvwuGAj8iyA+7E/lYpCcN16l+UAFuVna6VFPkU3qo
6Jhil1b5n9o3Dy8xw8OUb3VmDhLk2rQk8dn3iLS0xojlpqNRHZKeXXTFenmc3IhM
ulPSB8f0f5pSKGNuI3hMwZMQ0Ta6TFHihqinDJxqcG0afsNgpavaXmCkbyppNd7o
xsSv7OaMgmdl2NS0RCUdU5OiKX9lu5ZSgziaA3jfQAwkk+CX6WS+lsnfDC6mg2Zn
nok7kjovsZKgxC3x4VpkUPohSHJ8VpWM9T1Kh6rvd3Ch8ox17AoDB6eKoAWI/EDb
PEum2+ByX8LVoaEXBP+HIkqxvWESHzbwE4P7Pd5trxJN+Zt3cMYQyxBsxVpdZuj1
VChGrY2pEpQ87dgpmVcx4+6tglUZZhx5UVd/FZp0+x7Wmu+PV0EPXzjmrm6yxSKO
7+8i2PIHz/Oq5sP5tDBySEzpht0YvEkNf4jBAjiiPOPUiCKMaAinnWrIafUVK4U6
+6h0MWhsKJEG+TeB3XM4/x0wc7R/ZXsiuuYmsNPR3SK4xla9oGLW1k8IrLeUsszC
sgHDD/Kf9FlxvdoyRW/q8nc87thdo88U1+z22KPMfCoamKbIrPm87HR769m/YYYo
qu05hcEXlOqxxXF3MEeSGzQjz/0n7lUJi+HIA6mYRZS/SyERvBSXQZlQf/K1QTnr
Wvui863xXVIqcVIXnd1r9nySoT0pBh1sRZC13tX8G7/to69JrwBRi82QwR/wqWf3
sexlctS49HYY6Nwtl7zeItLBxwmQIzU4y4Kk22PqDQvdpE3MGTm71UBbbeOlPOz9
VBoIkYR2QUhKh8frWBJ9DuSIayxClRQH9W2zX/pMHjGDSmd8hip5iV7lTUFlBs38
yv2grazRkYWgayUGCyOYUqKRZUDNQQILZbYovfvx+qybYNtz7Hr8qrWOxLHhncgs
krNYCp/09uxBg4w+ygY84HaQqBzPMygWEQGNUj2LPGgHQzVM1iKEFLTzByTz+w4J
4s22TnLLS9BMJhKiAuFNPPd2DKgIoAjEMXszeovSsmHVntFbE0e6o2Gwtiyr6NEP
7b8wPqwRyXbofg4D2WDUqaAfnsR2iVh3sy21+vlLDGnfFqimulqKGtoquhOienPG
SHJPEeajFeDGqbodRx4ucSe9xD7PflnMvlw3oYk/sMCh0Za2ycgjITZ9X8A9vgD4
9Bqgud29qPZggvYJas1NDYz6dm1zE++Zy9s0Sb6v/MqF4nK/b5ugyiQ2FZupMq0S
RNdFY9bIxXcxKwfe1Ci/1LrGfoZyM64YQ0JiIYI6acG1Memr6f3jpyipEhnQx92Y
W0/O88ZiEP0jOJ5pDr/FEVqT5xjtkwLEwfdWKDgR70SOvZlnzPktjFGITrwggU4p
hvYnKf2s97uh5sJahsmngvjHx8P3sP+TeRFdlCQMur+Gd5S7Y2ePO1xm6ZqJG5tF
+Q187TNuEvvGWtwgBj5H/gE5Nsz71nah/QdHFXIQXpk+9hWmlwbUAtIQnJEclRJ7
vqyRY/Dz45EPmgkdGgxY79qU0kpHFXwldi0tH+FAaHSBxeFJ5A+cvPTDm2nx7IAm
pM8hCLsgpD5cEt9TAAWO75dvYtPAe9pfxfAbuCS5EAFUaq3eGmdbkHrFdJxS00zE
MyRXH2rosq/vP3TiPlxcz5YnHtgg2yD9Tillen+IB3pFhX1MFUh4m1gSKTDne6zR
oWnr+t6ElXZAMnQSdDM4h1jEPXkrMm5LgjSg6lcqTNZhzug9EBJNYZhOqxoEpVEJ
milAJGVvYyPEVfWb8aqa8LfkorA2vETVIKoRhmi7Q8uw6qmVlifqZXTKY1VNfcGg
CB8vssHiNPb8STqMBocuBuMMDWvq7fji5qey8yRUNfuo79dV2cpbJ92MJ482xeDF
TovWFAMPEjllGKBBjLA4IbOJ8n2FXmxMwdDUl94P3WYSMvEKjGgo/zndxEe1ILpw
rELx5sx+k83h3kfQQjVzWzQ+0zmTR0O0oTcrPbUpST1fmSRWNh2YxMVG78MUj8g5
Ouo9nU7zP6n9TPIpkGJD5jPUe4726+j6aTyMqI3mfS4zi1Apsb3Izut8PLXpkuVg
Askf9B+JmqXf3/CHzy4F3rXNoVeE5eZ7S4YCoICsJv4rSfsdOBjWSCJ9QaVMPX26
CfzdKvC0eFSx+DheFlcGnmXQyelrx6xW7v96WZaxoCkd5Vp0XRuEH1JK3xnDF+5+
aLT7QICKWSeiSj2dWq/7BHgUPQmiV6iVIzGiNriw6KKH9dRvR76DBsFy0rMo/DnI
HsHy9B7pNZPH9oefWCQVwgJMs1NN7flpUAtJ6cmI1ibhR2EkJWTAN1XhveNh3xi0
IFvnsWT0LLAMV+5gfqHRTHM9DORjCopXtV1m1+gbNDgcYrWmnO5C0VxjBdyp1uA0
9Jlq+5GUm5Y781uJ19Az1R96HKWnNF1+BAm4ryAyU3H9tHv9C5b7ffFA62v1gN/W
Y7IWu5oxVevR84cchIIMGkWpQK2gUMfj5xVLXPMNd/7ap79IO4j6+PbPpnzCvnOx
usiLtNKOzNS9i+CPYu+n7M54Bk0BRnEjMT5eFvqql4YR47MzlBft5gB/N7zl+YYV
I28arAZmisoKJ/TqmuOjRIIryH28YBNn+TlS2OX4h+HRDSAZzkg7auWb/FNS1QRW
bmumcEIc57jMd86TTIkRiCEuYwoooe7DS3723jFGx2PutY1mMVTomqVuIuZ8t/DQ
QqgJysBFOnWNPJDHO2xL2537xFvAHhAjxSyyJ+98bGs0/c5V9LLmlsmPHHjl3Bat
Mx9NayAfUGZ5OMjdHaSzrOx4P3ADTBiVbXRrgbF8/mNUZr5UxG3Aq0ZZF1Ziv2T3
fvuj8EG9sWaruy42aXzLveer4tmzF5onBwFPOMGg+8SHFmzLFW6Z73ezDSZ5IE8w
yK9rEnEPt5aesVFONhCNDz7eQEowsl4VDifVFOH1gdd6mnGvgG9R9BCRRNU7Nl3C
9uqprLCRQiA+ahRMZgwxOLlfs3db8nmg/315fNMp9viRmeNAEmvMrlZ5hBTyRBfc
tOufYFNazoot395XC7Yh3pkChXkZAwr8GejVoiwT71/iV3x7OMtIU1pEyZXGs3me
h0cdygmVEgXt135ReKwXiqFYSikgR36zblkQiJ4bwHZBtojY2ShpQBLALe84zhcH
jjPkGxKmRvGan7Mhz9fB7JNLsXhD0GUerkg8nkksF4RMuonhfhplMccy6GqzyyAy
eJ1/z+Hju9QKXO8EkGajyTc9cZgQJA8jZ9eSJEROz8k4+8V4nhizf3G3ccCQKWCe
sl5iZU1HhyBOshI2z8RLP+pb80WGgn/bgmaK+tbnMBVd1gP3Gxpb4pzSdqB74n3r
36YlatAnMdkWeoF80JBGrbzHWg1aXN3l19ROb/qs0oHi8tAjdCBozgAt0aT/9vUk
daxMVMqiMD52dqM9NJHOBcOXhjtvCkYYeDA7qIkqFwDaUGfQI7FA8eGjIM2UhA8G
eJcq3mBQm+yB17jFT3sA/bouF6xXMo0vf4bIA+p5CChBSHVJQeWMzXeToaApu0Ua
QPdhjmUiCJ4e/Z/Ee1XlFYqRut4U3F449BMYBn6q4uUav6bWnm/YMPRYz5Bq6gNA
DtQIB1VxrZK8ASbpXcqjS9LcM3oySUFBCYefrdHbplsuQRycnvuA3pmgAbtUNfe3
snJPclkTapDTGoVceJUh3t7as9nvGjVqIoL1wae0C2ox1vopFZlAbddTz5sVDSp5
ffDj+pBpfUYe1N7SPu7wfpzGCKf7hRG5ltz+JxVjDJma+GoeylV3Gs329Yye4Nu5
MGSZ1cChbN8pthyUN/Cnq0S73+DOmm13ieFCQwZRONVbEyA+PQ8n14QLmAp2jD47
u7/dEhFH/hG/JfVjIbV5ZzHz0HLaDmLQGbUVfCzvTYupO1eMSigSUGFuOGzYQbvw
FSyvzFmMfHQ4VBSnn1FWE0o+3VcqY6JZO+yCvKFpJkQ0ROkhZDvGR+rNTd+Icbwe
KQEAlGsZCheyPnyiCY5OZumIKxBLaE//Dq5eFMjJp4808/1KVeQOhnLGAM3kLdzM
pxOx3yQOWbSGsHL45k1Gu7dxdtIin1diSz1C1Bn7L4Z5zDX0grcKec06iKzPU0cD
wS7U506ysiOnN8o4J+YKpuZ9Ngv9rGEqvtm0WhPPpBe6rzwOXYZJyBePSpSvwzZ1
NxSX6s8dYLoN33jXh41+R7p7hDVtXr00Nh+uVB9PwY3PnLlMkGx9O5x+FfRkiRoz
5mGIqPGHdRVb+Ql6GhLfY2qrVK6wCtNH812YWafaTld719MzQe9kIshQx5LaO8Lu
ZhKVrdGTlKM+hr619DKU0ZOft8n4kcBaZzJ3LVja7SyU5SfaASCbT2/hV3m/mB2Z
FuFqWsXpZ5CmJ/iB4fnr6MKyLbfFCyx5jATalBGyJHj3xnMkAzH0eSEq4ZjRZxd9
xYLsciGDgSFKy96xxQUf5kHSC2UyzKSUuk9fflNiLbKY5mT3NFSfuaoYxRL9V0Gn
nf3pXLhXdGWxjc4N/TxEmyBi+0TO/QTsYmHcMCfnyIqmJR+kTrHq0sN3fCpvaDdv
wk7StJ3qGPqUbvR5y7Eg6kctAGd0RDmRePSIkv5sh0WyJx3MPHmKnD/AdK6B5EdO
aAuqsnvimk0cAngvxohFgvKdYktmwmhFZMMVTPyZWyYL3CYSjLuVeknptoLOH72R
etLz15mzDDOHRJZmxw9hj/nkk5AoKA1fAkzdeMqLzQMUN5LziKsjiKVmvuK5SRFA
xM+H+1njY/Ps4cuXM+z6IeKctaGhpWvngMJRM8pKj4G3uATeTpNOlsjLhxYhbcHw
ShSrOYrrl2q9E6nf5a1b5fQYAE4upg6640JaPNj7uRJaLHAMA6OY5jpsB5fBJ3KI
iRMneGoCWbp9qm3DXmkCBNKYui7E19AwRS03xCpwcCsC9bwtpejrRdrqWLzNaeJ0
MmMzlUZ5WRWJE3dSCwo49cm/CLwBQcHPz6OWtps7QWx+/S80kaKfhKDcpKpYZykC
vxtmko0827vSGemcz4oP3NcRWYP740Nhv2j1qhSkvoph/+6Qf8aoA7P9AuTxXmFx
Bq+yYUjAs1qPO3LaQx30lalOVyEHAUBI/iGpjDDkqPtX/cXqptIzk1VQnIfTGG/I
KCuzVo10lAnx4CKIpoEjhxSj0ibA1Sf0ppCedJa5xh+ro8fCZXExX+rrNWUVYUWo
UgACtePUF1yhmzP/V9ecAu/G671ZdKUXx0bICirYKOH6sF134ih5CijhvVO2oJVb
h4qZJ4dQ5ZLOyqykAv3VILySLgJa6/VfYeSSCxLcQLMK+MorEgn65ls/ph8YNDSo
0mzmKkOOma7aJe0AmvYpVxs4Xbp87pCmorqtEibg2pP1TEW5HBAaDgO66Whb0GHf
Psc6Gs9r8M7yc5GTx0uSrEqWUmaYaStEEEqCkCmW0GNwVbW0S9NppMGzWqynkVNj
4zFZLv2FEzk63KAw5J6suDigd/zoUdJyPmKCFg1MYedndX76RYKVHqY2kd+neDBx
BDXSfNIbaEVoFZfs8fKY/8WHbtvHIt9ZIGLSaFKHU2jKkkC19wGyp+b772il2za3
EdUu87/60Q07Bv0U2tqFMHpEnE8Ynvm4p9AS716DRQnOTtG0iF+Nipsrk4bFN9II
6DDwBh7Nin6oANQhyfB75VuIQoi9QYrsF42MSxFlZYvU+z/meaiN0+Z25PpR/1cv
oR1vABxZGJJOLYLRnSP7SpOcz68F0d4KzC9fVwz7qIEDr+VlVpvhiJSWckwabqu7
MziV2gZTW+abQeWJgofLB2f+oeAbTW9elYr1UZIrTmM3KgeJtW1m33XA/DnJ7ZNZ
V+sdQTJsSqyrDWDcu3pbg/6yeEYdQc0KAuXoZ7OILF1rC+UELHpx1FEKGGiIpxW8
dNpzLYy838CuFJoNtsJidHJIzZ0cZA9qZ7njK70TisD2bgX8kyK3iHZYtEp73dNI
kUkg/I7mpkgrAI4NC26FyMF7C2ZBJt2nt3A2mQ1T0xJy3gnL9QXMHw8IPkmuewxb
sJ/frBJfOFm19CLHTQRCC+hLnVsEScUn/NhwLEqQqOk+j7R8L0GYkn8NMTjDSOZI
Io7E4m9T83GMX5RCzn1JqELsuRvG+aOPvlcV6By5KrRkwaPRqPn4eOVrQXqJ3Bkk
RwWdv/T6EC2fUCWgsRcVlUgoE+U9f7FaHIu69RHCh4Q9yTbLe0g9Ko7fa44vJiTm
qHgYgKkg6ymYY7lB2YnP6oHugOXpKFLS9oB6me++Eob/IhkKsidFBMqthtkBb0Ds
1aMr8BYYBJsZVWhOuiYQdCzKVgjrpjC7ojM4MirM5fn253+y8Jc+iwMf2CX5dg3r
wRb8gE6EBtEqK/7zLpTunAzOujtdVhg7EZ6cLD6dcZhuiEfS7SH1uMTd5xnsUjoi
RlHySrw8XuG7xgjWxuC9TwK53CCSZ4EFHQku1Xf/UQCTp378CQgWQ3POeqnhoaeA
rot1kiDlzH9GBbCUKv504E8drn5y1t27gG/0tOdFSi3xuYIUhyDd2fhGyhpHWX+b
U7LitRB1OiloRN+Nb+f/9g6OWzKC8gSG0XmFyD+SmkKjtpAQztdp4vNrRArTpLWX
ZQWpbYJmCknnpMvWCoDm1d4JhRYhAWTauzXpkbLl6XIpmNR8iRIQ4tM7fIVTPRkj
lj6RPDCLWoIt+im5iLadP0aUJoBYOJwjNTjV8NMf4wYYLC4KPoEvMEKUViJUzgZs
Pg1b0PaXBVSHEPSxdCZNIuD3uqLVe/UVKvxmgj2TPISx2XZmLUJZj/e5IJTBMGLj
xUGVfc8/bM/CQjPXNnUOr4ZYFpyp2mLYjR5OqUJ7efD/x9bhfZINtTqakj9xCaAT
FV/Xo1PMJGI1WJXkN9FRyCTwGkNnXdNUKG/mapZthNz4QbW3f8RiLXfHRDEwF9mB
TxYgvrwusIroDwrb+e2hgl9YHuyl5gUT15280cvexzezvykDMxRMAYipexLoKQZ/
UKUqlNURPlqfJs6uksX8yvmpFGltsXHWJYCOZIliWYyu/xh+R0qmaKX6NEQjMGth
O1ZYY/ac0nrs3XjsKBarvga0frCNBjq6mw4KcGkJJmxMKDI+DWi+a52fZTRFCj4D
RQWNFpnboUjhiPCW5JQ9XkBe6QA5VwU8DXTfbkTsCF8Xa8fgni3m9gNMtFvuey0r
/YjejuavpJ1tSqGRnIovPgZ6qd7phJ3HL2xOqJhELFSymmo8VOwz9toKRxZEEGzC
UKFAUidrwiP4HnRSxUSODLMlcVZ8zn2B6KHcm3vth2tAsiJwqRIWkQI5x768Wndr
J3mqazj3Tdh4w8Svfr/TVuh1aoGiRYUlj+zauoR7KG0sR7ASXExULNWUYqsqdixf
cHqFwoOCc8vElW0ygusd4hTAy0Q1Gp7+nzQQK7f5LrYJU0pfGs0/Nt31uIGdRyak
Vo2vrS2UWyI7DCxQwXmPTbzXYYx9iIHZMQ418J1YHN3BGjo5J4Nbt9gC8sq+3F8W
n9quRe4SHZeP3wcBlmN2RJ/kZfqphZn79+H09GmoIIqyzbfEf5+Gfo+8S0J2Lj0g
InAhvdkw8zHZr9cMLH/27z32yn9vXQDqHIt1rUIaca1YdA55fygVaYwfqr83CiEM
kj3GwpKsT03Dq2sQhT6ezaK96FKrcblLUz+LzyFvw98QXLEjPC7ms8YwSEfud4yk
1xag8FStC8lJx3y7pDlFDonQWYh7sHSgvFrbikZsJ2hCuAG6yg3dWG7UIwFb34+y
Rq19LwHd9O888cfmXzIu4S9LIBJ4ZrWIxhxN/ga5Df/iZTRj7EWhu3NuArvhLhKD
VrfBywCH3JW5O/Q4eMgxODnnNtnn81ga2tG1KFx8MGSsMNUCgcN/NcrtqcZxn20o
VrQX08rl8umgLakQw4JKHRWwaRa14gP+pJn6GxJRDjq5yJ3ROnjwrIKtlOrwlplj
MWklYjNKw62siSjibxlVKzeVM1nyjVXYocL9/kSSn5FAG5EjQ8Ppkl3JTvjonesP
OCmc5zDCajhoCQn11+LTkINFsEsMPTfxIX4i06mkWoF4BzDsUT61llE/w2aE18H9
vVHcI0O2zdbySI9WYOUZBjaCoa49or1tm3i69coIWcjJolvVYAaaE8ak3D2n/UbA
ZeZRSNPH/S3GARgP2S/CxR3doy/WzS9Jm5UFf/oj4zzWQd1FqwE3Xar8mmX5+4Oc
ego3mvAQhExTBkkxJxuKh4ZIJ8XEsHhZM+ekSv3GwBQ7KTk1RScqyPPh67uAux+R
y8kO9uPhwcxsuTw511kyQAVB5SElhd++jc3HJtUmGGYqUTulS9/1VVe1EZ1+70R9
d2PaULkrGQ1oJG4anJ0XsW1E3eR07eSJiZCNG/gfoQ4FUrrE0wbWFoLblkoT00Mw
VxpqMZvpSk52DWPTQEQW6OnE7CNAz6F5DBaka8fY/cv6xNNz6HkovYojAS7GzAer
phylsGLHMOdTZObEHDFg08qnA0/pprF4mdU0j42TQJkoskePSrLhxCiHIFV/vFkD
11rjHI5FDjmMHEFxXJ80OJg5FdeBjYJTVXrt2NAYjCAx3hY39LT1mHrcjpxg2lAC
ntOBGlnNGWx+Hg0ZJ1nnFM9Bd7y2OKUDNaOK2UAavwJOn2p1QMMBQp+LIyXBqDJY
b1NWH8+11r0QCY0H/1j1UE1fr61Sa0Bo3e5dl+cXKd8bg2tSrcN9kDiQiiQ6/14u
tKxLuP65k5bxslkFkohi4kNFu3kCsU5F3bxZYDV7rcc7tZPfj9cEXJ3vtq4PjnoY
gd25db1gXZSVwN3GLF/qv8YIVNpwv+O4qCurxZ8c22WrHFNn0Pv71p5W4zRKKSMV
glqk4Aib3qGC4Xq7mbFhE4HjvFCfZYryIyPnAqcaVczG5HtiCe28PAP5He3sX+BO
Knv9MEvCo44qdAv2TJ3SJh6di2u+M+whQaT3ST2BMIsH/XNwtj49I9JPSsxae/8u
p6MQapFiqyG69jfVeQepQYm/ADdmSd3It7/ZvVmS/Rq4Xgy/NJav3vvKjPq4E6Dt
AGH/XM0rLcIDjj7CbWVpUgbjiEgbSbolrY6cx27vhlkWcxusNnrnNh6E7pPbBqy/
fesVg9VLwWAtEUPPeE4GNlZXXN21G5xsmuzJwcs5yFRBQqAJT6nhziLZf/jNvro3
a/CsicIC3GKbWSM6FjhPzuXZkR64TFAuC6DP2HqMK1a29rJ0KfkZSS31QhroUTn4
L8Dp0uRgDdgYziuT5P/TxwoPmW+YiRi/zVtQrURPiXCmaB4U58SaLfbdUWhAh0L6
JC0NXnSux1sBsQ30a9pkk+zgpxa8al0Rw2WqsDO4AW+hUDXAimfyKmkgsnlYCDw8
seqAxnFNW0/qJDKFtJXm2XmF0Y02O7S55OcdK1nAv5x1+l7OdHCzH+0nElOoYHPM
kNVj2xPqHbzE82BvgsFJupvQrlWINlFC4LzhtdqCVe2Snmp4b5QTncd4w661w8fA
aThrhQ14Ogdvi4um/rfIHzderUk8ocmOaGlUqqtyxEg6PMSykb0CayhANjlA1zeG
bkfqq8ChSXpB6bdao4gdnl0YqMMy2Krz1s/93r0N2KfA3RTNsOt/+ke4FNZIx1eq
OPOKKjYjiM7SCv62SLAK7HoXtNkT6riX/gaiP+W94dBYectDwnXsgilp65Fu5Fy9
OwsRAlilQj4zssGTutD9pJKAzo8B+o4eHVnRmS/HUIAkUHJtmvbG8S8pSbltP+pk
Y+2UmrECjwe+VYxJbXDT7To0kDwgCQNxMT4YqF/vW3Nz5cmZBU6AtOClJpOM5/el
sTAdB71xZPjpai+1U60SxG1Xf7DEp4r6NTHdh49TFO1F3HYdjvK9MoMo3oH+exa2
5bVmjTBeBzXdrPBd2fHr/lxS02jYL4Z4gpkYEYPleNUVfj9OxQyhc47A3pa/Sso5
EBhmjevvOlDLwu5arYXQXqPQSo+U0dHvGJRuwbeWTEYjXVovJrDVfCpd7wSVzeRS
88i3bnhaJYMY583vFiB8JFVG2gj6GbnMtr8qwImwJ4HCpRZkBagk/UfazWeQxPC8
U5zZ0S/CmMG+vK+70HZtzkUYrYcZVWcJp5jJ3SnR/V7UqIynupbf48MK7W0O+jQW
J6mdhZL/yYEUkSMJFNfAddiuq3/+wSFtCmxEQN2rQg9TfqJqRnA1aG+Il13Yf0l/
01rpmZrrd/dAlmj3g0OJSWIFV3m980HY+SlR6oC67GFiba4spokjoromfEiN+klt
M7oWth91a2NUW05dm7z7nWyWFGHvF+cGAQqS1kb9voULIlKnSR2nV2Gkcf5wnu5N
1nxUhOAGfAxVdrauAnI/Ykp/qXNwaAcpTzBs7QVDIJGPfGP/LpvLVzEeP2lev0y6
kRYnQLpdsA9K37aSClgZr79VvAMK5L0UMNZDW/L819sW/jYpTa8PPZKIQMid1pWq
iqtVm8Yp7H5ePoGbU5h7rTVYnBEdZhcOGzGO8QX7+XUgJMmT8U3UCnDX163UC7CC
ihMyFCtTzyFBQ1Ejd2dHWo4kfX/mi229N/XCdPDxrBzhJeY+XrA3shxDpr25I7W8
FYfCjKL5VVcAn0qZBU9zTx4NXF+zWe79FTvdJyOfU2CkL0rHlZ+WT1XH+wyz56yu
MSUj4UqNntwvbm7UjrSe0OnF5EXg7CArKIqMEaWmKYxyD3GfPlchMaZuAmw6ylmh
s5o8JLrb2oodl8XIGJVgZxFSDiNijkfiuJ5oyJqjv7M+2DL0GqAtiSQ2LF8CY4Oi
MMD2eHVxxspUBdPvKAYA1kKWlxtaDAkzdjt+087iYq/SF5WxOGrgVkZwIXk5SSLc
rW7zNpX8sIyFr7koqUiU6NbBPtYZgjmcA+e5aZYgS/2mDAR4x3tw53gwx1IKkN6V
JgZ8cQ44LIi5WvH5/oVHwAZj6VwVQD6StafoHB6PYxP5Pnu94V76XRMoE4hAtPV6
GpXO+e4MeE5mEV8mLswutQsobxPyyAmPuRXhenjLYbQlMdxSh52/kdED62C7EeMO
23r0s90BK4r+KOHhPh2Pt37mSmi494yhnKQmGloql8Rm8krFs+7bQNRs4Hu2RFjU
IBqWYeQaFUiiNjfJ5by3kQsybHwGgFKEQcFxgRZO87qBtyHsGCPaCX2Uf8pcpwMy
SchYYkllEXTpfh7Nn+46c1mIBencgnjlGv46HdFscgfK/RxFZg3XnZsEiL7vbzTq
O4qWLb9Z75Vp6g4vVqU3xssEqMA1h+bNsXplsPkPOEIWPf1TnLI0GHdICfcb9lbV
Z8h3ymtezNwRLChoHoV//hHdGHQ6PNOvM03EXixBggvuo5HXmlI4E8qT5D746dES
ul7bBAZa6CWGbn5+3seqYvctw/U/M6Z7cb5XooO8FpsPa37yCMMWhc+GzUBDB0KF
iY170Ik/ysrDVg98qXkPWZn36sH/o8g2wB6hhU7pp8ecWS8u9+B3c41MDdCqcmeQ
Re9Nx899q0lD07iCMFTOBEMgeslRQniwibzgMVXO8k1/JNwuUVIuqLS8yB7NyfkJ
rnh2k5SeO2Hb73NNWbTdOOS74Yhvv91f3SrdaiVUqdmE40CJDHWaGzodaoqp7Z0W
gqdx9T4XpIMA003e7/KMAxc2yfElhHgqiIO/8tkQFLd5LF5fk1+zSR+ddR3er5Tm
d7CFn8hegy+uDbKdD3hHv8xDnUPgNXf8ei5VSv7Rq7gNqhwBq43ww2i6YnWTn0Jh
d+XAlk7XIUy9IvHoTwmdTriAQOEDmemdWSHM3/9PGQLOAf3ls9RWszBwec1jZMUA
UkESf/Jp/7Wf5NdqnGOq9ePptZRLEGdc7gDQq5AMYi7D4B7/7Dw+k+Ij6Q89fQhf
G2MWEiY2/XOGTBdg8Nvn9SrVHSlL3RUZ9KjII7lhWGsx0RSrwJlLdOV8uGuVqIje
FKj5Cf0dF/YX9hXCXxQ7BC0WbEcePoQj0r6Mtf6IqLRTMxuhs/1t/0nhu2u1ut+q
eW7yZGFTq1LKbOQZqs/pboKcPWDb/4WknC/IuPg3z9ZHLuuxHOLlfVqEnDKUwe6M
AFWmJMgBUAQWkUx7IkKq4wHyVa1AxK0JPTN7Riyr1SrBnMNmbaghZCetUWfX8wGx
Kgcckzff8JF4Eeya/Xfc5Ukrtlvcozs2dCZbhIHesIZqsu1U5Hzil5Za5tTmasP0
xAi6KtUmj49Ar7nV9p6jbMUFc7ha3neSuXOZwRnBzUCloPkjb6mg0sH7Hl0NUclX
sTYfTaCSOtrQEx+NQAMa8FXXLaJJySlEzs10kwK6NQQQzBEc9ZisfkmJUsnWo8Kz
mXhZCkk4tT1+kMUjaKoDC7Moe2eyq6NKhu52jmpxwKJo5D+8gtAAs42rAkG8OWH+
f0JsHC4rRCiDfgKjtcBeNufacPo3YWo6GPqh7rLnNCBx/G39wWCO1W+CcbbZelYa
rDnX9dGbUZa5r7IvoWC8MfVLHmdfVAvatvOSvRxxcN7Lf3jHc+qSjcuYDDv69vGQ
2HeWaoBjr+jyCbyB/HMm3zgW/axcNpdNOVqBZgtOXk+0Rc8ww9eSTWGTutbjye/x
yVN2eu79wWiLTrS/SoyH2gAKu5LIXcMPFpde0OI0BgD8n4risaEDb5QSqZ+TAF0m
qwlK0FhlDK1Sw02df1VZhvgAgeLFYUEBIOJd6vbjJiH+fS8rV3LfRXuHz8VWHLyf
Q1+suu9IyKwUSfOn4YQ23xfKwEZKTgbETJwuI7NB5wuf2J97PXu4GxEeKyj2LJRZ
H3mhcWF2slOmOFUyVMzwbjB7SyyLPHe+w5/QCr5QcmQm2FBhGxn6cqm3mzhBjDO7
qkMJ92V4GdA2nThuI8aDaoqxatuFzuzUmEfg5IHId53LquMQMWM2WZAZ2iBPeZ45
ClPoycoALUfOFB9ebxFbNYqV/eX5m0nI5fgf4MnYdoaUtZ3N+iPgaCIDlXJsO0k4
FFU1lrGu4yuycDra1V3WcBsxK2muzzMXnpoycTV23Isv9qCZPCaia2rUpsl8vjyr
pyo2oYpGo/gjvSXMhJphdC+nnMQ3ANk4YhIGtaW6zWytbmI0hXiMPw544TYQCDXq
YJ0aty6ka96kdM5iwW1/4E7upsALUQlYBJbD6e1DIHxqDiAOFOu+Y/lKvj/pAFiz
B77NdZEgYiu6SwqfHSx+XUmM7RyVQxeKnyDx72on1OhaXkpTUbix6HcwO4WiRTSV
xU7lKmuBYNwN+7KOFXz3B/eonEQyilnAtvJ7U1RyZUIll8+U+iFexsoKzajLBB50
7BFgCnT+1CwBNajEFIH/IU4bal0DbrlOeodQRAEtO7jej78lo+wYs4w1UZoQ4vT8
YloobTKtjwzY18dwRTN7weSUbqvoQFgudqo9KAQ1/S+YlH5YRTg+y9vR4oRsOM6B
HPPeYzPqRrsIokUCFinmBnBxKogfZtKz6JG3ZOWKysbr1rG/H96NRXCw27RN2MrJ
QwZxUBVRl71DbZixiVFOvOUtu95XVVG6s3pE8gxPyBC56yN5OG4LIztDpv4u+JBN
B3jPFqp+wpZaXqfXOB7TgKXWTo4LG95SoZBKsy5/NqaY/BMEFcbq8uFX15BrnwnS
PKPz4ttUC/CsrW6AiaWZqsOQqrmqOSDxDsUNfpc35KHaS00I2BFx8ddkdfFmdKxJ
EdE+0N4YMjptXsfMXco63Lkur7umtMpDgTR3TvEhicnrsUtGyOTJ/EqGG0/MXKxU
qw0iCPFI7sXxK7xWaffgmk4SU7djrzEksSSlQEY3uOap+VBPwdQNsPMQDI9pvKgf
S3bCsmxfkzWlANqxXEQqhKCUg4QeKHLL/12tCAhsASA/nalsYffz17xmrk+N1XWf
lC0+ZN22ZshFOkJdLc8gswvSXJ4Yc7mbKXAnOqxLiYmGeGhCApW7HCxF4hXL+M86
oz2INki9hBeBXrVY+NK4N0t7ndG+pT1YsRwjYx43/eg5Q2FOJ+BYEXLg+w5HO542
RTkonqJD6TuDfVPcI59rX6T4YqHmRoMLcvd1UORx+G6aDiSYwqlf48XP5qUkJ5XY
ApeujmwbU6jaSNrnBbSJUj5gAwDhneS6iCkB0RPz7aUqai5WTuhNEjTydMkmXoxI
5qnuYIgJmk4eaMLZVjkKu+fmt5VMR+/92lBAnb1ADePdMQ7k4z2OdlkwuAftmj74
vQV3E8sN3X+W8ICTxFGtT4r2PoPPKs0T59MUszKMhcTogQYRpaUNC7dxAsVpWjG0
aYnU1Q8fIyjNVSODgGW5p+6i5XJLtpXmkX3hQLPiJqticLb72FAlJRK4YmRf4+zg
106Ym7bMaJQNsyCsB/fR5q8w+Go+4oBbdvD4aLoX++skD3O4YDBMtZzqLo+Mvwi6
6C+oLHgLHvyDWu6PnFLzvjeGm2tbTzokfK+MErEqISv6hAhQSE1We8BlpOZfk5F5
+y/1U1Xj5rNLqI3tmv4IGINh3mqSEOg0Bfsy0+GVcJKGZUiQlAiwN+QxtOBEClaG
L/hsQDJznxFyTonAQ23GL9Y5AfbVdmWOyKg5TDnX9xf7WKDpM8qqsVv10wP0K6Gy
WF+Ext2SgT9OxWT+SV/EMrKZLdrcbi5n4uCYHF7VB4MMhSR/2QheCP+9gyVAy3wq
ORchoqECfHiw4jwIUURJwp997FOfqqEHopit/LcjMtLfXEiPjcU9iJCN8BpO6Nt0
nvo+8fRZiPJksEyNatdRG0NJHQK2aXa6tls1H98ImkJZ4Hh7v3HB5Or0VGcTsbbR
QDNisSii0E25ntcGeulR8aUDjpgJs2gbnLkvf8G8uHyLsgF7eZad34K8hp7qlsoe
S9R2CBVUK5FF4K/YOPgNEryvzEAotM9MPySbj3GxI0wgghcTbEpIAd1wVPiroBuz
isf1TAl/wnjvOBuEnEiveWvasBWL860oHxqD4D72O+gl0vTJUc/SC6Jx7vbbFzRR
rYYtgfdbDELiCJmrSL0G4jqNuzcPdoN5pheYwnUkPfHscuY2hZfqOmSzwPQHaYun
4pGzlCy/8+kY37JlDeDBwMq1bFzAMzH1xK4OvnSpp3bqYsw2cpefzNaFr2hl2pOP
c5ncAnrN61W3Jc3SOEn0eG1uky8CzhnEFBqTqx/aRJGxJqEpaNI/BJyaNuPsNJO7
GtmLda1Bh20BKDmPTUp9JZJL3BqaK70Bg5sudaniwWAqRjcF2rKFSkA2aYc8NiaI
psn6lGZKAncfyjVX0pFbyN5PG8yZ9VCZZViWgJphE4Fot510b7lqHM5atBRo28i2
VimQWTK4/gJ0ISzNEcRnbvw6wVNrfPvuVGahuSn+oW2JkMvxtLBpywxDFzQDu5X9
fDqz0lPhDEXgCL9iE6uBH2kdvzm5TW6awToyw23IRKiclml/WKHb64aBXT6/A2Yd
yVRCcRVThmUk78DQAwpmD2xLMB0O9daFrXrlNN2dWccO89LjgzNyXENuAPYWVWxC
+dJ0OXFWKPTMlbmDZzELIO9UDlGg33LHecwk68CeOQIHNWYZ153KsYRXLHNLPMaf
ibWsZVhJjnr1OzWU+o+u3S0kBfYcks8mkNxO467kJSidBydmB5DAdRPOgSczLoHS
Knx3v/ETaW1dHjmNNahW+0toJk7vccPSL20RTPQUVJ+0rMJxADv2dIqwWJ8KdJ/n
uQnlWanZzU/sPMnHKuJw6oDzA4Tq06hJvw0Gi3DXwDh5I8zQjtHmPZ2S6q9Fzmjy
poEfW0sQohl9Rq7CliHbLm4eILfE4l1rkkwoC75vgcOr0RqGkWTM0xA07HKGe2/N
puykkW1O5PNFEuPpTFbQY4vci+VjnjDBuMflWuKq0O1wLhlLPzoPJGRBr9czryjN
/GlqH3RbSKUGvhvZ9+qN0SuBHLy5N8lzGUwVfK1veFgPexP5vwOFlmhoa0kOZ4TG
Kp9ganpzn0QZbiHBoy/Oum7qqqXWK/Ln2cLEuGX/45TozACKjpI7ld93iiyhLNlR
XG5jbsTIO8W1xNJx+CFhbSSUNeD8rx/m6wHiAc+R+FOIvtBIfqlHAT2Qg2hPKLzd
Q7zSUhsFx4GaGptT3z3TARwOKbtck1gnBdzOD6/vxezz6QTGuWUsE5qczCvrAl/p
TQv84AYbpfFNDQwqiETaC6I8TTOf9RvtHrDMUflVCys2SSsbANhpFdRVnGuhytUw
UOmnk1FwzQDRuo8Y+CDkSl/ZTVNZ8iF5HyhGbBeYvisEba8WWcqxspb/cANIl8sM
73LNoLAu5WxQDJBPlKD7JN2xuqqB3DrafI3bqkfiE9YSd7bi+L2W8z5LfArOl2wg
hGrnl3mpW6U1BeDh/EZ0dO88bV61n4Ri6JquERMg69hIRe7G3PYaRWD/btO/WExv
XU52Xu7I1DVc2p0V6t9Zb73K2SxHkeKVyKHe9xTGwp0KrhlHNECtN4SG3PbVGtkn
/QvF/EnpnbRQ/RI1YPxDd5BXn4Jp5BotMk4so7lmuU0Wj6UtCYxF8IsP87KqBSQq
nBl25O7rYBZywWaq6So7WEy54xqS1uiWSD/w+P4qTfIIbNl6IBL+OIdke0uykCVh
KO8kJ1cqd1irP/BpX0opmwQ67bqlNDvudIZffxoKiVbDHpTemjDbkB9pt/rvcxfL
UxEWx4bUIk9K7jrE/GETMUDy1UGQGgK1NM1Y8B1uhTL5kiiRPL6DEquaz9Vf/jyg
6PNFwxV5fSNYB4yu1z8t1vkDbXoI+EilcUuxNPkliswdIBse2ON3jiaXzwBZgegU
RA0B6X+gNqoq0pasMs8C2Uj3pDVFI30+vz82z0GkdkYr2owumYXsVVRsdAivd6y4
ub72qUowUXM0XN7DZttvOBGTJAjFMEty8SfaASwcZfNlndTvl3hnMKedf6Gb+5+7
sSmLPkCL1mfpK0xPnYsBFt3wSwD+nwAmMTDTcmfPM3cY3WJK45UOt9lZZCbyzdno
lo2SvRPWLfJRjjVJC6UguZ4/qHV1teBEaIEvq+UZe/RfbQn0cJXCNHJftOBrb4Jm
xSUBnQqQP+jNDXIzEL7qXtMT4rHyXZrhkn/ii/n5m5HUhmwg2+kSjY1L7o23/q19
IUY2HybKUVVxKceldwpLc1leyW4hoxeaqHlwZIjpRCM9fAzRrca++rKe5iwU2j+V
Uzhoyc+Re6ZpCopcw26nT8WGKJC9lGrDf5aNPLVODPy/Wb58YmlJaYdVxgGhn+4F
THtHkri4uWffBT2DqTYNev5TjQtUtl2M8U/E4IEdBNAxMM7iZKgepc2j6WAEBQav
mJ7/21DEQCzctmiUV6dJKtLXJpoKaA8rXRkkGQsZ7QArIoKCcq956zeTN/oZT/oc
VgxfnpCOk9c00+Xg/mOSD4yTOPkWV1J0gtQyPWvuEqA1S6nL7gXQ9AyFN9s6CYYM
+31BgF3efxqbr3ydwGlbwK16ej/LiB+Mz1KsAuB6fEVOuohS7jdBRr5kBfcNNaLw
3zVpFAMGb0MBBhKW0//KKX9nnZJnHkHU7DGgFpSCUWScx9bIR+AjWS9wRlidOMB+
rZ2cok3thpXeOvcG53Ar60H+ytx3+wVQDr4SR00/eEJof8X2cRZkcsD/WepPwhlZ
PgZoR/tcT+mlxQSG92LcsU7CNK2CdDhkRAu/dQODf4+z+JkLI7O7vQ7Jx4pLK96l
OYGPDhE0eyrUXg00pzXeDYyLR/gucyxRl9zDm4T/TKr5+ENYw3rNmaVcnhiYkuKb
Qf2ZMgB+vEc/EFfCRbYv34yPCdCJ/JAlNLrD+gI8DqbAIBP7O0oFZIijt1cgy7zt
6SQ2598vNFAFLuqQv0gz7TvA0F+LXjEfBZLaW66XHJ1Mqzv1zIKxRJDYlrZqVq/D
TanYJuXwk5ujswtWsSlRip2QGIKrU67Mfn7BYIYpJwClYEBPsvl4MG4D6Zq8a1JS
6lXZrpkUchbQGTe9hXTQubmz3NgaAGiFFi8hq2Xulk4PZkaEarS4WriKSkxEaQqS
lQgUiekExKrhzYciNp+Gu6HgDjfUIQhdlECieKDiJxsrDdnYEMn3nC+e7pMK2SIb
6Jjh1Hzngb/ljiVm0ojEm1Nw/enMHJn8BKk/8lMK6pwWtAtErWpJu3piolaYE5Mj
dWFA6ncbwpkfAARbEkkeQpcE8b6YXYwATzUWXMcdlbvShA7pJz+lGxEo//oAgGN5
SPMtGWfP57VLecjinT/97wsTdj3p+f4EhuwxH9L7fXhBWWvnoD3nRSXUU5kJcHS8
MdhQbQv/WrYzPMOGlmjEKunUEoQGu7iwVUUofvadFhoTh6N6d4NokFo6FxlmxMAY
FDXkqrQxo6v7IE/IEClvc9xQoEaZmdXUPxyhTXkOnS3GxcKo7Bh1KKG0zqcdj4FK
UMwUlsdr+vGbFV0lSuyKj1P7o4rHaU5QueQugr6LRTHV0F0skgt31Asg8ELxPQX5
giIC51f045QNhxcMq/zw/DlHu1MPkGn/P48ktGQC4aGGglBuiYDrgFXtbokIGTWB
6gLMJ9Bor6wQb2f/mLyuwd1N9YjtBtxaWDZ3aP/7aEB6wdaUj11nWGiO6K7gy5IS
DAN4MezuagZh/Y70Sc7dqAddEMIiM4R+Ea2+ZBFH1LDhL1GEAyxBPVFmuJNBJb6O
oSTpkCQrYC7vizDBmzf3BS0AAELn/X+mY0cbZBbqTRjmv9jR9SQkJaz4ZL+HYUtX
AgmmiaQ8TfGqCGPi9xAv1kdjn4nstW87nCfjBdy4gaULZQqP0IMd/HyogAeU2X0V
X2aRBaq+bGzEtWEfBC3mW6dWejSAVrTZ9fgXjOc2TsUzl4a5AAptAbi5hQ0R+6gb
phCJGemPOacmTpxKcbN9ekDtbBGmSGk7AV6Rb2M+fpOp6QC5N0beOiDthxkQcvS0
bd6fBgWBbFjel2KtdPPYuPhznNwLKQIcMihAE52ELbYrqQrVSUNzHW7qfCHGjWWR
JrQbbNNecMfZDzyRaSfIHCds6SL6DrvXGZIyOeS0rQ/dK26c5S0l+Gv5XrZpXzoV
Tj1d3EXXn07iuZT3GDLgDIb76v/iuBOQO6FLMS/OVS04KuFKtucm/afB6U66d3pj
likn1M2J4E0FTa3wX9nE79Yd0XJMRax99a7imYAKHQw0PqDMw5Z1id0Woavcc/XS
BGqMe0aEoHi7d3t3Qta8xkpPU6chTc/pmuHQeLjTXsP68gKL1BIRXUjrEv8ciZkr
bjWCgcMPjsZdYewNkYegf2dUpkOeF+eaB4jjggDEiwlR858y2JgrA+9MKHRpm+Rd
PYko1UReyETm52sYMtC6wDxLV4YG1R8fIIe/W6TR73OePvXcNmYgrFRn+3VnwCaD
Cgqdka49yGlSZpSNaYGjLLl2yGLsuJV5bqwvLnQPUCZFTkkHI2u0+HSPzp58eg+N
ApT8j0HgGPcWGKle1GOuhaoiRmGPWU5DEFPskeg2BJDDtxEqG1CKJLseqMw2qLnl
0B+Ilg7/zNhUtTFJuUC15MXZu86xJetzLCGDDrBYjOCE5rCxoJ4H3AD9GPEfGd4M
+uAyCwVeBqNgmF1mh71iV41fmWGi3QDRCfqq5/RGxbYTxwbAvR0UC+aEI4j0hh9F
ixA025a+CQqpsWToZTZ/qWDoBff5+FpLsWKdcGssKQCdrZC7sHZntDW7Z6KhPtMC
xnQGCF/+I6Ub2ygo3LFxcVa1BFEgX3deS0reIjR8cDg3hLj/g48fb2CDDZwM8u4O
3t8NM943NI/cFqWg3ioPLfOY21IIyK9Hyrf/ptCRH0n34ee1/ftPoEeQP1Msc5Ip
Qh9ej7H8ZImSqDTwxhtqLP23s6Eg6/h2Tg1qnbOSY0F+RbOrZ0iaDo3mV7qaWBex
8hEFQQ0blGZdggvYEWgCGWI1wx6cjPkiCTZOIu4VN3vg/7L7fr+o6rzt++7rAllq
I8sxNEigxYpPGi7yNDZ71xuibCodNZ9iOhl0lXTvoJ9XB0SfpkOq3/CxNxfUMiRz
UQECBvK4w8Dq4fYtl2Yr8oUfAH8IMCRJhvV8G6S/c7/VAqCziNF8DJ6CYQ8ved8t
hQmk2/stCUe3+JbXQUS2FJyZIk9sERDM5lx8sBnFy7nurX9twnAaO4SDb+4SGfdO
ctblzZT3VqvFTQtDQKyBNZpGv1/ck+lvSgpjueMbO02S9s/GgD//85LtlMjNSGSU
BX5U1RXxjP7K2QyJTAnfjVLk0Ut9i2pAaoX6Q/FbFK/AroqzTus6uh9R52ktaGyc
sxZk6p32F1LOOnbXNxyrYzmg76uIE1RIkpP8jydJ4s1UWxJdwSJIpHUb/Iam/J7y
pKIVIwMRBSYpNU2OnRZv4+3lRQPYEXDMAyxO8C8Aypwt5GiMnU/1oqOV5uJMyjMz
8INZhTTYrugWBed1UibsjmybHyA+s8CvsFfQGCpH6C3cmExM2OZt3Dkibkide28d
MntNLdh8EVuH66VLqeY82rcIjodd2yAYTJz9JRVwg1B684uVcohy46cA4FsPbYiD
XRTmhkSeZsm/Kmc4mTGcpnrHrzclmB6TnWVVjXEifChiUFyca6Trejqhnzs0KCv7
QJzZ1eMVKmO0TOeGNP6myBF1Ja0CizDeUdxOkVLz/oM0Jej3v0buYRSmo6Rf7UAo
/oXpmwnp+a6nwzImwQN6HkEEUmI7cTyGadii6NCsPfsmpFEZxk5C+Ea18DCDS2eF
r5m1CLvqYk8QkAzBzG/KqZSzLrkCckOQfIvCTABneGfh9/s4P/2WGutbO4NmzT5u
MQ3b28QkaNlVnKnIzyiga6szegVQS+ZIGCOznvQNB79X8oCTSOI7+aMheH7v6Sg0
9iGmVLTUVtIW7xAeDdj0gPvS2qXzWC86UMzb7zJv1WwDdmC7TdvHLVcHVq/SsFem
aS1G/MfnOnXcbYFWC8y9hUhAmomb4NeLfGX8fVXYeanWctBCgneHUfBJ5HJXZAtp
XjEcbIeArQfV3UtiDEgfw+HBWCw4tAvl6wZdtsbV46+oBMHZZM7Q5eK/rvNejtql
pCssGIocC+yLM/er7OSN/maFyDrGhFW2IK1gP/zoxt2EPBr/n/04J4N3lPIZW3VA
ESuAHoXBQSVOW1mHGrjycxEIQZv0zhmR04EsoFCMfqx4QlXXekZ9+/6fVUqRZEr3
8xMM+Vja41Lvpka2U8TBvzydsEGfIQTpnWCOc/a0+dsDqMjHlU/TXQ31ulxTm9PB
SAsvV5Z0sriVmoaIQPyPOj8QOaVrQie8K9jTIYjEAmdzFHTXcfTpfoPs8JrBqoZ4
Ydn96lT1Zo6GW+UKI5i3ADKleTLp672/0EdW77i9ZDLzS0N0k2ASj2KnrKXlY00k
vac9Nit2Lr2TlQC1K5U462gIDPI+jwtU3oAerhc2Pffv7hjcH/fMjJoDTtnljCzh
DK0uwdEFz8HAvP/lkv65ZkR/6lz/FSE+KRtuh8JUf/7FlFTQqHm5/rp6+DqJLRv6
jldKvf3D4cIo1K1s5Mz2FItaqRjqOhU2eRfAeiqs2MuOftSKoa4aibm9tuII1v7+
FCQ53o6gJiZkEiJFsAFEkBHVf8Ce4rYYolBjoggsxXAUR2hQtQgUas52FXTkh0rQ
w0io1/bjl58EQQzrFBL+mzkgl8KSVadRRf0A2sDlxdeP7VnV05EkwTl2HY+5V2F9
kW287GhW5U4UGNt+HvRWRcVVoF186gX9xzm0EB6H6tkDgsWZwlLOAp8s27UhGfo3
kRwfl6yK0bY1BHBLHri+O7NiUm8Z3DKndfFCny2X77tYk5B9KBCmtPU2ns3dkRVH
0ocdemB/OLRolHrbEJwLnuXvkEHfqAUZl0/BkrQW2sehfeOWbfcHwmaH/HmCgoxr
XzNsq1bKo21OBRcxphBEpaP2Ck0n/bL93mQTmWdsawUwuCdbQhZIUbQ6RUlgZBM6
PIUk8TlYSsia6InJskAyiyIfIBgcCuMuckHv7OJggbuUrp4ESRtziFA2LMMp7Nls
4NI+arKVwwaejrBB8CFvyeb+tCIpLkk8bPpDrnkDAR8flkKZs41LUoOUHyrIDtRT
+PEsMfLZYIxbGk5cGuYELFvBa8wZ4WFTkoam19PduDWaaN+ljHpRv+hpOKiR6UPA
qxgqTSg/GXZNnyCq/ybo5apKlxcD9JCYH+mMVuqnF4jn3nXIdxWB5MhrP20orFSZ
5bWDKzL9McE6TymWIawG6l3ztwR3+Kcu4pigfLOmd4OBSX8q+jlcmp2urkBrVimo
qDdPrNzmwnl0td5Xnx7pwFTQEHikeknR5IqVzSwluHg6HHw010JTXF2eSnX8jUvK
JItN2S8486Y6M5m64kH05HsA2lrtq0tgpnXUM178M5L4R4bqZhRsizA64dUHV8EL
k2XjR4QjcOmI6a9tRRE7IdKD0KqzCsw/0KgZfK7d3yel5bN3RDOXfNlu5ijMcwTs
+dWdAxxmCAXOrMcGjYc8lunfePDWn3S4QnJvkDx5WdX0z5+dpcggFyaz1GEYDNdl
zulQSm4ZUtgUvKcHV5Ija8XyKG5x7vDvWZrOC3SqaFway63kG9Hgto3jnptW5x0w
daRH5BXX/UHzEWdUr1Dnl2u3Alo2OhPEfwcNP7FIgt+Gj+5iZM8BriZSxYh828EB
wSbrIvrqWLt+ieMkdoe+6CdSni1yM0lCaB2pFl4JeIncSFL8viLgw/DJSLQ0zZbQ
mWLVsRnXLKYZmX/Xe9k5TZn5tX1BTvFoz5hB/8hEecKskWiZTh2N0fm7BEgOQiKs
88p8l2loV/9DwjClSrNlaSVdbL0V9o9+3tt/vIeoVWlILyU9omMpJCbxyOLKJ1Fi
TgvriSnd0AV9UQCEgD1JZkpR9O10R9ZdADIlE0D43SxtXOCbhiKWIjxsqaVfP/6/
0fRTvI+jGPt8KwdfbQ+1NeG+vSW+j6LiZqPQnxtV+pxorWOw5XcS3vJIPXkk9e6q
ij0g7/GRgtTWucdGQE2Pw7q/uOhwNKqnczVlaWdDviQbQ/kmbO4l5uhoRo42GQ+M
SjyS0A5wEy/mdER1P1F8BVDTKLkeMkLyvwW1uUEIaH1RGMfIYRfWa1gyUrztNUdK
A+27C0c0wXy4GgoNi9FRBrwtMZZSImheCYaox0hi9ghUSpDGfHBnIIntEkfOO+94
tM/5Lj7EsYFVzrFJNOiHkPJKpA3W9Dk0Yv8hzsU/8jChLOvviQ0X/03VnkKZy9Af
WxutcQ/IXAhu/EUFAQNW4W28suwQPBhJ9VxLukP4BSQ1vzQwd7ry2uVF+jGUr2aG
d5nnmAeBephluYns3hMFdOT2aZbnDiJHT0WifVjLIdFBpRtmdmD8AT4QzFA/80aN
P2P19sPxi7vewsaWYxQiL+wuWwNV+ih8ktv3CpoLl8MDyWjNzZS3LtN61sUhZy9V
fJ7/PHIyCNM3FrisCG3uJNR76up5ULY9ERy+YEFrvQiUg7DzIdkZ5aJgy7jBnIIj
YTr2lHHXuwuyoC9at2N676W6cPjdbxoTjIsNN39d4nu4eMtsQbOdLbL3D3laAs/U
1Ql9UNOcvtbfGFoewEDmDhUiBzgSRP6ubAZUok/K/ZW4q+G1MMTHbKeK3xVBwvpS
i0uskg/MfEPSQ7fRGTaaWrnAZ6VibMzUJafIsF+WKH6PmbFU8571nrKI3gxsJU0D
WJkyTmf2kFIgD93P630z9xfa2AIxoA7JTNJfSNUiWQq4KLylfW0xTAjIFQ/QX+Up
p0WR6wV5YjOZaXTG2HJNJH+vRGHBOF0SfciiwWRkR+Fwow/lpf6b1UKEhtVx4cQP
UzkL0SC2Owgpv/uZP6k++7CONUddgxVq8xjy4Pufz48fsizXvsmZm03e/oo9kwd/
A2NjgL7H/VZgwheke4AEd/hwG3QTUW3sybO1QCuurWfVpAR8VPJg8WCPmuEgwZUm
ea6F+a59pwl1j/tzacaMHZamzQ/jPmNU7f5IoEb6Gweo+qjHmrgGS+uhxXPzYmzD
mbCMe1pxNyvgCm1g1DiolHNcRNJtDVenDSsO+FY7bNuaeWueIrrYcXEkiiwtn8Zh
xY5Zho9aCXWfoY++P3fSXB+I/hqefe6j31RHNM/BuVcJs9HPIw2kR2C8GG9gqtmN
mG9uE0dO5/iyRCOhGRxoOxlrWbBxos9sr5YgWn5v5rb1Q5nPTQDqBT8KKRC15CAI
gpW9B+ZobRHPOty7WRsQF8ff1XTW30cbfmSfpEb5glSBF1SWwlTpJDWQCOOyuS5t
7SJv1ziBMxvSeva31+TX0e4NVLO4oxufELyqHQhOrdkzFLvPA3RVSgkohCdHht5X
1Vvb9wW4QoHc4C7qwUgKsjypPF05/K4ZZNbp2Wg2VoZFNEjzCYo3+STOjRDEiy++
HpWGRV+U5t8cOhobcK2F40EqKHl3Oir44SMfQq85H9hhDhlwBdPVnp6yUYBszEn8
SSOuWcZE0RZ0tTZySqFOikCq+QF9Hm45H5AmGj4c7c3XTlXd7c4HE+QFygJVLYMA
wIQI6Uwq365AW3eX+km8QfVgvlgT6Ji6nV6EPiI4EG2mQ0PFSlxl1wZmN7+Actok
pZv2lnIn6+uRXv8vDZ8B8D0uHnNyRlRk6h0t39DXpKYlzWO3CR16HqvyHeXK+HbX
dcp3+NUQgXRwfS/ovsfWZWkPJUpVZVrscWpwRLXqIUipjpuTJdNo8UhOyQg1Tvvm
DXTfMUJUXyyTwscLis6LxoJOLW7RylZz/walTbmlpk8V+TRdsrkSAGaa9n8iFJ8a
x57b2cghhK3Ayu6ZARWRMEdqqnv53UqeeFmMFD+8q2fP8V0Z4ynBauIKC78Ryg58
XzOcjorsPR9zibnARMoB8dZBd0XV+hxFg9FeoaK5pKtHW79BHgiteU6YzLN2LqP6
9EMg/wWfWNYrWoLiAVwA8kQ1nqrt6v/RCEB160SVgqmZ3GmQzKzgVsDvPie8aR11
Qz+727cjCPUk+GIxrbIg3S81BgfAt7xVQRJeORUwCJPeiCYImqJgs2i+kd3nX9bu
nCkvylahLYWLOJ5JLcZwLhCNbjXBJ3yLG5lYx5bmEG44VvoYkDPjdohpxSUN6WUI
ocXJUEtfrvEW4+d7YF8LUrV4O23GC4l9LXv0xq5g1SieT3mNLxY0r8ZLkqiee/rG
JlAoa/+xHKr3obZQMZoGyjH/UGWJmpVRugJCAaXATwHdSfZxKd5pmqxV5uQDwcQ+
2bqX5S130oQMxqNMS6Adk+IxuBC9ymb59SlesUTPdtAsrebQpwlaD/1RuoIhROmR
foYvBgSR2NNemCF7ufs6s8YVOQWD/5IuuQhSt4rCDVraeMcMz3fHdVPTJSmDq63b
Pjqgn8hG0wNsnNY5iljRY8tKZWk/G0Pbxmuie32kmBuCRL0E+KESQx+DGWNy9Yhz
fb/U4dABIrIrsNuvcKuB6+TFwl6SZVrZfV65O9V4ML+hYUMS9SVwXbU9LMtoP9x1
y6Myt/Iuf626Uol3JSYmcp+vchtqLkzOxYCoLq1mQXHY9E+muOkt86VMruFhKVxN
XAOzXtWX5/f8jx7q7t/dCaN2+GiwzwzSXSAhmudtcXN+pO+uiDfT0dQ7yEWSJ3UD
n1x0zWGOy77QfZBLPwqdqyAD6+qaKAR2L265zko3V7d/nbCTSIj7vEai95+Rt9Hq
OxcHjFWW5tjMuAd1S8CEc1lr2yXES8K59L8tByqC3psz3dQw1MTnaMcXwMyI7zxE
llLn0NHOS4ZyW43CDtNjbNYUuSh6TyOo2s2ViV4YYiBPYtwmrrBB46eGrnUO6scB
b7ZiCuyBmGbg5AoSvUZxDggzx1Xl4ap75Q69qhRsFwIhv+f8XSFh0ibT910TARQb
tAu6w9cpHDImotyVf/1pJvs8A6w+w3W7HnD/xzYrqnATk/JXDxpyu5oHUNZGAcIH
s6vR2Abf6/W3g/ze+j4P8ASPfCrYGk+odZMW0NpNPGu0LlIEaHrLMJvqQ4Gni4EH
xy2aqjIIcnrRkCaanPvwzYzkXoBKZsYZiKyd5EOk4Egzj9HI0JwAy0NQcY9QOGKx
0CIOLe/Ad4DuowJBlOJ4BURBNiYbsVUp3xE8YtqwckkRmGwRtZpVbSzNmtpc/V1R
+p6MLSKfYwtvNkQ7exDdAaGfcN+joxblE8oIUSvudFeUlbYCVU9bTSY7N1NqdaAs
XL0mUPmQTkXfvU/fUdjppESHWRfhFrTXW3AcfrZpVLSC5gyza+Kneuzs4XvAC6XW
P5UYQTJhJHLlz+Y5zDwW1oJ2HJv4KQafLUGPSh3U4/c9riHjUwyhupOiJLJDjjvd
IV7ihj++jmnF6Qpj9aYdKBjiN9cR5kW+TBFCbSSwqgRFcm/1H6/c1HhYHrezbBz8
B26PSYwNUSknseAg1oGTfmXM0KlhsuaLzqoF7kdER5ZbfToK1z068T4pr3ZR5Fps
NiiCOJZCNU4dUSVZg34HKLK8VJTnS2q1vydHXNIhDLnl2SBjJiL6Qu9Miwl20FMi
8xTVBaQpOOdot1MPD1OA6RnpBGx37ne8hezbNAmcBtwqEvQOOMqUDIGryShBdAc/
93YQvNrjo/A7h4a4L0ZL8NbuCzqz/4C7lVK9LUfBASTJ0evWxHY93swwONQutN4+
ftaeCknDDmAdrPkkxCV8rlP6/VsCK4I07QCuZy0qqXA+9n3dB6VDYc41wqtIdYR6
3MOuRyYFgRRXCFfQzXdN1RhLUIxptxxM8GOXI5zss1hklPJLhC6ldMwisvBbshZm
h8k3893JzdtzhGCMhj060jF9mR6fSckQmgkRFXNSeLRWljdpAB5QVt2oeiifbPBC
vVde2mCZ8HaNdgw3pdG+wJD2PsPwR77wX9h3/i2fUFqjqFezsu0qNXFdNAiRqu3Z
jFwPe0mFTQt97yok6yrj8ee1is8jc+X1NuN0/fcUiKDdUNdaxWQyj99CbsrZswVE
qxnr0s+FG1EN6hg0NCRRvhqYrfnl+QFCkQ5NoCuNqAy90NETSh9iFE7rksYRm9Yb
gk9xaXPN/Rl365xXrZ2+XA3677k6147OxSY/GVVPDmlY4aVk1pbekg7LIkCvLTza
5bKdsB2Em+iBvXEtEo5rS6a12JEC4/8hZH02PkawdH5zNRPly/6f5VRSGwQJBHgg
C9GVEW8KxY39XHF4Jp760+xBITIxS1zdjSbIJMlZkGyIDwNTCNEnXQMOoNuyTT/V
GS45b5vzXUCBz78wEv7ihrG21PlZaPQ2hYu9DZDZ4HC/7ZrHYDZnc+EfU23viSjZ
S2SfYHYMqecQxaPOYZTW9bGzKx5Ub5rRodsWhBSCN2hHopQt5s1Gh0u7kVf/uiAI
HcfLeE4719LlCj/dHtbmxE39H2/NEnfPA4aS4RFewCVOhUcaum3zDXLHLSuGeRc4
xB2dxVyewYdiijMjnQHfktajZe1/o3BKNLP/H/MtD2RbmWIOX8gHjm1vqxhP+KXC
VP1AlAk2kIPj/1MOagKJpNjvcraCcy8m9XPXiBLuZ/FMBAQYOvWyk3rsYTOsgUVc
GxgwZ/QxfcMG7Wo6rH0pBNyh6DgiKcUyJ9Gd07dcrpfhCic7gvePqaDuds/+fVWD
XsOe6w+g5dj8rWpgVEr6nslMagvL2sJEoE3MA3dkQFsq6Ofr9LthdeBNhB5hma7t
UA6scKUDmACuh/WTv3si9UCtULX2C1jfSKBPlkK5w71ahA+K4oHYxBdKhB1pVoZI
5XXftUIF9E/63Y4lgPgk+f3bSm3ToV0Dwcv1XyA9dXI/agKeTx9i7pUflM+H+EiK
XRTYBHeARq/5G51rFYf4j9D6CUriAc67UpyJwXe66a7w7oWq9jv+vHqhXV4k9+fW
NyN/vtueAdE+q6GfaWDECXvmSBjkVc4tGxifW2Ls3GZjo9SW7jd3C9nTPjm3HSat
RftTT6hhCIcq5Io4poGLhkXxSHnRO+O6n0r7Xr/PrjFUFV4rY4SRTU0cRUko/J/y
nYIf7geql3zJl2380/hX5N5NkW5Vw7+rH6ytMs5rvacz3gC5zQFZasCHwDy/+Pcf
baTq3GWHoOzhWSkF81kcNFM87/nrgZFoYpCO2cwl2p2GHuD1coCmY2dwknbDvSTS
kqn1abzgsfYloEsIHdEKe1fyQHTeTbhVL8HjGS2c+YOZlxu4kVA84y1Jy7eHG9wz
ASYJRqNnHTgi5iomVWNUNOVnhOn7l/+PYHXtFvYzDcCMR45BLo0oUxTO6h121zzf
4Jw9jZpDPoJUnU31C/FBXYmfCWrFI8GHlQBKLl3d1Jcf7jd0iFDfwRSDZEGdvywh
CPgFGQzv2AeCZDkjagdL8EFFj3waABCIIeQLEA0aagHMdAJnbXBtlrt44xLl1gNh
jZu+lkwRIK22TfdX9gmiF7lZNab90AKYtMURX2m0zcIkXerQvijm0TJ1KFuphR6c
nk9a2ntNL6pWP3snZiB7dQoMbE+B3Y2ChrfSYvISQMRO97gxtfy8SXskwoGrPuxy
Mxiz3K70F510h8sWRxEMmZ1VZ2SbKP+nxuyS/0NPCQYVOTY/qX6DYft0+kVKCmGN
gNas2CW23rgj+Ha3kwUECkFUHeSKmLUL95mbfa/MCjahLtFHqPnmSf3E59SoON+Y
NZEklIxyTxB+Acwk+cPRQVHv7KDfguAYlQA2zT2QQBrTd1jk0Z8fllVqjuT+QMSs
AHx+kn4OiV6WPrgFFNTS2VbRuNbfUB+012itfYDaxzjBkQ9QhkoVdzDwsRTkKOyI
tSG/0Yfj2crzknB+wMEwh3j4fhfcORmToegaqxcqAmVnfqXzGlGTCL6qCU4K3ws4
rcdBU8KmNlmj/AhVqE5W0FQw9gBqmP+YxIpgYmrJ0EH7vQNpT/7wlG4wau1IgaNC
BYBJEhoYwtcNHQ/eZnbWBvwHgt1NuosBF++3iySfO9V+taW55ggHTHt/8GJnje7P
zIi73mEI5WPMXsBEvvgMl3fabLEZKCWa7STLPzY+FwvSdjNT+8m8G5Y5wGJf3Nva
6Pj+6W/fbuuXzgOsjmvgImsj4Md06aEFCmODoO5fQYQU2tEAOjwAAhv4vlFTnGqs
24jiwr0Fr2A0RSNHeW84LD7uJVMv0l0cYQMK/IuyC11THXEkeYDz6Xunxaf9oasq
GyDgw1hOdnoGzKENpjfhnsEkWpwnPIrnQsDZXXy8g2QIKWlW39DXBNsqGoRyowQM
xE2YbRiGIPIt74gs5aSZHYxaxmVSWfjc90SG2FR6jv9Gb2oizekjvoLzd3MaxzjZ
szL4TwWD5nfnpIw41wVwwczjiDl/yJjJJpI3taZD3UokSf12FpPrMLcjX7nAoYra
bUtfj2wtn2qsuwyyQx0EiJ9xe45fyOBfCH5pDJV1TCKw9SFcUMOHWYkSbXiaj/r8
CJ3CUgPV+deaaq7wrenUBUq6fP7DBVnKX3BJ20pIgJWXOI2g8OeQpV29mp6y9tsJ
UAeDI/5MV+RR6bGXTXFZnjphZNZA4lnDuuFo05Xh6dekP1mD3YeuhfFrjMwUIOe5
gmYG+6trReE+1c2mZke4rPOzgeynZPcVpOAGh+bmHzUtIvLV2eWx0VETOY55GgWj
1vxeQzPhMvAhF52gjXdBVE93o2adff+I9ahbLyY2fWM3v/EXRzLkzjnr47BEDpk7
Yy6oqnIl1Rsgfq78uzH4LTIh/Ibx5RyTt1ZG6Ic+pVvub0a9o8Pgi8s1V4l0CBBY
D0BFMFv82Pl43jGsJHNma3JYX84mtTX+5U4UcZI1iRQMUqq6N5j9ntVZwuQHXAH0
OuzSlU+pcfjZlGNl/ec1pgydx1s4TQmdAGbL1nSVLsoR5V8l3NlRNokO+0jbvKe/
5CbIBc7J7YD9JZRqf7SbB/ykwnN9FgBZlGBY9rMma7CBrBj8yStc1zI0DAean6eM
H/2Srwg8B340d5Tzo2AP0Mg3BO45dNuSDwNcmqgH5SB4RCapiVCitlLkwZhDXF+F
J6Byr8BOuL1NQUhP0eCe/dE10gx+f7zexqtatoXsFxBp2wV4+CjwJ9f30zb5rkYE
GiBp5IQOZ8XV0cmbkJqbErKIVPpC6Wp6rybPm+vBCQtQDBUeuyD4fFgTIW24Q9Fa
Sf4LeU8rRhJTUSHvm/lDGrzMJT1GGGPDcH587FHA47w2QtkXjOsesbHs5COIJzqS
2/qNRv8Wal6lqKW1422n8ZjtiSheqblSS9szTR7MBWetcXOPos4ZeCoSRKYGDknB
J92wqjx/nbqD2CpVSo2OH0ghxa21WRYZRFBQbt0MHVRbo5eY5gpthf7zy84jeyOt
Mp+OPZm21V1CvNEMzZ8amraC83cWCWcNLDMIC7qaiG9K4ETYvVf2el/W49lCiudD
3/HAFTrAApGq5qvk3kanZpU4bFToywgUzWB8243CLNflCJIoZJsacKgv5jaTcmxv
SUnB7ZQzAMTbCrFHhW0u3sHxp2s6GJdYILMktX/YxIwt3lB1RVgpuJWqlUerNlYe
fbkGRGB6SEnK0pivjlpvHjUO8TNTW+MzdvNWjdil9EQK1MaeyF1zacVBjookcc4E
Z7IvRg/W0nST7UVR9IxO1X95DSTGMfmdRC/4bUvLnvCcZlFT8j5CHKd4MXvDkcJ0
JaxoA//JxL+IHxCL8lXoyTHDEnChYsiqdZsNCk50tw4PKWGGdcwEB2xcxgisjVY9
M/AKwk0vfDSmVp1zzgKLmkvpulwzDezoymzkDJJaT0VD9cnoHAdSMeY79Lm/vecs
FYF+8k2fZjsos+MOFEMhmzbQT8pVAjKN0wy01tbBKu1IwoPSp+PUYj2EqO4Pdisj
lb9oR/NkpYy2PfIE3W4lgItsVAeT0z4An4Ab6clzhLFSm4cOjiLrCwyzuI6ynLHD
hfhbXmWjSIrfimoUPCag6msrXF1Pe9erYaQUXfFY9cyef98zV092E7amSr1f/yhV
i8BxLXz/7/CkjZx1ATnJCeIXXCWEzlQDcgDuy3OBorQ4GT8vEmyh0pu3i3gvg/K2
8eyccH7ppzte7pVTg+QPqXXkGbWCULHimYA/eCzeTEYIq54hkcQ29arrhUY6rhsi
YpGn9QlqPQyN4Mbko7MBowfji0ti8agzycG3W5Lar/TDBZ0zRCYFic6kTt3eO5vN
GEtnAqReGdZmQG6cW5wNvVCY/mDwieERRMtPThmJyVGX5CttJtTzRE5hMjfWujod
HozT4DkAD1mRe1q0eT77Etignc3BxVUVh2daot+mc8da1HG2/BnMlZlYTHDy9vGG
tvhYfiRdX4av6BQcuJfut5BSojcoskQwVysyW+B2MxAkKP7krleCxw5t2RrSpzLa
ZOcqva/H7oyHo2R3oqPAtFfwN5DNQuAMHxzOTL1B0cVL61K/VypfwYASazvTnE20
ANk+fIrT2/085qBOM1tagfIqlujWwZt1auz9bDt0HkZ85r+bjl1VLw7RekbTFhW7
cVcJDvyBjbLmfCBmmKs07lL64jFJDrPdMkPbzbEwX/sfw8Yi6VtRJtuxRjffuQYX
YVjyXzusrloGYJk4JAu2270ruZvCBAcMPWUU4NbXxdZGX1MekMAC7nmYj/ufw+P4
yicsL+hW+dg80r4BpeirpCm+34L2mrE+o8CnFNzi0ru7QPhtsfuNoQlRdA+am3gB
MnlUsPfyiacllDXol99NuMEHK0Wrw5a8LL/Jh22ymaI9QP840Hb9Zg+A4jO3n9ao
5vgAOnVBIhxTzIbYJ8b8Jd77m0wSIxCgzc2+HoLumVtygVKP470jlmiAAwnmGKt5
MMS8IuUm5Bk1Oh51pXQEhJSOmj+6YaJTNjfOcNaGYiK/LSVzl52MO8KRMRLa1U3i
GqQJVwONhgGeMnnFy6RzDLhypGs1ZEb/MtuwqLcMqTEoO2oFODHjrRZ058VJPUKw
2HKkG4bmmS8Ydpl3Y9O8CR5yMC1jncJzV9J7pIZZx22FqES3Am4IqSaB75IL+awJ
LbKOmZzLweC7Oi/HDE4hCrQTpPrq45qwWU+Ac+aHE1NFcUfD8c+sc+OVRd0x7nEJ
ElEG4WH5Wo2ppKYKxd8YXaYsxesslpXaxSOb3rzcnCV0yGuXD4oPhhNS5fjrLXrc
SE1v0KmT6A3/TTPiH6wpTYYmbZ3/N4cKXav+Pkn3Y0z5POFG/sLNkRmnoEbXBL+n
VzcXh3jxcvEo657FPAT5+yrnRp4DINoKWVxcn5TZ4VUptedE7sSighiJxICAHYh7
a2kI9r8zbQwSW6ar3qdjUSPcQJTyOjrZGe2T+lKV5tL83Ye9aCeloVMKZq5UZEHO
GtiR2fDWotOsnwoW+a22MNhHQW2esaildZvIzj5HZBCtWbbRX7P7w+T1/8y1m2b+
Y4PvDtBtMdvLdy02eE0sQAi09WjgQBeJ1XoUJ0K0aetNdykdb+xViLV4NmMqs/Nx
dwnIpTQw1i3mJRIgst0oQkvLN5FOEYdch6aP/8II982FHIfBn2BDK18ZyPyvCEB7
Dxn+/fXMUM52rXjC37LP6cdMdkciDCL7cQCw8MEmeABuf9R6Ad38hli4hBMHYJl2
0O2u9V8mQ3pzOvTmx6cjPzULlKm5vqOdArkHMWAoJq3CDCJKKPn9qPP/io8QVAjc
h03eO3iiobQoskLu4mebRwMes68EOToCEhfm0EE7SkD+CrFCysgbx+5M02yweZgO
pne/LfZTeDhPw4wjQwpKoKbIbr1ZvH+7/y3Wd/pCF1Va/I5sJFJKIZ9iG40iMBcC
EgD64RQdGsP0Y0DOMDBuEwAoytNwddsJfw5US86uMm1vXJLMdNJ0aXaRx1p8PIbK
eQhLHCzO1Mnp5gf6+6B9cgffBJeKxpzz1yJGxQGePzhq+At87QSEUuv9raAoIW+1
kTfkIHAkLthKB6zM0LEgYefnOVsxRCXHQBz6eHr3TqntPHS3s9apeQLNGCFSSQ4w
o+nETjKqudp1IdTcmzLpERawsZOGBZsg4A36IrPwv9mbOLaBcqvVDCL9WMFvkIwF
4jtbTkxJZMWGKIhBP9re1kWqVbgLTJ0SABI1rm4zc03MRjmTrfDzM6Ua5st7lV0f
o0n/l88bC/VytOkZ7rxajWMJDpjEumRjUmq15UgpSxs2unmxAx/VtLAOOdzVcrVA
qhWTRNkvQ8pvxBZxbdb4dlVNNqqJugA0qRLxokC666AksGhi8rpLqclu5GmjI+9A
kJZs7eIMU03MP17ZMv+Ac4F0LLgftfZUTf7H7yXlmSohfzOZJauI0naxPxPm6crD
i0ziUQxzl21XJ4+kD/m2Rk3G1KU/0yg35l7UVLcGtDBut5MGL6t9Zk/dYkHOydT4
Yrbay0Uwmoy2oiT7cfGJrfK4OcaRc61ygLkkPQ1MH11/SMsxJUnu5xyhHOTDoEWy
izlYs0Zey5h+pr5MbrJ3+Wm2Q5iift6qk12HsTAqRaVfS2lIMhw+2KSiGz/CJaVe
ylK5+fRYwlFr6pmThkoDF0B3NcC3bo/SS13YJinRTzatH0n0y1vvTqwkr7vDue4z
BPkefEllazUEeiKbHgsrCtnu44PSYQKGnWCY4yBAX2s6B+yC1kSGdlIroOQs6Xvn
juDwVH6/XcDKdTPdIdAYs2QB5zBVQlN5BSQleIJKMv2PnLBZ2gQjJXCpk44+McKa
eyYkEb/7zgYeYJDkY2HWAEOP42hFuPtu9+XaA/KsQ2ppilZgTaMZlO+O0sCqAuZ6
rrc6untYGWffJ/kxMUHfJFuSUbMOgi7+iEmA2tL0wFDmpBfE4/J1iWabcPzJ6ZDI
NQ8yMtkpWqykxq6/DjP6xxlZFU1s1YOt1o/2dAp6EZO/zwYopTGUd3HE8XvsHKYb
4knhmtK5KDqRoTwvjYasH+XKj2tmME9I+oQ4jxZUIn8uF2IT33+wHB7HkMSNfVYx
OaNyDG6u+6k2ZVb2SzdWL3qU0jjqpg9MvcBRxd0AplieqGnOiJ6DBXYyI3m6clSg
Tq1UgbCCDhI/pGQu48g7CVHJKV/IAzEBb8yM+4Qtp95dA+gRz5EDd+b8f4lYYswH
BrSnryxbbr350a6opIHvxwgL/OFYW/puS/FisOGT51m4ws3P+xvjfRI6feU6wC5Z
ltzStyRc+2XT6463vV7JaGuWROQ1uG51riG9ghzfIoUxPgxpWi6RyqmJPrf0qh56
vAXuR+J2W+VGmJoAM5GCjdrLH8Iys26KoC1baarZ/3J0yTI/gZmypmXByy4kvVPj
b1Tw3UYbI33ClHsxA89KCF9+BQRU8vSB0Qk/dWOej+vPqcsBhVE7JFClJp2oHZ0l
NFdtWLg4mkstwwItqBeHzAQQapHtAHYSbrBBbCTdBVNfAt9RZRbqWd4WpDwUpq8y
WIFa/kePkTM5Zm+Z8LMYSaiVu5IWhWKrJnWcDN1ILhXrQba7AsrCQ7l3NoaFf798
j9abWuDqlbfeAwRPi+OMQdOJO+9b5hh9PMk44xg8F05LVTy6OMSsW/RoO/5jLiDP
Q4i+VAPBpo1qF9b/yHo67veDYZ1VnS+nVtSCZbYg4MFQbVrRXsPhO12E9RSJvtmW
d77gWEdYVQhLXjQu1r3e3ictXhYDBdHUOaanaA/LwYKvqGrv4IuavNw/ivHsdTTL
qhMIgOVLQCm7bGYA99k402jgRP2cAEI/Ut3WH9qnaj2whX4u8ulpp49jn8q6J/7Y
T5XCl+zg1zoUTkSVjlbHlmFGL1U+VNxgebYnrvbMGgVHOjUtWnn98fthi2xt/DaN
PLoWFvoZLHb89cMAd8nwxWgxmbRdV/YltXBkTGhFj+EJXo/u6cDljYX1sqVtoTGJ
20lUIEakyi+jvp1DmU+TRJkPbPkdgo8UyPK42YXjJbuPpfGqYpxsj2O6fMehzZvf
dFd/YAeWvvibdei6uIfZyFeqJe8w4aCw90u3QK0VGsBL3k7kCZGI7RdM/KjAXH7P
sh/0OtgABiaOtyFm2t6ZCG57f2BHDCP4iJ56dHriXeawvWA8/CZxVyUljHTg3pEs
14RTpv6lbHPDJ08xZtRmdxHooTu68gt/iUDXOZzyybLo/6yQjTjC+KmlmRtfpNzB
WsBqxTRd5Sq+CfkMJS2dWPKQ+ym9vS0IwRmBv6zfTQPyMfVLE6CGCb/YJja2SZ2T
fz8eH6b3lHBAvxH7jYTzlifPYlE+Ep/FYX79tx5dOL84rPNUpcSMb5BAveqTVhkj
lQIozenrlQ/zE8obq0B5Q6dWhAVezIMBoWnV74W+daDeOXoriAD5oE73cgohhlNG
Afv4lRK+zeuzuhYrbZ9ynPJZ8Kx7TZ7o7e2WdzGqOVwlbeOuywdtMvPOUVPB25X9
gDliaRhn560NL5l8vrgZ1+gTs2Vdi75HwSBtw8wl1iQV7dhJbqJ32z147ogF7P+j
MvbKj7h8gqiv/z2UxsWe8zj8MZDAI6fqE0liwEiD1TcqzntNwxTlzyn8UVk5+t+1
q9k665oG+ZfXJ+xmTuftRx7enJVUJBsE1nz67i4v8kiqXOgoMyecLMPeYF/Tlu+f
OJ8RXUfV19bXRQ4m/LMdvFbHMgw+h4qWLjs0WMS8cp7EnWIywp5xGd0H3DzKrn9s
XyF29Sz14r5Ya0az1iyhqTYqsYQhr6xgjqLRXuKxWhz2dc97ysTIKNOqdBEPWeSS
Tg7qKZj9NJVXUO6E07iB9yWBvKujeHnb4DC2DPuCCjstUyaB3PVnPrJh3K2n7qJL
Jkzt+kAOKTUaC+WciTQw9vow6WJm9Eu3huoJ7WqnG6Zo/qPOGORH2r4w6mqPmGt8
muyNgje8BzzUWwNwMig802VykDfWBELmIMI4sc9TyuqjmZmCcYbeTSTDNMV7VdLE
DLU+Hpb36TtlwFyJ/D1HlsHMs3oYvhhINHC3IskNlRUW+X99Amn7JLCoBx9EL7Uw
3PwFakw/PNCjrJxHHBO1BxRQ85ZSisRWhU1xTIfdY9sTwT8Dg23F5J18PDY3LTTP
37JUwbR7zL6xUQRBUaUNAqtsojuYRUVn2V2usef7iJ5oodUDhMfcGsLcwHgEBQDn
44+wJxixdd7iSxOFeYyH7UyHQRHfikzwR5KJkIk9zSWgALtxQwqN7eNTyL9jx7rb
3AN2cpV6RpJPryKYDB/1KQEO1jYc360qlU1S3HZTrDjcWXw/9Mb3lFe0WQyvxlF7
LYo0p59jfqx2qI3N41eGqOT0xEeCSl4xsvOKMPDnvPO6/pLTLPaG9iEJNX5/3Lp5
LJ6zhYMEzbXPjcZNsGzKEWTknwlGz6iEqPxBNMb8v8TYXZJTfwaBxMZPaBRA6vPA
HirdSTuT76touDym8SyyIqAOiZC7CqE10Hc9dVxm1gM078xQXgcLPd5Tl9cOQSW6
MeuaKu4qagf7dmPNQ7O4Li4uO1zNxPiIp8kYJ2tWa9EwMGB33KP+jzIJ0OuNi2uA
ncRyB05ENWlnELm+cbLdqcMU+ETVWKosaiRD8NrxlnFyUxe2l3oyt51O2wQKaEIk
gdi3uCNi4r9Oo+GEE9Z0Xd//XY0NvQ/r4bR8R94kR8kXgu5YvFeTV4RsEt+ts0G3
+vIwd8/a+SgqRH6keMDq7hPpgjVau/iq0ry7uW4JqRcxcIV3/CSqAmAD8CLiLsAf
qnh0nc4akvSF7fjaQQFfdu9Z4Cjx8TMqAaMJB02YRT5vbKZGzuk17MkbVocJ6I8N
AXu8cpgfdlnwJ35bFqPrD2R1J6bn6k/Xe9S6UAKUwpiQ1v7SQyBM4vFTSovVNMQl
PwCPkUf+k9dnp0C1z2LH5sHMvE97NmBmUNsgdgSB/kzrkZyGE4j/EMTCi3rnhaSQ
tyuQc9tH9SziSTsmqEwXudj0sHc+yY9FQuA4pVlYzUJbUASflcKUNa6hDXHZiFSD
H2dSOXZ2ey/vOR2p1S5UZZuyEX/OfI7CZlqYLofMFpQfUdXTrCH0YcZPXGvh1vWy
3Bh3LPfGZUK3qmck3YRJEXeGvOjWSl2KJZ14IablCD5ZQjQViE//Un97kHq6ZBSe
GKB7Wmk1UlZAETgRkdTZNSPNVFsqy+W9X8/FTLFAaX/mRJePbQvGkRG3g7+tXi03
rwohV85Dq+LQo075Bu+oj5BB/+/s9f0X2YcneMuul+BURK+j9k3gOfp9pJgmLmg0
W58iCuXcN0JB9x0Co/sFGZTxhS/BzLYeHf66RQJoDRqsqAXiJIFXIMDGqBKkMMyU
DH9kkTRadNY/v0xwp26wAbWczUeG8WcjTLTieoIKqe5VfBw4JKWPcNxdXPU0eICl
bEyDooiPLYIChkNDmdcc0hSu5DIjC3Xs+cLbK6vRWKg9OHK7G7R61u33u0orXO+X
RA/6E9OsAq8MtjpjIqmNOGyGi637WpAvsH8rpI6E7J1weZh1ro32vIPzK+7MMt7o
zJjhfitJ71QGbvEK2jtDtWFFlZNyhyXIidNVsyPK4Zohg+DKRGD2X4d+fpTYLHL1
PIT7XXMPVeFp6uus0mbxOyPU2j++jbSdaOcc8PMbVsiWTOyvt/3wg1aKd2lt+sbJ
joLFCezDE8qWqRkzGXXQSfhn1Eu4NwMdewP9qlWSD0z8UfZIJpQUxHTd8CbNtnqQ
DJlE9ho/FUmOpyKlc7cdbhvGCLfd+dRml+QzBq9/PA7UPR3AVuUoKS2qa47bLfSj
f/88FcWl586541X5bKsXjrlLql662F9GbR0z9ERZs+1mfpLWqL5aeTsCsqjO5i66
Vs5GeuNQW4ZxF9/8SsG81uuAYCaCdfbjnrShGFR+aCBo5L/kO680VWrPRkj1JL8M
h6C12atOwG/hcNrr8zBsz9sWubEWSQfz7U3dk9lGaqwLMGctlVqfHQYDtcoeiwRV
i2+KPa42LbC6ZquICZjA3zr03xq/MxIvO5+3AY3bZ2WfO8bLWVYlhkBfN6gtG41M
9dQqBdVMeZC0i6xsaDDxYk72GbzHt7apwSpwu9zwi6Ro4VqybNs2LWdffI7nMdhn
+RhntYM/ZNQpI3tp+WEC2rTUUeVeZr1i+MHcrsRs2FNRJYEop1RRXUUvuFuTDPzM
w6ON0qiFi94dqf4Maat1RE1FTCq/IGjIhES/yXVhqffoXftY/33hz6HucKJkyxmq
TURuYSG6b9bOIoMrKSZttcX8Pu2WCGhWwWwKSZv1DizMYDXiY862z9eYcNnetqKo
aYp/t8fi7dGtgeJ/Q/GDCv53XTWuZWt20cEKi+fs0qgTY6bXA5DJgtjMHZZr+EG6
6Mz5LrkMjL8vz7Fu5y41dxL0MZtcFdpydfTK5Xh4NdOTfDB1mbJda9eMVG8XqDHk
fMqdlw16xYeyUPcSCVPrhZsz+B8/Cgk1BOy1+Mz20tuuCBQj8H/dBvhcDRJBQQXJ
1TIQocybKPnJy1kvuwHSHJaTl8xx5JBuKgv55QpsP2Wt5AreUP4jDe2n7ddoD2wP
jDVHOCLCOtJ2mogsl5uj9fMvhCIHtMD2JeFGZKnj++/4jZfzuF7aG90XUlgTXp33
NTiGIzUu7KvC5v1f5rUjaTiYgIWrTM1rgAzvy6pbxu/YqUUMFB7kAPBHgWDtyNLs
BTjMceSldm77FDFYNG6wSR0PXnnPfTKXMhsjiLsQ2UNqHrKG515cI+Usrmfkk0bZ
rrrOFMiuF3uzkW1lAZ7ETSmbwEAgVaSIWrS3gJHhNUdsIEylzPd2VW99bpjUDR/o
QdzzUlA5O3zO5zizSMF+nV3YnrO2EgK2cdJkqUPmgKAY5ZT3Mit1bVs6PsVR9ogV
ZieDQP6MC1FIxcBGmraYr21fN07VPmEZRrHFqLQepu34PM/QcQfyfpN0I6XbZYCk
9+G1rWzfYBo5jd4rogiX6ikJ6a8rhrZESmmW5tamSLacVlO/9K7AHtxWxPiwgL+1
fr6d29K57UN9XVAeiNpdHYpZA98PkY91m9YzeBP4QOoLqQ3HhwOCOMN/rhkjDFuF
+iq85oP4nOW9aJoELjrm5/On8VGlu4SkCniQRGUn+dTIp90FK10AgaELj8HalWwT
X8RKF9vxwjSoTEyhC/y3lKsgGBGpPp9ag0jh7UNIHxgBOfqdvzSTsAV342q0xv/k
4cWB1QV6GK1N1bSM8SCXaDwFaFRodQfy6cbie8n+tie0p5EXBKIC43VcFRajFdOP
+JUVrI3YVA8V8K70neQsD2w9qBeCxqwqUlWTRtLSVqpeyA3fWd+IxTsUxlVr94Jb
b68+e2kRjYeK1ML9jzqcQD2nVIMsLXAY5oxEO5six6SjtGsFkl3hFqt1h8wKnwAj
Mg+Sx4G3GsH2e8Lb483MGY8dxcBOuFBOF8FuEb7muJ87qsUrk0ANJGKIhIvj6TAj
ZpHlfv5/3SY6eusEASA5GeBsz/gttYLaRF0B6yEijnnZbsNVXh4FJKik8DytcvBU
VFDc7UWc1K+pgYJhEKpymUbIt9xw26Ds0Wzov+n9tRnFFPuCjz5/vo2AQTfSnFtN
fIdNd0h8tPLMS482w7K8AJbABrNGi07zus3swzltvrkepX0XlpeHuzTy3/WEus/i
CKop7ZD6QB4t9Aq7zEHsCqOddEnsClacbTlHJM4eKdlWILyGl9XP55HNtvWzdFpn
2gE00AyS+x+FXQ97gKylhIfqERQybhrvMVd7kqMH2bW58dDWfLjVy3LDFTjjI+u4
FsHEncVWv8rdexD4txTgVp+odxY9diEdsE3k6lNmtW71HsRI3glBvR654k/8veLz
5dPksTh2xPIlwBsUV5OcbrcCChYMXeyV3BYycgD+JyyVV0PO1zJx2Q5w8a0lYdKi
lOJwbPndJn5u8RBUY3RnQmW6wVqH7upg1f2P6PQU8msYpQAbjbv5BWPeQSYmFSIw
6iRWVHLsncZOOBPzIwFyABtQc5ZUiA/sUbW7pzhPDhGVJs4M5qGrQRSXrTNqGFYg
7Ynv/lId2E9C3si3ytGHoepT++kBzLIi2wisV4Xi+hIWY6DYoIT2yFLHbf+aHNf1
keTyRCky7V2uMKCCJK8+LMrYbz1foMUpANJhnXRrlz5UO0B4MV4hb5NqowPD0DsT
pMNl4XTIWFJInFlmegRqwaLkOgICACku70dnopz9kQ05biF8+RDkG6SopETuLSDU
Q6XaM52z9+ZVDEhzkJNwO72yhHSHqJDlVpjNmGI5ursyONle+BDKEWr8ChYiO0o3
sypmJ6iIxtFloTvHiuFz6LJe78D0cbjWCQkJWJEjBlC89krrwlH4ph+KBDdkXwvF
WsAg/IPaJAq+CUHxtNWAZgi4MK93vHtRauXUAQ4nqRh2370hqnbHMBxGLAaaSd3g
7tSM0tUrpw9gQ4WH7oTxXNKf1fjD4SqPJOuYfv3qAEaMN2knpoV3cphbB3AQkBmv
x6W02vJG8/6LmFLvS0+HUFlihuON69L+Flgd5hvvX9IQt5Mz3vROtdopDK/wj5My
y50VeJ9mf5IeboIxD3NS3xZH2551k1hVFHiDUXEjSqI310CmuxDidqPZ7ihK1R22
G6sx7H9s1OGA7oP0aKZ8zmCZtSoH6ttA1FPVpOcl1E36uFvk2rMWlQ/YsfqF4ZHB
eWvw5BW0brSRIOq2unxbGCBSl/gFfbfNGtvh8KR63XsXxzf4P0qwNrhp3ohXNuPc
qAKo4gjH38jTZysXsPVHwtQ6gggEDIHwF0nRXRs8Q8eLFAH7hhWbJXMim3XJLoQd
bayO6WJuWws4go6C/38GcrrZYGUtb8ST+7NqzOZqy1gszmgXLvIiF4YPGLntQK1c
ZHtoWUYW2t6ohe2AeuAO8UwuJg5RgWfhew1IKsudxDZDhTyhkTT+dwqRcAzz/kYn
6pFAjX8yxjRwSc2Hy8pz4F/5Me1BLMxiVgJ3W7/lRIIDQZSIrXfdscniReZuPdir
oVPsGascbGMIaS0S113R4l5mtEiDifCbspBzg7CVDPPjkOh1STxrTIQU2sTXwdQ6
TnU7DIlUsbvHHMxHrb28DHIKKSvMUfd0XuLxnFrrzElO4/LQgEfObHYxFbCMM9He
mQt+fn/hi/1cq2rX0UlLxZQtf36OofHdQLDHvTOyntJO/bhe3Pyoz9ZMgdd3+oQl
Ro9bWVwoFLy4ADH0hBOpSj3d6WAckh4n5W2oaAO8xg18msHfEpSRzX7RMgKcxvv+
sMfPI0qzAryBKUhCsu5beZ/avEcFphd8mHWWUDF1hg2hjaxfJF3jlmeg8S9JOihE
TEveNI3xa0rs1OG2eUlTjJQ1XNHNIfWnxEzzzd72CroGG/7n0XS9XNwvOxUVvczC
04vBQzf3zdFDQJ72lg7uHNj6NKD1xaJK5go5WcdDRgHouNpWbQ8ECB4LHIiUybTM
lPIHqSoDPdQ1ALuCMJTfHrqolJP9EDv+S9CnJQmWXkPXYHwG5IGf73G7QT3h6GWS
24Id1lT1dciBIEI39T7HwuWsQXXHei3fY0mDI4mH7LaMU5L7/eY/hPAUHukxh8/Y
oy5c5mNLAwJRt8fkcf2UkKHP4CVdDEemS+L2g7LJI5hg4zv0d6Dd/Im4D38qwCrx
neUARpv7mVr73nIyGbxDVOP6LX/Jbht+gS7tmrt3Z2BCCrpz3qfj2BtJ8iD90GK3
LnBPQHvo9K8KCSRvSaxvOKqgohO3118Nc9omXkLVDa4U12fPMQgd8eAX6p0NM6D8
iNcvIeCdAY5gdcB1oWLWjR1bW8ioJQrhXwoT2nfC2Wk1aa4/xh7NS8LPAWZ3UtKF
VUxdG2S0IHMZYB6H02gjzlxGM/9C7XI5jWTxUcXnUPv/KTnPGHz1g2O0LGNtSxj8
7H9F3Serhq6D9ft6m85dzWjouvisTpSd2AZbrWAj8sEDEWJ6kovw5o2f1LFYzoVh
lUXAO4qtQRTSdemmhjyxu7yCgq2kN2XMBAhVmrCCQlLfG2JPkrIreqXRIx7j86In
FLBg3MOoiLaOHBtU5+HxkFcGLR9NyEbhD9eN6QSS6cQhnn94ryVElfLODSOgIcMe
k3IPkpeAFnqYwYvngMpbf/iLY9IerXLlyyDly5F4Z0uygSlUWqdvM+UUY8q6VX83
z4km6ziR5EusV6GbA3M3nyHw/dywxrJyc8RdI8SCFPBuYQDvuSpcjz4VMHYQQh/3
FwShPacsfKBVn1ClVYGfdEX6fFx/LqNwyx6xHLAxvRV81QprYI9kyqELXtt0201/
x1jzTe1V6rqa5LSkGeJNx/2w5ON+auC6RG8rNJbElO5q4O/1iK+oFANeIGVYfYkO
z0YWW0IPe4iT8nd8x5j1VcLrKQZamu2zYzu9lZjy3hhBvusq0GMPoO4y3S5biUyl
q6xSkm6UpQIWnqrduGJAzfE0b9ZWSubm4fqrbbY1RvABzaGx6Q5QY2M7ENWx/Y9D
Jum4uL6nUVe+0o+y7KApQRC/CAmPTo2YwW3wRuDdTpUCVo8we7SwPQx7ECeY/yWz
f7qVU4XXV8RDp0twwybCgNT6KOZDHXcRACjPLXD/ZNm1kInSLvb+pCbBfIdJB4eZ
7ijxV/BEI95JBh93fsPY8oDi5KQdmpS7yTkki0nZhouW7ozT9RqtrN6ffQLEQkR0
vrBj3OuTvVP5euBZCoiP8EwSmrcmidEqpqc8bT7kAPELiIhtprsXXIBav7OkVLmv
a5G+vHA1KhmRQuS/rZVQ10Aub1W2mYQfkbO3dZPe7SGu01dRPqr3PK1CyahsK+Ff
X38v6CFpM0EKZY4hRCB/g1tV94i+EHu4KP79erXre5QXH5XKe/Wbxk8wu8Fs10dp
QOQ8CPOXrBqxhgtT0y3Zt7c7o3+1LNskQ0CtwnbcQEQB+XnfrE5/aPGE7ObWNfuJ
xLtoDb1TfQ0utf8pYaeD2nAQAQ1o+0OdLGyCZ11BWTfoDNvxF7Igq2z/Cc4N+gi+
6wIrCnhFCv3GPGp0a4hzRKqoIvmCfDQZq+t5zgYV7hjGDgx2TvNCmrFs1flrbF4u
5bJRfsZcN3NRg4zfL1dl46OeX1f/CSdopP26i3iDPUmPSaje4f0pMGa9tHtW17js
03UzlEeZcDwtmiqFPvWshoQ2aUgP1J2cgzbUr2mj7AD+xJWISDCieHL92ZnkZksn
Mai8zjVGxdZhsVfy6ENK2SgpQ591NiNMKb96FBRO7KMCMGYzWj7C9nG4IjTkvWnN
WaRbk9gX8pHRcnPEwREr9Tfz26gqYWgtZez4siFO3P2r0sSxsjvPQPS110bVHAt5
mTandtJe5weTzs1froPUm6+BI2Ml1gMlYb4ppYj/z36AFJzWmhACoNHaDzCG681M
exRsmGbPjju2nhSrm3G2hcxLYN/Lw6Fw2CppjbJoUQtpCtqO4I+2UzcOedjVh4+t
3EPQj/iuBwpy3NS/ypauxVoY+oAVRp4Jx4wSraEI2CeeGynDNMGgBeE4t6K2Kf49
pZnfk9gyVlMOR4uklsEkscVpJwuou6BpNd5RILbsvzsAQtgn7Abm66nMi9noEUtJ
80yxhYACozGnP0OLdpA8XZ1doa094CHeyNW32X4tIh/taBEEJoqcXmWd4hO5fe/U
1FmOYLNkHVi9DYxoq7j9YYSzBHo4DhIM2eGdCSYZsGM5BDbMqa66s7yursQIR/pw
4S5rz/O8mnmIOft+P2MxZ9BIJ094sfDDNSIpi+onOxr70uKHAafKFjiMZsl75nBy
4pyBBWFv5MgTU3rgp0yPA3/iNjTTaI43i9ZsVsLsMQ+Q31S/KbAzLSo0MowgZYw7
FlB7F7kN9NKrACh0UH9t/eN3SMSqu9JZOJ7k7+1g0MB0RPEZQk40dcdWwGD4DrjV
sneYRAvLdYYb2dSTXgsU/mLqo9C+2rXJszDkOoPe7fNld+l4pXWlxLqC+fap3ajX
6vxktX+wlGYlbgHeHwgOmtzrfIGBfkvGz2kDWO5uIUgWpO8y3yA5OOaDlxvBqOUL
N2krpXf9bvfkxDqa4XMG4Zc0Ix1O/NS+yyYBX6AiFEdSRXkiwQpe2IPspAzqeujh
6BU2ihfCRffJMnbmjug3SB9g/OnZWxSkAF7dcCS9TCT4otRAL4qX3PP89LBXX+7X
wvDPhnOZBLGfVEj7lsBDyadB/arkb7JHGJYzfeG2b/dZjuvSHqVPKXyeb/F4Xn09
Hodg47YsVRGj44NNaKzDiEW22CgJsV9RRaxp8jU6vAYLNqJVX4sFm9EiILpzVaJ7
JMxyV8Gw/YBNG0mnWF1P6GsUwjwktvSK1F/Mv/6ZGddLBcEpQ/tK5xyShPXQ1pXa
Ul8IjofypgTTuMkvToDbV/F541VW95AXpDipBvo/5pEw8U2EqdoOJR1ez4NDJY8F
HAbbHsOdVShwW06tCjL6Y+6xDuVx5j7vxWmV/NofdQ/piiRYnXef4KCbrOt62H+B
+O/xEXAmZdjseUUWiwdSmYZT9MW+TGV3ujnNdTwpGon1KrlRLPSzZHq3+/IYlejc
SwKzSVFgMfwBowHDJRnts3nb9u2xm7bA+3yAGMsbq3abPGzvKsl2dTqI0qQAwYzR
gMYHf1nP3ejfIGfaUhquWkllDva/A+FJI2FHw1QRXgNNJrCLGRY6/tjXZiMURATN
CKl5A8yawYQ8C+R2fDRixNQhyGVA2EQ2KA1quhrE2qQM3ttM1VytMw4Z/XW6IvCZ
h/ACBAo1R3MsRujidRtPF5T5X4lRLyG2JSSDRUawnt7nPQ5hrVllZeUSmMvvGqK7
50tGQ2K77zii2MuTse3grEZB+aaJQwDDlk8w4ON2rYIjZUdi9jCwdmrHOdV4kxEe
2hP1ebBBJOg6iBxRqHxwyI93eR2mjoqpdOVM+pf9HRIExonYM3UiQpnBqYr/N0Qb
R8yBX/9i7FtxhxFPfsaIZwOI1M8N6riz9atO9fjj4SrcxUKqOk3S4zbKNCSWAsBZ
AbDYDPbrpdDKBhtgktVWqVOKoyOV17w095Q0lAXYI1SVYRsFBtIv6gMYtv6IsK5U
+z1S73zBnumKwKMBykVSlUzrZHjVyySCOSm1V01Aubd7cFDAacqYNcFzVNz+xMMy
ftRQYut0sbv0ReInvUkNtwxAjn1cOd7dS+0jpgOO5xgImkTcOwCKmiOe0pw8+x3W
jz+fUAYAmhbPuG3ZqMvDMyMNBX2ZKxnumPojKAqoSxulkvmQIMFAIJCmcn04e2Cs
qxlNr9zAdPaIEK/gG2WTAqWx5NBUBzQ5Ovq42a1BRJtJEEtb3hAZEnjI7lbVNr8H
iT2J8iWMyCFCFOmBnAcM8XuxxIY3dNvrbfpI8QKSBnov1X4ffLNj0VY3CnCrS4PH
lGCCxByE1CfvOcCiSCxURbZHUbX1rcQkwsLZcr815t3o179NOlZ3RyG0wmnbrJum
+VDz/gfBDZfWPAdnXS0ksbZBTeOyopmUXlpJv75CZTQnK1b0wJy1EKgDHs12jOxP
DhIDJ3EL6RbAQwnDOCSJ0PSAODxxKHE8sw5QdMzsZALxXPd2jEI4oQiBJFQtOGde
3G5G15ze2vNsKW3jwO988cuF3lBl9Wajs6eBVY/Gfdfuf/XwIvQZO+z1DWE4aet9
q85X38DazO5sNErzR6jx6Rtb3jwtaLljcemBqD8kN/odC1aK6SeUhWs1su5jOGs1
nMjNK3QjSSz08wzMS/FI+L3b5K0aIoyMTQ8zM7S5IwJ926pck8kdO4tV6RNpk2L3
gRuJr5rkVFzFpRRTdYQxWYOYUVLEZg3KU0Rfx/OIWewI9n6pL24VX9ICTxk3qy29
eo4zFOD/V5qwU47c/RNBBt0EWI0mgfUSsk3dXqtDTUNj+Vf0iil+0Lrksf37oPMH
HpZ97LK+xZBvhKfDGUU0COV6b97l3XuaGpo3sihnX1gIsfqm74YYDoN2UWxhfGX3
YHU3uwkAWevZk2zJY5hLAVG0KRVdHQvRaNxbYR8uZ+9JwQeq3hHALmCNmb8cYyio
BobWAj+hdIV+mA4xSLEun0nWd0OikYuS2fZfJ/cliCIP0IG3HIvRtFauLICSOl/0
LKjcxl/VOJtmCNVTLmaTLMU8f7s4glDLfYpwYhvCdq9fDbJu8lC+YkIywCUFlcJe
qVQGXiPSm/BD8fjTdPMGrSV3lYAl63M8J6NMAe7Bhe9PUHxORTeXoCf1ekd7Szwn
TU1D0fvGEvESzGwmvIXQVyHlNaombG5VzLrymxOM+bB4a1b7E1QQAJRJHTb5/gi1
6sWX1zMYdRSHlkAGJqQgvKGrst6J0bczTJEMfNQaKGXU7hDVJS/8+ppNwYphaaYG
KYCdDZZPvld0zxClVO+C3q0qsJASVakfChxiyctcOY9wV8mjfo5WNpJiBxWzVd6S
7lTq7hpBAkTl9ZN6NJsOwEF8MJZ8usa0lTOIaEAcYsAV2jaFfBN9FwUswetXpqBo
54CSQZ93va8XLe3//3oIKgjSN1zzpQd33IeoIa9u95fMMUcxiKHLB2Ln5KAw2Hy3
sCOt+5Zys4CXdA3e/F3yrMFhTdsbgpxwlHp93YDJ0mu6yQZwm9TwpvJwi0cHxJWU
13cJLybF7WU0rk2fc54KopYf9a4zvEWi9031aw7YkxpORo2XMSvw4g2lPaY9QoZe
Eevd6nu1QMe/V8pN4qjdVZL6s6SK4lPUY2Lr+vr57AQINp9RiEJgEgCc5H9zyw8H
0ectNWOj2zhTHKPqLnNFPu+c4XBzC4vGqI9bs+01MkCtQBsH2YmImQAGyTkWpNFn
Zv3WsEa+FKDbnVvt6BdBKOX600G8b3TTzbQtpOH0TwDZOplwhAkgbKfFq96zaBL0
lrK9clV9V7XpYGoOlrslbcU/WXVxUgA8PhMrmUHOrQkXivr+w4wXmeg6Q6Aqd+CZ
kTp6rHkxqLe6XKP7SjrlR7YTpwrDFQFLSh8mebp2AswbYVDHHZ77mMBeDbIuheZs
vmzelRkfbopoOX77pIuu8R63Ukgg9jsAEMQJKalYb3HZ21XojlGBqwqxLadEMH1t
QnNtKgRH0fLGqgXlvQaEGABzB3N+RBlzdShP/7TVBhRnHa1fliDYa1krXDNepbuW
AejAT7LOlAa7rZHzMEVggvzuzBLLdhRhWmLad1BhfyDysqzst70n6KXJo48sKjar
9koYp582Z8Fwk5oNTQ9ldq5tPvQaOcBldDJd+xKB8+f0rN3lI0WMMVh3gg5GipvI
6gs5EqCsvD4tnqfIAM9Vg20YNHiwGYHnYMia/4N34rjpH/BUDk1hMRPVy0OTUMsz
CJ+X1sdJ3NjndFw6uGQp2yeCnHw14FXqCsd05/i0oo5UoVxeQuO8gDZ+tjkDDccA
/Nd7hkcoN81V/gqhqyXvc6Km8Hrjugm3AdMtrQBhySIQ4r+QYdJOyAhekYi997gS
SiMC8btutosyss9X8WiqRAw/DyFuO5a/dDovZWwqn+Ezvu1UdrnrEMmiRhMOQgDP
7CwLwHg8Nw7Jg26Al6Qp8FK92OJCXV8/RkmX9tAflTGbYjUvOi2CKc0ttdcwNyJ9
XqkbzKDc8fMK9BI99hUiraIICv4CztRwohiPqPZW72VDxb+RSjjRRIskOJCgKTdj
FzflicqlmlhTHkaD0Xwi8n+hWgkdO9JHTbTG82PueCAvUsPJQHGSwhW32AgCVMsN
zYOiD9qZ2ccwr8acTC2+1HkgXmNi+F/uZdwtJFPbjsKrPgm4OhjEru/dYkFjlblF
6g8EphUg9gIF8Az/p1ZlfPl3WTiAKGZz43CJgTXY7EAwiWet+HT8ZPnMP5FqMaAl
GIuV2c5VPI8wGT8BMYAN3mTnLnQ23CgD8/99VHiQSuzcbyNuoyjfO52HfW3yZwoF
5LmKagNVDDhzVlX+G7ZsghB9+J1dzKPGnjtVpDJaQ9Hc4gNiV9W5n5VgFaPZrzYJ
F/fKbBRVN/eTV2NiASPo5z6kutjLAOS2z33qr1c2pf4P1+g4K27ceTabP+Px5AkG
IC1UCDA/KuM7eP3wphJvtlkNjtjbdPKvT8+Ef0OdwC8LEtMxI7vQdkAt+Eeg184g
Gr1Fn0XE5btAhGu8XjxsipsksQ5EswWHTE2ArBObAQJjBMKFbgvCweKv2s1Js6fq
cWmgq/xX1T+h3g+xsdMwlca1cP0NFx1DA/NDqiiHZsx4ZxA5K3+ZqawmgQpAdp5/
eKKMRnLEB1esxbE0AgBDEqGHpvx/bEnguGgqqI2c5jqNOjAFGvlLlaaBYDIPo2q3
hmKpQlZrCjaAjfQSKUBkSFlLKViqn4vz0thYQ0OfonRCu0aXsiyS6hQPP892xQgd
nncggW1tBBbP6mLTvEjk1oie5MhRSanRVYfm50cedGCI2fg5oYUb2Gi68QO/D3v2
YwYhy2E0ODhXsm9DE80Mty4Z29JoIryHtNH2qkvJXe5nqE8BVmAMI5XVol1jXwuX
9bW+0zkN6FH5s9mBSom+uVVwXfNmJYubbTVuVox8g2lxAA+AOxbXAWx5EBYoGfR7
pBoIG3eD5NuvRqPXX/j/fLLlVr3z2SZ+QZ84Hae3AVtIuKcd4HcC3YDPD27civb7
uDSEUhSPlngsKaJfRmIvhIrmtTuNarAIjzmyiRsohksCzf/e03yYE0YqBTDSPary
zcE0mVklTiuocrIPTsIxtBEK7Zwu+KlgO3UQejy5EjqQJBI7S01jc85rbfdrzrw1
d2JDTF6fjmAZ5Sk5mw/BKIADJtNrMqgyCZbQ+wn9PW0+cIygkKchCcQOn+i367yl
yPQ9ewpdiisCWP0ewirk9fgL4HDhuwjZ6jagmPdr74V/K8k+/g5I6oJXhcbE1jGU
uls6dFo5WIp5WbtrBqdAAezXLY2ajxSWdXmfzm7Lo27KKZeXAzqmIrfVwkXE5+NC
sXHejw+6OXoZiJQMDIl2U2q2ZLsQSQbPNcVLcscQS4REYWsASkmrdKwxdbZks11E
wQm4rUiVSPzzuvFeELiIUmHLOtp6pWG9oSJu1FDhzEPwJ9hHoyj1XoiDDqAYDjA9
Q2H8Di8i6B6zbb6Y6zzNF13dIi48y5CpDqLmBTPJYz2LGn1N56opXeHBo/jG1NnA
i17JG/1QEFUQvNgZrv2yBHFY69dk+dHEMGBmlzhQztijM4J0XmVnmDInPJIubbtd
+QjWURDkMzCGOHLQmbspUHeVCdOi77SG70v5rsf4Rr6qFrCQHcGDQeB1mrnCOukR
gDzvPb3Hb5nwIbUIo9szj/4mvy2PZUNm3VvKtva3a3vH2dSeifUpGdTduRVPkjnU
S8k0Gt7LxsWosZEW5tGPjBfCb2D4da4LScFRUopxW22iouY8qdf0YdWgt0Mu3s1v
A3C5hjXcvgrZaqXrb8KTrCO1ZigGq4bORrVnag3wUFmOYpwl4CX5rstRNfxW+Hr/
tmPdShMkFGvPf0xuirDTnMs/sW2noS5IXPJVkWKrsICiHDrxZqKTKaE/7tmul7Xp
MGGBjQ11RHRg+VE+Ldh6QwaKqxIYK0X7OllFxi50YMm6CQRDBiskTiToy1+RQWnY
cRi7K29Z81G8zOSZVmrwkPCAR/Gydviis+GD0G+qll6OhrItz4iBC/XeYS96zz43
Z9xjijPztahVxTSleZs6H1e3o0KGajCSCDu5SM/cXl/XbGxhmtjvQ3lKbEG8H9tG
TytH86kU6oS90JnSnQA1xW+kewrf1/c/tK1V4e6d3k34908CF9lJOx3/RK1OF1r6
2gaRQtEq17OSjGNJML2BAHagYnxtRrdFegryVVtLF/vdicdCMtC103jR9p2JjgJa
vK326F/EmGnaNP52eoYzvfLYF8CASsjTkTzYVzdE3vhJDzjpY4RDjG0MfWzipze8
LFBIBsmFw0TzyjabWTebsMSCP0ayCuZKROGEPIGJ7OZmu8qmhuXpuU6o3xqKzMBS
2vglgab4JcAZdDsrO8e+vslRDcEKMPUiEw0mTbj/lTBCOjzwHhuLrzDdQKPhbtYc
PGJUgtHPtaOp3GIfUKYQa5+tMP4F1nRZ9I9KlmQCvL1WCCJiuQ4TP9pWXW2J/+Wn
wPQo3NR+WfBbH17bUqVwNuE07uN1b2/woBnpF2/GjIYN9Pi1xInp2Xs4cphmGeuW
34y6tXSgWNXAjRBEzxGnuqfUj3ZYHcZkiqla21D9U26+xvvZ23bYaI3FdIwEzRYs
NlxoAW+2Kwcajm97OKAR3aZN5zg30VqsPTevUqQP91+SYD0txm/0Z6lQ3B7BhLzK
CAfuqGTP4nD+XYe8SeKkLXK6NHaCcPAqg6QN2rvBesfxS7gKYJE5pPziuwDZ4RBT
PrRT6MHrC+0U2zhErIRpDjKWX4IHAnK6QkrJlFlah8smtXjogBsNQLjXjOnffriq
XsImnMuAaUQxLT2s5AMxdP/qzaM+rs0LiHIWsYhtGKnniC4aczidmhfZvB1XTRuB
ANsQheT+aoRilk3kFebsfqwlIgl+GxODi5EEnnVnu/5Qblrbo0f3vC/pXHmB2RFf
q8PLdwMp03q25y0TFdc3zujCGBZ4m1QbSZZKlBWiZ5C+2FD5i93LfCPUSSZmo6xY
2LJ4CgdQsJyZMbeDfQ9EO0rYWOvsrQFfKPn94JsOfysgAvW5u8TeDga1z4u5yGnB
iD24yKXWUnAVH91UpdA2OFqATdyt966+jU22REOFvOZJft9rTijybLV6fxjJj2CQ
9cQIgA4KadfQFMvJZSR6UAxuxPuJ+J+eIhD7fPiwx/Qzv/X+eyH00cyZaDYg9uHh
uxUfC2RhTiZGRaaOpT9qi/hNyUtydXZIyXal3Cll0GZeQ33s6a7YBU9n+s5bakU6
1zUwAobrfD2Eqiat5rSZcfIpEpQsjFDMKyNwh86aGX/Ob3qne/7VOgD7rp80mKkz
tEjYMtUSBHthzvDuHAiDKZhliXdU05SxSAHgt1MbMhifU/CdO3/GSqMMPu9cDPwE
8YuvU+WzUqyo2Wjn3f1cvwEkYBFJDPvcwnT3sfUI3EXarvXRYf93imq8qqnXJnGk
6W6sxILEiXDQ+t8uEcAFJRRcvOM8ElsiStkeWsRAEXssrZd04zYnx3dSRyFNdE23
fXC5t5gRl1Ysep/Z8oLO5T5tlkKFze+OZRAW1K4MFqIR9EGxIW2kplIaDrxY0s0j
R2IuHALWaI722dUodtYGD1OUkxVyRz/jUO1nSm6N4t/Qb+APfq8FYeqTzJh330wg
cmelXT79Ba72J4sefKHufIPcIYg5iGzxr44phkr2j/HQQ0XfIZqBkq8ZshzHYfO0
PuNsLpnqk8qg+eDY5ZZsKWzKxqoRLvWj9Wup5aD9v52RUcdL9XavZV2w/EV+9rdJ
1mCwK1CECV9jTeviWHupOgrjdaLn/Dfj6sSeEVZcHH9bdQrS5bQRFuHSI9H+i/fG
Ps85XN16kBLBp66PklLl51GrFW/4CHprtgN1nmGyFhOigHyW/pe3KN0Mvrlg+fqu
KOxbfoMi3qXzrbPEqkvDOy5QnzwCBNMfQ0HLfbAQxA3ZhCzryMaZaHgQzVhZvOvm
4eC2YVnWWYyMlqYnazL2iG7F4lRN7ooyz4A9azrXSmqlrHw2cpzlHqxPolfeyYL5
bFAGstIGRqLK4bhLzaJ9mxX39ZoAx8O4vsjzyoFvyl9Uw2KXcFCanDasmOzXyD0K
40OKX8g9n9xc9fB2Q0XOTiL0PYYorPScIw/DmagGVE0NA9rN6VWhlOZZhraa/NWa
ojaFN3+7T/8ER92mhK3hYVdsCsRXl8hkXZaZ/6wnVidBlQnrqkqPN6oNmp3tsJpI
2oAV19GqfK/FAGxYdfk2zeRLcxoGmiAh2U4OWyves77c8Ikl0LYeff86odH3H35a
EPVeShnN9nHlHbyKM/jtwx27iJ0/glHe0KC8rjlA0IFMrHAWjRbYSkyeaubziuwu
Vs0SWLCSwp8iMpfKkMSE9Zq3VfodD7tJ39TRI2m5J0yNk7zzB++obM3z8gUmeraR
G5m5XX8YOx5Ym1q4eY8xjoDryyEN1tf9Yp0T3Ad1r3ViKtdXEjrEpEj0dGsL9zp3
0FCy/2B4yT4oo3RyrVGKcM6ifq9/skZ3V6i7XELhuN/y0gmn/GhES0ouyT8HiLLx
rT2clBCZgiTwSJQvq8Kzl9wUOwsR+ZT7sYY7KmSdwUdDGd0E0T3sKT3AL/A9sWG7
xr7ddFG8cjLjReOZ08rtC3euO3zxW7/SHXa++nKO+7F737yrZp7ElfRORyWYx21G
7NCKTB2N42T2onsAZuYGZLTpEDvkTOqI2HdKBV04iPvi2V7246PlWa0MhCVBPhRF
EptSxk4RITlY2MqBC1Y1OMly+157x/SU+lVRy/p2G56He44mL3iEuWECeN8MpuF0
BQr8b0E9sh/pAvooEvwfw0HtHTgRameYIiQqCFUoIUIZbETzheISX1opK6lp5Mbd
9j03W3//4/k/mCJJDtQyYqYIhG/xKU1azxK4mRoQMHaw5oKChsWbee5pWLn8P/lF
wZuuQqQS5z5yIAPuNUgJSfIEvcJKPdu0Y9wXeNaQwVrozcg/Un6piZXIVBwO1I2v
g2C5AXQzN4S8/ulc+S/G9R1AAuIsXNBMzCtoB3mn0a0FRrlTzjmj9uMqsnqAsjJ9
LzAxD9P5ChCrtVH+DHFPQsanLmnftxo2c5FMJUs7stoFzTbTcly3rFONZn9stoLW
UMd4+2MK5e8orTkC5dp4Kpa8+OC5hyC8jInLyA2aLIRe3F6lfOp71nLMvF8q2roe
PpHYr3wlRuVbja0S8eMXxX8Jep2yLFpHX5Nw+DxfbF/oEt5wQM5FUreKyhBHIyg8
N7620xqrn0P0w+d83AJTIYns32bD0srjjEPK8vJPQRW3fhGHq79gavuukwuhm5wF
cbY1Lnfwdzhcn37afUUjiqHMyR/ipdcb7a6Q+6yo/hgDyWWYDquP1d/rXxs1/4QM
7y8UHbDwZiulsHvZitBSLDnpMWwlm9sFMnD+OBHR7VL3UWCqU0mBHCTo0zmUWwdW
f2GiAC4ZRMKZU07OiyPZOl7wpqePwlqIxGOqX3MxAzOw5kD0NjN7H/Hnhip3xxMT
JaBNTai1csb9joaIvjS/LGVXVSZGv6feACJLBfRTTMHhhAoaV1lDsY3+IJ35XA9/
TXBkEKqX9PFDGLKuJ8Y3DWw79r8zj6SgZzuZaRMWPEaR1tci8CrBrdyJvqYrQnsQ
q3nj1t3dpS23KbMvpTzQF1Z43ouvzdYop3sw1aZzuIIPdTfT9EkHirT2CklOp7SB
iRc9dJNwNEIBoHU7pgsiWd1CzWdjnOsa0mkx+9ODaTHIRycwXWllPuIjUarpFlgt
/KN3nTvtEd97j3WDCyJ9JQviKnfWS4KtCvxw5HmMoA5qNGR75eX6+RkoxwZmRWYj
X8qCggEJV8mWx9qhfMYLssTzWA2WUodEgvKVIKES14UJaDuFSNkYduMIykxzYIGs
e6EZ2gKGfS6w+ZGVlD/GQlkylLdLt4eoCJ7e8MpGeoI+qZ2ZdDHffG3M5JhfSxTz
AHfEOfzm7EDb+jSbsPtgcqumx/io3JfDndv3x5G2mmXCtLGmEkke0tq7WW2dRnvH
acbyqVyhCrgqt4iDXuTC0tcAhsR2gjnOAXLOyFisV9blleI8tLvn64yJTndlGqGd
Ces8SRn9Bo+/ve0gZzBeYohITr3BGXLyAiU6h6pArO5eSAWeg8KuxsmI+8zIBRhM
u1JC9P/IubU1rUj8+NTGbiyHCYUZRUL6i0ppi37Fd1YlqvwK7ipOyNa+U47kgKKR
qwPYWQh+AGTYUadT+6qjp4l/PlgtXcuZRLMBNRSTrfez1HPEH43W+LgJZ+5a98AD
oD3RikDj4rt8irNLw6G///8OnTQi6VNsyUlSYEY1T/BwCO6nGWAatF6dMNaSNeSp
dtNE0wEvwgis3UcfeZcbPW4xYk5FM2xzJf+C1tP4NKkvHy7V025nv3q/r6PqjEUI
k5su+yBE80GCPFCMg1F+FJVDTJzYJq+37hqOGn0hXIixAyMK7Gg7nPulxlpP6IYv
FVe0TJLraqaf8nMLTk+nSSNjXUGULxFxc4Uh3+5aSmi9RyKoTnl7j6dGhqrzhtND
4d4+4jWHcSGuklmI+gsVMiikhl5aHDgXRvKXUii4BD6DpCdDVbEf9a5NX0yibNas
zv/HJihw9v8WDDk0A/nlTvzzxMYDeoh6sIj0mfRN9pICdxucN9A3U0lONBFF01ei
x5hUIh0+nLe3i+ytE3xrW8i+lBBKrumxrGZlC1PTqhH/jiyMllOGRgg3gXAphCRg
cl3Xsq3rdkwPCpwXD5IkAHkhCJGiKqoex/Z7zRO+NhFJCLTzcZlCKM27UcsYka+u
cUgYx7i65blwJTl55rusNdRVLS/bi17S2oCYKvC4EUfUklFTbjswRkHUdxVO3wnz
ATHupiHJxR+/zLDUtOAUhdmV8hoJ8TmUm6wlQgDrxoNq/0iya7IXrCkbGWw0o7L9
vE0vzOarJGF9wmbZWYLoSC7ziVQDyVQEcfhRjka8A81lDLHGegyXkbNdqT4dntMG
4SEwXYeWZ9uCbCEouwiA53+Wq9nQ8Ly3ZmY88pfdz0oOdl6n/VdgtYfuarl/EGyE
v3MW7GxiZdL/6zN49YeX1EdjMi0wkM8eefBC9mqlh0g3HCvfMb0hoPp7EByFwIwM
1MWsDVLuCWedAEviMlx8Tz+xydsAyJzXInun7WqJ5S+Wi1DSyRVsp3K/+OGmDn7a
ZtC7dRBrZjjV9QtlJeSYS/c5YKXmWnIi2Fn/bSGLQLMXDUueILZBQ01B8HXiL6zh
CY/GAH7ZYFWFnoDS/V8Qd7uFN6XWhdeKnM3noNl5wCcCJt1YTnSXb0n9BWaWs10p
`pragma protect end_protected
