`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qcguZKqgSNLIxpzVBvWQ/uy3ekCzPXejDizKAk1M+s9AX3TdjIVUi3OEuBZ+yN6h
Gjl0UHGmdaDhqZgmVwEkO6LKSacVB01rq5gWPR+EPtHJHXa3HruAubXKYQv/aGRq
k7MUUWNICzmV42r2HgWAZSWlb+A+y12DigHul0qVyyY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4784)
pxZbLdomvBZRO/aWLkBH3jZUZCOSnNCxWo1+VN4UXE7IOHpwZpdIL9jdM3zlltDr
RwZ0uTuYSNkQDaAm/bE9RosBlsAX1ufWqHnGv0kuLWA8R7KsCKttmjVWQ+kVwpgo
vJHz5oncXg1sYK+sq41cy4C0bhCD/Bi5cjdksKpetmrz7GxTDBpLsX9NBLQoVt6D
GYOyb4eDQRld/mL+oDS4BplYaXZg+I5G98HxxrugQDxy5qN77S428nz7+s1mTaOV
eCUC2HrE7UzjctgDKP1RvIm9zFAlpCG4x356x2K/odzvECkD8MaGVkA8ruktisp0
JAGLJIvn6h/pjukQxGNa33F/mZMSKVAAQqMIrsNhJNLO2V3hx1/BU7rh3ZwLnRWc
+hbtIceqoJJLjTu4N642un/DD5iY8NLNVQIyFdPBgDMBaTQlzecrn71nd9RQXpzo
lsCINFkhZjXlOND/2J95YldQgyMMvb40jnq42ZSGlQfqoPdFH8oDSjMRN7yNt0no
v7sdB7dQgjUoNz9vP6nHHknvvg9jVCAmQbC0VfdqwEstCBzdXAPP0iZyxEbwOiXx
ejLeMtzE2Q4a7KCnYX47OYPHHkzz5kXF8FCQIcgr96jH3z/ttYlanOoreuKM7OUi
HA5JZ6WBiMmHBbcDuo56n6U6Ydd0ruaf7FRtcGy6R/1mNmJtnsfasPvRvldww2M0
arBMDo1pBx6tSor/EgV3sJFEf3JInVomleHDOxDQuI23tywhWFFv1J6v0k/ro6iR
k8FxhOSUOWDf6jgfmSGhsJHBeRwmnvksvrvNMVYAn+/4/6jHNzaHo6GuCS24WyqX
TYqsvtuKJLtqF88vTSRPBshsjrleTwnDojlHjabh6+Vgic9RXA22whpU4Zl+XL1S
OV9nTNaBgOiQHS4w5EiVwVHJ5gxytg4pv0JQLR2QLMdwX8QjnsO67vz6hDlRX7BU
HjCihIiu0+eGfBfYDeVhNhSGBpiqy5wydNNVvTGGiOv8r18tWN9QLH5Qnv/GaQ4+
/LPmc0iG+FlZPWI11GbayiByodjgLjqaV3wyWWAUM9ZGf6oq3hAtG2XZpNzPejQz
V9OLYSuQIAATQgQPF4Z3CvWllsuCIvv7eI0vc4JTPgzkNyXltyDIEFzVBRlsHx+x
/2SjWADADtzWEUUdK9XUHPjQsLaZ4/XL4L7SLYyIt5tOSkUwG76gtNLtDVtTvjfk
ohXND0Sq4EYNiHErS8Ampl0BmOSWKI+YwJq6UKPU9YPY107u2Xe8CfIQj897Aszs
tk3XXdicTgFhRYI6pAvAjSwwy1XO2hKoi8o/azNku4OgegVsO/Gx46hbHUgwujRN
yWx9yU/4PAQIEne/trVYgF6JSSWtlSxONdz5cSfjfIy9GYFKzz0zqk6woj3e8mzk
6c1Zzi/6DD31l/rWMkKxQGQadoiBX6cuNABbDcm9oaIqY6BfBrlxU6LUNEwIdgZ7
KUqbCgNuBAeLHKeVNjv1Kq9ioY+pwiv2CCGFxygB+Ycs7bJQnjZeBU/FvrQmwEHW
K5JVeLmCc4Bij3G1sMudkez8AouQfvl47BtuO7FilJ9VZnjTHRZU1jWr4AzWQIvD
YRu830ghfbEU6eQAILhdPaUIIoUsNinzuf+iajrC9q/+hm6TNqdKyFgSEIDrsSha
Trmgl+4wrAKbjdO31QOCg+jpz4wR/9J+itzWNsdkMy7pyuZQoWzydK7x7GY8ECp1
ca3CRQfxCufpqw47L9qBgpXPQ/6yU+q9CHrAwYiwlUjJHpq0n0W9fz5EMgoUaJA8
3e+4keaWuWFW37nr8jAOU1ONTX4wBTViaiCIbIY0xkcw3P24c5nN78WMOap+BcQH
ULSSPNRebR6K0VIgJ4iRJ1Oq8yP0dqE7IokkLFAlyG2hNleQE5/2G3jUEHpV4W8N
WElJXd4Y/GaMbkppTy625tV/v9yPxJkA4CGkFIpdGCSh25ecx21BaI4HBeMZb9E9
X8n5SKOSNfUMVPyG2PvN1P+NLP6Tdp10WtXatogJCZ4xb8GnyDSZL1c3nvNpkmMk
AtE5nQYy+542z5F7Qf/ln0gjyuXp+B6chm+4Bc7tYKXAbehwOs0aXT6WkoqCM7Yr
uYL47cvd4GgSixSdY9O5GCqHY//AeFZ85gLbbIuTETieX5uLlxhg3OlLL+o2YIgD
aVSeP5ycbRELcpm+zJXXMmG1HlKG5ReHSp+5vK3vTvZIQdmlUK5Vh3sRRzVJ1DMX
I5HJk60uhVUNCNmfIXsgpyQH8lB7KFI5X/6TeH6wFx1QaUAFgL0UOsxBnSjzzuID
r+VNZju6vdNiaSoMqKmFDCcoN5JhBztU0zGvNBUkSC4wip8Q3s4i5M1hsei6WiLs
BFF1x6C7M6mV55TlbmgTNXO70A+tKk1Nb5vqAe1HGutKQiOmeO/qndi/tJ7zmcsW
6JxgyaXKVq1IjPEbwMxqBzETakb6SColEM6L3I1hIrIZhK40R4Wbe8mk60x2Iw7Y
6butcM4iTLD7tq8bi/C1UGz7vnDWxL0wwnZN9JlNFX+SsAbM2BmM/Iyx4WkOsISg
GhoPPfVzpbCEDVrX0F/cZtaTnTtxLvfEHSBfRLdSlaRq9KtMYRldoc3+rJ7/eSCm
4uVWyvnOEQUGL62YbKNCDvhV6z2+HVPKlk8vpsDJy6S9HW1OkHN2qggDypAg916w
TmWXeNUuEcW4tMKoCVpNIf+mcHP6SLtNgStMNFonKj0R25mwGhfNK8DCjLAo/8fl
vQmVi9IcxNp/rgtv0xS7mRl9gimSsNLK0mHG+2VM9lMtPBE/5TiNYyWzDjK4zsni
ZwpPp24Sv7W4Dw2toyUTzbl6EPMgpznHkWcjLKZ21G5B38AFTzlIhd1PzQILIIGk
kashj/yLZZlCFZeuTAXlAXcwUIbzPGRFepyZMiynTfJRsIxk3VYm8AB5rLCAB4Aw
QDNA96f83tEAqllb0A31S/l/tft49O/Hgf1//ekrK0VBhgDupcdgEcV8FTHTaDiU
IhGH6ZsPCT/FJSX7eVhsQF7o+8MXbq6AnTfF4DBh8DsKZlCEhE6saahcV13W2m22
ZI+b4xlJ6PaPrHXVGeo1BTv9FT0A+/fPPCFxUpAVOBVIx7FEyUj6c+DcPfhb+7dp
rWfmUF5CSAb0+UCpe/q9O0n/MzQhp6TnddMTPjm+alVppFp1YH1Aw9NxEsaH76Iy
6S2Pb3JxcHyp88C0W21FzshAx0ZaBTucCdMnxKD937MH+CzbTYWq06BiDCl9xENG
WlEzSNFiQcky0v9Eu3mgYQKGt8iPrTZA9kh3GgyxtfxKWNtrdX7KI4ChP4nTOvI/
YU7wbE/57dBm//a/BntXmiPpmJalABnAFugIhgRsKfPw3PlLlu4nxHsj8osff/w1
P45TVGv77dtNHQylSMJ1lgm+CjvLAFW0tZlJnUnTNtxTt8YpM4feEYzbTGQwBj6q
WS20jE+7+qnueK+9rgYnfHMOX8g4vmoS8Z7+ixeyMijpQKzeifugmDrzYZriXOGO
YpCK8Q8FuMFdW8gjnq5YWXdsZi/7MyVXXwyNXfIaHhUA8gbDhWnR54j/o5L7Rq/Z
bEMUovVumMFqiUe+QdaAq2u2W78+KXFJoHE676sxmbnvxT8EnjV0EuPJT+uWMuXK
S8jvDaTkC0CJDlq0SBoZ+DTD0TsI0XpiCR9Pf7rD5j9dDo5aZYv904yJYfRIKqd6
G3JC7sxSHJRiaj30jXWig7/bnnB9HNFOD/ZSgxHr/GY1Fnitxo2FW+R7HyrKFp6f
yuSf2EVlDnXbrZoWyp/BUGZQfRdTLPYxvV7Ztv+z491WFtxAFqoEsCX9wHZu4MO0
FMkA7XAznQwR7C8PCNd2x6KXJOiNwTmr+H2TTUzymrwFeq4q83H2mmYv3QS3Stpm
kNL2xbNMxGAQYDAZCdcrz5pG+pusnPlj+DjsttC3KPkhNq1B4308kDjwQlbieKiJ
/CJOk9VTTOrHvyMpuVqgPzXZEYLIpSje/S3qUIq19aWW4RIXq8NT7WczsbdGe/ei
egZ5HTp0ily64gf/u4YuEj0edu1b4YN0V2aVXCDpSOF12j5GvVDuEKuIrtkQbix2
r3oyqQrZitH/y94wQpI3fu+5YATUgOuAwqbOkIrbSTAl1jIiqUgF3YUr3fD3Emij
dsd64Fp0o+4pIELg7nYfXItSCpAkvpjDPyQEaap/t1BNEOhUfyDq+jyeOtC9jHq1
BtWdE0vMk7FfUmUQ6OkusCKh9gt6i35HPrKpV1QXQBHoJFBJReLgWWREIuyasJqh
ndItYBAUucT6QFQVGpFXIgkHfB2okaN8hLmJOlhewO8v2rK6K7ARKUPcNkCSt4XA
cHRYk8tB81bbmuGECRE189iU+u9BnADFbAmHDaZ6G7tSB6m6cGReF+4VDx2IR2oJ
QtQ40LxRrGmok1OnXPmyQwmZF5m0Xjv03Fx2L7EBjzwKSyhR4uVisBQvCnd3iudD
UdIrrQU3ZYT0b0Pv+MRfz7uMVOVs/xidlUAWnfNNCNrKt5M8dgeHArrCMjBs4GMN
ocBrzoJmp6+Mb7g/ZHd1TSPQIMFmzV9hTPwJuELdusfNNVgubAmdeSf63YyZB9Pk
GfLw1F0VMK/TwALmqVVIIasdG+ivAdqvonSXEMp5t8TV7jq6M1w6wdWtfMrG2Y3f
fv6+YRNOnF/OBdFu/CVCgGsia+20Jwj2cmJUXx8JdAG2VhzQbVqvdNl9eDg0a/59
1h+ZgiW9WyVIn0AU8FEV3TRKIZo3A7o8VJEQIuWtqNUKfTAp5I7Miw4LGR3PSTyH
16JntqipaB5h70lDzTxqR4NIDjto+Au80CDu9LG4BA3EhQ8dnSK8GtPkYy9B6hLg
UGGLeqgKrZRlkfWkwgC3UnzaHua0OY6ADd3AS8PBWGgXncSW8K8ELG4lcWsZV4IA
CRbLCrhWG811wQNfn6I/1L2+AF8Yw6Z7g4ybV2QhM8b1nrUyjWsl41bkCfqKYYlp
w9y19AHlyUBLHAwpjgfAJkDsbpN/B6U+IFkV4r2k6/Bz/i484BIEFAYFGduHx/dm
gb5vD3qRNEqjkMMNq2jV/dvtCwLd+WItmfYP35wpD2MZNmR4aEjMUWrVd+DmTqNP
1qDjUIoI3YzwzcY56mOu1E7eZ08PH92OFRt4QZpAOPJaR/o/27FnKP6zKRB3wvf2
mxt3+boOI3ne/OP53B04QdmXeBv0Zl+gxpQnzPQwJ8av0Kbcosc1qQ0FKG1Mj7Hc
pxzwo84smv5Vqg4v5w3zcDWcpVxT9qpA2Djstc5WUN7ER0O9KYj7bvIZh2meeS/o
AAwALPqRZQbNPbbDwy4iCrLB+cOJ52hDc5QfrcniCo+FFL8ZJ7RzMKVFsyUw6KZR
sK7BN+YdEugZo/yekkGqNSu1qt4K/F0d7UedLZJXU2fbPe5syh5F054Xny4Mt1bC
sXA3d0wE2fpsenOP+NRDHT4T9ZUsTjQ8iJnl53UfO10UXo6fVNM1Tl82Usk7vW3K
zdvhFpe2hiGbwYMHvPjKJhnn0GkaZLdQ7YPS53QrF0/WPR6CGBD98gR8ZhCWDGjZ
+mrM5b8F+9kjIr52ZaxxhZdOfL4dYLXEdcPGJUyAG+oYT0HDi6J2ljDKGsWzzUjx
IWq1VjEh6pJ9ebPQdUqIdCM9Bt1ElKfL0syflhUP1zEUJ0B/QbmpoHunGlhtZlnp
O1rQr1uLYV4i7W0yNvyTFFu5CTgTGFzeFy6ydqlw/wwXjF2pyc2tQWvyWSUYdu+0
7npD8TXp0FpcMQsWbMR7aPpFHV9oGQaGKHXJRFojo0YlnLphPDOM2ZSqMcUgA9Yn
H8aYqPhVMMZ6M10ENHccP1izPnhudILmEAWr0dJQD/PIIaH//Lo2xG0qwGwnM8zl
EFZozzKLomxQ8l6gYO4K86GIRdxVpgS6eO7w9Xeg3tkO6M9M5uDkoy5wzKbDmOia
Y6Rr+Oao2IRO1pneDky83u6qP4AkfInSSVizc5gUN3UnLcE1MBjifqlii25oWqkv
IWcj84SWWYaEqy1zDDd796787eadqu3GpDvJs81W5vBDiq7J95SPIGt1WTHkflld
nqV6Es/+2/Y7D/KBAix2kzINzpdVEe6w3dIjGafmRoAR4x6XAS9lfVZVNHygM7j8
wWDTQOQQb+zt7PvY57ihJHv8WOEkUmVkAEhTYmqRqglvN7SfkKqCaCbq6JDqut56
PY6BiG6BFyr2I2o0YihrmgVx9JqBRWGN2Jex2d6gjo4R542AaL+Bw1eM3tkmcHL2
c6RDrVAQXbz6EpL3AUBx+JheC9OUgMfWI0kzGS7bXRYmrWMcV7gODglKQf9F2N1M
YIx4e+pGOOwOSEA1lStR4XMYkTr0T55aBsyEsG0EEH4=
`pragma protect end_protected
