`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l/TES3OShwy4kCeeKm+gK1OIbb9pQwAgWvMHag5c/KZGI9oPZfiAw4LoLN89K+aj
bMGtcrCIasHeqNUC/hjsyjRTcqPujHIoFOtlnwpGwGQpeAnR8ppCg7S6bw0d3cU7
jcMawz4Zk7DRFDBA71Y0384s4dpwUOrwwAHScelroGo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18368)
jkozqD86TkALambFMz2EhW6UmbOfn6mf+fnSg2fiDgzePdpESHAW3dNBSsU0PWqa
d+SFdN11IM8hmQWaYzWdPXqVk2gb2fcHM8g8Tzi/SSWSqdASzpmZuD9piEJnW387
zPAVEBHHcdfCl7ZlCCCDEK4detg5gAfzvt7Pnwwd6447qAIhRxrm8NgyMf+Ucvst
PibwsKsvzM9Qzyr6IfrXAhFxuwoBtW1xW+/7+R+4Yl7P4ihYQlFs0GTbuPY0kdgu
IX5GrVM1gs0Ig+OWUk/wargw5ApV7BN/1FYAL4vMb3qS9585uJbJkRvSx8KvkzlQ
DncfjaExAmQLz/vPpslPFyBCaf4VS3raMomValtEt02t/7diZ+rCWv4FERlS+0B4
7tJ5zoowSGgVYrcNzhe09JoRw30OV++AHItIlzKtXT6XlExBjKr+BcZa3P7Kjy6x
prhOgTfsAK6kbYFHngPcJpIQlsrQx9ekr1zEgk4+gDElc7ZBwqCrUYh1MAQwsmYz
432E0uDEMA1LZYrcOEcLAR/PP8MAHdAemlbBN8kI6M+1i7ncRVDh8SpEIHJxhu4b
9jE+LH82lfhc9y8GtJp6lZuuf5nMMHm+E8dIWuo7eN4GWUcUs/1hT87HVrUcqRU/
t295GUNLjJDzBGgpU6ADbO9vGp0YnlXTTF2ipQ71b94dvoUyaR6R1ioOUjFImB7D
QMen2UHdYWj5A+UQQ5ZFLMvzY+JUgPZiHkkazcXAvkVO8/yx+r0wy2BwwmKl/Up8
PIvFN5nSilSdrmu9P0pczz9z+gg9/M86dH9gO5JHrGI6aANEFHuKPnxi/KFnUv9A
XvJvpe868zzFHL4hgJ/cqrnvb74if8rcf1BS/90JdinLu0rE67wPROS4Mde4PBS3
Dp8w+yt493SaXrauStq8GG18KeZ+G1w52awogLCwgTRU5/DyQ2u+ZXYq/EE2Jt/u
1GHTQWj0B8FU/JMYuaBc0y/KQh4Bw0rQyZRCRIDY/4sgldF/E8b8dq7hPs59mG8V
2W4tmDgHuMQ90W6tsMSyohGz671nJBFfQUfnekJPSnv/UaD0A6fxgnJy6gqQbpLw
SUuvKa+jM+OIxf22GpXHaHHkVYv3hP1DmiJnKuwnc20GBRh+3vFE3vctHYs//DuC
J8e5R/qnDEvxGI3r2aubWJpmp8uKEKmEbMwbsYL9UzoH8YSMyLRnBw87c+/MuhjO
HVCdCZ2Unh3e3Ijb/8Ndbv7vBJhi33eU1XSKH0g47rAVeg6nJzj4i6Lny/sLakp3
SFTqn4gNw+1/MdIm0bWWGayJSvG+FzSLNyf0nzu/3PPTrRflgtnsd/koWJ4yS4BI
vj9FwwkObRlQvQ1oCgvgmDHkX6boKcZZ+PVRw6r5KG5BO+KKDFTRPdtmxIDQhDHA
ex1mvQ6K9+PE5GbptX7GM3vwlCjBWijpSDAa3qCfTfS4BRyAucdOVW31tYxJiYCb
8TeXs6OvcAk/LGXtrsG7F/wwd3fSllMuOTgqXfHumnc/pPCvkAIYE205YdaPCTYk
qHQkhJtMv9ABDiYzrfBXaaKD7Y5wXrpO3MC1WF4ePmvk69Wki6TGa+N0C60SG5SX
Y585J9gJ0rvY6LgjVUp8wuR/6aZkSoBGZdHMes1nZ1yrRuoX70uepZ2Gentk1lWB
L3PSx8N9vBNyQgBj/Vi0lwItAeRPSmpzfuiSzl4zlv1dawzjjtXC/eGWNsStbb9D
jIxk7HpOeVObvNzUl3zRaMnOG9kJsY5hmviUMZWG0G4D1A4tF48dI8sl/7TRFNEu
hNXebZyfYtyUhQ9zlOpEVozW/tefaPclPN5h6DKUyxQx4q5Qx/ZmPTIu2gyY5ja5
cjunK1GqXGih5g1LzhGD+aHXQMZC1qGyEDdC9kyrktCtNwZSGii96BB/ngqAMhd4
ybQJlvvhpGtfYq+Gh0HD8yMC68b84Q+r/UhZ3FNww/rWRDii73y6Si8jopSrUqp1
Po2OlUZzMwDssAg6ityG+z4pxzB33vQrC/13na/RIqcGXDeEWI6xng9rDPZvxnTk
bi3N65AHaBb86Dz3vDcYcn7MJfCbpUWEJd0sf7W6kq+gTZYFWs1Li9bmCOYx66zX
bhDLE1gRCGPIHJGkwbdy2uLC4T4AlaIiza6hlzGVyeMCedSfxmZE1ZOvsiQIe3xj
OEAj0QZRG4cOpaG3Gp4rMpGo7l3/kqxRhBRJe1B5Lc1+W77rcaXogozxmf7qF3BS
JJOKYWbl1HjxsaMtslgrH8spw8paajRoS4/KqHcrZXp+ad8/nCzNkj8Z6XkNzOdR
f3PW5ZjkAJw8Rqz/9OyBkufkGF5i2xIkk+Vhr15nYS3D56pcHpZpkxz0VbWcvCUm
ea6Eawf0BBp05IXhNDUcvZxcJc3itn7hjkVS3rHaI34lbmf9EYzSD5YlJESE01t+
Hidyxfxls4uTh0AIbJ0pwpvEhrI5VMXyocOk7sossOmzpCJDI+2nrdO3QfjhkASs
CtDNjztqSuzMgzPnollrnyJyK7Qsshu7anZldjvf0YNpzCpsXNwchIEl+DCtBtoJ
BMzsuUhYHFjX7DLY9GwOu3lwl8a27XRuHkkmtioT60lzCqYE9byfDEFY2yek1Pex
jTMhyEYzpyWH/NtXBe4MeZhP/ydwGhNMXWpV8+mBV6si69YoPciZRGaq41BieemO
5IB1w1SXaQjyQ8rrSjFh0PWz5Dg1rwNU4AkQdjYo3yjdXMzuCaDU5OkOuzqlmRMs
IZbMHA/68qJ3g33uXvm/5Hev5LUmD4qY8tPxfbwJGt/dSmuvnXvoPVFJJwA5d05O
NSaCSOXw9NqDfZZxz6Eemu1D+rvrK7YG2QFurZQFrJz4qh0lx0geLjLoiSvL1ljY
qhzlxvPz5S5DEcBJ/f6NicJV3WQF9uD4vAmzjlD0l4kXIw/TGqOynb3c2+N7NxLv
P384kFIVB+RY1G7m6gPCxiAfqCBoQutPqEz9ZqiRjWEZ6ESfAQIngmuGd1kt/h1L
uJU1zNo+2Fdov7VBh8VnuIIeQ4RFnVR4qmpHJR0LCzJxymBN25RaKshPdVhXvkpL
8OiGUBRNjY6Zqez1+MTdfnUS/zsmBcWsEnwwaPmeaZCIEQz9Bpd9lhl6aEJYit7G
BeCicxg7DvcnbhpOZuZtcimuB0F2oz/hb6b8dF30sGWy3GU3UwnpiXxJGw40j3ti
ObSbcYuGgWw71OnotRVC4mKgr5jWp05UMzZiPQyVUrzFqPz2qy+F4TNYgb9/NTMh
7vVdDsoRFEKw1zxMZNy49Wp4Llbp4oftgOHrk43sqzeMmBmWJRO397pYPb/6UfEF
f/8WimzSxgg2voJm4+wOIHJlwfme1zuBykpdOLWTgKfzW36I8guYGUmIQH9AZS35
5KI2+X97jgXWBObBq4X99rCn0t1XbDm5dzUldzAlI1OHqlldSbXAv920DL4ieZzy
SNJjW3P3GutPUYIPfSHBJeO1isHHgmOaGmNP+20EGhltNwzzZWiaACdaFMyWYo/w
veQ+zk3JCEhJ5rVA46vO662s3yijaXfrlxYmmvcQgFvEC5+io2nviyIL/6THioEG
5SxXM8pLEhD28rkTalmZHUCE+Fz/yv0kD8C6cr2pleKh7sjyYQNefYlFwV7csd3g
7KcVtawP/au6OyifgLcCv+Efn/F2kuwuDrYtXRlsI/c4YV9PqFb7j26k0FDYvTE8
wxICfiGvCuyVtp+fEBetH9RR3syjsfKZNaa6EAtdF2Cm+/oOXTTqhLLt9EkHRrdb
C0dtSMUk114K7s9kJ1A56e0nFVmgMbVWslBkWh2y+usRKI/iGtp9Lm6PRBDZ6C7v
5Dy07pPnZaYSzYJNUCY44P7Z0BENQrf5KsDFZeLfcHbOfUJdmhA/mrInJ537OXYY
64O4/8dcoCblLq7Yv5I/sWxX/qkcr3l5mtUXpaH3uIAkJULVU/DzT99k7rDRgATa
5GC0De2gPLT2aD+UybXjoWQE+oDR2niCRZqXErarJEEOvnvgzdtS6q3Nr3+HohKt
shavNWyNRSoHidxHHzrOYkAXCDaufADDDG0RZiJ+NnxDzWHtE3WGJFS/vQWuDKxj
IBOBALcp95LcODI6gwKRjuERB1ugfKhVjRIP+6g2CslrIeFL4S86lQRwhabMOlAW
IGc4O+cyoCtAdz1yfkmhNTJlvznF1+h8SFfRnNKBfl33vrPCl1CD+SVp9Vxn1SjW
bPoTtxtMCVtNpR+OJo83YVbJ6Wic05wPe7EfQMTvZJsxVZTnEO3LMVxzmRfeC0YU
FKD7LgjU9fIgIJz5vMKL4CeHditmHYDMCpjnqQyFJ2rag7NlyjdCHBqBdz8dRGs6
mp+Hx3yhly95HWttYG9Onbv2aWMp31DwTjg+HHXWZRhIEjuYIL5qI0qHf6+eWvY7
1uQcenctoZq4fRNIj7pCMd24fany3DkpCTHvItSv5MJQGRHhZl0ravJJMAOX8GbZ
HVbr5mJUuzFNAukroYy3bEe4Iv0muZdaTH3grCsApWd48ZEO9y9BqfwEddzsdTRs
H2dP11oi0HGnv7MHc7MyIV4Dv/eJgigjGe8OUpOZaS2JVl1fL2NUkbUsHVTTuA4h
OPvmBtmOCEZlbaXwNLIdUWCV4PG3/ol2O9n2wwopfOo1mceHdcKLDYa/hXL3xlGA
6lPHBgx+rKrwn7rT469tfOvPj7+rWvyBnXxTXrncXO+1vEXE229GC+K+E42RGPBL
+t8XbGa2VSdTgTPw5ya0cN6ZaJqBjxx0sSCHjeJlbl9RoJoB40YcVKBRc4QreLdN
EZlin8YLi0A8HrsZmIr9QkL7MF1e6V6Wv1cF+BDhYXiNA+4cFlvTG0Nv7RK1wdEe
JeWbEYFEiAi2JGEYmWVKaZ+JqhvC5k8XRQtnzeQoG8uxjDvT6hWAmGnPlg4pA9Lb
V0uaKUdvqpDZGogG6MopR8P8MZrUbzNsz4YpA2NFQ1RBolC0rXRaprggHJ9D8Td8
3EPs/ntKd0oVeYPoqJ0FLcnCAA5rh8ALfSNJiy2nhjV26a2/0Tl4l+a7XP8G+GHB
iFIfneE1hSgbtxHZ+KPt7ODQJlS4JYKE5THhKVrbluhrI6SFAvl2o6uJGshvLHJ3
3tbV1BTmH3C/Ia1rTvKAAecoPt2m+Jgko0wcRtA0jVUKwfvAvohAZSlaVy+NlIA9
WmnCjteuDZ/s2W6qYmkLL5mhTohsCGiw+zMQum3b2nbC+8Gp7QvUL7G35tf9aji9
znXGTyFJR0+7Ij3Hgf4XJt2dWsYMkiwry8+1nBAfaJ0KFqCa8AkqizyFu3dU0qPr
uDvHJt6+6xslDs+7Eq9BVW/UhDpYOnaLhThJj9bM/VziWfv6HcnqWB08q4hgcW47
/NulRmOBdQUbJyIrPNH9seuqlw4ksq7kdMTmBUNXEDhgGiNcBZwWPFvl3IgZaq2P
XkaThg+YyTxj4+1re3x0wXhIVv63mNL/aUQB/Ga8hEWS1dGV7Nu+INoUPU81htx+
D8RGImar7PNCYruBP6Lxn8K9Az5Wl+XCdDqOWyxqBsSirLRUVJCYUoo7vo8p9Q/Q
luxXwIbi5g3wcK8/7bw4yHDrCouMbuheEZKwzS0Etq4muI6K/f4twLIgNpF0eS1w
QPDcdkqqrjGUqvdnM13o4IcIsT+N2X9wgtwe6u1gdIK8S4SE8cymSzWbburcRa68
owFSaMACvl5+xbfXUg9+KoCTrMw6H3EVRV0tL113jfe4DeXny1Xrl7trxI0D4UYa
UK/5WWuSpyoSmck4KLo/MxG1dOfbMIReIbWApxBm06k55y710AWrVOeIqsQCXo5X
f/QWLUE5PDhng2mU2vXTY3bj/UVb6RMYnTwDqmPx46W9FNJKjSBC8OxoQQVCUzBk
47EfpzjLrDXrnk73fZOWD40WOYl+gYjrrv9IUk8LaRQSJZrlyb1E3gaYZqGJVnJg
XKzZblSTeQaiYg/pshMsEDyLvCl3IA6n1+hULnNOmfl4bA+BscL8BDo9T9mYMb7A
9a+3ApuOfcHKFnDtlDFHKilx362DG7P9TeToIaAOubvFxXP2Gj1ux2lGrYs6qLvr
0jzDqfO/xNJjldAcRNiD3+p5Z0VGBkyses4LIuJ1YfOpluoxWCqyuSExODDuSMij
02q6u12XwV9SIERXbO4hG2aHhXAAi00s0KvZUE6p5gqggPfduWepNYY0xyhAQyhR
GPtwlWKaDauMUQLhw0Y2AhBOkCbfw+kgKuKneqJtQQl7CDub4leUyv7KxCGtDBTc
8OVkYxbiTiyqDrlcKNBGT3TSJAn2RHnsvaL7OAjC0BJIjk+5QlPnaFWzqhgsa+sH
FuAITvGDVhOVF2wm4EY0VI57REtPHlbfBk+GzGDArDNdX3PxSCbdMSOp7kWm3k4K
v7GvtriMhEhIXGXl7W6ZQvhn1Q5Ccvuu4EpsnFC3lzaXEY7GC+aA0l/W7gULlNkw
n5NYihAil6GZQTywKdHxd+y1Eu7a/J7mpZbJw32QZ/6BX3VoN80Iv6/YwgcRbtRI
bJHJ6WH7ruqoSKTFaF0Pgv8o47HAC5Ym2gtT2Z76EHVEzkekgxvuJgwT4Y5f+Qec
pcJjslMF6OCxzwKAIkjYeWg1On7OrhBN49YM/4pu3o04P4Pxp7pZfLKyZfA7f9TB
sBR2rc9xGmJxfMHWYYI4sWe8b6MBbA11nEBrvF3EapM7qk8UGPgBhyowW/f5LVVs
B8lTEv9ikCCHsdjTiR4ROooyJ5HeIR3R9CoW8UMA9Ot0Z+uJb1PMRYwAZxBaasLV
tIcnSzvvB2HZ1e4hxFr2RxGUcf1Eq2D7dGiKuX6u0EPBoND70paLP+J+ufqpF4LD
hz9598kyhK60CO3F7XHzubImBcVeHiv9de8BTKMiSmjDEp9sxGI8xkGNvEAUa72N
RI4wDWzBBovOR/mrlYSQyC3hvXOuvVHjDCj8V3W3+H2Nm+XQwWbK3hy9yYFM5I25
Gtz/YyvUpcxm9JmQdqEk0LEJycqcN5R1efqqZjH742xq7+Q94L1vveHkaj2A1Kuy
q0rV5Js6+8FJhrXoUljUgR6r9B2jExRjFI/luLQLja0F3myoKyhoDe6BCppzL9aw
MWs96US6dtFReaoJUSDH6hkjzannNT4xPIjCRXTGuW76Q/uUYH0JhCpcQ+U2GFDS
n6UUU5xNDC8Mytdr53NPlD1QhdziYSW41E6oX+h3fADQr00LX4NLGU9zw9XYgoma
g7TgmsuvXyW3sKof2wTpOawLDD7oDuvPQOGdj8TL+PUQHMFjm1t4cLUzHuEoSnLS
Ps36ES7O3B0IW0Yh2BuM6a1hq2v1q0Y3m9SzjBx1RD6jn1NHYT/QNfe1r0A21xpU
DNiDNTMJ6ZeCrrvj29ju5x7E1M4iFjVP4uxjqSRzgbMAnbW8zRWTgD3M5fdkWVtj
VZE6GkesdLOQY7sJTri/COabiS2810QhoTxJtnT5HuDhHd80o4SVuzHnxylp3E6b
LPwSMM2/saoqtLZC4EYYnFVUfcZkmgPvawQLjsqPrPgM9U9gDcr2HdK2JAfCgKFh
G/wUAaIJi7Z1nU9YBm+5ONLXv5U0St9/06VxGrBU5ydtx3h0Xo8hjpicHiParBHC
Pz47fTzzmPRvxXVLvZnQdUB8+Ps/XM+n/dEj/C3/umauqeA/GEaohc6kFFiFwR/H
YvZTBBrKz76hwS+ftcdSoBUOSWTHo8wm9Lwocb15lktRh0LQW2UBjHOEUB73Ec7+
Kh+Cq1DPcTIjJkmR2ROFMdBL1sjGda4qnR8QBGHRtiVsOyVnREDvorZJCQpYQHV/
8YqWc1jBA6tcAkSs9eKZF+yxd4iUZTlnuoKI1Gn3FW8sOIOEtL7yNzBDFZmwF3Pu
nYQDNvl+1wuDBX/FMySiX3k4dc+VqPHXmLzuoPnY8MZ2M/TM4aFyrbIDoXDq5C7l
6bdL2CMGRFL+ZXWzKqi/AtoHq7pvLmLip5JBkmQYJsSxrrbUPQxVpjwohckEAS4j
Gln6+lRxInfWTZeIhFmBzWTXdkrV/LFLgmmAwz/S1M6sUkIcSLw1Of6K+cgs21Xk
wCGRXG0rWT1/SjNBvOXLnV9mO5zdLDeTio9cS/5Cc/vA9z06K5kS7f8wtx6MnQzC
XTiUswf+8h12Y8emUrc02L4syzxzq8MeyBe9d99qNTQxMeR3zElnEtPyQDlTifBG
bti4nQNma7rD+mJgya+GsaVFrNc5f9KngOoCBgLMOVc8CVtkaeCPp6zwiaqSCwrA
5Zezd2POom2pM3Qkbscy+/EAJWdRRgtu1vrRnvaTKcvaPL2YrPwPmx9863tNi7gg
Fp+CW7KjAA+Bfx7DnAL+FlSyLQP1vRjBDtsiysivWv3JETQsa6LOPe21tiT81iTp
SB86FQeg74f+MZn4mC1ghT0ZV1D7W9373SkXTQeKJSOIbf3JuEb+OFXGvBjhIxHR
+kow/2MBMMvsjmxDLzDydVIvfxN0KjHK+6roUR/npSQbUs8hPx2ofuc0j4dMno2I
MLnqPamczrajQmCShh5TGAQzpAbuzMp8DV3vK70lsvOfD65mCv1wUdytDKL1fNV0
Wp/+dA3oQzLEnlRMtB7W8MAr1IryatJsLPO4zoTve91o++hsXI2fcIUYx2xJFyJp
H/t9cZ0Ik8cPXCMiM7kuS3mubZCMwG4YA2o1bs9IZcjRkuZh77THpM1tBnm2CVxf
4Kj35q43PkGHjMZj5opqilTrm0638AdCUOh1q+t9FEy06/R6rnUvZSdaMcUdS/c1
Vf801QZrxYADEaeDj9rbk9bUkMFtwNJGpIpx/9g0C2OVgYc8MAq2UFq5bzJ0Xjvh
1vPdgwadOKzy8VOYKHTFvbqG60nChUy9zALz/3S/xI+ni2zAGmIeLoN86pur39+g
fcopH1wAC72Qe9kmuEwknracxir55108S3xusCFeZTiBloMQqb0HQd49V/smfekX
cPHRmmCzGxU2jE2cVCGicZIBt9mi9t6ikXaKnYZl+gRUGZasax9k+HU0OP3JMc58
zgzW6IuZce53NEbEYx266EE+CDCEBzbrGZn7z1KZo08Rb0B0n8nKWtu7OKBb11tF
ZThRZCzrOB15OuWYqSkJgGe3aDmindVUHZzRC2jAoM3edN+6UW/uMy3+08hniIzd
vgXS7bsoRR+JBehU8l3E3Uw0Y1CS139lVZVN+LXuLpzWQP14RGMArWndEMya8TFt
bEocr9j5JzkrdIuUKQSMJGLVAN0ReRkBRuP/IyHRSrTbAFeBYEOomtYU2s4UlbsU
t8wzZ2AtMQXGrL2yoLqPECrKlnyFHtZ7SsM1825hvhGhAi5+MVBhXlsT6wp17ZPH
pQfO+seGmFM26PffD5rrJTjm9F3PB3UEdP9rCUbPqTkNVJV56wgb7wxAF5z9ieUN
uxbNASzPuKtgkNVhvUEfIy97i3q8Jn3sKbceVL0QKFtZ4zDUBNzqT8CXmpFqimoA
/h+kzIjbidn+r3lcyEsZgZgpeWLUlYTu2eCJKvxzK1R1E1YEThneveIl7le6RxY0
s5YPwgZT/wpC3p64nT07OsnyBrHNaTGsJL3neJv/pliIu3ar1kQ0fHOdjVDrfQAl
diyTB9WIGoFSmoqbzK88rTsPoJX9ISh+qg4GPXnrGqqlwdBFdplhh5S/0/pFNvGe
+NlEBC+HeKprZZxIFgw8mnVIGLcGwY5gPxUhVjeA6TocbGDtLlmp4L1TzTjEvTd8
EX3/a41k7FWvLCWRLavvi77biwW52YZrPOmEaJcf5LG7xf3/BRZsl5Hu5SamJY+4
vnQwfNaWUF/wy1v3JK9/6rV9MJFL8cbX8+IJgitX+6Gz3k4jQHUGmhIf691gL4De
7GYbsjFHXKIRDOk4mK9zeKSM78uz97eHGE8L2bjvfRjR6kcmFTTAoSZKHfo3hjWy
3aQjE89YZfU0jNb7MmtF43f1BZSiZmQxd23rwt6Ay6zaKfUpPuS9qeTBrbWskAoG
URIqg14eZ8I0sn6jXvO3VMWRXak4pTqu9YWG/weoPn/SonapwxAtzJewAFRn4Qz3
t5ltFAk0y95z/FIBUctzeXBalXodF99uFPRiWp39VynV8Gw0wu04hhNxYYDVf7zy
usJB5Fq5yybG2yYU3aUwOooGkTvXpgZB4TlHCwo4EiN6ItcnDbq1qIH6m7Y90RwN
Y/FpkBL4d3YmfdcmTTfI7KI/AygwAc79XbVefp0rFrMLLOVaZGSgUPWG2EScdzQF
+tDfKoOZnEHXjCUxXOGKyPAGY61I4jFRXKFirmE4Q2VBnRU4WYpICqQR70Uwxq63
BjpVNjktpTGbvSSeThiPjsp+Tacj0RQmzjOgzqnZDaOPl/h0eTVZ8FBW4i+43ABi
+lCHYLtLxAUsLHpPtoJKR9QPp1I3FfqmIKNC0hPrx+RVcQ0AS/Un0bU0D6+TamtP
nmXfILE05Zen10pVXRn5HXmWhh+UXvOaSCFPt/1SBgbP7rqfR7drm4SerZ3mMjO0
qLeZhVPqzrtqGged0QoDnwgZtJtKr6/ula/Ws3/oPZReOXOgV9VO6j1520yAT6TO
ViBxcfa9+nbpoywGBM1eln5cZ3fz/tedMyLIIH7OcPkiuRGqQOFMJfK2r2yb25nw
rBbqnNarqKvnWtTQ+uwHasqan0IQDEAjsFKe2l3zvEhN7DoI+AoFjjB3tisSNs+Z
HZYBwmpB7YxJtuZmC+yK9Lzt4L2rhdIW/y9CpK4tJ8UO3R+8dHapGV7Xh+n3at4Q
mAmgKFQnZGaRj36yNq1QJDn+v1nZWP0IWhcXAGvHjr+fdAlrFRlT3LSfoKen3cTl
qB0mv+nzRUfzU5W9HbssgSQ4Fv6susUYN2tclGnZUFZsqgrDxlTZ8Fnx64IA9zQl
kzu9wXc5DeOfbr+CNt8XnGvAIpllxZZ8/aHqqdbSATV33U33I09tZJFQucKkaB/q
6qw7Wyd1JPU6V4iWVG62Lg0RZfySkr/pol/IMvCH15fXdrK9EgCz9sz8oay08RsL
ad9C666J1qbmSI9zTdRbzGoosw8Nr3HVAhTQ/tcy3V4BQN3YZvNqUErWrF7rqUaZ
KVRjLGTSKDjTFCwfhBD/YHuVh99Nq682EfTzBvTqs+yjp47aEz55kSNWSBAI+y0M
DNn5IFDFwYav/o8EE20ITTnksPxG34wirM6fA79joC1p5b8keGo4nzlZwt36AEdz
7iAuvTtExnE+sNSwN02PMpmA4429/dXq53tjV2ahjjgmJFU+lFZzgKNv3lD2aSZk
mSP5Rk1OrKfLgutFUDHNA80ktn82UoE3meb+ttaFt7K2V6Ax0wUvuQ7f2KivxjtD
GOUmnX/sQZLCot0thEiLOzAg47QNj6HyuJrGzg8yBUAA7dk8PRzu6GMmM57bEtOs
OBD0DJYvowqWEBsuozpl+toILdsxEulPTnw/TjpoSyjzLBwTwShBibAeH5NfAP9m
xLzh4skP6VQrKl62FRyN4d8ury4+DWXl6yn75s3Vw3RUtBuJYeBJGvGhYOZl+Pi6
XCCB4f2QKgFCGwvUKiUsIX2hLVBYM2ft/JfCxSCo2WX7DBM1F9MY/BenMYCJwUsY
/dW6x/9q2h7KgvZNbKbJJSb+roLXG+i5r/WvAH5Oe8fcOKgxaJfG9F+aT9tyTGHC
3YN/C53OWv/WNYhNb9sAMlBcLcJYX03p1l2MzMEfkKN9e4orDPgQsJnJl/roJGJy
Hks1PVt/RPL9gSGIdUHEeYCyOdUtMT6+FvM/bg2Hf3hA7BeYx0vowCbmVPNhXkbJ
0IDV9Iq+LoXBdjCNjVp9Z5OLFjw2knRGBepajGA8OHpjSxHPnLSRzxTBF7t4A68f
AD75FV4EWkJZH31BQUqfmh5c3C3ZRSeqUnIt09Dxz1S+a96Y3Jk8hNnLQSEKtkCh
ua26KlZDulOUu9do87lNzghxVWFRSf7lV4R/SlNKAn2n/kICA+9mpCv0zwxHglEa
sWiScwn6GP23TwSYhX2/M7OvLxd3lAOIV26jzft2Oz4PI8gHek1TVJjrgdDRX/n4
LiY/yM1QQPhpvobYmkd0/TXJCeJqFLCbNmkMCIcyV5qMhW85EZCnAuyaV5/1oN91
e0uLg7AEiwSSh2Dsgi47Ia/7QAPJGhD3ckkn/0EMkr1ltw2kU2J8gwGNfCZO+eYi
B5OF9elg+6I6iYwkzuEQ/H2Qdb2yntY3NDYNzV7D7dhXbGqBtqJFZRp9v6fv3WY+
ig73CXOfZZK7e1ggFgcXbEzXuBQScBMhUofpzOfWfU68MWv48HFxaWVijWrkhGxu
VEs3HIpHtjgBJ64cZJeL40Q5LTf2IZrwRWqaz03RU4jU8NpaJo2N+JKMgsB4kyaJ
66bgUGt+2Lv7noj/SwZpHeYbunDDuMs5Baw9qQoMwEpGgWtcCZdi7RDlBqFFDvDI
RaoDgT+k53eWLt7tkgWweiLj0nVxtFZc4GLFUzQiiin9Ho9tECz2i2+1cNl8jZCE
LxLNCmQfT0Dw1usIWO8fiiPaILO3YGpv1GtiJACC7CMneveH1NeIKHnQJqrX7/cm
HEgMklk7he0Xg8FR01jX8Gl1n6R9znprr2XhHbQXnjzG8KetQBfTazAYMjlHZ5kJ
3iNqNT3zT45YivW2L/j13Tz8OQMDWvmty0cYhPpzCkOi2qrEPyj9NrNcziSoVzKu
kAfLVLzKdzUXYqsfDzOwVQYU1iGjApJqYeL0MWIyLKS1hPEmn8yyOTrzUXlDCxhx
+6ghfnY84uhwxJNEkq+O+qFiXkuwpFv4n0uaGae7zytvqvg0psWSK9qnm4m+y+HC
/NhuQNK7okXBN+6sZMMIDpiDx+9VB1Zr5C2fwQ04SBd7n+iaJmXwDiHXGeIDyALr
nX1GG2u6Fg7rhjDjpBvQBSg7FBNo49L4rYX3BJBYyWLSXQ/dl5iQ0bpqxzm8197O
5327dACE/dZwkhLoRtXo3XRd7kDe3TucgTCcejUVZ7J0HZQhcO0UPzpUs/LvTbf2
2ncttpZ3nGzjpo67zhuTyefFloLJera3MY87zDtvlH3Q6id5bax3LXqEg/ZgO5ST
1S6C+trvQZ3Kp4JWm9PmkrN8sS7noGIxG1wMHL2WZKh+YgiR/OPbDFDjbT8NBnQw
spDxK2RBFctR36xrksf9jzzAa157TVMYUdRB/ykPsJhEcPKBBD2H/aFTl/xa6rD5
0hl0ny41Nka01kQyJbEZbsNdzT1vJGwzfdxyqyJUfeDl8dDRzGKG/rMKk+yAbjUk
qX9PjHoO6PrCONjLfsbQ8MFofY5ZEB5Q3mE0PjHBwWQxDhoqoiClfDMcRH7U57nB
yIpl9Od/EicZ3M8ow5NdMXrzElJvmE53zd4kKc49u/NuBgCxXg9y4Ly/7vyQRkct
iSXATlcFWOF6TSyn0vvZ356l9lmGj1sxHW6vDwB8+xwEIw7A0Yjuhef2Ag7JSptB
+u++OPkR8bbxwfhwBLnD4N2zpmGk2mZwvxVMQvs8LI57JcH6lcvMe6BG9O7S/wv4
D2fkbgV0O7etu4mqDgFKv6jDF8Q7HZ4JthTGz45vFVPaalw0ED5Zca7rpn7mpYkb
FccIr2Obthvvn+MVCOBoGwo5G9xUFGqgw+OnstmUZuP6l7Kdv8RrVR23mJQAoBi2
8ai2kWgTtmFJDYiOWHbZn0SI/q1tZblFeKOUYg/cSp5hwPyJCe4GDSw9rZk8PcEp
g3LsCE8cVrffK6SLoXFSItud0tfnwc/k4IyOdyrcMnxYjPgU5TXkfGU2Yis2Bh+/
ZmwexzUMmuDKefppVmu5ITnh7t5dxnWbs/QeMfEBlwUMCeJ8hEekvJ1TKiaj8r4x
OWGayzW8ysDI3e6+sc3WqLA4v8QLyBW143E88iIMhVdUGGBbabu18JhjV9muxrXs
p426+vAxgTGsQOItdbX5LYRk5CoRvrABVPa5/M+u5iZvDjVOtzvpiMYc+XJ7sn8x
kWgfaKHyNjDjpGWA7II7NktCsjG4CmvtNWj0Oa11vN3oF+8U9ArAML8WLuww5gYn
rpXt2d2IMbiD3S+zMQEIK9MhAkGDTcV/HOGHkY47W7uQdxZvlG5dT81ZAQuiFIOH
mk4dP/3SkmCX/22VXa/uYH9fpItCX8k6Y7LqeXGwYdcxwrKFMAtvO/5vXniImUTz
90HMlTVVnhbBVTBKOy6vTveoabkMmcfAjwzHifqAZYbM05UE4q0STNjw1lGeVYWb
0ZF4DZ4NuczDHon9gWNo4HQ9A2sQeO4yyVhFgnZpWjoaIYb/9bvPEDVYt+uOEIJp
EW4jInATUDHnSUDm7mfbCZlIMnXXPeJqFuYsaAE1qURN5UPdrsXW03fuMA9QdcMW
gK3feDhIZ8lSYqUKglrcYoa/isSiTLhqZrZsxcKyfK9VBQEvHC/S7Lo17tqQpOtL
wrtNCKztbOhoGH5R56gCuUIy8hq6L5dVtgCBKI6k84dxx0n/TbVCDSr8T53dCEcv
hCCBzYYJA+NXNua3CuIlytZ7yPBe5FPhdy4/UQJAwgFS8EKUSFDBxJ7ZoCPHnB3o
R5PKVuoSQxyuFw52MAMXnW1ysmVUGexMpOYL+C7AJ3aDgSTXfmOmFxeHmZ64bG5L
58G0AsOVrNtg4VGgUr3aDpE3SPDKT0GtqjqKlAtluO2D+QhBdfTN15bf1VK1+nSm
06EQrtZkSpcf8zTajfIO00+lDRzB6v/OEx6cWpRb5pM8gOJTD0PGmdYfYdNaa2CD
U8oUTBR+0HzQfT0JhjZZAjh7BcmSrRk4QV7BMNqaoZLWejK4ZbxWAmC8siCjvnJA
QOjdpzj6f24hN3zkEAQfDZspzqmSun3k337f/SuSSZEkC05rxCgg29Iqwd7QCTB3
M5/vcYFCUv4ETM3CE67OD6QWV1huZBmmlRe1RmrjNKudMpx48i4o9AjwfUkViUAF
11y00pWzdptx13Bon1wErLp/Ry0Q+RqiQ099I0ob4t8x8wQa/Rchr/GjscRhkEgN
XvsX/pkduF8RW4eIy6F0kWdI9BhtkVSjHqjUlDRHZI+cfdOJQLRdz0UtuKDrEHtk
U6T/SoGhrauHJKpyK3kzMhhhmJ7THTWM+Ndk6XhNifhr4COhYCvHCFCNNvLDRlIO
GYZum+LrPFQXsQsZFdDamBfz6LIvvZz0mX1T9RWMth4sPsdEQqPDtsastPQIturJ
9M5OhQo7b/i8s5n6ymwZFm5Ww2in8HYIhaxykeEJeuXzbaqu96hVx8wDUPC6Bwjf
D+srxjAKQ4tLhtdnDXv1G1vuKoypnaVy6ga//5Blu0yitjXO3UR9SV7/VAazR8jE
SWGa6UZo/1U6KSs/0OVlmcRWNIBzPx6/CL61AVd70n7xqzn7Oig11EH9jCKTnBsK
5lY6KYtvYW4OV7hbogHXYfFBmAd1XjHimAS5p9FEVcjwHVTlsXmMIX0aTiTndUdJ
83Fm8OPzhf0aFFy7Y0MqhoG0P0SczNZPm1KP2n0MZfKz4tKM+cCegrbecf73YgS1
MCRvBOhio3eeH9D1bKlHnXDQNBj+hEqENwEM+Hiu9wXXBSJLFpWqL05BzVFHya5K
q/F9T9zUbI6MzXM49gftyiA2E3LoGB1lgzSeBCuSpXqPc4ip731Ir9lyj/188Kz5
uDjkJz+LxX8JtHWlzbUFx7iq23dmDH4vUaknwb5kxWFeysFFjZho8sZB3x0jIY64
CkvXDq/Zh5yeCHL/ZkEF2NVhqZOIvxj+HLuUa1yw5HxtCaiZLSyRuvvfd8YkdRhh
cXaEeJwJL9oIE0C7fq1gFT3snBoJrJHAxqG9YYUHZUgjf6vjeTAYg9f6JyWFiZV0
QkOCUCeSzVNZAIIkhVxpuq8CKVjpY6PYSO+gxJkoPx93ydS/IPkiHngRBvlkAkN1
vJXppCrsD2/bjmil9tvGrWy6Ciqy6AwZvY9+gr4IgShhMIVoc9nqj8EsJdsm5BsD
xWzIxbwaM+l6nPSWh/3NUvbhQxJLeGn83s9aiHRGFd186RLb96cYkb8tZ3qfJ4Gc
J0cNMig6l3ws+snfawCF4r+RW+yE2SGl8vNj3Zg8OhV5hnKo8ywg+qsJQ3TFLRRU
+nAafYOgKNEGXPWnf5QEDgPwSaLzl6R+IbpvnOyJDniNIHRONx5A+3lGWL9KYJ9o
O5iKywKTTISxnjxycI1Vmj4K42Oxq06lJFrAEFjT3ilpVD4+As8quztitRpxHSIJ
RKAVqeXcDdrP3eW7Iz7jnU++ch5fMBuibG6TalFgP0l+KGcIAAaLOfjj8DQ6HvoO
cXfOo55veph9fbJmBuDWbIqlALpiT4JR5XhwK0x2M8BDGzp3YcZpm+Ehib/v0rJr
0ncVqsHGERN9MR39gSeUattJRzOLfAC/plDv5MJ/MktQAbdH3P7Byrfv2UyjekCG
wkXNE2z0obFc9zbXssNovHowPzcEhxCFpH9ua+zWZD1VdfaDFNWjOK1O9sV5k6RE
Rk/ZB1kf6SpKRWJlHs72QFFgTbqu0/DOG1YToe1fH2J3DBXTZn3hzM+wlz3XxiUX
dkgxqWFKIv7DWxmrCAComxKIClPP5JKyckjmn8gUPBHjrYlLa6UtUQ7P5kwOyGi4
DTSEJ5mNzkEH3cfzlUxjn91CCQyKW6ddCsz9HsZCmZgjjEjKwOmBC/XIK3HN8kmP
j2UgseUXLVZR2gaBi5Dw18jkRpUI/YS2h+l+BgDyQxqRSarHjmuGZZ9OzVzALSYL
lMSQOvgdD2JNmuF2raIkt2kn5WnuvPuR0QYb0dKajbmmJOtL8tVIWrQPgaLl8RN6
CDL0kRuMXROiedac9buRzweaXfdtiRa9VUGs3vOhlm0L3k9NbeEB3CrxJmF44nkI
Q2NsAAP7Fxf5fyZMHoO0fakrRLitBH53dJz9XUIzdILIzEiFsiih+W/4wLkQUm+u
bWXr23FW/etTqg5CpUha3r7B9hVw9ks+KNTSI5BnB0SB8+Z25EacfgfXx8uc/sgV
US0cijG9ASlc4K3F3F2Q8C1DG070RpGF5PA3UjuI2xVpZRycAn+7zurtT/OH+3dd
Od8qphX5/qH0+16/GNQJbnNEsxrtdYDyXkacKDzArNG9kfJvp0aFdt2ibTa4Wak/
etHGXcBO7V1yr8mHGCCOz0yNYJiSYH1SGsnRGmFTZMaGDMGZK4vhoNMILfgmiOU1
LWEWJtuc6xhpcjj3f2Gxyj6Rkom5l1Hd4aPglmKtMmTYuwRehDGtzY8ohRMnv4we
3+WYAuUtz5fG2UFAN8H/sjPvuRZM0pOCgHbokcVUXFHYZx/CP7+NBPYeF4qjLnQM
UYcYzQ3G6bmO25GdDGYo79MmrH9GEgmiEa6QTeMDUFVZsNZ2APH5gKslZlOBweri
0e6TrLmZYT4oMwsNik9eSGTAIMG0c0FAqVX7DeyVkurkZg/j3vizRBvoyIcRwqBS
dFcf+KbsqehoZWjftZdaMBsUHLcgx0roOzc6cQCo7287GFf+Kkfz3T6kH3TMLlj5
GZ43uVVyq/JrNhWuq6QpuAOVPKU99xtZzndDvxjM3azPFvaU2afuPHqku3Xp/ty/
1kogWWOijuY5hW7qfP1fCJNe3AyKcvd9JzSaP6cEVQZJAsWKkrE7unsA6m/KLoMQ
kGIc1FtyClvk7P5Wq2gxFMbUJjf27V9ExSeLQfYhQMw7X2JRuqscbWKnBTNnPa2K
1dzv4eYVaq7S42Iakutn6YPux7qMkF7jSNFUPJYPUjOQfp0Jabbc+mvonmBg3rXU
9tEkpwORVgmbYZQGhBllBajK66BfB1tlkVtRi9oyt8UF8WWkg2I1uOM7RbigXOiB
OpnASo090mIPQXyLUaSHfQUgUACCFtBSd+2QV3Do+FyZicdoE4hiMykA0c4Mn4zh
+7yfn7aArpe3RbyvothLf48u/ANoAgMe8hoz4FDtMBaiRV3BlQdP2YLTjvMLd/If
V0QJPBJAcntI6lLtwfX92Ll54F+WEe5DH1jvTeINbLmgVL6D4PhofTov9L4zFEH2
eXRZGgcTLjtqJt+jOp6Ov4gZKCytjZeleAVbJ+C10Fw7fNowylqq8S8PfCyNf3WX
ptYMP1fyxnzA83W7aXsc0q6MXukHhodTssqBajfO8sgB6NEeTVulWNIoH0de2QLQ
nS99/nwa/hjq5EBPmIazI5gA0vYINx6gcF0uPIq83Lt+9WqIRY+1yGV9/U6ch6LN
p4QihIUiPS4QLxGZSaxhCsOw4elZ+vbKTHavpXHWcNC7gqzdgRmxhG9P/oRSTfUT
ePFfzdT7lrBwFM4P529IVByMmTfILM4PG0kXMJ1qcBNI/Fg9jbKrKb2BIVdNo6O7
DGPicOqT75w6UeXH7TGQcxQb/+qPuMHSrPadDCW7m8C4QMqTyUha3jjETTY938B1
g/jXe8sa8j3meqHKeuR6fqYlsMd9ZxrS7S2s76HEWAQhWal6/SyvViEejmjW9J3X
5f3N+1aziwv4swMUrpfrjCYJlP5z7VpdYq7waZZ1UTBI9EEKyllJRwMZbMkdyUwp
HjgGoKF0hJHTeIq6qwWnu7HQBVWMig5AZR+sj5kx1DzW1qhmuOZ2thOpvRVzf5iX
hCr30oELx+ysAGQXgUWedaMGDhJWJ3I6P4tVxQdLvsqs87ZYw7Jd/sG7nQanvFcZ
hY8/cRbIxO0XKV4i8YKyXCRbAr/SCLfx+R+qBEUpTtQbMCi9IKVesuKoFuAXeJ2M
M3/gSB+4x6PR5pfJiOX9N2FHvcUJ1fQ+ZGhrAvHPwat4hODLUiqbm3Cmow7vaiND
shd7d7K9xF4wlbYvxLT96G58A3Tica+oXlK4bGCyM7BRC8IQRwpW3rSXWfDGI8t+
dJJv9tzE6tSyFJnZuWDnfieqdQKfGDUcQD81kNiSrzgj0O3pG+4u+E6O/MgOA6BN
JGRnObBM9oeL+KShMx5nH2S5ErPtjusJSRML6FckGZdjKOMdywVg0ezrvHG+0h+k
Uc7b8ZJwTKxxRhclZAQ1s2B/HrVWaZ07tK5TRh2awB7G/ifh9ByLg55Amyve7E1I
dm22sp5C2N0wtvBVa4NiUNHs/PCWIqdfregwuwTWloeD1/iaBfb+hq6PInCjI7Nv
N5FRSVNUKO0XrRCvoj4opdEtRMtjJvOHnJEKYEiEaAKA39AuI52fOYrBr/DwW+Rf
LuRMmxfcaD17Ne1Liu2TSi0uEggrIDlwIPs02OxGuXTm2dyWNxkFaStI0T6B2XZW
4bgKCd/Fb6UJBoK8ghBYXEnTKmg3LYPbmb3u5PRbV84qVSiLwCdB8MrXUNznMNck
WWa65x7tXVP/6iQflWzMPriw4TyOcL37t1bD2xkycDz2oCTJRwodiKpIt/sXrvp/
cTuZCnlJXlqEAX31C3+W6Xj4E/KFobIwK0hgA/uVxcVw76/CtaLkXI6q1m02WfqV
Wim6kSEs9gEYGDBEX5ASnxTvZSnw8ERpYxzRadaMCrXYuseh7JLOhjGhgsgmxQNg
33FtK8Sqdvjcoi6J64spxuQJIXrpiDLTU7t2vNhqW978BzUHv8uK91/8+60ockYK
/wQlRlcqheBrhIZ9gyv15FA94kI7RP2z7EIkqFXdG8VGq1YFycao/9OzQ1r3TZng
fjHdCwDr5dONo1bXlT0RhdVjyi05etK/6RlfBOybS4N1aw7dR6nelE8Ud6u2ClSi
veVltcij/sKYDkfWxEFbN6ebSijD379BpRYdrSE8awT6f1Hv+thQDYaqpQPGmgXe
egQaetRDXQBF3Rb0u5SNnli1CCoft0s87kKk2z7VrnX7DztK3ZgHL1G3XK5J/ymv
6tQLzNc4v+l8vd5TTrZRZcxVmGnAWoK2G4FoEZG5ZTLYf9GiQzygOnb3QzClEabO
NJcsAZWBNXl+5uvMhmn2DCUWR1Jgq3+PT/hO9iqr/xpZhT/g+XQLrEIA6pK/DZrg
YjFfL5qLwULJvFzRS/Kjatznp1ZYzivhzHPrAjps7TktkCK9CzXYC2AejasRKxkD
IqxDz+YnBqMHe1hpkLpP3hi+qLkc60Vo3Ayuz08qJDnBQDiEwNSKX4Q3aBhyBGT7
5H7lH1B1euonMnMxJqvgcvHcBRa2nhuFL8Be5pv3xdoilkKrDH2SxcKlaZY/LU5F
5UYW/Xm+MeQ9eim9GO3GszqSfK1ZtdF6NLfKkuLfmGt+4zZ9Uyv6S6U0goMNOz3g
Cp+pNXVE4+/ppB7cHm7lEjUbQa1ElxpzIZWezwupEWXpF8w4+TXNq9YbUWJWSpK9
u87aIyF1BgeqOBToIGDaHLoe0Qh7mqjZp8X4XFfCDFAABHjcsIHyCFZ3xDvuzDDP
T9r5dhiPlF6kGEUoS6VsMewFGQvpDjV9GbX/squjEft6wBXjijylmIB2F5lDPef3
pGZXwJ++xhXSpoNjTGggF2x1o3GQpGsyCpLd60Jcj8XiUoG/Lxp3eQDiHVbTvV54
PkSQi2wnNYO7IMA4H1rBYdZ7EGtgpBVOXd9vuVl0VyaObVQtI1vE4+qh6fFaLMAi
hI6Ym04Q60ZEa7kUqtV5uxavlKxbMXQrzaD+cEwcs1dkUxUO1aDxkb2vH78wKRJW
2AtmLmYv8xSY3yxooJdWHHPARzN2IGnNWHGWTp5jmbFTggK2UAX17VsJzT21R/vk
lIFYOVH4/coisv/XWArUOg3CUWza0OxazNgrhHzi4Wh29zV3s+IsuuPj5zYvKGkF
COh6+YnsQnIHKj7b9d6svNtzplY+dIpW/50pbh4+yIBKg6UPgskIc+T9+ikgaPXH
iHnU1gBUpX5zy3Eb+2Bs377KeA409UeNC8+W05tPk7A3UdOfyLNDlRlXjW9aLF3d
rsKZIYtyOa3UY314pEvZHz62cKcSzwgkTyhp4fvwPzNbYkcxDG54XSd8A4xW118Z
4UWW1FDie6MLoyQzhWY9EblWRApqz/vjoZRxt4yRitg3w3us+QVvQVU3jUkiDeKI
Y2oYAw1ZNrap/SvMxl1pVFTleDtmgjhT65lsGHag7R8SAtzHFFCYXBg+SK6hCzFB
bj58MxuoRpyTOOGztcTe6SW2QemeNbvBaqyPKILseY32yXODdpjvrP/UDC9nMlVg
ZeDQeeGkZfMoWbtfPZykDJxGdZB3W9vbGx6Bauh+y2ho8I3B0jf6phSKreFdNksH
1nHiu0DN4+EcCbfDOxGn6KVBQIN57p4GfAl0iSyG84LnfH745Kn5r3zggTc9eM7i
ze1mKj3Yrg40IsDlXTK9OTGnrVnRJdT8eWg3zJ6w2ecuW3Res6LC58SkfWD9VrK3
NpjXzTIQJ9vxq0l/G4llBW4GoDMnD2I4oZmtvR2OLbocH3Zzz5TLhIxYZAUmE/pJ
oQBUUmOpqlUJnb5wiBwulYa51/gPB1/9z9lrI4D3jLFMdyyFI+34ENXQG+9bHK/I
+QMUzR1MPkC8TVul+1rwVtjz9eCq2z+sQWja6dThWdJoFiWd+iO4e4UvFgQcZm2m
L9WYUaqITQ7mROm4mlqJ9ikBPdxLV+kLwLJMZxrD71d47ckSTQ6ltAivM8ofuhro
tkF/eeO+l9bznahWfoIimOjljJN/Jk56z+4DA3MQsBz3lquGmPad2rl/c7FK94W4
VjfRYAt+Yh+7IPNQqC03J0pyPjOeIYrUe/F9XGOAn3T1YQ890W9/SJQFvb/lfhT9
uJtGxyMv3owLu4YFbi4tqV4gsz5RTFi4Dyo6NJWWv/O0WECfMqo8kvxKCSU2Vrnd
Fh3fqCDMqC1ijiDPRyfzxImCARAK8+QS2MwMVrR8hv7Mbf4NwHuCzpgs0bSVYmGB
Of7Nypr6S/TdOAqU9vlzXaJ5RNQCTgXJVJZGb3H7fXTxk5fmlSnY0JK0RLz0fjyp
t7nDfHZwA0dQvP3RUjzQcmcGmgk/zvCvK+up9nAWLleZL/IWkZnRlvMRvUrXHc2T
rGknmQjfB4EwV06TR/EpmJSYOJYh8w+qT/1eunY+YEy4h4279CxC6kROUhs/s78E
6Wi5SpXdRYUP3hCNAvWqbieemcqGks9TTIbBeO52QonjMSRvBm9N/4DsC1pBBBQv
vJyzCr39PDVKD/UdoeWjKVr+k6VXfSMb3z1hzQ9VUZdCj+brd/vBrQ/w7Ei+L7xs
8fQGlRX0mv218t7xYBzklc6WTtf8wE1Bmfs1oSXyymLjiVyn2jBQD+ijRKyqAkvG
7N9OjpYAgHsidUAGfIeUnpvgiS5g+hIPi30r0xguv0xxIU3gX8wS8CI5aWtkWGBh
doBMSuG2k+sQ7En7yIPIaMYroIDQdoHW5Jf/N7AxJ1jF2fz6LdZNUpHI/hTEvmwL
2XrIO6MQabkMXOnm0YmAY0CKXW54aMbHR9kmAgOEgHfB4RlnigSV/g+RfDqyPb2N
9MZAUqHFEIVdHqqOqCxU33ErRN0Hf5uDBtb0yMHL91oJFmmNMBUygaRtGWwYVp8l
AnZHHlPTWQqtjHlfuTD3wnAwqTxNLFpCQ1unlqRFzmzbX4FreHVYPcpmyRrpjOlY
6xBvJg+N82vEW+QriXYlfGXrwaoqxYl5m0jCQTtrF8eziHuD4R2/Gi5fni0rmuW0
L49wHUxBXT+lBOfxQ3nWjqRl9Xh2JnJG5z7ChV+syFpxEznzEDxLIoervir2yzVL
0/QRcJwiXEtPe1dmNTGTVL240ifq7HT6zxDuNUVpu3Lp2QVz1Qo4Hgov2z4gHMTY
a36WWqtQ2DEOv5m4GOONF/N/UoR8WwgLIUEF9VWesoIOUObuHfb3DHvI48ByPauU
q5wdgI1jQCuW/o1dAOd6tMLpDftyLbx5tQzkJlOJ2GS7i8zxN43DwXaAl3hi6iOy
ybPYAFHd6+R9ZFpB/k/giK1rgKUq541Pnm1S9OLw6vhQhthjvFmlOedkLBzE7vJP
zEcLUuRCmJvDxPTNMFwThvThV25EZ0NHYZc0texdQRP39rPqU2kur3d6IYcbXNGQ
vXLfeJFd/Gsw2sSnlvDW23ECNfmFKqQtmEMA+6Uk4MRkp5mxhcod8xpQTVc3ztY5
9LaRZIDqGl/Nax4CzlKoNTZM+xsBwqzWq17W4hwqCEqQswEpGinoKYCdeWj3vADM
kUtoegBIxxtTwKKIdtoAS+XFQ75Rbhz9vl4aRx3O3UtWz4kKLODqG+GhGOUAy+nH
guPORv9+ssvZbxh89DnTPt5UPSLw2OQvPjb/6G4CWglMjxI+inJ0QujHFqGRBVdy
R0HbRMm+fEp2qUH+IRfWa2JYGF+ftNVEjVDGHkez0RmhcwxnzFB6BeOJyuWU8V1r
JjK5vyCXnHnJfEvUw1YlzYfIu/PM2T+vanXiylklj680WfLpmaD0/+bNGxR6OMaj
Q58eNJCvlSdLgy4oNfyzb8FgwNWyjCVKlP01osjVeK+CHtixUU/KX4fLVFcORodx
l7a7KlXe5eQGMxvxg6SPK+dGQWO/d5tsijZBE22is89C56zeZ5TnHCTNo39oHu2y
0FyevWObL+YWoxwr/AZosoGkQ2/9hEde39b6QmRPs3+pZH80K4vf0BKafZ5Ol0Li
xQgHnQb9pHdmaYblEFaxZfbwWtEhpKVqXTBEKo8RmlEFmwd0sLMa59vtu/FR3qhD
BYqeGF4E8/VSoxVH+VI9waIxhLSa0LNkId6wZvXYJ64n0w6WSIqqRdIlj4CdvPFS
dm6bza5VXTvYAefH56gPdVV0wbvHCvyTXege7kgiiqUgChBk59+CGLIjUHRfGCXy
AAYjSw6eLNJNbHq7l9zE1tWl/ZSGQHSBIAy2966OV15G2w6aNqR9aShjYgf1CBl8
2hvp2bcTRklOL2zNVbhPn7seMmoVrKwNXJhylVe16Iy1l/k6Zc/QvQG2E1yF/zcD
nwXv0gxAAjzFwowHeqaTSHFfdsOTGWhQz8zmWPZm9Bur/zuif2C48ihyxR/2aimY
KHPx493nIIcuCPpYWPYJ8AQVMgwJGg5eO4kc7/5rWRf7/i1NNPb5xpfSmF3GvzW3
WKkgBBprNplMUjbU+tW7Uw8HfSy1Dz6BqbRsLaiNVU4li2ndwbXMvP8pyDkETvy9
4dkLZw7pEyG+1mL0i/80NY0/gc81dDurNengoknmIZSvEW6lkyzT+9UitYXO45ZF
7QiAR30Sn/AFnkWT8pLRG7rnFffDgp6OuCGuks5o0WIwVJ6AjVk8/9qDGGH4NQkU
l1OMXzDRt6rwAnUgkN9SLthVY+m1SSDSP+X2XF3JCkNkY3gbTURJhYolWRP1J5J/
pWXJbG5qY5C+oPJRwUmkus+i9UtHuuoe4e37DTOKm7eQmTsBM2Xeof5npUjHXcrg
TDfGh0qLpy8hIycNvUvG4jB2kT9cMV7XA5O0OoI6DCJKIZBXNWLE9/Z6r7RYQv1E
ygc4RYLKAC1B+KXX5qNOlhuTjs8QCKYIKRkGqBf8O1jNKFiwrY0aYF71KXRjUxzK
2iOW52ZdOG2GUA/BT2JCN9R9bVN0oGj+64yYjE2i93iaHot+HygUXBgeea1QrgYo
tkiaGTD++Y4y3V5vs8dKv9oYI5bp0cmMdQbOzKL3z4A=
`pragma protect end_protected
