`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SbL9+glm6hhM832hnwKHOs93nAo9W1wpWQpz9usI/buE8Ly+xfJBEj06YcM1jkF/
tDU26CCXxJ2Vw/d1Iu+v2vqOTKXMdj8BWxw6gXNxLNymGgO2tVeUYWtrh4kYAVvV
lr37VAWy7Ekyxy+U5rVI/DreqwrDS4qRca76A9rLDJE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
60MYd4KxeQO6UEijxOMxbL4Ov1XkR99t2T6VBmz1jyOo4Nc4thEtIJggb9AfTnB3
Y8sQorWCAqkeTPV5AW4DjRqHhR5R61iapXn1/keoZe4U5LUEoPVM9F1ueXJI5ZNe
GIdGXuFkHq+CRLYInpm47h6Pdr8nZxH+06QS0znDJwOx6Xpkr6opzISuwPiR2Ueu
QaiptpFdWPYJVt1EcKaXMDLDj1qgk29BSLa+qm0rwHuUXEhzusDSWJJMVtKmPzjq
UBGhDy8xbLrDaUDuK5m7kVKsJHSPKcG+J0NYZttK4qR0t4ZYNuFsj7gaNqQblgSB
NibR8KWhq/Ed923A7BwnxHsSnVNfMSWqox8X83pzXY0iZDVcs/7sRhUk62fcP1y0
uvsq5D5aodYwEYjtf76Y/8wKEW1ccIV/ktxxJnoA5It9tdhE+xtesqH8UYkJuuoY
jUAs1L1g2Y7AYzKuehkYC9brOEhFJ52z1awbGDVBZwEIDk2rKLRxlRhq8/fVpsD5
psAFfp3XHWheGsj1n/GSTKUyy2oq9MnBo79bQfpZnX/hjYi3VXrNYXbN0OCEZehr
6jPqfcoTRoaLuX6s+pqimiWB05JaJ/DdgTy3MFit8S5piRBCgnbpzFVZU4+QR9MJ
/HZFUKFolEDJUz91UaYdnugYruKp11TOSf05CB/xAjsvlBVEjcHhDGSWL2L15+SU
u4bQQJ3VSHMHolJC23krxrYW8Kv6UXvECYEj28Xh8A7V+XjA9zg6zplIlcMwddhE
6ctkQjsB1iJD1K558giWJ/kQx8Ku1HkCRV7h5Sw4bBeNyNtrqtgswPcWnqFS7FdG
olBsvEu4i8L7R6BZdeydoDQnfxrRCbQQIyAhSd/xfwKHqMOtHHN7y2e+hvHlPy+S
6NFybkYgOIrD6JcVWOEu45e9b1pvSEtsotPtBSe60TU5074Tv5pKfWKX+AC1bAE/
Z0vL/CKNdhXVzE+ZKqxIu0fkuS8L2TwpasrSPmaJyCPYaKMdjHzxDPchYd8cQPD8
uv+N8cW4wOsooPxeSUpBEsf/2VDGxjZvOIqLM2Xrfx4Xi2+yf2ZAPKiHA97zQlbZ
/hZGRam6mgIYB5iS8YUwJULkKzjwt7amq6SYXmbLezUItspKvMD6mu9wa93Dgz0u
8uB0hmBr3aBwTaQLvnx9gqOoc3RI2qBzj6RJmAy+t3AHa7h3xnzdz66FT+ffKlKh
H0oX0dx4fkr57+39vOH2QijfHsnNvNWgQl935Wuh0COV89OpI65LbSfhahP+CSGD
0QBaJw/xKt65EwLwhLMpeYeNGE64vyTGeeO5vwADqSFcU4IqkhY3SO+REkBmZ38e
2hhkDZMZlBODpFLg8EXEEijLqUJjHQD3jOqFO8G9hiaUKUthQz+eUuTd6itH4wuN
1js81OGS0CLfgA/8S3UhOR7QlxhNXrwHuaeIyBpqhg2ye74nbvjXo8mK7qlTRn6t
B509YO5ht/ofGfm0RVOY+ayMH3wz8g/ajUXVPplrkZF6/X6bHWyIgOfsvIgR0V68
lsuf4USamKoWhyv/Ynrweug5Yc0F9H0Td2AiwzduXrmrAKxkEQLNcOC+9uYtLlTM
DdrWWPWeMKXSJrgKdN7e5J2HXQcMp5GLK0xE/ge0P46ylIZN/0fuNNJzmG0po0Te
a9RzaAiZ/3/T87Na2WojOBupVxr2lNeo+yZF+OMX39+zcTTBsX2txHuxOjbRsUVM
1byjOiJtAoAptPDhOQrhh9r/DWgA/gjHLPv1yyAR7gCd+46xzDhmfFLb52DL7H9A
6C/CgjbId9kbFsBX5+uB5LyQI1WAGiM/1tr7VEEbjNNH138jOCOh61gsEH6HJnqS
2S9zMl25czqQvXI0My/DqTBDSQmiKHvgiWhpG16tlRRO2pyMbjm19YSqrX+JrQ8V
kZTGMTh/paKQh3e7Jw98NoTQfNUrrg6sVbv7JqA/x6v7VwaTGimCpwQjbpCYugZZ
7zO45yz0qXG8OzI9ZxiuNxhbkOAlyKDxtQ5zQ0AcGFeDRDu1ErAZ9eJA1LqSXZ70
Mm39h2QFkhOaOUo2p04JRlsRPYKdm0K2bFngRP7zwqpg13JvdhmEmJAwoGYPUrs+
dzianmrX6OkO2zLEcnGB04zGc2hcEx/Xvyiv3LnIZWO6VYkLa7opoGeFxHT7z+uc
2Kz9TuDtE+JM6iqJ7dhAAVumjTO36SZyHMYbgyOJB0G/6GlkcNLYLrZ4cln8IqFM
MioyvVSLNckccHQZcSpcEKQ+mbB0rJX1SppbLQRJB70C9rc0iDwhYvXUCMO80pWt
awH+BCkDTqO2Jvbx3HwJoNPF36DGPyJ8wK30FwNUtAviAdwFOz1e4j9zgIFX7bvw
Pn3dnuu298XOnPPq6Hkuo0i/nszmnyu0wCKlH0QbQzaD4QjOuuKWxNF1l41+5eZN
F6c1VsK6ADZG5NZ5D01lz6oBjuMF9YxbyuLxI9BowswEBcIfmr+WUJ3KcP/awTTh
q9JctQspjtGvpueSJhhPxHJw5ntverpY8WwAkvVU+vbqYS/ZNCy/B7OcMlIolgWd
WXKa68QInd7Ufdqb8aI8jpILnhlf4CpQ7xHFs85CG+OTTfPlVos4qEZKAeI/QkXs
Chdd/ah6YNOoblHBHsYfOn+tZTr0FM7XqcyFgPNVWYVhVnc26FsRZbEoSZZrCDUP
wYnVJBaVmoS7Iz5IAvK5PcSmALnv5NKPnsfi4ZsfPQ4zaYdtTtNV2nT4rJqbgNzc
qUhbRhi32X0/YTXTD0TsiQnMI7DPaJgKf7AaTcvQlMvkr5svpQVfQ+Nw1LTO7ONd
Dy72+kEwRJxvDs6IyVr3m1s421aaSB2tJtgcZZcIHsQqHd2CpZ8kL4tYD1jfDWz3
2EBTSLrG/B4GoWpOW6b0/q3KINycdXTBGUkHumox14IUw6bqQ71yXO6RiTAXhPac
vC/vif8SljSBZ+nLVAiKztFJbfLwsMTgq7q0ZEPWpTRKYtxljCvAmgksp61HcFPL
EKs8W9f4KAoQ0TntBkHQYeO3iDQ5oiNP7ZZTEPBegGJvwtZl2QUPAVgFicxW6i8d
e5P6bf6QJsvuFysbsMwxXzKZ2E2Nl5UQ343P65HCxJdVAf+QTBac9lZwF3q37uZb
xUwzrI0FBgkDfqAk1XDv1OMNfu2VaFbqyh0YDRWaZ3nuXowpttcmnFRJbiKPxT/9
pHmBFiEcjoj/ExdIlngYfbVHJRc6RywQvb3rYZppVw9HsL1a1Z814Hbo1OUL8N//
3sH/WQBuvJP8uJLZhMn88XcOaDyocePX0PAUF/OROS+hnlaTTC90xlhijzhfWH/X
DqhD3S3dUO+3nAnhiGQGgGhEDMQmGovlTH5+h5LRMsQIxXEZx3Mvv7gqw3HoeI+k
tWLqnaXeHqqBjvl42gArGff9PM90j1jJBenUgIj1Vgx7oihxqNpRXff4VLK9rq4s
TNpSHs5tiILq6u7GNOlcjn8prwf+0EUW2uwzWOrcgrgd4XfIJm3sj9MJPECZKzdD
Xoun0oCiP7AKR0/HgtyCAHdLJZh1wyMPZChfxxFYYYBs9Pxyaxd6PsLj7UqWG/qV
imn2eIYshmTX9a27kO8pZpbLMQr3gwgk8mkOzoLklEHyfvfzil/Y1N31y6salZEv
CSyIUiWOCAaaq61qiQs+dhtxp/t+cxkooQ2DIfgoP5v/cLZ+IEmzUghYMpDYhUXS
uIBcHGjMT2TixkmQsQ1nT/iElpk5Lh/NHXLm4tXv0YroRGsyGJLdfgjK4hQKkvMj
d2V1K6ixs1TA6ErQoBUAYHswAsxOh8P4lwGhDSZGyvojVHfjEtsO9qF3fgYfGnVh
+8xxBIcQn79VVYwdFEctK6BHCJPzSQgapoAx/laqC6X0vrWLT38ucpDRNR88o2uo
HsGkSLZzw398ZMTMTpzHNs1wyJSR8pLjcohs6lELH2jO4OkQuHWKOJKMSNF6ofv9
MpObuMcJtc7qBb8LRCZ4vcsR17+jI5x2DWlLAZD3Dz1S0DAPiIO88Guc6VNfSocM
puLDDcHnQxsT1s+9jKM6e6C5XjsZA0seWSx2XROiwfeWI3t9ZmPTV6g3fP1cv8XO
4gMAmZgR4TBgHE+jlIOruhv/DtfPPD5v0QKmcwnMEduerOlIDBwW4XYOr6W9mEM/
rXa+VWe4qkk+IvaSd+sb/tGfxHRKUnM4VG7/VhE2tAr9yQeY2hAZ7ysXdAy6cXA1
zk8fN+hQ1yZXSYqD8AQj8P5jNWJzHyh/TczdC9MwC63cxJ66DgAxTwY6xXutv/5z
RI13hw2x2DemYyiWXHj6kp+otR8XNlYq63DlzEDwVAp2MrLPzvxnVTE7REx28bz4
uAnMi/RC3pRySXtr1y7NHkOVNmT5aSH42QD8B7ECTrwBAzv1Jvd6wyCQapdcHBWn
B6cdqCX7n1iIHmKi8Z+ps51GyF3Jt6B+LYMvkrcLjXMTmkG0X6GVG/1wJnlR71/4
8e+YZTJVVy75wbY13FX6sN2zx5rj2pGTZlOaouPmY+4QLkU7uodhT9kJsdTOcrPb
2wOKxsPUJZpb6xWqmaWI0uzwbxVYS4Q7TpeDjK08GYSFwum+Jku1A60/qSwaHKaa
6sz/fdAui3Boxy3SQlnnuneVuNy2oulyPF/QGfc43tvTITBHOojhRm8GV9BmBjCX
Fe24GDGE5A+xHIXTO5gD8rry40EVstoqFnNRC/nB/xq6KtmhLfbDh3v0o5dNvvEb
4RD1AJzr3tq2r5Qk2bafYq0Y7YA89P2E5fSnYLRVU6FNUEbtLIMVz2Vwm0OfU6uF
KQ2R1vynVNM23HF4RrsQgUjHMSK9DRLm+bwCVvIgSRyyuj+sfqFKF+Cay1HhApv/
+K2kMD43SwGbZkJM4Z9WxcYkOk1MTSyiIm3dIGbgSD/TOWQMz9gew1NbLivnodwu
J+uU52IacGws9uat5aZRIUxw0+IIlXQP1WCrR8lKaBAejVP6oyOmXfc8VNteEE7T
ev1NqOd1XjZ38H6LTr50bsnw5W2s6H6U0eFCPGJ/2DWP3Wb8JDAu3zdEA0/leihG
E9HH+6WqJpR032Hz8fGw7g+zbWtqNXvbBzqAwRKxseRAjUsof3GVYcQC7UtFzRkC
8Du8gS2QDskyppK7Uzq2zxMYOCRnQyRwVptMsUQ++6ZWfZGsyP0GX46hkSVt1+Be
u8ShVkD7vFBMouqBsYDoz4NXau3vPOveumFXLVno287ulsFiZPn6HwxV1G2koISU
qjei98mSUkc/53fhIXSaArmRIcEDPeCphcBN9ZUF3ZuStXXsi7AGszxdQdRzYtPh
YDNWdNblj/3PeivY9EKOO94dhQ0yHAG6lvhH5o4Lylb2uGPAFptNQ985ZMtgaM7z
jiGQ8kBYyNNR8QC1vOcZJiNL7BJ/RL5HWBUHw5+qVrK7uMOB1Q+GEntRwWAPFvqZ
IOIJRpA1hS+o6zGef8/5Xo2KnjCWpknThX1U/47W5tFqq9YVJ43qUMzgK2LLQzar
hRdvBCaO9wL51MDzXgTTCnSZrwFm5wGOeww/uKas8JebhMqI/XqOsSzPR9r7ACQp
BN13ZYt6kLQvwl4SQ8Tef7aunpm8Rv3Mb9sNX7GL8EysyTd09vLq6bJG7UFE+nBF
FxXH5PFxvQVhe21wrDIeWZA5qfrdGGhjRISjJQIpiXS/7wn6Wklz1TNThHvCjNjC
FAR468z31uV6o2tO2B3sTI0UpnUo3Gt01Gq2+cHT+emtVYieBSpLkOcPQW0fJPV/
mGsncXEPvOgpAWmf1aiKLX0+LmZN8W2pbC4K5HuRDDStYUAJX/s2rkzcPUpEihug
QlBGfa18q90dvm3n6Xx6GjqWT2bpJDOdvFyKJTQ0CiQkfyT88f4TzG1xH/W9Zuta
kxq2YQ5eRAoziDH0JL8XhepYPgRVACuBL5Y59qWZTYyEkwK0I8uJ4PLInvmHgmzE
tcIQXg8MYtgHDuvAbGkwTQYaG4FtG0FbQ7MEeH6ji9G5SJazAFKe1PQnbmQ66hsJ
5fqSAKbLGVFMhK2YKQ96wwfAWnNg2/G/VPm/MuW08fxqib7FIMkRz68axbImXZp+
QkQFjx4k8ym05BMKYLXVoSzkVoHYEsepzPPitO+o7JPzs2+hmWXltmOz/iXQq1jZ
1Ss0BDMTm5nuD54vn/Npz4tCtQIGFGlY1Xb387P/ED3+r2OqZrSJTjGrSDqcKVrS
oqy0cPaJF4OB0+ZYcUtWJ9HQXphz2dgumqG4MSzEo+uh4YwICuBPNyMOzZHhaKk/
pYPb5HLcSPG57v9/FOdvlnuPTtFTWJxgSRGDGfKs/Y2bM7OK0CT6VBQsdU02IKag
NDyo118cH8I/Oj4m+CmAq4CFd8thIcHILYRluOG/LNaiVvS9+f/sH6ooSdPlwAlc
lkXd3ECIRjSQuj2fHkGqNpGam781yRdZIscRku1KcgpHx0w+18PyF/xvOXEC+xEw
rE6YrEh5I9K9aNC/ryLUHDG5xoCgRrzEKhNyrWY2ANb5re/8ym8KcKJAdz1mMsbq
jv8O3vvdP7rocVmf3cVYT2w/jSdrRGCC/vq3xhd7hEvR1mPcC/nlb1Y1WCA2E6kt
7Nd2ThEdkMPCvOVANog/Ux2tWZ6uqXVXfAaV9x8yFqLqrge0dH7lUMLl/R3jj/zD
UPnDTwp5s0pNLOUh45IEadlBn32huxG4+iR2cJa0FqYL+xzI5p+wbW5L8va86X7B
dD5bgFRTnKFs/9PzRw0NWWs04QYmP5gkc5JSrtI25j+unJOnmExGEFmx9w4DeLdN
Ay0JkP3uoBcrxfrjoqmDSQ52MmBERm4ZNN6AUEQy1JOck4m2WKl/9L88iOb64dqs
X+vHRXDkTkXIM2ZochML3iWIOHhEAKqeLLGzXmeay3Buw34yQ/AQa66TRVHUb6AV
50QESs916lF5jue54PDEkXlyEio3ajR4N9NmQ0eQWJwVkqFn5dwztKDfN5dyDloF
rR4RKtJUmMPo9FgoAaoHttjGq29ASt+DmSbi2oZ2J1jHmjlhP+f6Z+sedvkir2Sa
wTpTSon8h5gjmuVHB2Bsf8GP3QAXbwx6dk7IoTRKq1EFByj3rnXyl2HYIuUSbTYh
9QJ554ZiqVFk4LiZuGa9xTjYsa7Y0C3nMFOWiePOZv21OqlFe4pedvk3Jh84gj0J
a69Ttn/WRsV0U6panuPU70Gim+wTbzL7FNzwy7yN9NAzNmbeoCfKDzxe7tI5uNH/
JVaattNsfKJXnZDsG3APJaUOtW6D1QySOgTn8Ep0Wn+NVb2YM1vAFuUu8UDVKDbp
AzK/fM+5o/Ol8hIHokAtIRiBzTZISxZRaAdZrbvJcc46LHtY4ae7Wb7pTH7LAGGk
kZkjlXeh1YSKmBADOgIicfWuBq7YyB2jSzqnVEJysZc3mMt6A1CBgrx2AFgQC+eH
C8QxxbzwgBLK6T6kTa8dIASJv3v04vdJLocXZNQtDcx4dz2vpvnSWoQ+lmNqlyAO
q0ycpeeRgm2llZV7atQHuvW+CbGu/U9SFcLeUARuhw5My9ixaKJcPiWGt9fMegIl
b2FTEh5J1tfbWRX+yXKOhjnMPAykJQffalq4VhQOCZLFfDavMPIHk88i2Rd5IprH
BEeQzPlOAB57cI1DlrS83g==
`pragma protect end_protected
