`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bje2dWY1hVrMzBNeiTzNCfUBPS6sZJ1DtrH46mR4k9vcQwvvgZDsmeOBnt5JATlg
Bl8tQVjUxeY/aL8E8VBDpUFzblf98fCdmjri6gzjHltF+MC+0fEKc+oGkg88yR5q
tDHSszcjc/4QVUSGKrVew6xQrxwrCL9uwzrAaNuLVtQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
x0IByhZosowe9mWIe4nLWIl/Qk2asgq0G2jUWIBmBTxrgzgceYt4ZMKIs5zwXRQ4
l4fY7mfjD/wMt1U7IeT1LYrlyA9VfpsvXl0AKUMovgV1GYQsCFiJSC3YjJ0eQxFT
mwZp5nLc8KXVYe/VXkM56fj9tMQiUzSghshIwEUMtPKD0T5WWSqYBPCUPItrp6Al
t8jJoYQ7ZZtmj/8aLErXdW9WKQeOJaS9/2R58W+hDCMLktD49YY3lgUYUxm5wMKN
Bo5eBVZj17Af5gYRxLDAWlIkpmrDWyAWOvZaiX/6qx6TUD75r0+GTF1o/aAFbgvy
Y+cJMkxnhFQjIT5u29V1hyq6Dee1GVH7iSCkNDRkU5wYCcvbFV6PG0ftHzq2nWX7
3ILT+Tx32atMowkX91ex2aQvxT/TusFIiMlIJoH5cpfgi23iwz5wNTE8iAK1kdT4
+CcwOv56zwkLl2VGkn4HtsUxndFITnsy+UswNU4Uu2CUs8bakt87BG/Jyekk/se+
Ozw95Z2xYeMHsyd+wL7JARu1hE3UkHsln6Anjhk+COgvCOex5BqVyZLFoMowC3fW
e1IHvwQ/iUTSFW70HECLwXwy0Bb4VaiSmvsFqOxg9dfkr1Ah4Z98yYX94djpdv7m
9GKHvb3owbvT0JHVONFfHx/2G1iRGRxY4kZEYb5jE50RMTV4ShoGLgVj/AzIPk/E
5hrPC6YMfpPwFTHm0NnJ54338Hrq05KxzS+hGVE4mJpHFciQGaIKmONqtQOnDR2K
1fukRbU3ml2oi3xiBV/NHHQCyELcKG6xrAcAryDtZq/Psr5/NGw8QAAbKOa7KQSX
SdtkGjm0zo8KmhoEWXUipe8xMKt4jEJbFBtAf2G/XGNbwbCjzjUoss3CSKmZhxQ2
3522mSzt/rXj7ejQFiUb/nwkXwk43KebAbqNkjR7LzVKwQl9oY/6Tcz7i2bW7F81
4a1MTIhTzGPlEWFiXypksKySm8RGVXM6GHrxot7gtMvSS7Da1+CISGHgIv40Iin3
ScbJTcnrGTsrf99uO6Caq0mViUZwEHUDtpmnMfKkMlaQ0J/UR+SpTZdunm0d4erP
Ut2boDyLcVd/UYlps/aIC/gfujBBNwnra4kp6CwudrQ6YoPBfXcdH6Wx5QMU9jC9
tq2H2HYTefAhXUHXI6uz+WOHCpvrRgX/hLH0shDBPFDG4NwXvoH2aUlIORG6IEav
p+IV7vI397d1Ecn38r+BwljqIBxCXxEH3dElmvCxVzRCLdO2HuFDCRXMiiw0pPEj
rIHQKpmmoCZmfzqC9z51z4KZk3v6x98B66L+BMOtMSdx95C5aF1zhs+juMJeldPu
iBIyWO6Hg5v08n30kh3X7n9GnKEnIhpWod26XiMXmTPRATP+MAM+VBAax0zXg/4m
9Dbyx7ieQSSeq3dSUeyupPMnanTcCxmBkSy3Vw4j5jc/h51RbpFXF8+YjNYcdcsM
wsP0F+u9SaWxAsID98tl8a0zpfc9KeRzbkAkgpU5vjDJsvL+LW4LurXt5jC9KrZj
bLxG2dXwB7jINnvw4TBRsOcfdcJ2Y64HB8uL1lTWrodsyFVlpgvoODxj4F1IY+F4
fshnFM6RFHvdaSNztd75QqX1KfHMARF0yi3IuFTCpIeO0X5vZxn12+Pxce1jTuvG
c0dKPDozDiD78uH2ofhHNgdHuPc1h+x4TTsBSIok4akPUEefC05HTk7hJLztWLIt
3y0zDRO9GmsjIPQmqcVNIahpjI5l6WdaID+Og9Sq+BwAzGZ4kVnEnxh3JnKqsJ8H
k7cSinA4eHBfc9XM5NqM6/AtQik3qoXYS9j+T69vco88Z24jt9BZJuxa6n86gMGB
vtWCEJpCH/EmdLmeJPGwOCGA58CsT5HAsRUDlihFl8a9m45Ro+0Ey1GcYlEBk230
neBJ8CaR2sQ+B9uG0KaE/ATgsQjO3XhQFOdT+qJG4fHqIFAx4TS4c8EV8pzHeGF1
ngYVxsled1mPx1Vg2D9Mg832Z8ekQeMnMu2MjERuLPMbH2t/uuRARLuwRcBz8c+c
Af4+aaLhm+F4BPJqTw1bVPL3GCcVWXa/1+XqU39nVBSV9aOt0bQPRHMONny1juG/
ijHS0EJwPOwJfcBjTnWN5cWidWYSQBuMRZTMvX34HenJnqIzYorKnHgCUrfqLETX
T89jJOnGzoNrLbBDTZxiO5V8BgV3RSEV1K7VBfEfau79H6vTOnSklSZ0NqZ/31gs
/L31RbLVrix8ANHSrjeyheh+j8c7Lhu80wUDstUM8E3UWQEYF9piYbX8mUFd+eQ8
+SSNxr0a/0Loh/5i2ZcR0B07NLXwnP38bNbyJ/K9VpVbawblJ6U0erabF5J0paOS
Rp+DkneLg77iVxGnbuv2+aN6ZbupvGc0L5UqrNavw0PyA86yesD9MNUbMJkmPnOv
J5b+yfrzFw8Kfkp77FJbGyKFmRgPbTzFqVWQqJ/ZdUF8zFR0uUaKhHrNE3HhyxH/
1xKb7gvjv7GllhlWtam2AylYZEAIdaMq0XQZWm41aT/EJMRoAGshh2fseZtzdyns
5FUJ32GaXsY1atpPXRzPOF8ySvVyvof/I14qKMTFgt+z9slWhe7W3Vn3AbOkORZN
E6BijPEwAFX6Qz9C9Fb/lDZ7DbplZCzh/hJyyc37FbG1REckKV35vih82+XOcfzU
9nwLk/ruBd0pPVdcu+fn4OpDBjVYHuJwpC1MgpAEleKrf+Uz4YXCqmZH2xL+1+3/
73/6gK6hk4oQ5Pzq5aHeZDnhLVbC0z/6B5eD1cvddZhiv7++kSdJtXdtOePr3g3u
2ktmSuvi6Y/QWHkTm7/MyT/PqTaWgI+QQJTGB/7LvW39nWoMaafPDx9tzkHlAmkk
AhqK5zni8PfIA22TmGLon/gaOfrzILKPcGVon7wni+2CJe+YK4y2Hc6LYg9cVcTe
fwjd3dG9ywacnnxDnNIM5eoV+lkCe1RSHRvuI1Ztj9CVjad1Y990fvvPugtwnzLz
uX+QDxCRsUPnLqaMQlkW+7mOVnG12DkdP+JnVjJ6oS4boGgY2VMAk+wOSknbaqWy
Y9CBmwFcJrMwJoYymRI/vjCVHXycPFG3V4R2aakvLSgfVyeSzTDtBntsAGGrqqBe
rJNIUKo9kYgEecP+X7paEDVgznk8j1LDD3cCypxxZZULXEGC7CIPP1phOsEmBdTR
3nHCEIqkHJgjvSUR38a/jd9yVRIr5RM6K+rhws2E4JK2PwCIbaX7pusQutNCMw/x
xn5M2KW2jTjmMAiLy4nbOWhusrdSoMsKN4ot37Wllqti7nevSUyFNs/Msm3Zuja5
kFGEDRTDMSPj7fDqTL59z4SxWRnXGNQ2Yr+0TPc/IPnndGqGH2rGFc+EKMNpPug2
4gws0AT4a75Oqwe19BIlHIuHQ2FeBZwEn1SslqTSm9gEjH6Ol8TaxAlEKsHUZIeJ
Dn3IMeAfFkgz5uCdcoIN6JBEZgYUe4xq2q9LCyzG/tE5BObP6UCohF6j9MnB2gl/
e7QqAmr8b9iptZ7mIIasuXi22wi+9P5mq036lul3/4bHyzzBHBDKdWIKAlbLeDb/
1o+D3yFaJ71sP77+IGiwrufEtSeIEvU+6PmEoDqSBGTg3rFiFvePeULxiPNRhaHA
LJorzyYlpDfDeA813r/GRyQKwuLQDKnfk+Qt20UezPGw8wVcPEnH3rngIVKtljJY
ZpwteFxVtS+F3UABom5QnavcHWxeWjD8CHkeivWcWxUgJYYUcc/Hht+U5RVdtGxF
nDDdFQjPP33V25AfDNdd+P0Gt2hiyk8pl/YFfV2ecwcKlZyfee479gzZGtVzAaBi
wh093YbuUKuSow74Y2X9A3PJ89TVCjpWCiY6aD80hKlkZzXzY3C9VEpOLWI5T7aN
vetL54arJ92yo4o+GiBrOJLSVpYtGM63dB/lZBb5RNc/zUJwNgvBj2ZgP2ArWMsq
pz8/iUnHVYArcldhdIjlMjPMqmvKYBREBg6gvbkJPavD348zQdh0s00RZpfzqexc
v38xSvcpvz+E4NXlO8A7kCeI41c+fgXN7DKdo7wswaO3qI1n4DKnMz76/J9Z+nBu
gSstosdOu9qgrLOcLZIXbmw4EnR4JtSxkA29pjhnZqpFhnE9cyqyogCkNY/GVZyp
9B2Js8kafejx8B5krYlGMRnXB85LFGh4xIlLnwl15exrbZUyekarM+K/ktRcNp4U
bXF0F7bN4EGk4hTozdXuJvoIkbovakqp8nKYWpOhIxWG9Yqs4mN9OJoqBTnhVVCZ
ztBg9du0bpoj8J7Lh82jyPnIM9YuN4PR2+cTHdcJkcNEYTke8+bvNvZ6Mv+hVbDG
iVavAXCRFx3bjLewvTlnkhziuEXvzI3dhgsf99VP8azWCV9Cm/udMa7kfCOko9LQ
QMz/XjJobj4fGVMhgdHbbqkVPW/b39OT4wU5y0wP6xuReBAjH+f+WzDZiyO651ZI
B3IvJC2xSgXa5bb5bLc99Af0jY1H6jqxBv00UL/5UcVOmv8t/HYkIj+Y+lFi+FSP
LA0nehLlE+hWQbnc+cZAP5awCzeQ69A7fqP2dC7R0OlF+sK2tGsmvtu0YkzILXi6
a8nha4QRQRMbh9aBQrAxRgTagCKMNslmQxmITLJc2i+dAQh5I4fnIklQd74VD9yc
hCx1jmipOjMqS2MhirvkbO91ztYG2Y5/s/v7ylXcculsBfXrsVCThiBA9PF7nlrE
Wz5Q0EbXqWWN7Vr0ANNTvyMz7D/N8wnjD5jCk4CfGO1TIrBZSvApIhkaTBiYWHdb
r6L1xgcp6r1PmgpHpdvGy6WsmEN5uNoT/ojorE1nwY00dqRfJDpjU5kMf6IEe6fD
cgSPicqnWzMNXhA/wFD70TS3dD5GA1NwscVbE3AVZ95yMLSiI8WQZs2XMc3Lzect
GuDofc39jk1c80ZYdQj7a8tOo/zFGixHM4NTNpwmZg/YnrKQpk7GyjZg5NzjhOap
MRBQ5Z2D41rGE4yLSe6NIL5EiHKtrjLRPY2K22Nb0cYx6+uqsPValnrcoOKLmXgm
0rqW5S6U9D2wL4JO7c8pSJ0uT1zDiYbn30/r0A2LWLQ3qZ3+qpKW7NZxpcYC+f0O
poK5gD27VS5+vb1p4B85XGwlD/eGYwVlunp0DTyFCGujsjxo++EzflQpPvZ0Sj/E
RfuUMGdExxE/OyVbAnyGFCn5SIzI3vCvnzsMgn2Z2S9e8k9BBKUKC+9lDd0d9jsH
lEzdhtxY0cWQ1STZFol2bBOYZUaZd/znez2zihZdrW6GK+CK2O6h8Sf0ZLEnCGoj
W9hwIXIxmAG6HQOO9Tc95tp/9/LSU4H87/2tkMXGnaOGv7arKPHS8rA8Z415B78C
jTl03+r+ii0Ol8ymtc+p8tv34eimg5v3lMoyiNIjI3Ia3RlkEbE9ZCVlaHbxjvGc
bZzsvLHQmKa9ry8YVqXcAWn//Lzi6ZWVGWMwajZ09WPg0gEInRNc9t125wYLiWxP
ApPeyEnpBchOjrtNHl9LyvO15ebTdvhoeQmKkY+Lmk8Gem53bTnlLywvJkivHLrd
EXia0As8mGHHz83f4vxiX6tVIhYKJHwFBS4GhzC2B3KVKnOZIxhBe1/+TjUi4cSD
edc8q9SWAbxIE56BJs7JJrFmfSNT2lBjb0i46OM8c934vJS5EcuMft+3+Gbqhnr3
GFzvVCvFTQ/clI0e+LNH3VHL+vZVgQYks7Bz+YqZ+IdOIQDnvLldMKP0qDMJFGQh
YrpQxGc56V29ehBQcRnOrA5dpdUovQn76RN0vGm848sabk4B6/fVY1sC1Fu7JY/u
OHFy2Sd5L2+hoHUcKoZyi5ZrUIHH1lCUCg3YPzvb85bMVA94ogO39Cn8rxVUVOEp
H9OT4VRDIt5jL5CCMAtvysEViLvD8J2AOuJthDhqobTjxpJRcYCXH7y/A9sk4nzj
2mkwE3NcLG+mN5ASxpTubaseeoYs7sN8gXJR/woXLMEKk74qgW9cN6EJTOKq/kQ9
hvUJod4b2kAFwZZOLcS/XeQhexjxVk2gGzN2lXcZYNSSaOq/gmfPLUv5x5NMf14/
Hf5NRmejX+qAUcNYZWUPMcoHhakT0CRXsmxwzKsjHYIb82mlAN5vL/Nb4YshUDa6
bA4u+geGdRdx68LUpMoJ/LiBvezRoeQS6zITEFJV13Y3BMSLa35xY2rT24yJr76q
XnR/7YhXB0RhgvkBcljW0ZU5nYzKGxwm2mIB9COkVgz1IVL0t+DnTFPo80Gj+jjU
O1DVicBM6t8Qy1WJPph1UWAKC4n+4OUKhUzSZcGXPGg2CJGG2jOm9Vc3zbfpsE7K
Y6/ljN94zaS8xwxJ3geE11mUGYry4Tht3tGeRudJR+EIrx37nI3+7HizvLpUxDTN
/eLlY/EeNi9b4qg4SaGANGwnMKjYfhjFrC4yHUnntXiqQ4MW50Y8FwTieC9FiaAW
ahvVGQpBH7lkVuR/huJuaEJg/+Z9z60QSPrvNHYM/wpMwGTOHuP9DkJdu8lZj2vQ
Sw13dPpizlLP4KAw68l36Fc96HXHRUlXu2AkMxeL5BoMhqk1UrK6XD0fs1YKADxv
75h8ppd5T2cXr0ZGr9SGIVNkL1ZPvu0wI9vLKFXqw0GJN9vG8tcsHMMqk/tWiF/q
9BN0f8OJGHkvwt/A4XHgUiJvet8TE7q9au91nm/ZH7chg+AVxiyhZQcYOMHB1od5
VHZz6KfRnSOMjd6eZHXLuhD/GctHwO/+DMS89K5EmtuOmctgtO6td6TTNbTt+dqR
Is+USO+mAy5QkGSSaLcT39619T5zx6saxCZvaIhQBdpB/ZyykVnXd0RR6Gm1yAUl
qagS6szRkp8cOz1JVEjjMcHA3C8ahmhbzfYiAJmTH69JnYy71gj8PraIkfwzfw3G
wEr2UtS+aIrXWJXCdv/Xg19z1b54KZsnwYZ9BMz7BmzQ4Jux5AeEUR/cvve3HaE9
BOpJstQIJpDt8DVxj1Z1mBoQnMMnnaxuqAP32gZsb1oLJhGnfynEIila4nv0WX+I
olTpSjhdZMu8IZkY0ZLRA0cmU0Yb3b1EpINIvFev5O3IOCKpOIU2Euy5Fb1igrPY
SvdH4MXhssSTzv1uLojStBZadrdKtgFSmTbjrN13zcPuno4cEUMKsx9kaDv6Tbyb
EW0MrfGZGIa18IA2Dir/BGl0XA3voU45D7rG/RQPVZwfcUgZ8dcWI9/Hg2W3JbjD
2xLrB8XiakRd7HUdwmQLaVWoC1GGyu/aOGsf2zh8Rq/BFXVABAzxNfnm7kzAZBbu
75bAOfdvt92nCJx7f+J0UbftzistXYhRFKyBTkulRNlwBZNTJ40YE8dHlMExFaMB
SE9UH5Iu1bCDf4boQS+HGbNMBS8DcdxHPX8w8abS0x2aC7xlxByggL2ea/zewfbA
jZuWHq/ubfSMCMRQzgBuPBirR14HLKwu48UrOaKrxIxDi0rsrbBKN1lM3yyQTLyq
t9ehIixgvGnZdYVJ1SX3KXuG+EG9wLLR6A/g6w2BcY7tAYoFekoqYbfI33MyA6t4
vn/tK0kEjSooy3hOgG4QzKKaigf0AZrlEuIM1xK1cCHP51QEvOssF7hwkb28fNv6
Je+m5Nl9jjsM4XojSHlHpz2HitJdo/1QNGGrcVFD2TcQyFQFTHRkgbOF0pfhZ1OM
7w+E7qMCaUJs+nWVrpO8eM3mWb4TEMY6hr7wI4kSMKnWJUzdAgZ3L9EOVmipesb4
cMTeVUSD85qUhu7n+XUQ9SS3ayCyGI/KQ0vvFvTYM0k=
`pragma protect end_protected
