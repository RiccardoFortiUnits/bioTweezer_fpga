-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KqBOgLed8Qlp3L4ZE6O9MZxYbsiCLMoUodp46JTN2cGg4RRmPE1yAPD9Rk/QcpTk8CyIDZu40plM
kted8dldS+isTnTPsrqJbrjkce7vIfA1RbWTvel92PNx3HNZmx4WVHuJNQ8pVG+E58HJbN404h8h
WZiMNFNmaYxz2nFr8DG98plJ87Ork4r3UEWcg7cpyGCXcn7iQDb7T/gDyG6ASvsHuCz2sBDazBC/
7GTUcw8orwmV+D3RX786SjV7JhWdcWS3YRcUSkF7FTpPZboHz9sTxcLgmLX3qBbnnnhPLMfaRvHD
DsUSwCNLtybqVmVENQoWKQxvpQeieRrhLaeWGw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6512)
`protect data_block
+aZ6+GmsOIp2SiP/YWZGtzwr+L2Fo9QQXGfNzKya/UVPwuP2mwSUI9CZe7B59Xiy9EgDmfpjqqxY
T280LiiMdM9G7d9kI/WY99iX4mHGVsB0f4SBAU8vljdP6tC9lBU7ydd/dDd9vY/3DCRjGp+ikRA8
P2cIbBORrnQpQDM/9B+MrIS+pOLxfFcu1s5fxaGFcYi3V+Kq4CsDRRdWPy+LazPM+Zsg91svfHZr
PjiIqS2DnNSEDcmMfVS6rWatcZ3miEdbm1HduIGmvlACI1mk7gvleN91Y2SXT5qZbQEfPg9bCjDW
9reGPmBGMOU4ppQzEKUQDPxklioulJ86pL1vrNutN4l6TSQ+VoalGBzZYm5n7W+mlK355GitjdUY
WDi9nopsqLsO4gX79b2ucPg0EyXucSm4xv+Ypzf7U7JBij/Ay7UHDqAMEJxlQ8QmB0cEyvRW+EfR
S/U68t387vzWeazVgdJ9kQFH36FYcGf8G4367ABXN4Cs19qRr2RRUnM1ttjBJ9gTJ0c/wnb8suJf
UC/6rTLtijN2rCUeMYsGGJzhKWczRGH3wjhvU1crEVtUZ2e9okf/uOuu9nFaXU2WYrwObwlLfJX9
jKcM3JZgESoP8Vb+i1d2edVLVOr/vaOjFgiihxLClWNl1Q5xRHQqbcbpFzQF5GGRFFsnhVsYiZs/
PB316wAH0W5n0V/L8JUmY2NF4BA9oQIm6y4dzXLJ2kAP0T8L7K3H8lM5xFWr2V4B95eVXibccaqE
y4uGfZ3zaPBA4Blg9VGTl68Pn6i+skJp66gsPY1L7sShzEBnb5xYcEPs0Cv0q1Kel0YHyqMG0Anu
VdNdD3FZY3UWR2EbSt8MZrTtCDFlA+glOtaNbDhltd6ulYFPvhrXrckHGAkXOPzXBV+Ko5aB61BP
3DShEwFoj6D7CSeWH719+jbAj6SEcHLMlnyjYUbYpUMBYKqTBzTx29SEkhhnrf91OOjrLbtpWM8R
mIQD1C9ZmUIjlxANgJY6HbW6ZMCWF+kcJlnCARhFSLiFIYXhr9NrschAfSCcquovIq8Cwqaahq6u
XvBnXpnBTGaZjpS+J7fataY6ttJgYt71qRQP3PFWTt8OBRTIQGP5OB4MTjE9SzbtOhC5K+UUvlX1
5r/S5zF79zFf3Y1IZoAYRXNSP80uBvRnuy2m+u4jeHfQc+iSrkjiwm0Rao39+eMxN+5NKvJKGND9
k2yUinBLcE19SesL3eJoyqp3DPcxo8ImQkYrEbtvGxNx74dRwOhc5l7YqCbZxyd422fv84+Ih29f
dWE9FKTwLBvCpSvFgFNTgVNNBUyCSvGtE0VStVECYU2aWUzHNTeaUKblOTFnOs9uBqUwIAkPDbgu
qrAPJuFMnZ9E+fdcgUXWscVvS3VrxZzEmngEBMluVIzZmRNZcItt828+LbQl7MZ9JlmQfXsIQIGF
M7EipoIulHc2a9b0bTRl64S+oqdcP9QHD7HnURKePCu8GoHTDQ5MF60HasvlqrluOHjx/FkSJWo+
JM1UmhYSSvzQzup7YlZBwJKN5iUtd/ThcXXggNUm+FPTGPGrEaJDQf4jPft1lyeQJxEV3YXRSbqt
p8l10XqcBG1D2k1hvUJRAEsWSn+ncQx3JH9Eu9txnPy3SmDu1bWTR7+zm/aJrGb+2+OwTTCIjW6m
vkbsRtICpTPKckg40ecQNoA5xhCWkJNJKud4cNuGD8t3+TnInZhnQARvsgBq2IGkatruh9Hhu3HM
6fHt70cbAbIC6wF9I/jqQq/2AJNyum1OPgTXmApoBQFXxXACO2M2KtWsG+9KVojKzHqj3BIYXuYJ
jNPBPerzm7xWG2Kd0FqyOcEOKeiklL27EnCCrHdz/E9KqEdmNPeByfB7woAs0sZaF24nptV3WwgP
JLAWq76kEioHH69CLVbsRZBhiGAnxNrPYEdxVIJm1gV9j+mfm5yNBsXYc/yTDd2JLgH9z0rkJLpW
A0n6IhTbX19HSt3jXwrL/5vpFm25vSLyjALec3qz6eX3IFMOIppZzpnG1bzwpK/4dwzV10nygXhE
A7oZgTsv8zh55mEFQDk+eNAS80reGYWz27Z2kcOnf4/vIOD56Hx3o2+bbVgIfBgzfgxO8rttQVA+
n8JjapQbpdP9+jbn51vC6NTVZOFfLE6uB8Qb69AkALzpXbfH2Hh9Dv7mNaej94jM6xBzWBL5bAaI
AVfVbA3TpjsfhPbwcZNRyrsDveYss52O618BezWKc1g1pSzxPyIXFaA+6gBKCutb6S7l7EiHIrYh
+33cs+JGDIIcCaV9ptcIRYk9m7eYRWNvfk8c05Wpv/O8UjDyBb/zf+APa91CzNxVr5gkqOTM7bqp
g/j0oS9LopwRyl7zes5vdEReo3O+tyWO4DQ3Cjg/RXWaUIXNkaMTt1iKvHvrlys30P1RfXJIg5VE
9Y1dGlOlwoZ/BB3WCjm68Z0IVq92DOlFCb9C0QQtls4w4w9s3FBaO9boWGF4YCAPwq97KLH0I5O5
YL2lU1sOYm4NTzM4jZof84q7rqwv1gJWY/cRK8UOifNzWX/rb2bElNP1lO5SbL2AY96nPtoewMhC
NTj7A0HFU4Nqn2wUTvi8xO1h8pQRLgCYb3anz7wP7t6jdo/sUNMC3Dv8/6nAy8cg2tXO5PeroT41
ls2wJ0CQMvCEdpjqQTMnHL5tWfnp0zFmZW60SF8sChNsK6fq04663sfG2lMeEjUvYfikmUj4auoc
S0jD0JQ1zUyMvnGratY0WKFFqYelFn/yDtCqMYZtzAnEqfPmVrZUGkzjcHANq+CI7RQDeaEZXbkt
RoG/z31nd9jM1diIizWQ1nW/h/ricUx6KRpv0C1d4G0ZyMnwy0qrtNzJHtfhITVES0fTwyw7JCt2
JeR2kfapnujCje2cLCa6RjmQcIcsbUQ5Mpso9PSK/g6xzCSarP3oXlw//v1JlLKlJFW9CpBoO3fj
0jy/tt3OKOjDgClaKbX7iLW61kfBte8VDqE6jZS7FT6LB7LR0TxRBKct774nitHcwcNLmmS1Km6n
6OWNhGKvu4zPhJp8GwlPLNjCfhuQcnbTDJu9aIHhZIB+boQuSCDTNbZjjELq7oKbGKubqfAO3jeI
vxBAJtV699toRNVedt3JUVeMBSM+M1twPvCx4yVuku0qmxtPeJrq96T4ad/HuzZ4AV2TFgwDwYnK
Uh07nWHaZMF2Zy7BgHMmJyQP6d5dlCoC+IvF5C3FTkuIBlKXWQs9D4QCNT51zVFf2z+iz9PATQ3g
9svqF2PmRMKHOd7ZRyHsvGZlzdZQi9Se+ZZpwS4ejbFYUbga4ueO4NVDY6pUuVAppG++Lr2mPIQQ
XWPz62X0hXdbI4jKNukE1FCm+GGo4EFhvs3Mu4lu7DHOGk4/cNMZOzdb0dzkXAuwhvcWwoaS1fW7
h9H/6g2TmOo9+rQflw4xofZKRYTckmvqe5PU8gKsRehc/M8l5B0QnUTrkJMlkvXLLRgiRRgC18bW
Oi0j371sS5uw7Pz3N2GfhPYtQQkHbRs3awS5HPw9cJwY4lvwLxwv5bnZ3PoyzLfMwtdtoCbGjucW
hTdp9GFC7wV+r5mDyrjkIIDRRlwfEbpjJd4u5R6Cv8QctEoZc1kJs/YTl+M1/a2tdoaOdKRwlOO5
bbjLe3nnCIGminHV9Y/MaTqSSQgyoAg/TxMSfEc4MufFswr5OJtyoTMOFoPeaqrK+nWH2Imghsue
rdO0nIv/YknmWiz69DIWEkJo/755KPTr/G3bEP7J34VBs7wFfS0DsBx7bLEm9wXlGa1DYxsQYQtI
EO4OyuMS6wXRxPz1Rc21hrTmmCoU9YyBzwtvsa8ETN24HdO0PuQ7TjMV8KPttVmJ+GEQhFzSusHe
PgJWZShVrr5Qbwdhgc70K+/Zjggbr3ZjED81lCrGjOx4Xp0Rq9u+xuCppRHU7y3WY9TGvKbCa62E
bYuoOdidMbeU/fndzDSVURgLHnX+NXav92fe9Dmrhvii8272M1/bHFprnsuuy2ciBx7g64eqacTP
RNvpyVrrIRr0xfO/PepYHPcxbaU9qHEkDeqb8iPMEQSj5TqHUjD2IjNurxsLffR7b8e1oEXiOo0A
ro0I0LIIAJUwXelVJ+vUV2GD+BK9vqNoFeFqJ6aSbb/CE6oocM+HceHJ4Tmpf8Dzlk3XplQIqE8U
khLSqhwIs+iI2XPbYdWLIhpdM6ig4HzxaG9ieCBELOG8c5kGusjGC3RM4X0xyvD69abyLyUfUPTp
hE/0ncLvaDMpsyVKfNEV8wwVk5aOe60z2IJZl4EDVO1tscyrI2qV7TbCRhCIABLnBVgcCFoS8wJi
cKJSgHtVbrpuHnZ7LzFPz3qV6+rGwHiQdH5qfcBBzPdgk0KIv624h0j/llBFyjMwLnH4AbersD68
jXAHsQRvgAehN6huPR5oxCQ4ddxfybATF90RZNgwIcBbigygZcKHH0QxXwtv4PeoRTzHUo3XmZRI
CU0V9zvIpApMwo6YDzL8qpbIIGfg3QO1D/iECNphHttzGEUVG9qCzJ07pEUl8TcKGShDxbOa4ULj
kq1T2U7WhXlEXqIkbGTjP9IfrQ2MheehONF2dFvsEWpO9rFuXDvqADPBbYkU+wy9EbMKfETLcytP
cvqhbA0XOoAUv6XCIY7z+qmGsW2o/ZbhsvDm585fU4iuyu4JW54+4ITX4tPmLq+TB281rMi48Wdi
2sQwPmnT+IXo4F8X/wHMD5DbGtg3k+XXMtXuUKYMbCjtWI/yfJ2KP6k8yy/XVuVZLA9ZyXwpgRab
Hals0tHOeiHWlWC7VHXhYdOb0/T8ioX1ZApg0lplzSUE/JXITjuz+dK9QFWxqBrMZ0J+2+FVBy6B
WyoVeRo+rTwAml+B48kTVnHWjwRCzKo3X9rspBskVEV5ACql/oTmHWIiBgdaPwGkh8UgnKq0NGT4
g5ECJkurBwaBUmO6ThLA94av/alYW3PaEoUNfKiFy3A+0Dr6um6pWsOXNwf/Ot0Oc0NEojUMgTff
0mjUPZ0YGYZKHEX6JKFKHggY+sw1/GkbU3Faey1wztouAeeiqY2qxY+YP5OPVKh9ctrTxBr3hf0S
+yQARKTAzEPTHIumClOSofFauBE/FgF4tIv1RZDPWSnoRYiyyA3s4S3COWlubTn9ifAkoQrvDoFf
Q13tp1XnEUoc6IWyga1bHJ81EGwzHH4um9B3j+HCakOq4XgpTgM0r6WY1Qla0ml96Pu9v6ady6uF
YjGk7vSfHDUNItHjp1cVr6ukd8/0AV5pT8gwirBWzAQw1+/scFTlgaZNZrzAGUptpcSkrjWO9NIs
yuhiHxW/PbYM0SbRmxqg+s4WAhmr6YzBZ+aTiUMquTnpuX3K/sUqZ5pq3PFWkGkYEp2WSs/sp3m3
fd7EZpLDTGyd6pzd4rMjA9KztzQuPkpiXIwDrVSdo01sltnpgkpI3ls7c+EKMG19mPmFBms/Ed+Y
9ZwH/zxihM00ZYyT3X5hwrFJ8JW48Nd+Qkh9rK+1JsZ4G9jsjxUrOY+v8aV4dVgCBEcCL7+T9hGf
tm6xu3flfdZN8MjktxSziUsuwIUmJw2BTj0qGbkePeOc9bF4OATjoCvF+SzLXf+0baswXZIAoM6C
MGDV51u21jYf9C50WiSTCR9xIHCmampwSs/LF4SB5kk40FaDtTtuhBMJC9Yl9Z8f+CFgYRJN3h2Q
afnk899Vd0qheO38OIwmB3lu9q+eN90CZJ3x3y7cyK+RrlFLMr2qKpFKbcD8w63Jc4rZNZhst7Wj
gp2VGF1skSXaKR6wtpdv9YJgnvXKgsuhvcOeXx+NfsbVVkpEdQAdyG6V8VMmbBdlJQ3Q6LpLJt2x
GYXmrycKccWqhyPFICZW1AID2ZegRG9rT5iSbw9nY972wsjtR/l4ul1m5M0azD6/luxCZQlE9SbT
djs994v2juqqAgxJkfgZcvxC/3BIvPRBhLU18yByFqYizcf2KGsY3ruhNM4lAsKnmgALEb/ggFu8
g2vbMlW6xYlkzhrDVehVzq6nZ55mNvdt2kzYzn/UaDP8SLUeoWGPtCDi8b6itgIKsj/4xn0MH6Aq
jLB5TsDixBFYKFU77RkW89mM555kC0E7qnrmb/oFU3pYUiQYLQurlhINdN7/Fqx6CmXtVGXAdTiM
kLg/xk4qriZiR1X1sylMFXOLAOy2RT1jsid6TcZT0Kw6Z4PAlJ2+EJA2M4rXrA2zhz/sPyS5VjES
CIivGRi+qkO1yTKhPAcn16oJ4LrJqOQNnR9oTb5AXBlM9pNxqvyyhmIqTMuCFaRTXnkjndX8PECo
MFumxZvBjQpY/AbGXR3yONkO/NpC0JIyjh36UBvnKs9dO8kO1yhkIiUIOphXVEvKTknycIDprzAU
xahXU7e2FcB+ZHn48kgqzP9R5KPWrsyNanA4UxEJVK031XA3bVKKU2L/hXO19JHucKvyLr3IvW0s
sMPicYNy9O7MbBSlC+R7h+XuVBFUGWZOfjKwYPiphoFQNYbwjHzu1G1yjt1BKABF0DTOdBiZ08vm
ViRNVimSAovFWIl1dqrR6Ls/ossyWJP2qfaJHz9D9wppnPDKDFBn62zf/uZRCRZYhGK3hqyf9FWL
E/AMg5NNFJVIJMPdZqtO7Cuuvvt6J93Ey5oybkv5S9Tlzub+ivKEj6rCS0dbglIlTcyO9c/Zg3w1
ZW52L4vDvJVq1qG6mkYmbQl9F4gO2vP0oFZ0PPQ4qYVhLUMpBppq1EKgvD0wI81695ag4y+oSCvG
iCnyucKgk7Z7hTfggucD8k40eWLwflh8JIF/WYjoxjQgv4fPduohx0SliiVUP6BqNws+OH4EdngO
ZU6hZjZzGJ1B3PCLXHZU2XYuNDApVDVjYVMeTrTJGn/9k36q+eEJgq0GDH9EmQTPGL8Pzv059Z3d
9Fcx4H2sWYG6Dkv8F3QPz0lekx5lgCKoXA0nJLMakOiH9RXlchJqUrD/kFB0iETjFsMAb6BsORiB
osSeRH73nDYbwiWZPbiFWo+D/ipG8DMSnMWr8h2Z7/zhREmB/zwCamXDn+lGwgWlNcyU/9HLVrsF
c2WbYFchtaPr65uFbeZ5hr0czTvfNLzQpyy32P7pSyx0XjKheCXAKcdwVuws1Y+kLPsABh1gyDiH
WE+dKnwY5+jsLg7kE5TCeyinPLK1e2kVv2+OzsJaXeushcuIytC+aFVbYJpXazKuqZ7IjGOm4o7c
7RwwbwPlzPf9xzrzTihl+lkGDUEeKZ5ozJPfOHHag/mM9KnrVtr6TbSmDs98ZtqPakQ4yMvZY8Hj
zLB9SV53W5lk3IjDPgcr340nIDA06bjGnBQab8nVbjvFBZRDTL8/iMmO9vjmfHQo5Fsa+7OnsiY8
9aqbkyey2ZcWp5/B9NIlvKZGGk1vcYfJC1hCAMiNNHfs77YgeJSAvbWcNQqZAWaTKoVdJgV8VC8M
ZDL5wpSJKIijpTPTL3xjiMsUSLf/yOUsaI9D6Iag/LaLrk/o0+/2xHhbnc3BBaZo7lXiiVqc0/lS
HmsgPH9HiMCj6zKDWhzU4V1lyq3bawoy1ObdHERnCHIg3kM9laYs8e9ODF3aztp03iSZb1XC0adf
REOI0WtspjzN4JwU8R2BbtSVpPkvFcbgPHn70eC/XDAEMSnGkYfrJ0dYRfIHF15uPKzBW0xzvReE
7I8jwcGLl8O5yVHEE2VtkI2hLKKnf+DlQz36/2nrn+UB9l+Be+fRobYZ03X4NLvo6mSuKvLLY7ZE
UC8qfwe7GYMugqhCS/yLh3IwwO4vxyMg8NBLu4SR7skNW/ywc0FrjQgOlRRImXfOVWoSREeqd9A4
ubyyGwXhuJRD6e4aoOHqPmukf6DfsfD1YcLUdgvmGXF6AoBfhmdbCRy3HSWrfk90paCIKrTgfMn3
AnsZZwmFwYiY8PCAmB3spbJAL8yDCoHAGHCAP30s9hVzLvyZaveCS/rngjNxkfO46KB49zV/Vnhg
ActfmZBI1Qlh7XFvMddsUt0H/rN6MZDEz+DMJk206HRhr9CrSBuiKgOI73uPjHT6tdhgHe4iCrwy
9QVJyf4nPbcxEb4g/+EIJcU3o7RXnPThSO/g6RK+wOAoUT+2FE2sKE8Kp79HR+nzu8skV8NauM7n
UAzhSl0wHte3KKY+7EXASXdD7ASW1vVB5Ob9dy6l4PNVqDocS5rD+DxwBCTSfkoXskZOxrapgDBp
7sEXS5ykhNd9/WZ6Ytvx6MErw6woA8HCVJKcXh1DCccMKP/kRGvUA8h1Ewri5lybSeQzB9gQB1ri
hLJhXifJDYHVshonNbqsg+0mcmsT8Jw7fjJzNDFLKiP54IBDmta0BrMQ6yRRwKQA9EGEwr2TukWF
7FannFgTPjK+I4Ect7baaG7YSV2CSMQaPIMvukVdCF4hP/DHt+43LIPPOdEwqM3ZXBoQ2qJbSvpY
zmD6TTJqExj3iQQqcuTv/KY2CUbA02LjvqB0oQ1wMgn58AnSCdrGDOoNOtk7sTgHA3y6lemXJVYM
RWyVZNDLXN220h5Ss7G47mTIrnm4tP+4ar/nwVfkltIRJiBE2yzBFa2/VCwlFkkFe8VSByDTx5ZZ
SK5hxDGHpUS8rCzGVnMSecYpnLY31PugrvOC0Atw8o4PuvKZyj36ItXgSvFMDZhAXGn53w70q7TQ
kTU5ZbjoGubS6TBoxVo=
`protect end_protected
