`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eJI8QyX8gT5aht2tGVzniRRd08S17a6mlONjbl7U8pP8DESsDgPOCp+5AhT1VbYu
6j5tpMJGsYljTWoQ8JqyWfi+whD1Qt48kbKAV4RdN4TV9VeLrpN9DlrIY24Juest
FXVbLIs4xR0ONn1yeBRRAA6U+A2QppoNMrDVXgmjKkI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4192)
hw/8dsKo4R0zFEwCRMPlF28tQwXybVU/YdAaarcdcoHlNlswyZXrU8PYE55BIVaV
VYMKetRCU2Qc17VRxbIL+a7HbuXnFTGpG2bKgbYYM8B/EgfcIMJSP3t5ntcEwECW
xCCEp7470O9cCYbX2YbVgOE1WE5YStGiK/NUS894xPZJUwkQg6Oy0CqAawe1D5vT
tUmYBGCqRJumLVUwwYyUDxvXSxSgBxEGRZEB5Ovq6nFUWqoUAi0cOd2mXhreIyMN
JVNWuqAOBqUGjLT6+zfai4SemyLnR46tT3BiBEuxAZHIc7oDxR35XQnbv2uFMdyn
7Ql5teAGrgb11DyIJqnUJZ+JHBYqvN8U25SWqomwHLJe6WFPRd2JPK2G9DdeI6lz
nd4xYDz87XAoPFA8I2QSPAxxkPSJ99gDaB8UineLAu4mtkMW7qzPbz/0DJW7t8dv
Vb0c4plL9A2OOVN8QCIzNNQJTCZlp5qzlTeVfx0LdBtGSkLw2LZmdR4JnApRId9T
IJQmdi0ndgge1tPFKahzBgh8fUkfB25GthWbgSrDE7xaVhxOV/zz5WHCnN9zLaJV
ZORDgsa9DwBPV8V3eX0UDHskOTQljsKrvkDDziM4kqNc0G8ar7bjX4pDG02vvbzm
jJvViv4mwNL66WOOjzZUtsJMltGPIce7fHqNJjigCGC5EgztOO3equ3BJZvjrFPe
cYAdDCeWf32RhFY6qD95no/D5nFSL8tpecrBsRJWE4HThN51mo5FHiJRr5seg98e
kzxQ7yQaw8ot/HV72MbaDKUPrvJ57KV4MfYScO+mDaBYIbzPw49Wvm0JDGNlHgVC
qhHzjp5LKwMaRt/D/1uhsCwXJuGLfP3S/QXsZmshoY/UDVpajIjjutsF8BBxw/dy
hUCCSlW8c7tU9J4gcMu/J2d+L8VtAph1eP6Hmg5D/j3j+edogqJ9YJJKeavLOn0v
8D5tD3A/SuLQKTMhAmnFBm6wnnkWunIX6Maj/BvgFInG3riV9MuAMm/xgoG+8An8
BJPz6y3m9kFujA9uNi7i6XpDEmIr1acqfKEaQSDZT9oT73beR+Uz03bRqfh8ssLm
eTwsUmUp93/QgNSehOTjqhw33hLOD9kocKZNGMx3Sj4yMuwhwAODHp1YmFiZNba9
Dkipb1AK6JESH7vCcJD5Yrcip0yoUkdm+h85Vj/+pzAN/0dAzAQJT7Oy1W8/oBTr
8H9MtX/+C9FPx6LtmZpCCT8k8e1tNoCoLruJODBX755aKZKNDMFJhdjflLJ6IvYB
0lyRK6mdOOyrkO9hXsxyPJboYDbwyFHhk08UE3iadEPa0giIjC8+zkVt83jMcTxM
JzHhsxwS5CYQZD/MWzgl9wV0F4MteUmw+NGN8unDkYfurzpp2oFe4g6zf+QRnluA
4BO5ZA7cypUd8s/p0avC0YU4SAAplm/4siJC5WBgjYFAH7s6BJeWHBCvwpnAsZnS
xFgdUEkA6wJv3y8lCrZpJZ+zFasYD9nOdvY0ZZXhtpZj3bUJA2ZomE6mNEuBvUpb
jgGKiUvr7hS2rmVsbX2SkUsnFCg0C3br+TakBeDmLt6DaH8iROYlIRxmKHURUuD2
AEioLgR4c8mTMczpH2KYg+NsCSjDE4vNva6b1AQ18OOT8wgyq8uaBB/WOumIRPXY
bvZusZ0HmTYr9mnU9PSdLYZHKXbGFZIF34ASB6/p1a6w/l4qntlyZ/SnVhUPApS3
u4i3xVCqodc7bRs4JvHHKCGEnLWOc29pKxcBOdSy4XZrHSZaG3s1kxMIN5K7WlwJ
sZPQ2avbYG57K9s4mSHo7zRPqjDeytYCbyruBQomQOfehumGlZgZBpkGQ5+pPod1
GjVCss4Awlfvlje1Am81zB/wo3B88i5cAH1cJYtVUl6pqQxuBLCfroSQOdHFP74q
+B9K+7S0iuDXGvssN6gm9XmOaw7IoxFyX9wuHRpDJH/KJRO50sXK+BDuhOvovhV2
JjPmRoOpmQga5GImKY4NCShbBsAlq2OkkCCAF9BSBItRz+i2+vMvMIC2vcM2SKZ9
1j50IOYd+I39ZCbPt9KFz1lXw4jhvcK5tZHxiyKxA3CeUDWSGeDcMm6SsyZSz1Zc
DyvMgPh5t2sEWQYgxTKOgtTHjS8IfMdNxnwj/L/wwbxZiU5Ujq+D7oA5Qs9cBiRC
P/K3mhTIswFUZTk0JgAEzrKvVycBxyoPWoA97x6Lf9ckf7WBZdEDWQX8/r6rnftb
w1KECfP/yctcqTCfjZTM20jplz5bPyuFscweaRW6qx7veJTEnJTgUCJCUIApu4Ko
NpuT91uf+LSwhY/KYlC6s24U/tN4etlgnV0HyavF5UNHTC55KC52bumXY3OIzm0z
B36Le175cwQsUpKwDfwhWBAB7CLSpdt8j11Xgw+UMC1yVeTlUg7rWVJAjLfY4mzP
pYhpBSTFjuSdJJ+b2AkTzGYmDAOQ8SOApBqU77c+PXjxpBsyA3D+4u6QghW6gip4
ExdbfBHxEIAQx0yo/1Nb+vm9Rg3wikcCdUQCiX+yIujBn7yPnj92A4B7d2ah7ZZ4
QFJrGzb8IIrJDUuZsbp2EQaoa+tA/ZutsutmB0n08yiXA1IA3BSleiPS3HV5D7GZ
IZYnvcYr8T1BnWxDk1sJaKmv3r2bi6XISqf3FrgPN/4a/iMAOn8lKyzilfPbesEt
97GfMc97vBUjPAmyHoIlecGaXPYS92hCInMgsTQVEpu1L6wLl9nW3htcsDSuq5rd
l/immxPSKVTSdIbkH6N67tsNJg2VPKrT0ss4aloQODSgfqOiVA4fXIVpnR3Gg3UA
osOfJ5sH2wyswUJ03vk0v4/uBEEiPKx9dYv0HcqB8dRQRS7hdz2MAJfgoaURjDJt
9w/m2gPr/4mFphkB0EJJLpOKv6C2cDmopIkRbDo70qTq3xtqYvSAQwnkoSAMfCVR
fqlgrjHidvA9841yAhX+c7VLh72oCuPI1yfJyXJ4BumNe1cx385sC91sXwdEcodM
AksjfPxAqiO9lssbNshMZl8wVLK0Df96Q2g2XUK8d3QZtAL5RnGYENSFmEeffIkV
lo0liHiQ/icq+cn/rJgfWXYvMeECR54IvZ84qbDtozHB+GVbfRcMWirGn+AfmLyC
ryj1Or49CKibjk1sCdoeTezpNa6+EFtO450K3SO31VqTrLVBmAkIHQgSHJTjZGDh
WhlKZm5nhkAPuwcyrjdLBCdk//2RNG6dOI6OgdzVW5qgOCjL/s/YqqH3EGCJwhCN
M0X2gKkpkrNWeJ8y1LdBdPkd9siTcD3r584rxJS0KGrnoeJD2J6UV4DIW723TLjZ
2t5KDEI4Fh9zhyHQ62CzwBP89eSV2mcA4LSH9H5Nvxc8N5RM0kf4lj2U+Oryr0Ja
GZ1w+/Eg6OttE8hOk93qaywApbRAbuBJbnU801gVoF/yJWHWgROzdjl6iS04pmEm
XvsOBSLi4y52exRBzouWEu5sYhgs6B9FvTgQHVnJH+vjC3O0Z0usJFqQsd93DTmd
HmwqE7bvkRF39nM2eMEVKNOgfWmKLACQQzyhzKkcKb91Rnh7xZCGq0CThVUSZCUv
LT40yuHqd2KYdcYXg1+Z1Q64B2J9+ZSW6/nHhOkcP/blT2DkkP76daxxL/xOM9vf
ib7ju2VoP0LpQizDxq9JdRNc0DzzZe8JMMGXv62Z1UCDQ9Bw3YOdXgx0LAavCVit
1vhAbC5PW/mL/9CQClYYEW9OZQ4Ka2CLdSfzmWyMUBTYVS4ORfgEyl0xpwLv4Am2
/1YW3NrFVcwFSodeg+qr8HnG/Oj4c4a87dEi/UZmavmgTX6t+7flOpfj7E+X1pDz
oldcbiGqnDT8eJumWj463cGIb27ljsnPnYfw/PGTxUprrezG60eH8L1dHfzBpVV+
O+kgAw6gfn9lWdwwv28FIoHBpnumN6YgGVoLJx2sP+IiiHU2ywtAy9P6dQ9dtId6
3eKFDj7CnIHVrk1RWS19kQgBWAtUHef/qjnyABlogNQ8S4FhyhmOpWaoU6UI8FUk
q5J4FiStg31rgDpzYGmf9GFHhKxyoK+sx7xuqGx0wIYpFeZM0z58/VZeILD/+NWp
VTujUmXG0rzTDRbvuigSUezUyyzHHjDV4n+3gig9QLZ9vnSTyiD1bdbLP2TwGp8W
oXsQyBqlubauO7VuWBnxUJUm+601sReV5Kfle9Oyxk55zRnZ2nu5XdX2t5XfIfzj
oijNAR8HRk9AODizpZRE+OpODqIUcgqI+N0sFe6ZcUcN0FdlBwy20HvdLjIlXstV
YM4vnL75JL9yPg4sccXgX0+Nggc72VMDFrSKdjLpUuXAlLYaTtlJkzMl7RdHYhVG
D/3h74J1NJLGi52MucKucmwBTVojwWliinvawgwAGvowe6Ns+XwSmDPtG/KXe7Zm
Vp2yhagC/cWLLdAkp0GBqOmK6lYyO+dpowgEPsuPk3AWBFKxI6mjCxONqsANn4gd
F3h3P1/T1HRbZdrGmjhiCRMmHBuia87UvkQKKJlnBi4CNAW5yvQvIf0Ycg7yO7Co
4XVnKhnDmYKdArSIYrsgQbQhhukSVITc3nMlmBms+h92FcxX4+cd1M6uxwn46Q4S
eXrMeRHQPiSEO01MB1EPBgQnnUZfbM6+F+9wXqzoXBs/y49ADB1AZh91ARKyUX5N
T4j4WeJG2PXwr2jMPU+2KDK48GuXaqD0a/ydQuIKNUsi3DxphNvVJSQvyzTbqkl7
xZa225g0DZwXrp1BMmSFXSGlv6K+7655FNuwpO+i0XTOhdeHl30GD73Gv6rswST+
nm8hZtAs2er08TyfRBsVsNZrTjGYt0aBkl4NOsLK2Oh0Utdn4ureGuZN1lBxG935
l7JsgQsyRoSHZR/47AQRB0yT+wGdUOVhytBtnp8IhAxXbAch4ZvWATweLnshtdh7
vycELt3OMghANvuI4XH6LO2eZvRmxzsm7hB4364mOJ/Kxtu2fnH7QAXZ+NdD+xR3
XUIIGfrO7nMgiYpvOukExUOZBDNo12+5eSO6FhWaP1pITW6XwjbE364LVOwRV0sP
OwtLQXd/m48eu4lQxacWze0j9+zXH2ERqRuDgLeUqPo6mmcEhFgeaDRilgTqvMVO
W+puuEqtgmRPccGm2lrAMNFnsWsebkG+BOeIM/R/DGNjajTbnIwGjyEtXlkOznFD
eTN/Zy8NbyIGAzV3JvuLUnY9IbHTNQT6NHciqpXNwP5NQ+bVVPDmU0CuuEkf1NpA
VFq5pjxcJgE7x4A1YEihK3dQGiTRDkXYC6DravXz7Mr99wWwZLVB+BE3+a62JkNt
eIt1jtawlbRla5ZsnourMj3ksu/ifRV8kNNji5e4ggLaRduHUNwyJlAH6XO2kOwm
+BDmy57kMucF9HSefk+rDzV00PObk+oOLGCe9Qf/igsxbUrezsinl9wSU8L2q6gG
GYGuPKbkeXQptLF8P1wi+M6yI8kK3SBuk7eeyTL6fcRtNfTyeQNxdWCkM5XdGd7F
OGylaKQ+gpRRG6bRegWhpPF2o5CCwPwr8tixDFST87WC33hlGn2Bv0QdD9fnfkfV
TVHzm6MbWHrEiTpd1flb5A==
`pragma protect end_protected
