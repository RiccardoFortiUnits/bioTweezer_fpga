`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rnvamzxp8WQyHKk2rSZwIeKi6x4ScwKl+zc3Cs5YfSZwnji6V9uffrOfcCsJMma9
l12NkDfY8iPYhRkVbG9und/q0anIEaf96/xhyk4Ki6+lyBhQrPvvbAm0HVxeddnh
68kNw5svoLyRzklHx2SmMnLGDE4R54yptRkssvQeXSE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28016)
kROWtefi4f31vXgV76MZ3aB3WIuBWPnsVSoxpG2iA6YKRvqr97VDWAZ4oz2rrTy5
EiLZ+7enELMy0NWB38BpcltfeY9i5rDvBrJwyIN84g7/BlCT2qiH4xTEuaFBZA4q
H8qps48ej2a5mZcY060qTs/p5COpk1LtePATr1lefVwOmBdqgeZizl78Uc6UIFpZ
dRQ3XQ5a98IflEGw2vAAYtx5sEmk88o/2S+5YzCZD0pWQEwRUAV30TjN0/fHDqZQ
3IGLJKwu6SlbVOj+FGXlQBGO5pV42hlTklaNs0BHJ3tb7U0+xh2Yn8xtWFeKpm6r
B5kg9XpYtRMG8AIoupvrnXV93RsQw+zyXgkmEV2KkgBs3QLW28OtQfWyR69CTNpg
NNlGUwCa2rz2UgosnaqUP04cgFdHEHkjs4lHxf3pxmSx9vA0zWTPtWGqgejgXrOV
7Lb3+DBnll8WFozn9Brh1dJY32cik/p50cy44IUb4fCRW3O0n7nr2agQ5aaDP7FT
a53/xh3va931j/fpwTrkqcr7aHYHRv+pDlUv0XCKnWddAd/y+orwKQehv8IDR7Ss
m1fBnm4kqZzqpwgqYYLpCXk5CCfmfigj/JDZTrjMyayKh1/m92K9k2HweSr17U+m
SKoAk6YRIID/VtTOMsVg+B3kalxHOx2UYBGroC0+0wkkdSnQgL38QQL3TNQfPkwn
F5T1mWO9q/iHNcm5oGRu7HG6zjQjn9jM5x0MowegONFUKdAXM/UbM8jRmPsL5izx
Dp24YhFwv7nzsK5cWea1P4ahV+Il1Rr/49Leru3L22A2YEECaGJIi1k3uA34zbTG
ualx7ljAIq+uVVLGuxmXlbCTYx2vTrA0yrGgLJ05bGZW7ZmbnJeletiFwoBLF06w
Ac8f8zMyQM2Ut7CqEeOXw9pUrRkep4RxBSGhTF2fGUP2hOHmQWMGNl/DmOqf3Zul
EhH8vKOn/gKPgqcLs6eUDXvhdKEbByPqzATagXEW+EtbzwRWEEpK0i1GhxhSxgKb
BtDGD6yOc0aPtIffJJn4FC853XVPxeONeYSy/NtrCVzQPvv5Rz0Y1NYX7K0YmY9I
ymr2wNYrkKUKgyY9TLQ2CBUOeIug6k89oRus8QqstU4v4PIh4k6yac+6MxtM3PST
v9ElUlhR2+O3NhFcYem+w8lbUUF2+91tHnKzCnvYb0X6yt52Yz3ICWlUrJcUd0OO
zsgRabamKXGoyesB7LrAM2U8bpHH7Sds9erhOy/zWK045LM8al2M4634bkbc4+xF
4OOVToeFQ9tg9nmYXG0wCAMIRCXkvb5NM0wJ4mC7mz0zug2B876dRLZ8u4ONc1VV
tXDRrgdef71+vkiUGbeceXigUiiHmGcAFkK/3z/1CHBKU8wxPwia0oPRGiOltZmt
WmeTpPEbpCqV5TuoKmePw2xChtdbhD1C9Dtxsy7trqZWlNIQjuOSnBrc+85JQt/6
+m+rckdibmd5QwFdPPmqwa+Q8n2zl5bh0CUmHFF6OvnlPo82YXtQBY+6ibFWub5r
8iW9BCJYle4lW10LQmM7KxYwOSV5f+cxOLLsAvp9F9RPQQQZcSh9ibwvnIlNNKbv
+m1P5FGPyUB/bph69xefrNpBhMzHjeras+gX+8a5bdOVU0R0zk1BnDGb0OD0UhOa
bJ0o4SNf3IMQAgWrminxP/feBYMavCoHpnr6k+QRdR/JwKhsWKxpk9QbSkQDO6sr
sw0l2PxradFYPI+1iQCkbGBPKbkV+uwdo9hgGCxb0KqTZBhUmtfY9z4ZF4TvBc1s
elysSXlbiC6yl7VbLOwrvhzmtHGjgFkoPQ2OuqOIpTIK+Icg815s35/wAeER04OI
+sJWrOyrZUPFRekAzlTxY5uv1UsPIQkB2LtVj9EQdKVDpNa5jmyq9DwIkatcmyOz
ypc7MV+g5u46nC97dChqP2j/8eGlSdkYNGHFuVxJd268ccJewVcDL9SozEJAP4Ka
VP8V+jbN0wWi+DzkRqP4/tL320EShGRWnudGwS0AgecUp9OJJs9PJPk9gfWKChF/
puK6R80L/+yvic2rmyebyb+lmz+W2p+D7J/gpulQPebeYe+3AjvMWGQWWyYGGK5o
w9GDRUddq94v9Fh/KA4L1jcCNsfq38sWf0zlZ28ot5yp1KFzo0LO1LSiAsG32IY9
H06Lx5QJcHsQ5NC8v1xZFnP6WLu2AnxABHAl1/EFSmEmN15RgqAn1Mc6ebXigPbU
nZH8knFk+kuArP3X7HA31BYiwhtjwOhJVjH6jdakf6ac5dht3paHcxn4jqCBKF/P
bLbNcyu2ynQZXsu8U15z+ozvSj+cdyA6niki9Cgi1jzn+egLAdaJeEGIhtwkByLs
yxhqD6iDaIA6mwnU6tZUxcM56xGfduBrVX8qM+dTgjaTIpMtrD0MrqNBDVcPRxF/
mv7u/HiQJvsdS9zDBdWxSfMONdgGBnOs+dKd5jTLHSdMK6U7RCrh+pnJJyYb+PsR
e8KWsz6l7+5GgG+kBK7lUpEJqogZZdhvhkPDp/PNxzNgBBxSdanY+Wi1ap1DDndQ
7/GdfOOTE1gVwaAuU2fHWIhOAoPQxQ65cp0E63EWC3RFxkf2R2X3W35QD2yY/G5w
0zClvY5ATITLeGSaTdf0xabaCRjHecvqDPvJo7XTR6p6CUuth/+BzfraSKu+djjQ
x9NCd2g64+jIn3BeJTkGdPT2soUTwzE7u+4tJ9OACcdZshKBiloImIP0q1wOlj1b
I5yI/dCbvGiHoVuXUU3QCluWU5Dz4brL2fnz1qL5Gj0lmz10K/OGKIjj7UyY1JV3
XKsccU8scKQSp2Jg6N3zBrPatebR/A8RGHI8RB8CVaG5RSrmeBRC1VDjKfPjLYx9
Xron6tCqFu1kSm718GO8TEVZu/+VZ1tPQDVT+0eFKuDpkybkvZoePCuIxoy/p79Y
a/zS/tzLVLP/HW6jm+Ct66uaFbfMr3fgPObmCI9G1ECqWPGKrsx1zkLM3LDFVWCH
afI5q9F5LINcEJ7O/NDYn75SiFtnC0QjxuUtzOZSjnVkfrbnaHkoJEow9YUL8PwT
mh9/lqHBGkynWn35kFeFRrXvKOkMaLpok9wtFj9SJJDLhhOkHyR8AHKx0p3UPGgv
TE2bOQZ/96G8G1fSzVo9hlSL1o8+FLEzTlVDnt0DGjQOOMrC0XonOksy+OVWDWe0
CrfgtCxm1/xEr9ItimAvRQ5+yhXUFgXuqLicwivfxrUAR7VyjbZmimIqFHCuvTHd
zaAdF0+UPGKeq2d8ixfvLzRmYqZGwa9nfmzaRNuaLY3W+7ZKj2HaHTMdyN7ivA5P
IX1IrlTAoQnti2TOb1cUX40tWRBPteS5lhs0h8wZ/EVMe9ngCjPoWg3uJcoKflWt
DhYC8MUf6jOJC3tt76YbAmVAqUCCnwcPbCsSjmrCF2Oi70se/6TrAyUKrGvU49wV
7CNsO+Fj2iDnc0hgLWllb4tKydBPJa6ARGFkwCMO7MWpOfTu3EuIb8IfDiBDk+L2
7uuugMwX1pJ4l46C/diPzYvnWLQSdMJH2mPg181DwvmTCVDpXwAEX5QqdOUIyWot
Z0IOs6pThEsECrwVNjy2ZOPH28+MlgqTNkJf6l8AmrXRe/VWoD8Zkn/eoSWIXUae
Jup4RSq8HvY90Sze8pEE5CWUABhkWumiZsvWjY50h+RiO9rxdGrvTIZTFeR4R7q9
S1csg6EhbKIbO4yBFU2kzFTJYCoaynLJ4qRiJlSakaLFRH+aLNL+lW/uq/CeKkHv
NkvBbudaEYoCk2oPyLu5vcXC0Aa/4tv2kwwNgynZciP/RuBwmGUTZDBo4VVmyuaO
Ae5lXGjiiaMn9IVmSINp6us/wf/inMYaehbKlJdPdLapX8Va/eWe7kQWAEvCbP3Z
pwH0sbYQVn0+kYIgajRZ6nDZN7xtf19y4FULz/NfdMRy7Z+WhVDfS4EcjFYdFxBI
FpQAVY6i4wx9/pFlUoIUrJ5G/BoTGBHcl130Jw8JOPAu0/i5IZE/Zb5MXtHFku+Y
fuG8UGXdo9APuJe48cYfKHYuunQXMopp6vvSFcfYcoWVUTu7mcQwUv89+QwSPQ9U
gLjeiqNZvAdQtRdWW5Chs8/fkegTFfbyfGzOWMJ15KxTQxyafsaqij9x08NIKmRe
i60qeKMSxLk8KUriyl2CyR9pYg58MCKl8S57tUebHspF82h4ssZA7x7kaCMj5pSV
FanpxYGCqfzmDSEtH36XBg/qFSuaiHC19qvHFAoISm5Kvubuy+qkvXXZgnn4eU+f
Ju8uoPVrK+2awvJPbYC9ZXiRerONC7gkvSW9SBzaguXei4yZooNRr0Ly3UAbKEVN
A1EHlC6sNY8rGSMXfroS1pILVugKcfGKVneONpDAZEcp14CLVXdI5XJm0er8gMV1
OktqDw2625GW8GZqx15UxWj3S8sMsiO6EdN8ptpc6GeTBmT9H4DtHQ8WW6YkXLfX
ae6eHSYNJqJ83Dj5O+2G4bTiG6Xt3iE+u41fnw7qff7gOGP5SU+xzBxexwONXEOU
CrZFXGfryk1ZU7xSSRd62gzS+ZayL+wt1vVBMt6yn8TxKs65orldJ9K3PkFAuj9d
iIqQ7MUJ2hBTBJ/E4pZY/IaarztQUsqGAvZ8i8fXrKesHuGTLNh3Nmqzi86ZNMJe
tnIcV3RFw6+xVBTzw+2Hry8EF3mmOnYiM6lvVvTHDI9tsdeAt0xM6wmOdgqotBZy
TG5CaCeIvJsU7+hpDBzo76+QyVZx00I0M4kMHYFyUlIYpdYjyja/cQr41M+nO2gM
9ACMrKRdPlzE3JfIQQQoruhUMr/YFNCklOsed7YZErovM3u2JAXSpWaADfAjCPA8
A4arGKReJaQR7iYnMzyNyoXx9wZ6BJNQ1NzGNfiXxHNhBHWXA5/jHs9lcV0QMijk
+qWMhklNPGXllJ88Y8iIsgItJawlSoUnQSLc7iiHrs+a0oZRFmzvO2pDk0xjP2BQ
q1NiK2GyC75BvmLuI3Pmt1lwa2k4gkN/UAiqW+9giTL3+mFsnmsy/oe8kY13bZiQ
wqL3N6zu0szUM4JYIUuhNs3fGZjoyZlZ3cAsGmHCI+lE2axYBDYh3ZaSVeEXthx1
+ZpNrX6wPd/GoEPC1mmvuHT5zmOkWcjffAvylI312S+HwffDgce/F7DOak3K3+lr
P+qJaJokBoANJW6aS2Vr2L0feVQPM+E87yJrYGKrf1lvTda4gHOE1v6vKSIQEoVu
FuPV2xFMPelaUfri7l+fQKKmwYR0YXSR39WRSBrlqOqL3LYJL+90LL8S+RREmqwq
TgnfYd95/fM2UBB02oBKNNsfTJs29g9/pbEjk27e97Jt/df5x5dTcKuo/5GJrQzD
xBKRtN/2gx8VIfmzBoL7WD6/W+EdrGZN5T8OCZrxh2X1V1YRmtFiTYWA0cuy2mLY
x6gg8RhjyEGW+xkSWN7wvObzDN14oSNZ8qe6Qe9AUm4fFizYgXuuxpV/4k3JIDfO
jUA0gFAqRyJWU11n/WX+/znSOziDdlUqq6Q/0alDJTqu1J/zOD9YFi5IQVkW0aWq
fl0EP3EqZvYmQE0UIOzZLOSxsuqJuCFmV0J6cmSWBQRQ/xyjAJ2j03ljjbPKzSr5
P6nwHsGplsiCiBWNPH32AXlNBjVvwLXLnSRc2n22yqq9e2ImdCaL1/U1Q6tY1EyN
EizqH4RvLs3SRvOVx5JFRIQ4RWS65n1nbaXxzrKHlFE/xmr+eG+4ern0aLWbax+v
+0KXhn2+RpkPUyQ6+Nw35WMIJuN6nbZ4hOkyNMBRNtoABNIsBJ48GbvgEJhskTQZ
ZEas4WJAVB0knLAOz6Mt5hfo8unRtQLL/eGwJ9urWsA/Lq4NQbtRQnxVLyFB+1lX
0AgtOkqGiYtCohlgVTehfgKhmkDrch9SPnEUHPVFPZRQ2E2uR7QAjBxrGLbod7eS
NeC5IyxwCldOxHNtOE5bTqHMkc9MhnRWgbdPOaHW8osof9AfU6z8bfb5qbX8P6zg
PoQtBP/3MZfqvfbC+pS7cHe3pn08/uAxKc2fUkajv4RwNG829S0ZVK1fO36VT0OD
r4+JkZ70xRaqedcfxbhl/5YTty1bzqKRdjrXh/G9Rq/l6UUPZg+vA3nuNQ9X1EyT
5OoFCv2utSET5wcFucc99m3yApcrvC+xi+4/Vg+OOMR2HVnBadT5AmHsJcE1GNfx
HttnmKpY9rkyBFv2A/sbN8akcdKqA+dvcUDul3x5yv6Hg9cAqgzafSob42hn6CBY
ZT8TkINCzRpHB/QQ2Mm642DlaMYCwzEnaV76ytOxVHf9vBhAZfxc10HRCLksqhHv
Sm7/XFW/qB1urQC7DXKLspKzlAGqPhSk8TdPWRNeb8+TcoEeIolYbj9KDtoLM9Ou
6PHh4NjVUmtPRKcPHlJoBqbBycUsFHZH0r7Tg5B8TRFc1jAPfJU/RVam7N1EHa9O
IgLYyH9MU8fLPYjIhsmaTgCu/GMm1qyamBxMR+lVEsBIr2+tRUBIm1+/NCOjvUSk
u3PR2+8EUgHU2yFiAmGHDjjQV0Cc52FB3VOLxd+xm6qrZgPZ2xC9LY0tFa/rdYFL
paDvCnk28igEkVAS/AYNFCRFl/Ea8P0EMR0T4lxombkebZD3UcMOR6470s6jZyjc
V2EO0KhzeZmArU1nLp/SYZ6AhSe9clQQ0PQc4mkd4LpXuCphWVhbV7UVEXCDyGem
TWa7S+r/F3rtgnqU1RGVv9Omkr41gV0jHbtNF3Jr32sYmCqlGaYXzHkl81pUuvAZ
3boD21U5/M9RvPZmCqiYeIv0otoeOzwE40v4LjrVqxuA5m6TiMzdK3CD/KYlTC69
j8eebn4uBuJknpasAMC3zJrpB9lwgiDQLrhMnXNZaoxUyfP4RHqhevt3I3rRJutz
AxWFu9ujcmIZoVCD6BBXJr1TYhZFEMr0INBb+2l7QH/qk6zVsMn0W/e4Ds+SW5n/
E1onHjOeVDAiXf/53D8boruqfqi/Zv1fq5Rid8vJlRR4sjaA2si811w+97u33Blu
uWl958YAjRdFT3IV8xuZx6f6KOAHLXzIW7rLT6QUZZ+bLzP9ZITwD5F2YRnR95mz
GZuwQ9dzvyZXol3GN4z/k99MclQ+T1JQA6pHYBjhyukqHxNroFhGiF8j0ijMgkGq
f6W5stuvyTTzllzMiXz8IgxQIdkQPD12iX7iO+mYhkW8nb0TrkFCmSNBbuTf6KEn
enK/XU7gAOkt332R8o8K24FnwlAEw9rKxCz5aQOzfsHD1OTSlAu6q+qmXnIcXjk9
5Fk09KEaNV8OOu5lbEQow4zeo3QE8cVSPVpHwpYCW7qHqzceylK/HEnELfFXkLlA
qPMlluI8vIHpyfrcoy8tyVP5aqdMp4FNwOCPm/oHX8bD7rLapYrja4XppLobd+pt
FFxR4hZyQ4xFbHGgQdfOXsM3ez5upBrdOOAhY9QnNQPPZhu1GfDFyi0ScVR2Xo85
PkgNNDTZkERGgnfFAGTX0eJE0xzkDBHYPVPirXlpEf2qn8CCzETAJ/8uywpJcvlr
ITl9U5sqIchdzY31WxFCXiWeW8WYL5hsktZ3Ogzv9gIhPeyiUAkP7GcFc0k37+PL
BE2Q1Xw159W/GafUpftI+e12r8YGfwH0vVNCGnnBj1v2mAt+5c8xgI+QuBh52mST
FYwdimbfEYwwvz7XQMnUq6ZQ7oljwGfXvx5PFsNmF2tADBCNWHLu92I9Tr6pm28m
5+lcf4+PNvn2N2rbS5kIT1mAz9bgFXR71FV0vr8Y4PlYTl+QhonsUVxCuJIx/64Y
/yDNQBQckuNyV+oGT+XCUd/IRfmNWmyiWK3jAiXPlt9XXAYZl1JtqgwEUsA8BP+u
oki+Hfi1Gg+gRC9IqY3XdloaEUn+eWxf7+GlJ0K2lL59QsGKfaDhf65xA7jqj9OK
gAioF6ItU6lraPyL/tRLy5X5bhNYtsXp0Jy1UYFQcE+XtncPDkjuDEBBH3Ee9NzW
O+M2ACskDrSVU+OGmR3Ds3UgldsooVtI3nc530nNxGJobf1pPGjxA5heEkIz/iMz
FUJJjCEvBz6LKJ2n8kEJg2YUTEvjP1mFxgQBWEYP+K4CavOa9id0KrIcgqkC3UxO
8HS6H0oLEp8btCq/2TfctuRyqUROpcolTFVIhHaGgPZ1HRSX8iKFrlWD7kKyW6m2
pPR0fGBlXBhQ6jXytSJM/FdhxpVcodh93PCHlJTeTy3IUPoBSAupMcaeWEG4f8N7
cGF8HcfLLxGhLMoEdi2UPzuMK/P5euA03S4/NBOooPiF8+4JD7Ly0RGdqX4EXKrU
ieFnx0bSnZwTo9mxeacr0RkVMqvDT3p84RoGO5ycQB8HqWnvU5LiNPe39gOcTpQH
ySncdt2c75B9qKHffBSVw7Fg3PAbVHspTMWlxVTl6jEKWFTHkLpHClh5OJk9Cecp
erwjb32a7l1xOOJZlorJgi1Cz272AU9gGZwgEBn6wIGSH76qXAIe7s2Yiv4JgloB
OhQzDtYajp9awn4fA+Aojos1YZGKB/DQ1NmRi3rV2HsQ3FiPle83LnCz6Y/vC7we
lVJNRjjxW0eWDy8Kz/PWBX95O/nUkha5iSUxeMmEJRAMJnMAAW65TCCRT0nvAI8H
v/+wAGo9CTMGmJltl3Qpvypff9fslbarIqX8ecJi8SWhNxN7w7ptYY9aRFqsv4EC
IGEFqABApGlExWPtVzig23UinWe44ifdG7uN1WZwM1TekZIxZGFyyx/IadVVLfh6
QkoajwiS9xxFgH7Y3OcrLtKkPvkL44CX1d3DwuU8oHMyp8Go0WOxCRyBx3tlk4ti
hKvCwXIsfzYbpjAdLXysiNkWKzSKbVeOmDExX6M4ms8t3l6WN6di+uDmvoup1QZH
rUndpPil47bqWRMgRomhYFdhXj5vaaRqbdT6nBdhpbR5kH3e+5wU7lC5xAIlF8Lf
W0PN4uPQAzHRpqD8uzAjmdSXNovRWKuXBuZns5oznTkRs8JorVh5wk16boZg6X3m
ixNl6p7+HwxNsZrfFMZ6f1kp/+NFbc/FlrMAxs0oHAPElsJEKsUQujqwVTBfcMSj
cI5thwb2U/Ww2H58hhQtPMurt8ZU3r9OA+Sdqdw4xyw5uy3pPTzbEToKBv7t56Sr
f20Dl6rtIpnjzlh99hDpnWgITrU7Y6ixSwHpJBGfRdRyoeaIERVOItnlZ/Z9WeWB
XAvM0EuFk0Lo8DSN1E/LnA0c1brc9/A2+FGDuEX2ipAC1pG9MZKm8f7sOKSh48Ae
ol4qX2bf2EHvTtt9UVsBuw/7w25LYzUX6myw7v8Ox/+LaNl8bHwChif3YdSgiBU6
Sg2I0Is+OgDV5SkdfDOHToO047+a+Pg6G5s27hkvIDD20cE6fw8mcvUcErg07h3R
8McWZi/SsGC0o1+EMq5i6p6rHZdyGpxr/Y9oKBoJrTsi5Bim9wPgITAnxbmqBAAM
oTkMGNU4X6d3gVikUx5HeXBCwJWQCqWN2MoveYfMGqEKUpRqRwS9xgDo+kphjAbc
67Mi3PbmZpQ4+tKZLCz2tUzPJLOjm0EqTHbYtOY4FgzP0afxukeyv2H5h3R6wM/H
nVGytxqGnH3UIDIET2sqFnuTzIbQ6Yy1NW/w0Ch8SUD5C2kLOjOwiYduwtZOlfYF
2zlWLIA6h9l1q+rXxnF5hMbW/6kJQGi9wWuSnEYj7eDKoS4IE3xTCsy++O62WED7
hTVmGuQtDw68uTL4t71oWtx9zo3n8akHVX2x0+E3O+SVJXfvdSYGp34t459qPjsv
zXwkrJmYYeINpN4ixY5dyhlx9fPB79uVUTu5R/9O0OPR/rUmLlvrQOpP4iSP+ja6
okCCJo8BIXO/qARV3AzKvYMXooZNWBQNywOncz57g/P2SoLCuXU5LF1hU/XQMrCI
SSZGI6hHH11jwQePz1qgwJd/TuRxVNVNm3TkQW2BpRWM5WnK6JdaRQMOW5c9qC93
9Ho0RbzsMFWoOps2AWM77PfXvkhrQkBGqoW5HIBH9B64EiqzFE82lgzA9kQNq+G/
u8OpMiRqT1rA0o7OlE//5djF9tkOjs+97Xr2WXFJuMnribotXkT7GxQ/n1RZ28af
LCrtMdnjnKFV9S4kh8c/Qzmyq/05N+j0cK38eBGmIqGshhumEyPiOu/4i0ocx3eN
Qm/hY2sn/dKp0Bw5ibOrPthWCiQKQcPgmzZwdX9K/B0RH6Y+pzRzFn8oT1kzVRZt
lE1qFzXx7TccACt/d6S/fximnamwnu/YRedbbZL0gp9xQuSKpWE/ESWKsSE8Qba4
oxa6zmgDhBD0ieYN42EROdSSC3kqdnuyWkaAOGA96hz5kHOJ0Dtnqut+p73tted/
SvRH/4mKYx2RKG3iW9Im828eizPWbBJ++ZGIQU9B4SF0C18yLf67ivnTZkgyKpGQ
u594XZr/6cm2fKEKGHqNiibndhFDnXt+dSQvBZmVB2jCEFG29brkB0r3nd1aQz8m
Akaf0+xgzhq/WIwauXMtgqojkv/RHBiMMx/ARtBKjifZ2C3vbsXbyu0kYAQ8XC+B
ffqVhlx78UqPaslZbvKsVRioUJDga/8dEQbRPgKDgqq1fh9sQGeUj86yiXbAUZdz
TUoHQ3eT6aWktBIeVRX6kwObKwKlAOimbPuFyBEmt3yUwSK3QWl10wIj/jnA5wcl
lwRSACzNDp2+2HvZ7wcUoFmh0WRJM9m6oUxcyYOGNc/TlbXn1LLqKyjPW9usi41X
F6k97L3SFYB80AoVeWwmGI2a6kHcJhXyl6fhlOpsgFTnLQURwAJl4mWRpuVR2n+i
VAFcMtEYc+ipVTE5rItXoZ5F0pULrZaTyEPcM6m/ctrkq9sPXIxioJADogKu2FfG
UyBT49S7b3zSEo3+AXTcZ5SamFoaa6dVLjlzxkrkuGZoNcuQ1kII9hXVqcmKRayB
9Qs59z/QKa0AsUuD2ZvRlKP50n1zwa0pkNtR5/HcKM+luMqq+gMPsvYVDdvqCZFP
1gQxmCKo6GHJbgXYqiEdh+vo8RbW0m/S17ITh+S23lvN65qa9f/n7mtBhGbMrLSB
4yG5h74uRnBIaBs8QccBLOiPhoG3SYGWL7bLwgQUksRljF0tIn19Noq0SvqQ5emj
HffK6hevdyhefAP8RK6LXnaCGWXZ1KqLQpnROueNsrkrUtjb84wB2GmpkKGl3gsD
nx9qmeNuaua72hSGCT3T4Z7ectQLHs7SSFRXXiBpKJROaesLsWRM9rvGUHbggXnR
pv3Sneodiyqdsh8XCvQcFPBAZ3E4V1N8VkrRDEECcnPTcvV7BHXScCvIUfyseSXw
Leqh7wkKug2VPK+lQna8dV1H0IOLQ7NAkzKQMG1qXueOJBzqnwcWnX30XRkqizrT
6DFpwdiOXpuKfucc7/2Ru3j1UC+RaS/9J+Y1ZXwZltEFUzcv9DGeZjic/Ghd20rr
rAAANFtq7VzOgLlMGqoxMGfJvc78Pk7qJzLrTEKagIqdf/7h9sqgOtL8qvi3yUtD
4KFQSHnsewh4It/ma7pPU6xKIeYXWVSvMvy+/NRQ5fj6J+gi/RUU0bi+b36iT0jz
D+KQ9a2z122lfcdY2IMj5srOweRZZqtO+JGNr3EOvnE35IXL6/4XuUfWfDseOX6z
a3xHmywG09yI/N3xUNQcrfbP03Ms0ZfxQryFlnU7ynoed8pHnRvoZvfEYASmPZTP
wVbSfpKxcLC5U1/9CcFcO06MRji1tj8NgkkBXLfgPwyaT+PXvoaLg3cRqKiJENFU
nQZJbjGX//43myzUo4VEn7berHDXNqHLjkYxQQ/LwL1gJ4EO0HGs0ZukSYYP8hRI
X9Wk22GPQhXwb7fwys6xBbEhoiWciBt2U7eB8didGhty2BvvfJcHWEWCj1Z189YW
hKMdjlwlL/qjsrXO2nrjus3noPqg23TNPkBDwbIDyoc4ot8EZOe0OAk2NgE+mf59
UF08z2a/BrvnyHoh2LFuiSCgfNG1ru2X1aWeN3nsdwp+NCiAYZjUxzmiYd6/Bt+P
AmlNsJQtmg1TWCjZu8KFeRBi8tMY2NXOPBQTUw7pABmV9nvKbrBWKPp1DZoYI3lB
xs960TC/Ho8/XoUkFyA+X+XOTEoSEXHkJ94Az6o+E7WO/tUDlXro8WJ81GHy6EBi
EE8hWDKxG2S9/Pc2kKT7NslMaa6RJXr/QDpzM8stlCzuxICKfL3PP5lEQuYow8Q1
lUYyQPtEYEDISZm9VEQ0dFXnnPC/OKk17Jij6kgvKdpySXmZAsqjHNrelHjfxQmK
mcML4gHOu7a1yDz4v9Yn9jAKy9uKMm5oD45Q+Fp39eqhyP0hABJ6Quml9RJ/kiAC
F71O5BJPpYjqx5HZVjMcHNGTaruAK0mjscLXRXtiNmSNenjMzWiZ9xpYfO40XW7z
VUkSsQkDnUE6qq17QWjrIm4bnRvGMnySA7M19kmcl5m1QJk4N7Opv88EYkJFNOzO
Ksyk4NvWGs8wYCNLkIerq1ym8HK6nRnTPeVHgi2It9mfGrO9FKyKa5cMZK0j0wGp
F8/pOZUoLJdgLI4urCOHJiTMcnyJF9GnHjOYN2x8AtGhOzaTmeUrbupUNxRCM1B7
8BKZhdgUrba6E1hTGcPMWsPSZaX6Mc6XqscHfP6anKIunVZtFum+dk0M4GKYyP2Q
HOnmpqGfe0v5nQUlmipMWFSTkeOYQAfycBtty/KQWGYp0i9podXwdn+hWf/tDYjr
1WebKcBkMfhucAvOWWf4fAzQUb5Tkgyz1TF/pH3hKiOuQ++a/4XgDV5LtpmOQYt8
7tYlxDnzzEDwP73PQUr7cm6EG+BvlfjmO3WCJYvRkvp0olFrshtA/ZW2smuPoZWZ
V7CxTb3ESCodZrDtRUTzohYuG+Cm9ksM7QJn3u00Wcczg5Hr8p72Xd5PkgLeQ0Eu
p7jcv2oeRBLOtFC6ERhzJ/7KKv17DGsjKQWlSNapTJ7yaDaulsIYlhtgDUz5BP7V
8d1iTgUNpCWj7jrbZkbfWjA/clw4Ttq6yk0rNo77RqHZzpGpWU0BH8S4DK2Snd78
KIVL1zWl+b6BTYADMTjqgfmtOUbhCOeTl9kYRt/0q1IaeeFVyYUvcnbit8A5vSSY
/GeG5XNwx6Hihs/WbLZqNc3Um+XgfVFCOLCAZm2FaZtQg+wFA3ncDLcOkdx5dAqr
jiGKAS0jOG6gMUDWJGWK6Pn+yeE69o2guhgx6FY81Cj5dDy2ciUdJ1BylNyeNHSZ
D6YHb4KuABcWFB4Ng1vQqH0xQJlQjFJEKAAJotawYojKokbeC14b1RtCEtPNX5T/
9KrLaPcTn3rcJJRpFtwq9bwtyKnoGUL59wlvrIein35NOyEDmHRBps34epUp7udk
dppyuqtXlSh2jJSnEm7rxSt3fFSpQr8alFg+xwMAw7AkgiVQA3Y8dav30uXuBIO8
EvIsS6F/e5sMAJJXk/Qt676IpA3/FSQGaVb4TV/pJvwvK9scplaciEdoRrNnq2OS
1C7OSWYth8+80c7+MPsXnGYlk0Pry8JYRp98F61F9+WoIZEg8A7UtVcL420xE7aC
YUYOlAQQpOZISSKlRnckmG1pZR4FvR8b0yyufPJm4CkAWBop4jSF/tAqBZ2Yi059
Pmha0uuMkAZvzOec8fisi2A7xK4VJL63Rx4HZpJgYNnBOGJDMQpjHLrUuXnqE/6P
0r89q7Zwo5JodPn/mdOnvJszjkK/FlVC/cijw1GUr/LIbeXIbRsA0ePyks/U/iUV
5m6Zzs+4dOv3H8YbAJBqqn1trEuZHeNwtK2HPFRBiDOhXGuXsO2fu360r4S0aydq
vpwRxbtQ02wiZgDQn/ozGhGZ9LX3al6CMBsIg/fXsWtOItgYRV5yXHvZzELl/NNr
2ZW8OfVHAB6mkveMIbGv0kKn94ENa0btEKHEGdRO42EvpCKTXxUYo1RYludvS/BP
W7Y3FJiRuUIGTsX7Is9ngsRhfI7G6O/I/KpVVkjVvSVCvmxQHadoxGsr37ZDXq1W
S5okCWmy0WRrgFGzlSUJqncddgtVzKAHQQbRH696SgQWusC8G2xjULLtqBG93R5B
fx6YjjJqxSDP0gqC1EOEyngZ1jO0VrkYNiqg31Tj9A+VALFlKKXSph4fUb28o/2F
LDpkrpn5pEJ5WbrmzZxlcELWgR6GMEW3EUQgFJhlXYgWcFnBsiCKeH2X7L4Flyxp
i7bhSoFq7vCHSgRtvxLswrKIJgLDqAXqyfzOYOkx9mCfCKBKq23ueBrhsC4DtY/H
s6h7KgpQFoCzRBRSkGK18jWtB0ttojTo/UjAxPpUz3OakVVClg9gqygrP3isi/9C
Jb/La0wHcsqW+IW/NOan86TJxCJduskjtGAcLftVWf42geCKRxEY3mYKSIFMbbLN
gJw+PiZuPs5aLJpxoggeXx6yD6yzPhEUkAHD3Bv/iopdw/bEGVHMi2S/wf0UJS/F
dwvGL3+Q6spE3RoWikdYTpyJ6YkTRi9gK6VPHePUmqeJT/ClpVkeATEFS0nc5AvM
Ap7EKnlRJPMxUD5WnJ0Lb8RkraExy4XnmOutpf11+h8/mT9aQ7L4YkxGoRVxtG16
hbTRs8X22+kFLkDzjWb5NPst+6f2rqL9o7SkgcO8BctKomdiDKl53KadxINqKUb4
V3Xlqy4zih9C6Co6rlN0WQdh1gHqgPIbSDBBQXj60e7sOpViaMZNzKvTq8ScBAJQ
cNEKoYSztKLjubCPTYDQ8M0k9t3VoBm0u9xIqCxtJx9h8hKNnArLzDyiDh4WtnKD
1BSKHvAUAvT2GaP7pvrhHRp+/CYrXs4tTE9nZ+0HcZsfw0GDneUvxv+TIfaYM5W1
wFO4Vk1xb/fLXloOMz4U5F+XZdT2M0isup+FTyte25AJPy1dOxzAJyMRNqblAr6U
SSwr8JHNaBn18hEiyyKyl3K4ILFraPF97bZumcNMYTeMUM6ir/cbFenwmSxkoOYf
b2x584orkt6mL9p9db7xmN42uQfL0N+oyFkmkjRQSwQUmrl0nkHyb9UDYXXEkwqA
bahiZX4hwT7PRA8smw7Lm30eeJwbBMpFFGzWnf3sgsuMPD1eduN382VWyF0S0UJu
tra4DLzw57ncwGMAWYzT080uVUqCvgZh3RLjZyGfTWZugM7/ByZnJPyTRYWzo4OK
t/d9JoM9ZS/MdnPioHBaFLi/Kakqn7OwrJioCKQoYs75umFROGa2/TfssIQL8krw
ce3W/5K4nE5eKwm9K+Rdu84VaVm57rDOcpoTRSn/4DTL+zM/kBYGyNXC7T/XzW3J
hwXlUErGo188tAnkAEot2WXphcbZhIBpmO9TDMyHmUR0aC5f7bcwTCnuCgEE2M7l
BAKc0flPDV0Akvz5jTtWur7VuScwgtzzKl9XGA4jgA7bFKtZ8IY41b6Wce67eewY
v3bIGLkaMB9v1P99/P8VDSOsKLlxrCb/aY9LddYmwEAbZZbq0lPuKMQcaNo5sO8T
Zt3JGPBZZr3OlUyaUULDdb5ehxyyzSUVpcW7iaaggZA9BYDpHjez8wycSiNpzjk2
CR1hRDLaeZWPzu0QqGtCQDiBLY+nUDy55+ig9mPji0WIwttyTtzv6PPjWwFJ3iIZ
2lIjuTLfbvlYEo73u5j4poPhNt0/oCBQFywTZbdeOUWXuNVAcEB4TLfomlZVSUU0
v+z0KLgKZXo2QWKBTcXLY9LxjoEAQA0MFimBAGqQNCfrGKfm3mnEgqCYTR9SNdH7
AnEvhDK2YV+dZv7eyD28+yVUaOCdlkG5axh3c7H7+otYtPpFFMzk37yE5n9YPmbE
M4WU5Vguhn0qkcZKn0BUpfjOsVgBcUhOf4meB2BSos/L43dcEX1GOzippZ3L/Ivm
KMo71qw3fQ/dkyGkg72Fjcukpz0d9UoNhllf7+NLjU7w6Nu3vu0C/ZwM289esNUw
VYxdb9ainByqN49PuTjh8IT/GV8vZZBqX1cFtsLUKawzyHMDRv/CzObTnLOg/OA1
SaFlTNxOnIgxKfnN3J0h3CreIGGgp3nWTyoMt486auJuz2rPNNJA0HPt2zLnxKam
KMP2n2Fqz7LJP/6k5Tr3DaLSGkbU0k5KYx7CFfNM2pxpJTecZUYs83dxY7BvwUae
61aVnST7hutSiDFDvXsH/sm8cYAHWGGxGqIILxRthapKfEMet9tYQ2hUZr+t3DGo
BjYIw/JiVo2PqHbDlNZjQa2xp+WHJBLvc+X3muc2VWTQjaj9cWEa62CrNdUlirSm
3tJGJr0pqLG8xpB9JCeYZ6etv2t0mfSgVfn14GF81rp3tPXLtnj5idqrYFF2lGGp
4unbh+V4zEPc/CMKYRbNsGoiauEsYFqcc5fqOAJruWvKXwDlud4nx7WBBWgs42oQ
vMcRAOeY8+bcZ8x7NAQ2PiFU9a6ekab4l+QvscdzcABPIF/gredqkr7QrAHpSaJ0
Q1Ah3E1BpeSWdpILPQmPXVnKi1psXkr1QjXKYshoZ2oozlmiY66HEz5U0FrcuBZK
mIBdJ3l658np6tcXJFqYFglpNEm0HNmjVJcIio74O/tutvQvnADMl+h3EuU7593U
ZWKwCKkOtMDF17K6odM8lSzjVuL7cxJua+cihIqUAeiUeekhe6oxRuWk2zz6LJXD
MHeF/rFo9YbJf7DZgRx7uD8Hbcfb43gSoTE0DRZ9NsjZox24vjMjwDWbCdI/zguJ
FedvmT4gXoq6z8fT9he/1Q8HeqY7BZICb3+XlYqqB5gWdmPIvmnDgYREOXg0/qPW
LFMC1IWUDi3Yq++zh6ogaufneQT4M10Z804gUMzyTH1bQNVzFxXnIHEpyntLIXiz
7RjbeVumlT3/knyX2ypTztFkeBfJE+n3m1fB4oDSwa+WacMCaKwlVB+sjKt7e+Lx
thjibJdDlJmUmbC8gLaNmynqrVYr0u5esY6nV2Ff1BVOCkIIH4872gPOq/9jNfbi
sfupI9huY8inmvOO5oMoAqzExdmqC7rwH3aK81hcpWem7XXmG9UBlHgle/sd22yL
1BdCMhmZXDFqsV9fwdVrYwC5MkACnPxCDNzuVzkU7U/V/C7WrLzIHJxbhFdN2vcu
GIpM+kjIqpZcnpmXfyKC8WVMFFHxtjg5XZLiLFrxD3QY/wF8HlcYr9aPdMmJRLJP
2gEbqkvZOrhRPJw3EJxq5wfSH5+qIp0gQeydAaY0JumGeaQt/gtCYhU5NRrogvFS
aW/OCs3FozuPl+oVr+MfmeDjfYCnW/eDrrqYv//2sXnrED2gpE6g4H2T4ooZVoyQ
zdudvXCZOEZyclLvXCpDM0JNZIIE1ZQVFqt39aNHwHWipa6q4ZAtv6nzkL9yXpJJ
rDTpxeBFDz+BfzfYCwt8tWZT7RuPCM+jbgxRwnTRr9e/PAAfjo/TuqvyBHPxcGOt
j+5DTJEwhfFTa1uvl3+ADsDHU9uRlsNI9UGYirv8wIZWQK9STXecN474za9jvZ2A
3xCOc9xAXkTheLOFHoqzvmAoNZzFdzUs/vcyCwtAEjfSJfBGNka78uWylKP9FqXT
dImIyYWROdPkVqhjcx4o6PUlfhEuflAys+kujWF8xrEhuvV6FgvbRRoCpvXz1XA5
Qgt/WfCZcqVAHhXHuGlqf8NstrKUZUTvf00kRIVeICHx5Wo0XzN29lFQM0yZ9jHM
OwrcyRSXlTqVd3DKAFNrhoDBexWeZ/v/WkesIOZGuCitb7UfgG9mTPsQOGWEimdj
HDg8ImIOJ9E3EZaaUOjOY1RiXhJ0ehu9cKkBNmr38PWTOe8TIEFeaYp8+h4JB2wU
cAGagklgb1RDWzSWVC5zY922VRZn2k2mpMfNlQpYAsB3T4kb38T1g0iq65Blm0L7
qYEF1fp7xI21fMZDPZjtnuidUsT+XgpVKyrMLUSqr8OCi+V3ABABpYEU3NTmMnPi
EIXKx7tDCxOqRG1veJzNOB2nUIyCGZLRuc4XWMlsa+NQkokWeJxBIjDUsmP+X95k
FFfpThtP+8DoM60AMB5VxeBVeZ+nIXovbNatSH0qNtfnRABbPB+22XX5zDaX/CJv
CWDNqVaOM84+Z1imLOyMP0L3SkaOzuFUsldwut3ZRmycx8WJ1z5rKtKzzOyCV2yo
DUqVoAdsaLs29Vta2lpbnNkNNAz9iKuDudbubWjQOCInkhwJXtwOZyLu6bp4TOrq
sJVyGkVfnLXV+7R5u3x0ra0FRIJrkK4nQb0IuPMLhvXCWa6Fu7b1KeAvHo1U4JMA
BA6GU0VYBUWntd0xpyHGmgz5EzWJy0/4cf3V7qTiEyTaY1hA7duzn1sea0KRiDJn
3fIoU3i8Nj5Wque/PxJWsY0a7+ZemTfqp2tP99hHFqHp81bZVtSEb49Cq+s+VFXY
4hWmmnEAuvQUoYa+MhSql35Ky2M9OHvml9AZ7modDv9GvFsoakRLGXFsQdD86/JR
0vr4zMApTNcmNRR3FhctH0XFGfUVfCsKc3EnL9E6w0hNCc9XCuyMSIwnTa9MdBU3
IPDD7fyZhOplqmuzSKWzPzNR3lSq0YwGGt+TNJ3+CDegxkPChQSK4lhMZ3FeKBFO
R3fjAxHPALu/yXhi36EugIGuATWu2NAnTL5/7IDsE0lrv+ZCmkLRE18qTfc9dT5s
CsbpNzGpJwmOA7VoV5ItB8+GAS3Wg4DNRKVBkAhZ+cZxekFwzSFV7xOl/08vFs+M
cbfnxHXkFi74IRjLky7puUp8BwBSBLOYfJEmsjoHKvg7rFg/EREdl8e6oPGwyaoA
SihcfY7Anix9iYEGiXwVGuswfXv9YId0+n0iyna6X+xBDhgDtRyKVJVMiuTt6JmD
CfAKJA1FPvyiUWwWkZNEMw/EsqbUhx3lHhDhiMdElgPqdU4qjfDpQw8Tx/GFrn4P
AwslZ90vEEcNLzwfAUDkMuBVTdEkuG4eXBAucvEPTxuvmVj1xDk3jwk4xhzSXOxz
f7sjBynMT7xDcuwJw8AlsUJkBaP3y8UqcwW1WmJT8F/t2rNzcNLiK8HSzqR1oeYA
SKTypVBcTLr0a+7L1gzyFAX5wr9bNthw6n8ag+rCdzzq+jjRbz7sXElD8NrBBcy0
Ip17g7mhSoIpxshQSGjcBjLU6pypQ59u0XUJfGcahwfQz3OY292FtCwJyc1Wovwh
eqxpRVm37628jQEyBu7FGT2h7wwBqizu+aA3EzVS65JgOz+E87kpwgnONLxm3UUv
coR9R3yBnyw4LxiDvU4J5wDyK3OlUYVdU44TeCv0fL9I8J+cyyAzbZRYB1NzLpWM
RzPyr3nCNoTJiZpcnCYjH4tz2x2kZk2BWm4Zrh10vyTWpljB8JmVH7J2u9ezcKy8
C8brL7Ft3X/sC5j0/xqvKACJzDEgG6L+MAxcTITjLFnUQJU/zM76OBCZ8W4gM04a
LmrtWJXdKTJtVT144lQZCRZcCwAAIX8UpZLY2Dx+XQK71UAJ7ej6DVKueDSFPkeW
efqtfwV6MLvrZ0MehYkNaYqRq7Yn8AUOfuaaLyBMXhh2jbFpgxs9tbp837xmbfR4
ybKg/wJZ0hEQPgvZ/7W3RkYeHE83aP/CepVTc0rfzuupDikJh9k6wZLxG5vvNlVw
BnFdCsJ6QqdAQ6JVt8d08+GoW+JDnbq5iW8fCRQQseVtYF7Ha8tguIoaDACknbM6
MX7AGt5Q8t124JHtye3ck+YszR/CzGmZO2pFE96vDGXqxHLVtepVjv5TjMS8ZdRO
6Mo2xuvKw0ryix4U2vUOYfZaxlNxyc4OycRdNSwurd3Kv+6N7ZugqAbl3oFTxHrc
wj+PO8P65eg+Nkuw/AiH30h3CmguynuGfG/jav0icVe5ziUtHWF8itmxk1WPMC4f
pn5ws6pj/me/6oQUbOZmqEkOqqXD8eFYzoovOIyR6LsyGdVXQ2mSsiw26RVFxccy
bm2rvI/M78XAQtM+h4GseCowJfd3J2aD2EmB2G1EO2N4RSaxSTFxShizzZoF2qVM
pykmzzPRKyPJtJB59bzkbyER5joT4h0z+lpCHtuZhgQDk5iI5970xttw8gL+M6Fh
H+hZtEzc2pPhzc1Gl3jKuPsMPIdPFWyadzp9KpWtFLedclM0oM6ywlVnWMdp+w76
w5XrsqhG5YV7bA6JUvjdtXtKmKh2+attJBrdY7ScUVIfF8bLJiau0Tx1ZSRy6UzZ
RkPIvP8MTN3/gRzd+gbYdsiBy09ii5Kcy76L8YBMnnCXguCWd10lqdMOg64ktxlD
fUAv7qQ3mIjJHxdmSj4dhBbEfZ+aksXFMlR6winOx/SJdnTwhjfwcZDXoqSo2nV3
Zgw/0pmgKWBv6pQOonnpSfSGYxXVsnDDMjkIc2HYMNBFePZNyDfXs5NP3YR5iGP3
XBRd7y7Ckpf8ceB9ZWH08/1EkpjyKeh07zUpgg4PJ8ekXMwSxdGIaGTydNlRl9hc
iBuC0TesBdVCAlr2zVFqfAD3RdpjmJD9kln0XzS8RxW51fodtUal1hCHS/ICPlhj
CrQoTbYk0h+hCNZmpPeiUGWZ3E+kSyJZVXlXPdkdMRAucrNoiNHkN1Uh8Ei/WD8v
zAlf6hs9/Z6YhBZeTja3ABScVAebiRB2XF/TqXhtP38scioLC9h/KEG2NZB0MzRX
GmRCiglTlhsSzyXqGTC078aG7KH4QcrrEltoP0J9VYQeR8FLESjFFuknNlTYgv7w
MqMB+lJXwJYniv6ubPVDu+2Jer08IbDCpl7eYn+rxYLINimhF3K7qAnW++As2/Uy
eXubB6RvWVgphP+xuH5fPr85Gpue3wdieY4x17oxEL+nmR515+SwcdGiAX19dY9E
Szj9AQrZU9IxsuZW2lgCNzuZeYKNPD1R2JwK7JYbZS3b6HzoZTYdhbwvUlTng7mh
cu2Kdze5Gj82KC8jUHdb45NDOky5HiFAH5d+BodFcTITXxxqt4CEmJbLjptdn9Jh
LyiJMeZ48hb5++NFWBZjIr33yN23lRs3cEz7zvIk2HEfQOXsPk0PyAienUkFsBui
C7DvKtp1tD0j6NfM+uWN9wqplFci96cu+jgvSH+Z2dRm/bqatTatHvjSe+BsSe6t
epIgLOpIa8WuZxjJbarocAO1MLXkCPM5OFLc33Vs4VmmdPAXtGUMjiXm3I17nV4G
OjUlMZ9WMg3jIZ43ch8h/+VhAHh1xN4tKXLmCaJosZUDnzF0gJx7UdwMd78sR0eN
6aRUrO9DcUGD8NNiDMghyXDn39w/5Qp5NgaiKo41wDmEpzrI5Wgnfg1LecCz4S/j
lNCFhFKagqyRbUNJBIYTOQh4zUziFl+U/Jbj4CTw8fKtp91eLc6EqLXsBUVpHiCG
10gPGKes8GvfE9j7u0muvZqGtc/x3G41A//UqFBKS68+rQL70Lg8FsnMbyM/4Ae9
/ZVXWBnCZicZietyIcXs+i4jgGSxcZcozcJ4U10coRS04NQqxAVOeQj5E2bH0NK8
weWq2vDuD0g+KuL6onQ4Gmqd8hMgMN6Ejrxa4pFt5XGwO8sCPmghwLm7DcZOOxtW
tz9Bnhi1LKgFRoHcQPHy2rF0MHATLKHld6kBaUttsIeBqWMbqT7pOv8DzA8UzcLv
eG0mgiRQwnpn7T8QLrSivuBCZt27uV2BHC1XUS2llsV//mfI0GVCh2O7jgvDtAUB
PWk9bQTV4bDJpr2vJ0IXftdl/tyCFGHVj0MBoARyIm0MHVmm8xhuO6AvJxfvsTo1
bdNhbGCmqOS6utmko8HMkDuu/YVAYFkLlvWZ56bF/Q4sUjTqSit22pVeGcCD/0H6
lm8o8TFbksoT/YBlUJMWzdu/iNxYzSWPe50zPKmR532EN60q6BT14RI4npVViGeM
mhu1y6TUzkWGxkZ+IrbQa1V9+IWXrHkbqSINe49admTw2FZIlwV9ZdPm0aACHumD
NJwShk4ewEIOQ/jzcjAEkFOKpwOcgVI2RJgPtnINme9nJpAR3yRsbbR7N2P7VnF2
RocD03ykoe/vSCkbcELInEUHtqd0Ixp2/ysOJ1poUldIn4f6XnpTxT7bR0tbX0JP
yO/vXcFc75dbojAFKtqqf+DPLzxGfxHJXopVjik0HQElQi2zY97h+O3E2OdODq40
xfhgvygPb8vLVhKwFZ+6gbk+cG8CMUuS79xzuZbIGtFeIcuTDHxBkY7q8ZTOwC9w
ha7T5foKqE4InnezDWSBuQ6IuNP90PUTUP0ytGQi+5ska5ElWjR9a/C4Gti3/TPv
Gn30aOgc1hWsNyg7CinM4ZUIDX6IyxeMko9nGVF1iUv0smPMtxuLXQqMaBuylv+w
R+IFZmTcKmlRyf85b7dSkNTvFaMgo+yZBUyZ1f8U7hX7Yhy76rzInjPm2FBht/0e
Wx3/sNSupGKCZ7rbAdbQu6DNA0hhK8VcgbbGjNeAHgcN/ZQV2wIDAMNu4JO1Jpxi
7s7gw9e0u97+zYloi8NBTEUZ6lMshvqxtfO/WGnKYuAfEUCDd6jNWEk2phaK74eN
Sy/QQeZ4bbOFgtBh2hXkeEAaNDZsKftOBJYcYZJtrxedVCRSNgH8Ymn4+7QlCBOY
bZATpu7+6pVE9f5/pMSYzckpHxouKXr6QGbwPLbhVdPI3BJAuDJ+dzrRjRhAmsU3
q7pbIc5xo9eBMejviOCqlRxdymku/JlIx8sKmLqU7IQ11b9pRd7TD9CCdJepirXj
QsfxzzxE3fPB8mYithYL8NtxayL8UB+ZO7/fzpwnXAPsDAVDv4q8v6NPfIbL0MEK
ZF4YCKfxw1M1EPwrLJqNSn44AmnjrJSFjna7SYdUu6iGp6gAUNvW0qgtfQcFaby7
Bb7Ocp/Z/ItqK9hcQudTSyBdPMbnvvTUsaQZyNGgsq+4uaTBuRXSyDVWvy5k+/zj
8Dkz7ijUh6RzKEmF+hV6KbjpczduaXJqcU0wmgfA7+axNzaWHYNnwacRYBGkyapG
IhmQGJEYaPd8zc9+kPu5GLbRrz3S1wN/UsO6+i+gpF+NrGOH2xnG5o+ewFG9ynY1
RXO5uRfDjLYB7GD9MP/4p0AhhDvWeOVYCG0piyfmCY6jlTaL6TIDveLp0fvtxMwv
Q/x/ECMsem9y6xVh/Ts2hDRXZHRpCaOwSKui9SBQ9qare9z8TnI/tnWJgTD5A4SJ
j2Leq7ngceZ4Bt5XQX1TVGUYKoc8N5CP/nOn7qo9HsZLdGxpUg/+tN4lApcIUsCm
p8qRmq5+4VjxgWR7acLtBd4BFASrXmohdK08EAs9DqojC8cIR4PBoCBeVhfVKr6E
dA2KqFL588wZQ0JpUjswXCTgJi1E+FNbVVuQPoz4j6A/hWLAWTFTuznLQSRG0fNw
QBvvBo2/yY59SUDaxYG5hACFS6zNx81lG5JXP+OVq/RZerSEwgBMAAlJ5Zd+NVp3
Bbsl+G3F0xrv2XfpgI3CEAUg7baOjya3r4QnI8x5AeFWVecFwUv+VVyKqLFbkcKZ
W14s9BsOYiOXzEEyTf0OcJhXjlfJP6aAmvzlE9Njyu5GknGRrWgUc/w+Du+5a2z0
eF4ZsFzVRSyT3EFMeFZ/x8nivzsxRjiQkDy5E7idd4hm6x5QLi/epAP5WHJMLc4Z
3/CSK8JnCSQfcmOZltb69+qk5sQdDltCKCsaWQvIPCsdv+IWcuOaBp1HmE/7CsIA
OvbWObdg3T0JmxPtl6KCS/ud0bT3iyBww3lqltF2HZeVuvoKrlFnUETPAg8Uyp8R
z1pPpaKy79/PC4jQd1l+6RvG3m+WcZLZwR1XTTfZmL7Uoo7L6jU8DuiiopInsWpC
3ZHLmGFK50aPX2YPDG3GQd4NOO2Npkcj5KMZkfxSiQ9tOzo6mzkQrOog1cdvyiJx
fyP51at7YRvC/hjp7Lgids6jfRS5K7GibkNijjjBN8cPEb+GCjTrwU6ej3zliK/S
YCOoVY/n7F+2XfiXe8ZikGj0aqXfu/NYspuehTPZi8iRQKOsm7/IdPVOsvRCOjXL
HyIz6IZuVrja2N5HaNGChRzc1SQNsZRs/7spSmODMPWGZB0ADr8bDCgekGjaYAxZ
wXMN07DJadRGhz3xZaVNqO2j6lohsw795p/IuP83K2PeC0ZNEJKGi7r6I/iM/Aoo
zbXnAo5JwDeKY8Ili+zunAEFdRxZWExsDTmq4A03DCz1d6g5UBFZHAqaRAE5adIl
iROZR7JIH3VXwoSV38FBc6tn7WDuGxDQ7guwEVR3KYBjZBnn8IFLJhn1N366nNV0
PJoeK16anhc+9TLLAlLK4fL9ElrcD49C6sgucaxkcFQBc1ql//gCL0Y8YeBIVU/3
NFe09BI3gHlHNVHV0I6xNFCSFFlV1/kZyFtTl/sGxYonSwaUIPQY7ollNVqO8Gjj
dHiEDngCpGMyJBDoVoK3laXudND103YHmSmdImGF0ioUTlTCKqchRT8eABQfcUI1
S8uwkzyCf6cdikTrzz2aTxgGccj5a6PHRUpSE1t8KFzXFBZ/ZaVjWlk04nE5rN6C
xNEoErygjJ5lxOGTdCmYM67zZeTKSmLfXAEzw75Lbu0LJnh0dm/scdRzb7fydSnq
QBMGdGGSN1J77fO+5poCVj+xolUlydZ/Kys+3bNaXwwoYPnlYCUJvynXEKHt9YaO
75FSBOtgM7SGQBG6k6we3y+isc7cFl21bhgUVZqDCS0q3MVjWnlQLrdcJLagLnFz
Uaro8FROQ/sqHYsu8rynY5Qr4khXr6tfOjXyBMpgs6Z1mqgWPHe67Aepbf2xnH9b
dyEpPlohYk16EkE0matBeUKT94ozFH2K7S0EEicN3IVv0jzLGTh7n8FeKGXJhMW/
AGvw3FTVjfZu4SGAxsBS4snV9M/VDH8XZq7sduZuHI2CHIyuqTm6QDfRJqMnPgo5
loMPR3F7u9+1svg460xftPwrJuQ04+yAI49B0mJXhKH+AuEi+fo6wzYnHe4ABekk
BLxhMB9ChFvjtMAe0nOhBZ/d/uoKd2NZl18MBNR0tcX34akTB6AEJFxZj2DQn9Aj
tvJMSj+FaTFD0RIOz0FAzi7er5NUOkxlOStrzcxhrrb9TL6H0f2p7cAqaNhkHM7T
0QpTqg765i+BbCd9R0VKDhHEQK/8IJmTq0/23MwwUaqZws/z16ZSUZkAlZImmkb7
Dmly3bV4F2ZJEs2HRrlRI+wO9TT8dkPH4TezIalVvb8G1CmNcVchiO8LOlvD7/q5
amsVLDgc0yjmLablJXzWJ+k/WjYMhpq4fQLywK5kDH51lR7pseaTs730+rzh4amN
1XhinwnNA6/LQMf2RUQH9FI3rhnNfJ4jp5MdaMXQvQOIU89lwFvHORvcZMuqtM6R
oDPJ+kPoHX2uY0j5wohZUkYS38Zd4F8Z8LYDTfz7lNZP2gdRQtjwbUoK8JFggw6j
VkUBY9hNmLfYbNVcb/BNsgxr0LpP4Mg1K1S2tpxqEItLaO5NsPgi3WJKC1KOnnOk
lMeEB6ospO6aCGQ4mzb65rxKs8/NMv/XsA6L9T5ZV+f833d7CqYNBNCn/PpVR78N
QUdFEFORt3+Hcg8JsPYWMDtXxPxPdInzdsRqLfYg/RoG9pITigvwgwN7o5GIeet7
hcvZWjWGR1ZqrQIf9Knq8k1lARgmhiqQyxmV7mlnFwML/ro1+vou2ERBkbAyEqzu
AkGFYvdo0RzgmodFTmn2Xn1nM5LqEq/4UVfA1B7nYAvvGcin2pcMugD9HAbmXRNC
J8PugB1xuwbdkng1ujnzCLDbyWkz4/fdJve2J4Yq/R9Ngi+ljUe1IOAyGrHvVh10
skVZh2BfVxBdDr7iFw1LvnMwr083gsg1uxasv55XbvG9puQZdwjoAinSLnyQ7O1K
mPyRgETEz33heAsWE0DL0gtkz/Dc7T/DNLlNi7hyZ7S+PG6fPrFvCv04bakIpRE4
2v+c3s8hGUopOw+3QWOuN5rzstrU7jq1T9r97XizadSiaRbJIO9sUy6gOzlZIhZI
D4E+P6y2CleF2QnEyt8nbUVaeZsPjSvp7bvelp2/KSfpJOrxJamXJiWZqPrzkm+Y
9YWcYVb+WXQf6Rte4ftVd10d7yE8cnRWsxRD3Sds9gcBxm+59Kgc43pnOClH8qiD
TBeqPstoU6fq76RsBoJykrUDPWgbEZu84BaWYUmVxSDGcVjIfEMdOM29uEdgl2Rp
WPrJnwJFD5CuVbMNqEomT2umHRu5f1cUXW0lGDrnR316X6cuBHFpUpDSmVWtTLiM
ELcuNLxjJ48L2Vh++sFNrzok0od+Wxj+gB6jBx8mnFIYMW86kTRdHbW+Pkp00+/Y
WkIQjhjga5yMB4XTNip7uYwR76PeiJ0qQpSMNRzjlP+m04SMqCGkvVJwqWChDiia
9ZAfGj4y41hTtF/8eb4ouREzrIgpglf4ZXrrN7Sm++hg0Mc+QPimiRx3gSGClUQb
WmDmG3r40p5JaqZycq0DKSxhalVu+ze17+UqJqlbqjm42Vmyh4UF/z6qynjjqA8R
i3Cm+6mbAagsZduKVgzlk3kxY2XHUJzPo4szzFlSD4gezICchlhuiHuN593wft/R
SKietQaVI1ESwLSrjdqKaBBeWKnjXm7v4ZT0Lt2ggzGuVceedWw9fDMbwrwnhPlj
gbTK/xPpNvlgGuySFc475L8473hkzP65/CeNSdymjZxnKupJ+jTWMtmtx1hpulxd
LMMaSh7BgfU9G9+mXpciA4aWimpAb4xIWp+59mtRPbkYzMm7tkwcITW3sCjXChV6
GisnS/heMSDHmBHiZsc9D95jKOCK/wiHQGa9xnKBT0xIqo0W+VZf4bE5syEpF5Mb
vyg+KEZwJW41ofxPyeF6gP6jPhnZGu4BUynV7Y12j0muSJ1cp7ArfhncS/c2wZja
QNE8z5ptxyqLyjKSdrsmgRaDpJRGCO8cFdd/C+PYNiuLvYxjFxquJygJqBv0dTbo
6lBDhlxca9RTLBYEseeKeJEUErR4jWwIHoaN2SEFTTk6ukRsdeszA1tb50yDz+Th
Kdi/ehCbkSthG9alTJp00qZbw0qKLGvrq/cYidoT+VrGxeKPnsulJ6djpJXL9iDg
d+tZCWZ693OPWGsx4XeebOOQA89QbJgtO3FKk08oc2r/x6sEoIJ4IkhMgXGn2+Sm
/2jqBjWPkJqp2m4xsYnXz73wO/wjl9fsE/FkEevO0dRi4M2rdYyXP29qgejoRsBr
zJli0Xox1dPViqAJdU+hfgTmBAUOt2NxjtcYqPGLU3+HFJNXwgAncWPji+YRGCQF
Jv+kByAS5snSOUyUbFm9HNHTnzdcu7OZNh24nzAzTy1dlaeVA6+ziPCpXVAIXfqm
sqvuNJFUT2L+1SW8BHXI+IkqiiGVRAOKKurRsDiWJvGCeUnWxls+8ofACUi6zHek
t73KeyWfiAMujA7JIRhK3Xk3CWHbX0lV9qZ0jLUGqvxW5xA/0RpSj7Z4E27w51u5
roQnPrvr8ZcT5tXuwsUjhBFTYNkr+wiSi9Pe6ce41iyEET5LZ5cH6U6jFOQdv6Lu
PvMHrcwKRuNcikKqZlWIVRdKt575BXI0I80P8e9QSZ1t4kwnHhQHN7lyZUHPe+fn
G75iVjB+FY0oOIWM86/cN/ELrnhe+zrBs1PjERK+LvEqL8hoqWL2mt7tsyO82nYV
cWpeFzzAEkZrUGr25bcYWOfMwhNaG4Tk/3jDC1Rfq8d1ZgIPcJbTU9K/KeJ83CIr
6DIWdDU/sB4Ffl/QiZlNJ+cgH5NKqSq16JGxU8ML5tmnaM1NSRG/MV4w5EGZTNdh
NUbHb9LDJL/uY8rW/oHsiM3IfQyxPw188yKz5zok+ugH4yiIlhBMXesce1xBJdsH
vbRKIW7LmXtZcNPA+dEZIUBfl2u7hnA7VbmjVCoKdzTYQX8pq0hZTTDcXm7d2XxB
mVNys1uROeJcDyK71HmKFJjYESm7D8LkLcUzp+8KkV3oJxeaUop9xsMarQwqpARi
5hID2MxRf09NejpBcxkr5Y3PBvzY8xuvJj+gw3b+4luVksnic75xmVxTETQDBrHX
M+pgR5aP5NxE/1fR9OfJT40YBcTOhjttXD19HG0Czzzz8gP+FWO6ypKhDzrvcLlG
aMD/ZsapewZvBfjX6uVm5qDAaE4N8tuAwhDEuaFciQU4UECmbdUClxYGadRT3Swa
ghMSHfZRo2GDmNZxm69uwCZVvyfM78WGAlJbkAfLjyGdQBO2S1OaRxyIBpORohCZ
JC3vUpgBz828NobEfjg7FwCPDlJqzArk5hTh7PdtF3UhTdwpkwrkr8eM0tnUA+UN
Xavf9qoH6nN/jGfDWvbyvfL0U+4jkaU8pkCobqYrFL/Q4SXKbtU7ZRKL7FDO5LIk
j8brVrJm9qgCBsbpILwf0cIYTVOL7IROAWWDjbvu+TQZT4uTje2oYdWKeCniWISv
fsbd6mYL4E3Zmec5CDkFS54xzP6CP7MJPH0vyCTFhlR5sj1VAbLFlJDIUhNXxeCL
CMVNhHd0k7dsYivIWLWSmJmzIN34Gb1VCvyxeYx2gG01fDfZmy2GJYLHGd2VltnR
NvkTnfNIUKZ+lf6EWF1pRw6nKFl1DAU4nOOukCU+s0V183zg7bfoucGXK/nfjz6F
iMQxfm2Etgx3uuKo8K1buMkEtKZn2ah2FZvfwpy8rw/n76CtEPa9QeWbY/IC9PU1
V1JpgIF7i1nX5G7Ygrlxgq/kHG42ISw5Z6vjyKxOusOStM26bBhHiHlIOyuJkP6b
AkYyoc5pxvZ+d/xTq9AWYQabF8hwe30MpDi8pe/ig//B3tDr95tQMidcaTwlJLOJ
SfZydZ1rcSRp6cCuVMtZU28zkxbNpBQR4rtJXJ57M+noDKy9zwmrF7xA08oBUl4B
mOJAzd/7utFu3asHyR6XlEMn4lIke37vSTFD1xjdlRjgePFH+wNwW4Xd1Su3PgLI
SLsrv+h27OklGfb3uCXI6XIWuHMGk/amRN98RaK+yvl/TXr/Z5JFmadhpJWAdGvH
+W0z+muB8tjbIQlyT3o3X46t5kXT6t/YgCn0jGIL/BTVYRjGmrPfiEamIQysjzs2
Q3VssBH4sa+zOaAAztj14EI0KFlFzushp4ulWQrTToB0ULygqlSpSVIPAxzrN3WC
23HJMXDvW4Z/8/o9r1UzFQD7t8r70arN+ifAuZ+WCkAkMSYhL5GS61xVWgBEgw3I
bMwTdYkimeHMQXZ4GVyWHxvgGbWVmKrtTx10ma/AKyRxU1/41yk0MCqKcYsBnWdd
febcLD9WKAbjXpO9bCBYC3GUALgpmuqs5Xiw2Syec3Ti+A9+JlsN5qkXr2S735bc
OMI/aShO/LntyusynZAVLb8SmPu+Uzkn4Vre3TTAu84G5UeztowQFku7O/u7G0U4
Qys+AgvEOblI6FX0Ny5da1ugdOqCSSmLd3Xlq48zcE77Re7ZpaJZO4DZtu3ks7jI
Q4rC7nPRClhdkE0JAR3HfdRMq5GDahe6kvhM8F7UoYfbviVtY1zx98A4ymSIJvCc
aL9g3MV+nVbCrd/X2Vmjq6b2yOPtDdOoeGxgTtxhLkjZdE5lJ0wsZRfK4fpASNnN
pnXFaXItOAJCMSFMrIk6vnQS2/Gcd87/zq9AHXx7tBNX4XRi+j/2UIEQ97Plka3+
a73n7h28cIO3hMc3GRfCbtrspbNO+38+oiPAEsplKys1CFS1GkoNz60M2VWkAyEn
UbWioK5Jfi0I/xqk5SxNbea/4RhmGl94hQ8MT9bJRlW9xZMrjBmjMmkFAY3Sh077
w2pLzq9bZzBUO44AUGj/ETfABzFGsMfq1n8Ht09YK8Df6a9fqvBjCV2eaY5di6QD
ibwQLx+XRBr4rI/gV8ABl20kC+oHkUMXDdhYeXUs7uEFtkwZQkyPx0h60E/jeJ65
3+KCUf0cKxGADK77jtO/ubSOQC9MiY8vVF7JpxpFFsnqBJSjHcCloYfaTTI+uaR1
Zvrg8OvePQS9yzhHOyl28Fv1KP0zrRYA9yUVIJd42wB+Zlh9U9ijNWe4zxos0Wou
QBLNdVHol/vKPmm3EiHVw6lhldYhyEMbzQ4N01o8XvpyiZ70j4ZziglXGoDOxVOy
iCrwBXEJc268o8uLT07z5AY7wU1R5tXnm8eFiEunF1H07dBm+iRXCiljAMmCAv/g
wD+co1JePFwqSL12mXSegw8zb5RvQZDRX1vWdekkfHthw737qAwcbAS1EVYLJyCq
pVcnkclvwooycN79CGppQB4UExBFgIKu7OmX4Jbl75s2KoJTcvgTs3spImH007/J
OM/eTz5VezjoP5Q3lJwGV5FhZi/oWT51wxm36UpaLQZijQuwzTLo6kT2tXftazKR
9JvskmQLvtXT4HYWfTtpH4ODImRvh4a/LybaNArpkkg0mKk0WEzr/Swv2VqRj3er
G7VjFwnmHauIQ7HkIToiNAoqT+DF8eQDarh0dVBqgFiMf0B4wOK1tr/pxe9Mhleo
3Y8TTY320DDYx/AOtNiztNrklBBEbfkARt8n9FtglsuxRaNoBGPpwmGq6a3ZXg9m
f0zVAnYnPkcuQGcxHrLth87WufJ0QA2CeSasKi35VLD9EVGiasTSR5oIxQbZiYeY
YS+VuCX4Y9XxZxdCNwNkzf4aOPfA6QDflKzvdELW/CJoqlVbUcJlAnpR/C9UqHF1
3dkHPQp5ZIjAqCL9chqo3OIBsLbyw34WtuXNNxI0PRRapXSS3cN9eaF7jZxR08vs
KDaJcPsZq7GKaGycEFNdXCZHydkSx8oAtreaCMSbp9MMRZf+xWxq74wugyI2xBHg
nW2i5hMPFvntoFoFLvKrDJReXzEJlPffh2Yd7rU1wv6av3LGSbliJirEHd+TWZ7y
7G4Qzo4GpuYZhaYU7QN4laaoNryUskPEeKmcngtzl0RFIWp62QHohrmnEXaCj7tR
htFxIrcP57Enrm0mFiKpTPkq8/zz4gvg/AmB20sN48CAqJsLCVg21LpvnFxwHin0
uvRLX9aUlhRFOjPonQi2vZn4DI0HxYG5ylN7vQXvzlMxoqpV7ZNby0jZPX+86oN5
8PLcSVm6AXfbortXJ/J4d135zPHajwj2ELbRDYVc4ePkFErf1ltrEBLiWztD4fXp
ZReQ0TjebUUETgWL1gzWb617ec/B+TfNOZR+pscaN4Nf7th7VYyca+fED0dimraS
lv2G88O/q8QB0NtqL/O/5wopVNUJCw0NrR59RhetGkYblmj7lWYvLO1TNEVPqUB8
hTQHBGmUmQChVPBnS9T0R9sPcZrz10RSYiaIqYFKdKnA4kOmRS5+V5DgLNy1tmu+
2HJa5BuXBKIaBA/fRrrKIsdtY3atxEgShvwBB/jI7OVSoHYd2s1pAed62vpztsVy
/uSfijUPsOhUFnqMqlqF2r8HmTqcDLT0SqclNeaV+Qvcdkgz9QQuhpJbBgheV4wH
IfhMsfKUgyuxyrNYoc1GoPxw/EmqvjVQfxviqDWFYuHHfendni2u/BrPgpGqErU3
qXulBxMULTcqpkkYlxIZXHCQZTvwMlsfsbC1Ef6OHNonfbTsp4ClgliDf7F6MpCH
AZ1soVnnu1kEVD2bCT5SdkmFv9GWNWGbzo80hM2dETFxIq7+8oQ6H0xIjYSXMvfa
yztD4AZDlE6bOl0h8+6+vmInyWnMxjwBF0gKElJtQ561Oxe09n3sUqdvhxSHhGTj
2d/kbRvCAsy4dwtSSZ7JWTL/V/TY+f0VPcFQqunezSTvs/SB3hnnlf0HiaMIlL1A
YTm+OSJZp17qUsUvzbr/Uq6XuyiGhxN54iPlyE6qVtyDrYjV6H7xX6vTozc2Im+u
TgxLWchOGqrPIUcgyodXATRZnnhV9nE/xsPNIw9Kr17hHDBt7PK9+SmKnyzAesVe
KzL8BtifiZeIl72yA9qd1QWleizU4ZSCvxlJBG7LgHJ8u/V+MnzEK2SU6sSFtb2J
j7GBRK3XkiPcfsr/noN5QBHnOr9qq+DH9H2cptor642hXMW42sI9LKZVE+I8LN/9
E5wrZacM4XUxXXs1H0FecFsx88M6fvZmeBUvfsNai1cmUXAY3tssY7yKNuNz8vTF
XotsK4w9Iilb9DB9ha+NzSQvbnyk0pRNNRDj0KhqAIik69xXCmzLdmCP9XarPnWu
yMkP4Nf/KTdoQzNVkKXxJqsG/Afn9lDPSbdktjAT/cfXG8kZvpDCL19aqWeb+Ce3
CeRqFVCN8aCtMU9BAf5AhmCz45n1ZuFnPbnCjgiAM5zuOuZLNadYFFyen/OZaQZ1
cw0zB6pE45dO5Iw/jqiVxZfbNiVFT12M3cv5+qs9n2vmIyEnz8XjgMN2GGdvCirl
0vJrnkbdOTybVv/PZRfHO97Zoghu0wP2C/ZkAs/efUcRABZrSpzFmP8UgX1EY5o/
V/pF/3RhUfZP288O+RWHrSKMtqit9vrWJH0XPFD6MFYI5sDE7+Ygs1Bt7DvEo+FD
ey/kXXm7BE8+5hviaSaEzHdq5fFnktwTQ6CIh47YijLHxFvRhLXdygKzdRdAvOy9
vAbX7s/C52llJvMu50FD3pkQTg/b7bX0DoA1GMZfm8MNsUf8emrVvAr+VytXPVN8
33jvm2Zxz0Z3Ba7k8Iwi4fbfRuBw95eMBClMyhKqThYi60xzPYGDXNC+Hxn2EZl1
2LIBx21t4+nfxbTRFqTI+ezE+dLnOW4SrJU3jNMaDKEPXXYV/1KBxgfWDSi9Mx/p
TktBCOCzMYnaFFQNWOt77MAEWQr3QnUpE+maDjiIrkGlky2PeB0UyBuIBiAC21ev
Z644X4L91Baoq4t58RXh+abJkysHjDQxzTSpB/q8JHawSc3K0waMvYMr7w6vpL0+
LVZexmM1BGXd4coqeAKF8vvMqBes0c5Q4mLbOmdeeRsUS95fOpbDY90aal6M79Va
t3j9f8f1zkIent03TMoHg5e9W8QHPh2xDee/pLaVzJgPZBfQbH4WDoopCTcNNm6d
2z0xjyDvCRn3BGfYT7VIGKibz3x5kM+svnVfbxhFEdVzjwlKaE1OaDRYk1c7XDxL
v8SOFyGpcIk1MWbx8CXJc0RDasXJDYJeUCyWwf9zamLB+Vc5GqnfyIY7zN6N4Xsa
RpbfNogF0JE9uD1LiNr7FtafHeUlskUKq/9sWBhyAAPGnRuB/8CB1d8STUWqGPjc
MT38Sas23ETuPBI85EPNfFSLOA59yZENwQuqhmEBO9M5d1D2Q29kcuX8nwcnX78o
sZGxRG2yTfoq7KZVsMP8DQ4x/zV/c9LBSntNYP4127nVabmKYQH+pwJ6/WrWFhPu
lucz/KLkIQxEYnLG9s2EUOttSFRr/nFxym5nzQsCjDZk4KGkgkKaZkNf5EdSgv7O
GtpBzZqcH4NFfizHKyyq/somM0SC96mXgEaxkujtV/n3uEGSKgASeBGFLrQUzFrI
D9O5FQsE77r9PNm0icWrTXfXjyL+49c5z0DGTE1SifnaeStCGm01lqh9YhIOcmjb
78lNIVno2JL1EuesvQt2xjKrxJbrGaRJP9Xvz85xkUpove7RABasJwXnjCCe00Hi
BesdjUVsUSbwDTKHQIDqq1xCCfetnvx0/SjVGG7swshHwt1LRyymARbHClAgwGzN
iPbD8NNdX65H61k17/befTfHTuwk/Xw3PIABVTQxQ1m0VmmMVYomBtewqXckIPpS
2Pl9/6itRbnRoIyaQM0D4ets7MkO2doFCHkzkALiPi/f2ipQUfgYynlyho1U03I4
1CtV/tGYdkKl4myZ71/nTzxEcSAbIPWeZpE9G8ZiNNa61HHpXV2XiE6ZxT5qFphe
3krzMKGMjOIhduGdov0IQF7xMFfuvDMfnZv2QRnHL6wOj/4G/ah6kk/cYL+E2Nce
Pe+A+/DPi3pIrUVPifkIRBbwPc90COwZjSuRf6SBk1nrrrhcBNbgry0wd0L6odXW
Zb/ItzKQMTwadS0WKIX2+dFUMPXMGqs0ecuP+n12/Lh2Sqlmh3k/s+PG45IIgOL7
Av5U4vhRXANiqC2RDUTJ0xWIBoNR3sxoiK8wmtVHPEWNjV42CHb0d6AAo/Jf0H6Y
O7adOmSEWBPv064GtX0ULF/D+8/XNQUpBZrnmV1n1Myo5fRL96YdMybBUEBCq6di
LIAN9eqT8+VnOA5x+TbextZtNAenAthBjmmVL9O+Q+9HszmF7gQMfEW1F/ZVYF3W
EmOQfv9TbaO6+AvFaAcWtsCXJ6tjZuBesW7gTFt21rrdEHeQb3uNiqFjcq7bjfaR
Oi2b/n4iJ7EmzUmmQolJ7ZbU3r9qNcR8sR2nZrjLZCNEGMNtBKYrSbASl5wzuq3F
VMl5oA8X3jhYjOPyMlu2rN78sPGFZ4rLVOz5MequsV2VpSwCH8iG9ne0SzONrRkb
Bixmk4gRJ6NLCgyhBnVAKpb/TiK8Q6es6cL3sxD+y9MBGP4k4Dcw7ox58XJXGO6A
g+pq9CxUB7AKwpJz59umjfLVA3WNoW3U7D90M/T5t/iYHuQjauPHM/wXVVZMBI0R
hSu43JHaSTXLsMtey+qmzMXnY3ZZAPD4TcCeZgBM2xSAu51rkSWlhR3nbrQYK1+k
fmu+s43KEKRuvWY4gMnLKy3YY9SVR6TJRw/Tr04qsP+rm86UFbBHCxAHPUUq4SgQ
QAufRYs5fY3PsyHhq47r/sWAulXloTaJ+OhNYoHD/6JK588IhMgyPoAYEwcIwGVo
Q25qw+10hD2E4PHoHys40J12E9Hn7qrKk0lQZp+0BYNcepyY8DObIlnjNxH3AS0V
00ejaMVRza7Wu/c5eiaQ2hgZxSCWuM++SuWicyouOWSDIRVI4olkYkFrOpjxXOuM
f8qkJi0ZpXG2e+sarv8yd4QJc5j5Qp9oPXjLpOuxQjHRSwPq9ZcGYeZwXoDdk4it
OTtqyKRZiN9RW/fQYsm8rmJyTeu3dRS2gYbC6p9J20jXjwbL8hMU8ADfKky2F9Pg
DCPEbk7PVAW90nkyZYd3SOTyFrTe47GU7NfWvji0LWsQBOP6jT31+FuQBgIqEk1d
dcxquxGHUuUtIuotm8Byxe2VfTJyxv8TO8AuHk8F06xPy14rk/7NaYQm/ihAezpy
B23iANdordu+EvTHrzf4i699Vji0tQA512AgQhzslwln9ZV9Uxqltph+EpETLG0g
C6FGf7GF96eoiW4+z7otAyGjdyD+fQLcSZDdLwLs12fOxQoGQMoksEQd558aCr6J
wLwmacx1UEsRfQF+vnA/rSh+Jn/i7onmaq+sshpeCJ1ZiALFeuMEbYabL3I2CkMy
N/eTfQ8GOJKnh3/OUJM+LYplJRImL6Y8D71+/8aWCe3lmgR7Nywk2BRiiEYDyiS/
SB0kg/KZgd6mzUoMqp6nn6AUkba6t6aS3e8JQeKm/QPk+5SfJHkYlkMPWfp5GxTi
44AaWaXtEGB54py2pJr58hZ6A05209IHOrugR2ag/+9H2SVdn7phrTRz3gKL/sYz
JoH/mhv9Zbz2M1wjdAeJtFSfwyzgLBjnwjgxYKkz03/OqwGu1tomMhS1VhCddOpJ
alnnFsGOHMdvV+1nYPJJ+BZ18z+BJ9tscPH7qCjgyhH1QcENVn2PwAKMASQPc3oY
s2dqpPRuUl+d6B0d387QCGy9YhPn/wVKs6/tSSgEMwkyev8jqLe/RDMz3D2vKbyT
gBUGupCakRvhzvpHDUaIJzaeVG27Ci4hVMkb8Y0ZUqUgG/RULhOn4gn+CWyZLxim
K+gJjK2Qq4PMFOdmDPQAn9ArfyvS5z8MRs0SFLBu8NsULIFsAO/GZXRlw7n7l73G
6BSHd2yzGfDHZdyKgkZWRVQ+xIC7FrA7EDYS9ief26L0MKM93kychtVZfit0QbQ9
/cEK6XdVdRA6Cx9dakTBpjXSTA1cEsDJVhYVUhp+NCKyNla8vrUHvHnnNxFUeS7x
ddMoWmFPx1eY8mIdoHKdxvpgyvNfm4RUZpfu6Avtc8iwhCb9D8WkrOP57L2UQ5Dx
FNqJon9IR9MJIOTRXCKD2ajt9MeDqbjHe4tp5rLPN+weNd6aQOD1ciC8uBv8c+rW
0DAkAaKXGwT1eXjT8sRUfgpf/+1bqG6jq6awS7Rn1TZSCJhB7Qpf8BO22nuBHW+O
+J4Qq47w44bC3c0EPD2zajeSzBM+gXKa/KD2rU8qtom9oq6INmex1/tFd8tqnz2X
Jc65xhfvjmzcPBiX2WcDYS/3Q0R741Lip+PzHsvc+3jPBlGKaX2Eo3kJiwHkpAMv
C42ejiQx/uCSkGmVvZl9e9Zu+Kl550iZvFSG4vWiGPci3HZxcuEpiQbr/kuWCLIR
RH/dY1sXhE5wbqqX44g1wo3dzZUgYaKboznuXHrrh7dkH6jfloZwD0Z4pV4QOqDQ
gu2T9oz0uXqOQpLJuVZzt2vICbvZ8yNTtKH7ufdQSjDNR7fRiVnCLiLmmWfWbnsD
qCha2YFJczLJl1skXzWQ7sjQXI5TwK4FtHZWfUKqQeg+P+z4LB94jiD6GNbB5WiD
S1HgejXxoTXFwRkFV6TGZc9Ntq5/7mRogCaCoceFwIAatZaHeFSEJ6Qo0LyR7Cy/
Y4iDA5NUI0Vqfj8AHtlZQkbA09DRuUY+RmWgRPx+uST8aloOYOc5GZ4bEpyz0NhK
5IW2wvlC4LQnOI6CjZnDdusemOF9TMG2hHTuHASIM2z36AiYq5x0OwgRMkVz14Ke
VM36DJtiT3+n7Z2PDnRNSshKahkEHV41BHAIO5OjDey0iuqMtiTAdrL4Rca88+eb
DUX11C1+TOtsw3yTqSsbhLNYEtIRXBwXQwAjEKTLJlo0Q48e7caWUIUNOgO47AWj
FgIoT5WyeM/DeWnws8exqEYrqwcJoTlM5rDuuDMfRxq18U7s8vJsqI2ujIlm2XyH
7FsH9VpRmfqKa/T+mp9bjHFg/Sj3rqVE/+JtC2nqNwmG7exx8AUSC14mCRN442dY
ylL+/UjTuEY32oggYhNCytUOQSDKjj+muDq4Gt7Q0VdRNHxdoSa/AkDLMyhA/wrn
tit6eRjz3crAPWG8TD4NCcv2UfUh3/zI7OaayHSj+4IPFxcMm0dHs7wLWTZ4nTUj
dPLPaXVHpD8LgLqRtnLsMy3wbXQZFUrLfj8Bmkm+ZTZaYQvlV7p/YzjcpU5Snk7b
5zDurRsCT5lHMdyw+ZZriMfkDm0R/72vholHnfmRGem9cUxD+O96w8Ofmh93MCm5
08QWegkSLKtRanjBiwM4Uhsqh8wKLIKS1HazV/JxOHPZrkTOUYcLvAccFzylmQlD
M2HM0YvUrZPk/1Im3Ug3jVIDHK6JpwZYycdPhR4J20UWvb0KDbeH25l8v4MLROT9
vwu+8wLftJqRa2JjC+RIG95fEhShB+AYZKE+Ug1OjZMf+d7hon8D0Hmn+sJiZJ+e
s0T9haCJeamD14HCiKcdAVIB85luVt/XATawLQLaIDQ=
`pragma protect end_protected
