`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tpNzg8wlqoPbIcBx9bKogS5cnd2wfzt4FIc+RLeET06wi4XKl4DVUO6MlbugxY/N
nxHpWtr8iOmgVzCE28X/ZdHaphIBtTkX1ZHIWz4dVSKDxLi+FWywcrVR7q/U+RBU
lwMOBumfY5w6nVmkJfJaH4bzOxbnFk8Hs41p6X51i4k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21904)
NpC+ffj9z9rwbAh4qetBVzMr5Or/Nq/i1eF/ABkcx4QpVMrFE23TKAbM0LniQf6f
naPVQP11Rb+UtvrX5WD5WxcGZ6XUxYgWzSlJ6rYU77hZQUbUmDf1H121acHWb4Iv
zqLxBk+SEqOMCC1KOYD/b/wPdSFowvOIEnWD4opA9qQp+T6SfKfVPKsmpCTp/vn2
bEt4yeJs0Y43bZOFyFHQVJKnkwgRnOTaq4vp3IrQNCbepvRIF2w1LdjJ5xyMcrdv
X4GPSmmFtp47oXXx7qsIUxvJSFegCgpNJ6gUScQy0tRvEIFIehWW7IqwP3+fv/zp
AWSt5fLudRnYd5sX1ljy8k5XHjTCTBVRZTF5PQL9YajSa0JS/y4X4mHQ6QHoAzZG
j7O5cC1fF1/ONTTyhHAlqoEEY0GQ3VaKcdWg+nFJrAJPOyPwdAJcrwWFvEUHz0Kx
i7gd3YRtuAjZ4o/iHwcH7p95eqmBVCKuGVe+dwW/OkY5f6T5hftZT2ihl72snME1
gAd7Oo/LTUAEsyx0OlgO7KjF3LgsjweqMQ7yDVObplLaxDfi76GmXSev1n7KJ37t
O4EGEK6per54HV4uz1An+NbfN6vkMswGZCZuIsuspYAJTVSpIBbCv/stMnMUPNJe
6clGqMbR/HNYRIYw71d1wgW2krBB7jXigqDed7wBkzbKHHSQHu8TynJ0jNQse0/W
yoGbFt9PgBeydLfBa7MVZbkjAV3Qnh27KZdlTkG4AMGNYkgrpyoMqnLqm5+vKH5E
YiNGoHjz5RJQaU3GWU1drPWU0IQxew3oqhRZ7+4yBOq30Ok3L2h9cA7YNHLapKeo
e5CG4AuBRHEX0Y1g1EBZ8LJiEkyyaKGjFpkzJDjOzcFqybpPreuV+vAlPGCsjfd6
OY2S+GblJ95bB8dLMTAfMuwEIuZVTJd0HSrKj3Hm8xVsxCpEaTAlSHCWv9gnWaIj
eR+p6wdw2lwvEwR47xKpEjKPAFsbpJkdJEQPCh4Lp2W7t38YdxFs2Ho8wUmhAqUh
fHpPm1JZIGdK0oujpUxlLIdal2+ratSGzRGi5PmLh4MyFZuvJuODzQcHwwxZpZ/w
NKxxSgw/G+o4+HPXyrRQcFMwynk1OTNvlq0hMWq7NLNCQ7XNPDRwelm6wtAHUOTQ
5C/RpO19IeQTBCFLp4933Fm3Dg6fndQ1/ka4SLP7yG92RTiXQmboxA1T3BRQjray
LwR0UXOxd/BY1Pf0sjGu/Ft3JDmCr3XQMEFDyrlxg79Rt/BGSW0wPcv2uJkyrrdL
rmwwEMiQ6zBCZzNzoeIWw7rFsBtq5PwVRAQCFAtpfRH+LsS7KP2EkLWNtD1FSS3B
kyiIRSOhGxru0d6A3gNt9i3XZtPAABuffZD47x1335wswZrzZgemkRZRZykEFhy2
2SwFyA0xgE2YOLtD76e4gpWvsGBFtZPfizO/I1qTC0XHeVNoSnAuGx56kUZ+qlGv
SJUhhDfWakDj3ICF9A0ODRUCz4TIaAa8jSo4jVLszpkvFpoWT1uJ2ZSMU+mjupau
f/Db+xuDqpMvSgiPSbEo74MLWAChxlDAmL9yhqAgFNZAArcSISKc1wdlC2m7U3ZB
bnAUmDd1Hg/uC4yQVXt8N83sC+GZqLxa8Y3liYpezBug9u6+rVzPofTniwPstYgr
GqSl3WZMGmwQvd9Q4wJpJvbVLUfF8iHJoiabRhaGJ+kVx4utX0I1hlAedPW5Fpnt
WdoZS1+oaylAimEBxY2G3D0grKuVyA1NfrCXaLTMdVwAM+9LnUH1cY7tYRuGd0WP
/z9WNy55tEe1a6JdPgstG7aX9r/zLmCJSjWQ9iv581MjemmFIcXnfPSczUOWCoXs
9X5FIJa0USt3NSv6CM8B6vbedrT9mpqLgkDxJepuTIxYLCu57ZWfC77BMkUiGi6o
dAGOEg1kdU/mNzImIeauRcb57kNKjNFAqKl+VEJsenRZbCAehX8a0qXi8JCKjsTt
OI4iIxp4g9bobwO5xXN1XXUrfcy2SqNnbOxGBfe0Ca8W+QE1Sl+JQrUsCDlxwxYh
P/HZYo+vztNQc1r+XFnKF7YBK6UTVgpBxp5fvtLvYdZlY9MI5xemwL/KvzcgVtFo
S3GhyAn759XvThPImP25BXEUZmTbZE38MD5GVgnZF7VXvt7CsgKMELdsqIUWehKA
OPoEXnmhGICkMWfvbKaKhHrE7b6p4htwi91IUHYHp97kpdSywQn/1BOSYeOYMcYg
qxd6c79KaIu7PjaQq144fqUJe9pJ7ckCxs+sggT6TK6OHnfXvX+h6GUfV9elchYj
sXidjuaD8GmtNmkYXPAiVkqzpR0SNg/tfZXrpRmQf1xaL/rKJprlIyCm7+XWb07B
szWPglpRBfMdL1nWIrsb6e4lBHa6XaiAtzXGUbEYDFrcLTcAZMsExgxywEBK6E1r
g9kjWGaWgzGu4aCroVs3fjLzNNyY6x6b1E4ty0ors+ScOT8HDgx5GDlSUOfseZyI
sQu5wLxVR1/A4WXTx3a5SGP0ZPKcIpRex04CkwWEpfdLsZkNkjk8vnbHlWDOb845
2mGh/MbeskZ1wgkpzs3aLdaKdceDE6r2+vo/38eE05NX9EdBmx2zlfUBB/BTX5O/
0Gg4a97AqWVCh0zx2HPYEYa62pL+bFtrTjzBWK0MrizPPPeomu6B0lylDm3W2OSS
HJ/yWseVv/HD8tgwe4GeTrzPeHBk4aL5+OI1QsrRey6TQJMBf+4oovCtKotvnc9r
HRPtY5N+Qkh+iRQSCwhcW5MpB8aIdG/MLSg97wZUb+6g0IyKafgLRdTVfWRC1jFg
CuC4sqkroEJkdYYJWxFf/PeRn8qpl/q+4DMQYCvBiVjuE919tJXpCh/cEOQ5hFzz
h7V9kdcRebZwQBCiFWY9ys3PFyQFT5C574kIH1w1l47+7U7uRl8ZGGi/Y5li5fdh
CMN83prwfm3ObWrNW4Lp4Rvis1LSaWzhrb8GkLx7WLLVqJK6dhpYc24QLU0UwDcb
ViDT3r9xciEs58uDckET7biRPRpHF6mvEwEyPaku1uCsi+wGbvAijIjIt9k1zD3f
e9R8r/Q/rVp3oPZTpBtoZ49+EuBWXmMhNthHEUdTrGuHFLo6uOn0viHK3HdKlYD0
8866hG62fZTA4im1jkIrWta7YTyLQ6pH6fnQJ585QauY99/L9YpsqVKhzohGoFdH
7/4hJKZAHFTEMkfaPCR9QRE1/0JbP7AL6J4J+bOf6028r1lm5D+Ji824gt2WWjIg
xBYMX3QSY2Z/GmuCyd2jS3H5pded8Hcikc8GyL9YbPB0uXs7MczrRQfxCvM09t7O
4Nd95dJdPTQgDdg5zkgdciFU7oKBz2G6Caj5dJpISRTCpmtIobqQ/6hcv0IumioP
1Q1/lCSk+6fz54CdcOn+RkdNWJJ2MyGC2gvPskK+sbqu7OsOo9evr3uSr356yvvc
C8WYIpgRNMIIW7Oo/2EXKl9x3RChfDCq5kLxfGY2ojsWCYn/fO72nkOFsarW28m6
YZzl+RhtPxuexLTrWVyIgVetQv1LQrZgfs3eFJgUfZlXC/ovkWBuFSc8BvoRCd7e
zAuldrw75WrbkzinHclik0oxDlB9j5UqYWkBiDACtp1NutFF3IZRDN+pD461nsaj
stVFdJtsM7pAoZltfyk9/251LVbA9B8dzL8Gci7YY6uWcLZTEbtDhu8T0JHIHt7s
KqyFVq05eDv3dkOMMPzW1PqPhmvPzblYrSahi2Va3xaFntnpuc1X6RvtcF7yYI3d
g2lZJsRwiQYXcbhV0dtVCrVZiOOHriPbz+ji6YoiDPGjX8im5PQ8bu/aYfKv1xQK
6bJ3e3jAupL/dgp1JSLcGqBTN39uZR7dvq0VzOCDYLuVtPUDvZ4Jh25g+b235DCy
HjlCafHtSPcDaHU6BCB4FOE8SZaBLYDbbMztQuOu3qPr6R0ogO0TxC9Do+Bx1zzx
eSyjHYA0LDLgyGyDNQ2+pIOfzUlUhDRj0/mmuxZycdCJ9Z5PUl3ZSlIYQhM0Y7TL
k9SBXrMHe1Sk5tyRUogr5vKqL98BmUz9TDZzu+17wxj/RsFsk5yd2zQMcBiBKZxg
JAUYsPigD9C1QZZoWWR/E/IAAk5sK+Xns/yClrb1T9LqQqvUdL49a1sPXbvt9UsF
GZ1elbN7cllEdhqrqwLqeagR9bHL/vGL/WfkZUCLp7oRW+vKYBjD0wr5ovaZ1pPA
C9Acm6HiHHfqH+2NDYPyydX0u4wDL9KDqcuiHx0nm6INTEYss8MgbKpft+nnGb7j
i9wFmyXvYP0Nhi5QLXQk2FSTlUrTxQuJ0xVbeF1mEXxu4QFUt/1s8vp53rtL9IYf
KPygrKBqtwOZacyzfNvU41mfmkMC6N1g/YDhgTLDjpqgDnJzLpYGh98WUO6YWkRL
0l5N8b0zl0UT4NzqIOJP/piUAao9KAGnpM9iZ5KaGHhIt/e+eDDfOBc6bw4z0pfc
ji3VGIy6hz2bkX2mEGhMt0e20iKSW7/E7OXq8l4+v0CW2zTwjq12PyAJu5EDwm25
JkTwM/56Jnvxl6XKX/lHkP9ISFIPy9zpK8OYa0YWSeDC7feDdnhmss9wBOTSR0t8
C+0vbtqRbZ78SrUaVhIUUA/etQFC99l47wdHWYT0RkCAlDzV8HxNmHc8+DC/7pgQ
ZjtTQLjJLXZLiAIJ5Z6Nn9MwDpF5YIDnhqOSwPC4doiO95XOkuYbv9SKOtIlAC7w
7YEZFTJ4veqA1phJsgPnzsP6EkAdPY3p+RmTj0uWhGQXWNYwQGcLiH15HknIuoa8
aqxj2aS1wPHDfPlwqH0Sp2+sn5kUsXMCi4k6etQHGd1iGc0Lv9cEpNj7jsD8lMd6
b9PJG9aAT5ZxyMXZWkbWcCgM3xWiy388MCP9fAowTdGaiiqwBm8qTyrkkh4t1pCt
tyyXe2OaYa2SKUQCmOvLLXvoL2q13GYO5UHR2W0J+0Jgu4QZglF2cIP6ZWlw92Qb
GTKuPw4L6ubzHem4q2poghkq+JMP4SkwNQ+s0klRD4r/1XukbsaM5PV6286FcxoB
0AGPTGIRpZ/1zefjQ3OJAUqJ8w0xWl9yI5Fkq4ZM0DwS6bs2WRAdvYINUYW1HKf/
nT/dhqaqMLOs1zuRIP+PENl8niGKs8PkOuCjKSlLs2jbFQHxZwt0vfeU/I62VXx4
FnQEuI0RXYD19LeQ+v0DnRRARbVkLrG9D5SMWJanFODVWCtTQY6GhOOHvIceViBv
STITzHAaAPYxDgYGEBXmn6gWxftJtOd6BUQbzyAmyYUvmH9i1bYRxHH5u/PBXcI0
pldx6VNKzMHJSjJ2gmGnTtiW69fUBDriv2swKkI+DHu0AsEe35wg7Rj9PUY6q17I
HW8Q6tQjrtazgAaU2PRapNTCPZmFUCRJK9dV7keNDAkUrGifqER0TaIYbTeM+ol/
2wLmvP7ie9r6UDY72x8YDoeBPLiZ3NFKhcEsMF4A7il3MnrKRcISndw9odBq0oAH
hW8ep5LVkqvjyqQFS239oad3zS5Jh4BOIMTZxjXel6prv3LLSBASRM2J5QJ54UNl
arDbnYuB1nMJjeCMGmuk61rIuHnmOtmcIe+z4Uk7MdZR5mPM9EEaPNW5aKJLT6fI
+LCjSZxIKz0LcydBDUSsPyotAJ7Oq0sJSIyVHmJGcJNsLfLQZmnGadX4mWdywLad
rOF9F4S3katoy49RaTqGh4H+XfZQP2SqC4AmCyxMnRSrOm12uo7YWoYr0/SLxqRb
i/mhjiui58W9cGJA0zrckYLFCTOFAcQD/ljTiOlGjcZKJu9elYV2hMAqEjBMIBTK
G/5B7p+bUcJPUbQTHMzYQSLGVA7aCCJvbwnsd8jf9aqNGkMXY8AGKeVkYVBlvnBE
c02HVQATRiQbrDhfLv1foamOEy4DXT26mqqHV2IHgHAV0M9elm0wo8pIbszvHG1+
Q1cK5usalXN8jlWM/1YpRuGWF+hhFfI16CyR5uCDDgby7LbOGYkFtTQpBsJJ3wmq
9uJ2Xe/o7jxtPebc8LO30o/Nu93ZCQ4bbXCrBH82laT8QRGu6DkQoBQDwbb8Iwfv
epu9LU9IIscHVf/+notjFFzbJ5XXyHqqoIVid13nbnSYJQdlOlbapUuZvxj4NAh7
878WB3KgZE1I47sg6a409c44ASkQ+MUJ48A4p/dnGPyllrnIjPa/NyGtQSQnaqBE
4uZpjZWNtvEoJygWpiQx1K66jebvjvKpLLgt4tlpSnjLeBPKBIA3GhV1MqsIX3b1
rlciXN9dFbrhlLUwE1mZCkXedQ0QUEx6G5FtoHZaBxYl9ylUuZQovOiR7Od+h6zA
KlT3zkDK7PLimkcrUHgbWP8qLq13bLUFb+4VMfD0LrxbMcv5kfGFHrHIb6YvbpUy
QbvzWNtBWkvfBNhXzCnfK/7LYs7hpSIbgn4Q08vSZOp/YyWFFub6GUb8d6D4xlD8
hfDJQXoZuoJjQsd0FuYbmglias+iXQnTrMQHF4ZRHg3iUAXTYanQb95+2civ4M0M
ujvTmTsyjMPLAg+3msijnaoHJ8G5/XttT0DYqfmlAwbCBw5R+iN5ox/nDohmHUKD
o4fUdjvpIhUJCe6PQGCzE9VQvbsAHPZIWxcQwRZOS+rqMSG5zqnBwn8KyrIPSq7E
KcD72PauwSpG/qRCwifhhYP59cZW0RqyeBdESM6MQHVUqABTKCWqX3L54d4QT9Ck
DMdiIQFTJ75Y/mCpdXuOE0Ukoy9SMarPTV1YTobIPy/yNBxSNc4KJ0xo3oLt7bHk
oJ8uH/oTDN4oZrBAMosOlAroFzEcS4Dd/xiwxch7Ln+MszP5j97G6lijcskBpB33
GOpTzH7YnkArPDn3Kykycz82DaCtuGtg94RNDBpZ+klMGTFQtcbYDUYjd+oj/C1B
rUCUB/QR3It2vMhzmdZJB065nZmSKYRNqlVox8gq8cpA2QSFciJHUmpLfNvPZeaJ
4d4BtGhBS2tNU/0BMCiqlXSzg3VWcG01+LCQxtFIvw7Ynojf38oK9LMBFQk0euf4
VHRH9ZdNTEdNGXNdCpV/+A8PW0Qrbp/CSgHS6SG7Y8dFNYPRCfL8WC7sFZwx9G6G
lD4IWHTWWBcfwGaenUsqUgrC+zN5Zz+PzzfRV+2qkcsbrZGdTvWHYaBaEJwep9rl
OaV4+8/FCumL0P/Wt1BoDP90UQCFTtsMOZO0kqGCPQDlH1ASRRcB5En5/fUxiwjZ
cE3/lP3gJ0/HT2jY35muL6IcdSyYEMpgVk53LS1+bdc9PDGN7g/15wWwVN3cIUaV
e7jf10pTnSQ/ww+J2LbRtddAOgVeiG/WYMcfe8TkDKrjU/hmjTpXvzVz0HoSUCe7
1fw6UEFUhi3R28A5M20PuKWD4vq1og97XUeGoLXrehyX4hG6zS7fI5Vq5mHLWqT3
yrRJovAg1fe1koxV68xt0XLcyxkSyXk9n4OL3UZ0nBPXKDzcoH9qgllMzkP6JIbk
QM4hWnztMoc16kJLUnqRNetjibsqfJZiyKEOmMEPTJAnaxn+kFHsnCv6Plv+5eB5
pf9sfgTdFhM0BooQatvpdg7GOarjvcvzvVtrN998RlmOWBIS4nUYYIvJQ9nbJPDb
2l/8BwK0fnCrA7DzRTdA8ZNIGRrxFIv5NuJ+kgUp9dNXwtVn2dillivrSapKmfUo
IHYRXa7SfxWRQJaOlhMAHxfMO0K4pbDfs7Az90bdXfp286f8+r/k0cM5iq3UBDj8
uEiz5HA4d1DHK96CjD7W3RxklwVSF/jrkFAklx6gtfeXXCw8UJlqmGiRz4uOM1jK
1XxqkmzANwjVqJRP5VX4yoGXCqblBcaWKgpGNvlNFl0MbfvkLh07b6MeVJqlYUmr
pEm8oEGw6NmxYEkmKYXXNN2WgaNskKoALbOfAUfU+KFh4HSrEJi3toHyJhR8mKNV
rVgV3q7qVy6KWFW6Wju/D1nTabFb7Eww0N+vsGsDjddZAkMFwkaEQe73EvONqSq+
cInykcEzxgPteirjISU8xGnj4kQGvpRetIOsJLu6tXABgwrBVDNrD8yQVFi4KFrb
45UUA95jB63Fo5Ka4p1zhGPWlgYlsXuIjE5araMXKBvU6iTD1w/tdmRkWKFp9IJ4
THSmxPkuRvRz+6uwvvM3nmGzGMtuO3VIO0waUr6+R8ssf+k2EecTmWKUDVVKyfHq
IrQdofBMYvBQq3nUhLXRBdnyOmMKH3qoC98No7+aQxiRBERmJ/5nQ4kQB4rmGOW7
QuhwNPtmfyU2rBCrp63htXBlPVTTEsEnaT/c3ib8o8g0CrvnR09s9LtAa1TyWSSG
qh7LCgANIg8YurNHoMrFZ/eHjRKC8nxtdk3N7+HV4JvBd0ewzQgBwg5ctxbqYu6Q
RFpvjHzWv+4jH4CQulpokEXO3g/T3fXhoArg5i5cxGVktzgFKZAxlarAQJnLS+Ba
BFgTlv14W4WSKN6KNs1g/EeEmH9rtdx/puAAQCfWxgvQfekhhFmHKg9k4bmwH0va
k3Sl5pZjzA4Wm0mz3V+rfg1gweIziGMOfEnTrYqrFcWSIHrHYmIGYtWXowI0IM6X
KbiS5OA03lMLZ8dveiWEIIclf54cUrhu2qk9PJ/54NNsL1f4ml9d4hUNpc/y/jOk
l4pfYctdAT7Oy2OKk1i8QGtDyimXTzUOtyxOMl/Iu8UtVGVXH5z0V4GWBTIiEPy0
qAkp5NsPgiw1EBd9KU3E9jz9e1xSeIFpaoikVwl+VWHn4iJDhrK2qYtwwiYUFvUv
fJ6A1CqaeGBPqgnkcxqrJFtdgAHGcZJin0WBOztS/ZEqIZBOiK+wTLwIIG+AaHUY
/B7k+PmVyn7Q7V6HWOQW+hl4RNKo1fA2w/GLzQsogQa9Ax3iP4ITIsa7pq47OYBo
HIuPnZn7JYpNCdtLm6oDxzCpG01wnZX1N9N9aMmRmCNGoykRWfk4s3sa/zwdIgc8
Fabmr1DQYmoIiJErIDfK998GVyd7uClWh8SVTZptMTPI1vl6RJtLWMFXUpS5Zh50
PxB4Uja7Ju/k4L0ovXJPg0brgSXXxwQC4I9H6lSVNDI2MUJrHuHdA73VdLa0c9mo
apGwfmPafHjM9XvWsCB4QxGobKe/sSI49r//hGKu04BMbmy4Xb9oBwoCRaOVkxiN
UL4qUwaOux40cPJAdwgZ1MRKFgowYbK3ELUK5Rokj59K6/vXlK0UpWWTU/1KsAOF
jzlQLF3+jkLvNqOLwThxMb0SWLwl2xka00pTgmcGEkNR8Ux3GqDZxYd+/kmFhY1D
bAXwDVLlBh6bPHz2VkpPzrpIzjrNTMlgKZKaANL2Pk5vQvuJjX1tf7MPT/thOGtu
Zz57Wfxnd6E+kotLec7wGYyXNHTf6LdlhUIxtzXidVXI7s21eNDfBr5rA39GNU4a
6WZJALLSLhDpLPYSkDPbqXs+4kUnY14ABYHDvWmW7GIhzDB+XUSosjjqglR0gjTZ
myd4p8V158VDvgG7uOFbb20DCPUIoOrSU94i5e8Rxs0g4kYayEpuCvOeMmQ2l9PO
F5iOx+1jh3OI0W6gfnBNfJ7Fidu6MPuo1VvUyJky+Lf+geLwBaZct970naVVtwtv
E68eIk+zzqDDeKZb0E31yTv6B9DY6hLHHW59BMBJ76kV7vpS55sYThpQxm3jXsIj
V214xt3gyFdwwuQyiybpug0LSWHJ/wCg3guIkHnlOvdxkWm/a982taNoYvqCFkhC
pno8jt5uhYu+7SpIpMlH9lk0yALZ5bont+pruqYfa99x5UN40db67l/moqkSN+/P
N7KLbKCedLvKImRmZbKylPScc+a2mumeGERsbBAd7Rex5derf74rVcKpnPg1LFc4
FXotILdHpWjPvusw1XIpWRH8CNuYEYwibSoIldUpFZoWwMHSFOpWiry5Hw+kDKeD
+wq5jaoTbbk1lZx25RYS+OTtnRvKY4/fbjes6uyWvjlOWElSPTrjoOmK1ZYIiwpE
qJBF4idA7UzoRT2X2ShwZN86kAyNUMdYUQJx6HPnf9fWA0hNpbaFa66L2mSvKOdL
d5RfE1GnxW2rZoPK3AohcQq096Ta/qPWQqvbciyLa9ZONFCq97tDRPDTbM6qU8CZ
gnhZvWdcjojJAN8svtqqIiC9lK/as9b3pOZ7F8TJTwrO8QtiuI2Gw1qzfQ7sZxqZ
/RR9W5LvlE5odN+kVj8fhISVuVqXMySOeH5+uZNUW+cP4WfaeWENKywEMbg241mF
yuvSfv6s2MIzsQwqiFPB3s3urMGq5f95kYPfOSREcfN84Dpvvx7qzKghi7nclhtj
2J8rSKMhLVipgerbP99ALg7b6zjyyW8vGykj03biG9ZQpH1yiEb5dEuvejxEv1SZ
aWkuYkcfQg8Se6MpesjaZc0DRzQwyWkadcPciRy0QKFrYj2trToIy+ckqQGTdlRj
U+A3g94rXzTppTURv8uQi5Dg4ARXYRfWm9jRBo0BvK3QNatZMQ83+BtfWHEb3KQW
vD4hnVS7FuaoS091G4LGujD+EbfEQ7bD8pm+YDE9ac/YUdIJj/a7JsqHvdDPArWy
o8b5ZVJms2JjwIf0qg6cPcQXXJqMKgaDWEYU8H4MG+ljfoYM4rRlePRpY+BORSbL
Xsan+sYHoNqj7pPe+64BX3ozxgSAZzMDoLnMXNY+1BoTCqHewSva+/LahsQSwW3H
Z8uVWbnaYz/l2syGW26BorSCjV2CmFXvgU1i/UR6rnlOsUWBEG5cImwqeBaRSJca
v5MMN4OggD9zlVw/34yjLDcisN5A2tkjRdGKCFF2TASW1QWaGk0rocUM484rUwt6
71mJMlO5pmd6Y0awoMJorl139hSrgdHkDpun9nyRDdHjGlkUI6Wzd+gbC5lDXqgN
rNUqDVXzyipwh/qQ6iT6KsvHLvyWPw77Ad9XVSxiU6s/PTyF5b5bvKqLObXcHwvj
6+PiGkpxo9alVnKBtmBi9nxHdKSvi8GgkqIXrKPeWlwQVrIugkTUrmBc3FuG0PFc
D55UQJ1jDdNEGQbYQ+uoTg5wAWvX27l/ERrRg5a/xFZ2FsIYdBWT924CUMB3dvBQ
WJr1Mi9sCnon2Cl3ierhDmFbmDEI0AjA0EaTnK3A0O2rcEt82UkKEUDt8VfSY2YF
zUnaZ5eMy8WquDb/QyOghmhPBlTiQM+1r20bTw/GRscCSXgB4nTAcMI1rK0uwmXU
nsqrx14y1mvOBs//+9P81+01g2aanPQ0Oi9mgy6POryx3PrJT3RxkfgZs5Qn1+zM
Me7iBMpbnXCM7wHKGyBBqo/LA0UQa2DKM9Ot/bZOnX85DhAAdOf/UrjpWGcPqIw+
CXQ1sfZSPg76SdXwp4EN/Iimbgy4VIfVp5WZK0eoXawvjjVn/wqznltXkBno3f/p
y5X/YnD5f4andO6UrUufDE51SuasgduLDCuqnzacBjjI0Tg6+pLS26SvKbotaCiL
uA8ufpvqh/okLq4xSOrmxX7n6cLI2Oz6kvlLmB+xxJCgrlW/VHo6cOL/rDmTK9Gs
50zvwpQG0vpvCIzzqJKx71TYwdRgcDpRWpIC+9ZG0X30A1/Y8Vb/FYxEdJtz+MA7
1eW3QUo1b6lBuL1UXPky0kxM94O2sSS1ls/aoZNmczggvSWjB0D8+pqIwK0X/bGL
n7h/mYCyFy0YXUYFGtlYN5hBiGAqyfUGUt+zOGto3MMLghaVE6XvL5aOXnyUOygg
h70s3XExfrvL3Whgq/sYEpWP/Q7sEnwSzh7Bt8l2Hnl5v1dPjIpBvWWyuczj/7En
wfyfGCCLB/rcq6/fux98Pe4spuB1g2cirwWMFMHMdHQgQ7bURZ2MtL5bCYa1UyHK
CyFe1ed45BIFaYxRd8F9GvDGzTVb6EJDwJ+xrC21XlRtXBHiVlAHrNfE70Ekrv8G
q54ny08bHeUUpcfrvX69bskELE3ftbc8vWVGAYVd9Ki0ZDGFGbYCH2qsjkevolWF
Fqhi+5ud3rrkRDYcTaHKwhaCnSMRf+XzLPO0evufp9gF1XggFg6/jvvRL+mOZA9l
mb2dZX4j68pPM3RtKx3CFmflxI/crizdNc9oh5fSKcLtZCEZFQOFruQ/55YimJyl
cg6vTzUm5YsPBELisvZT97l13o13ekbjYUbdXOnyDRmiFZ7Q6Z82JO30dQdDth4F
VXuglkghoD5nlgnGPu4OK3trxBiVqxLFymLPem/t7Y7Z0rX1fmAzWk+546Wpq2+K
IhsCTtK4//FzfWdCcq9SL5bmZxY2REsak7470O/Bqk26lKl534xW+9guw+B039/t
jScAUWnSWyZB3p+aKKJtr1tc8G4sUjGQW034pQnep3/fIErqd22dvuU872xbpaIQ
LrTrb8TRni9YjJmA31riTEXtxeBlFbwhgz3gyMOE0SMyAJNxr9bx16sDNiOVrEEe
nCWiR23dNwB5epI6eZ16b1SO8kMtDqE9AWWYgXGN1ym2VV9hxZQtevYQxqcyCNl7
5mcIt6Jq8IQspLTewVl74HTj20HlIT9bzrpE7vV2dtz0KUWM+cftQP90sQwQBxJZ
2NxQo5kE8uTmmFfHiqB0TRmqz/qoYQFfmDzIlawDVA73hJ47Y5p69y1pKWvX3FlI
Flk2eW2j8qffpilapcwpU7l1hunkdLvPeV3DJzuDFwn3aRwg6Ve6S0oBGsKgvWMA
cpEHKCRJUaoSUKceXCTOU3ZyF5WkwihKAxrKR8dk3L/K55SzrOUWKX60aoqrKP6+
tUIwFWwg4z/+HxJpBtuZyTnYFSfetgG4spNlVgGNkxuvWii1BOYySrGmMKBhWfAC
haRHHDnKcECTQxyF/FD/Lh29BDhoJR4gKZtTT5J9MOXWGzMhLWBln88jky6/xla+
j/uZtNs5A9Zkq1NK+OpkMfKK1tLUGTSb8CDJBgFGyOXj/dzSXj9Ghse5tpdnSYgD
7+bTSenNopYpVqtG9tcW9IqWEcY++OtJNtTBKJCPXeSl28R0rVz/mWNfkdMSmHfi
vlAiJj6xF5bvEiF5J4ukXaRgxCz5pmAo18NhXhSgyShx2M0Hb/FsJmSOtJoipbXD
/nCrDAhf6xwsVdNJJIdB1X6PIQRnIqCTaWaFuJwlyILwJ8ozlz2kbtVFBFLLosUh
Yc6fllcSXNo+YpAfcUeWSKjypnaawmev0LCGQQNHfPhc9y7+KRXbsU7jGUpaCBaX
U68K2et5Qs6yPLq8mTNhl1+d3EwXmMbV5ofHGzUAsBqAc9+pQoSz/XKLRvbL+nXj
tBY1eSD9E3fnk3pLpBKER11us2OoEnssP1n7nlCHIToXTme9q3pym+68kpWX5xkS
JuKJF1tFg/bAxN3A6dz52N/XayAD+brwWnEscBAhAtYz/jz+Lnni3MbjKuhnSDLo
4tkCcHKmJHTqonDjIhq/qntXoJm2IBV/RQteF0tf1EN8BrhzraUolpz8xh8+uAnh
mkyKw2VfDVdEQbyKaqzzg5xcCqnVjH6ZvqWjGJb/qYopjJtu0U82U21H7sknVfE7
0Tax8afHtfuAp+vbQv2QzOkPQvKoXmiFrg9sAa8oY2aGXa0sj/Treg+ckNd86J+8
w7N4ZkIHoDc59gwZ5OLnRYOJy3/bvU82XqGbT4dgnNCaCdJmjqHr+TI7nGQF9uZh
/pHdQZq1/HTLG9OfMUxY3mLBTYZnvLxGZNpzkB2IGE3tdPeM6d1sPVT7Q0bCqqjW
2OLGauUFiB28kdonpaLov6k4Vb/cBwNWPBu1NXWa/MsgbXXwLXmgdf69y7P9dlRi
eAq6oPwFzslCBgSVi6XE1acukARBMVQpoFHbWvpTz0QKk2hWw3jKfj6yTWUI0fHe
Zxl1cwH0h7ZixFM1lNSqLSv4mUfvSgngO0m+QNmLy3XNXYrTVQOknc9S+rZCPLUx
Q1VeardQAK9g/d4BCfyGtz8KxzeTEgkb4unfrAQ4RjSbuzCvUHcRfAIN5SV4BoRZ
+d7RxHtl4O6oitcBID8xakvshJvZKxPmTukkeJu1+ePHAELeNg+mV96Y7ro8a8uF
gv58gJx1wUf/exsqx/U3PiJiX1cir9AUoe6eRFUXZg/w/OQ6ZkHGs+dbEunQTUVh
6prQx6aVd7vn+I6vT9Afp8qEgotDAsaWJjDS9PGanwazQgWCs+NA+P4FSYdxjhqK
HYVpBcS1yrph3kR6Pbrl6vyIqU4ehxHJ5XMYkmi3ZGY0tAm4zLAcEFQLM8cK84hL
EUCZVrUNtSv+FDTLrBw3X/xEWS4b4oCahZ/FNQoEpciFDuXERweO9VkyuthoEZ+A
TJLcaEIXIpy3OcdE3jKy94TUQJiEyGZe7U8DRrDtVsG7jv+7sel+U4o1/NqJiTmV
fjjBSEoLcDjcnoEM96MWjMsIf0Q/JfOY8LES9C1jgQ5AMjQZc6sD6GSfb3CRoDaT
IH/kENgiYBEtfu+dNEiYltyvyzvcZ0yqISukHODIfxKQLCW54pWUKC8hBxiRBzaW
16BNBgOyTwoCwbktKRijXLkWVllHL5Q+3+ONy5Lb1eNGoiwChn1th1JUU0Vgk+JG
41+ewB0Rm0EEdmBdrvRfcIIt09hmpyV4YpzKw5p4foHw3xzdDwUfqNiebBqSK2/y
WBCz7yHnXeau5fPiLP7lHlhZ5NxQCTrgt6bfhs1iVKNK9e6LV6qh3a3pIsOl9WBJ
lZ0Pcs8HxywxufWNhpAhfDSM8kW7ZhdWvEYUHg9oBgUmPa7/Es9YPCXJPn3PDMDo
7Qr08GaF2NOIrchn//D1pqPIJF7ki55Q3TnOR9it6dhd9r4S2KrcNJCWBeK4xASD
2CXo1YGv5BwC9qoVWLLAKSEdue30zO4XSp4R0JPmjFH9DsXhUyJZLRN+233XF78v
7fK9ImYxtcNwgRn/cWTu+W1aXpDNyZbobzk170MN/bC4gAyaLKdSWGOF6BHPwHwB
r50cnOppH0M7K+6o5WyUZdEBfeFqYhZaKproeJvDRpgbNhfINmwSKApl7G/jPCgv
yCXThlvtfaUs4uEuF+fxJ4U46mvti3ktlMPeUrDvHuvkTivle6/oGsv54BeC154Y
nfWF3Pf3DiKGUL1yVVsx0AG9ecJr/lm3rH4MM05thwejoay+b5xsnFvZb0Qx/BP6
myrUe60SCeyA/pfRtiHOjXsBUgMLNCQqd4gbILAuDwgMHhRO5xDKA1XOMfQY28nW
htYLo1D7nWElMjnfOfg8mUPrbxDv7O7c96rIlOp+EZcsf4w7t616ds76MKxNXSqY
DgkwYIMpP2KdhGc3lFqZgLv9SF4AhC2Vl8Zs9rEmTd2G9P9PbEaNBLGsAeDrq8K8
xG138+Mz+KCnSPN70hIQ/De3iyrsEkDbXqTlUrxQT2mBpqn5ptkbMoQzUpURn+un
urg+orS4gADoUhNny0dMzbqHkTzXBigrEmSFsm6UV8aiw/HWma5+VgIc1eX4EcT8
2invrh6UIhu6dAt+0r5X/d7Ye4n1JxfAtb5Kge+fJOM6d2yekocRwNc3q2wgqWdr
SJMhESB9Q9rJ8rhbPMGpfsdpK8/j7UpO/RCT3DWZXnsBMftrVUGzdu2ie4YM7jVY
kZpPwfpVsWewBwe6/ENmf/r9KAvyPHxAVJIk1g5SDarpiCTtHcgNYEnMYwXOWk/d
S17rlNNxnQDdMfiHC0JwNSGkDCVxLfLEdGNULV/wSnxVys4JdknhjCg4ixBQWVmr
lkXrAaIf1uykFG5ERY4tPJQhIJZeNpYPqSCML2Jz5WHrecWW+DyR29/bsBDRZUpc
ZeafdRS3r746wBnbF5EUnl6Icu7OBw7gBm17WtK7vobLu7ggYBgVoEBISMD+jelv
HTtYoAKcfhJVFGQknCD7AVy8E9m9cWXN2Lo0bht6CUvqdgqO687ufb70iw/NS6A0
t2wo2aPCEp8VEJ7uINTn5oF28oUVeE2hIyK7IYG9LCjkW6t0IOo4g8sBvQjSpsJi
205UPv26sjCcFizFIfZha1IWFWNUVnmsm9QDzRKQVZ+ryhM9S5JlHi0ddITljj03
6Su/w4+QPb+QP9CaoKE3xYixQJzf6+eTfafRiCairOxXDcPqfuwbOXtAmDXEtEe3
Gy+lb0K98CzPkkBBTDcaDI87ShSma5e8J3xw+Xs1tN0QEBaswCyLHda1PxhYWgZ7
+BQqDKvRGgCzyd4FN2iASJGCZ+IRHhh0VeUywOoxJlD3uCQi7vYK1eeKql4n5vmD
ESAfpJKS2zKhe8/o3oyp3F/zO/sEB9q5LvRnanjTev12JRbbrgLEH4runrlkTDED
ZTHe+3KG2O9M1uqOB3AjRQLuyCEqg8Ckj7nbWXtdDXp/1FpfM+daBHvRd9RFT7eJ
xjukXLm4NQ7ISkf5hec/FWs/P0IDdYH7JW8FXcipgNODe7WQUNbGtCS7YbYGJGuH
nlvisph4gpfYsZyZGw9ifpR7bq2D5IvXf7n7woT1cV72f4MRAoeBUnoJqCEvS8dn
CEpYmJFx6UIz7xwt/GmiInrCw7QUVCCsVr8qQp5ijqaE0WD3FmFOic3p/m1c+h6S
KeT2fDD9+l5sdta9JY0+9jXbdxvmVCOloHbBR6kMQZTc9heEHo4i5ZbirLmqSZ8O
1patQjN9oVqXvDNztvJ8TeFHdF1/lNiBE5tiPut4HN5BMPJkm+e8afARC4ZU4iuJ
wdF/QF8UC/jve3cVA0zl2z9+LhoVLzbYFaHBvUd1Dgyt2D2tPtVYrzUebBShy55e
kbjRzNX7XsbDKAluQ99vSCmWkzpnGFWyARIy/qW1a7DZHpVIZbBxHT1Bs0bJdXf+
pKlPJ+iEzqfwqZPXHZqXzGpX2Shb+Fm1YPVrRH9BLl3REi8jWvpQucDVR3XeqmJk
wqTWl1r7WmT8BfaeIHqS0c8WxVUb1DQbzgnE/lwdOqZVIwVsgCdXwmznK+DzkfwS
a9b+qYmmLRR6XCkORnhcpy24rKhO+VtRjyh1LvP0OVzbzzXXvVs2jMNchVVVsZ/t
vYo+l+VZumObH9daGxw8ZehRqaRd+8G3VbftTPywkBgHB2mUmogpAQ+zUt3Aq/KV
6havGPI3mvnysd2jKm14Po9PSUh4Kv2s+QZqi/zTLgLZPAOWBIdrORb/g7CMQWUH
wvgMUj7hLL7q3ILNzPN9GxDa34RlHhtMXA04EenJuFfJv3pJqL+hJgXjzXRinljw
EYEC95lsWkYuXJg5MAc0L4HuxB7lmn492bXjgHyXJN7ue5Wvy1hyE+SH/yOrli9H
sOQ9qn399N9W5hphuByO8qmgM89vCIOTeNdvLwEjhhxZ5KHEr+CTU6Cwuow4lJcW
hPj9v/F1ba6A64V7j5Rg0vXSnkNssiaKUYfdff/CLmwtFS+M729WnMz7owb9oFlI
FyNaxkjw/mEwU1AjN/QRG8Q+PXCsUMuZ3TX2ajvY+cevXmWCObQfUnsTDcP3e//E
v/Bzk7Ux9lez2KfbJOpznbhnRNP1GlMUXzHoeDhIc8aageTyalzx0iI9cRgoY+KN
h3Apc6pSOrMXCEMQfAAsM+BKXTb0+HYvIznCZLGMfUyR9/SSgrbn58AXFyxXAO3g
+cOD27caIHJZPh1q01HTsAbI9kGKa3s9Vefrb1rFS6oSe0ynQOcVxhOljLn55tC7
E0zovP2DuMi+12fDPCdIeSkSOL+5zug7ftq7YlFoR9d1rga8JjnlMjnQJdj6BTlw
MU2ybjDXmsulJaOFDRLY0L7YcD1DW62gNtw82qE/nWj4GCczIqhKXtysJrNo9urQ
pNkTlMv3jmkSN41KsBpWo+PGLQTLTPIl+l+c+Xv4T4rSp8ZicS6mUw3OraBWZ7ox
5N8iIsw57RPFKclkpS+/kWuP6f60g1lL10S8WaY8n4it37e/l4lKL3dG9RwYuIyh
uZyOhEBuCCQ/v04MwSgZve2joEMBVITw2jHMTxAXOJPcMfRZVBjK89PnTWl+Vcnx
TZEBuxWybTtiU/GgONfRebvsCs00HluSyL9ObQVvMh2iTGd4aM4BnXnwad8fxsLx
CdQG4b8qJepsymnlmwFkIHbDQ+t8me8d5IiiPuyxqn4lJep7Z5BGGZg3I4xV5mfq
Irc22bM9J6pt5iUm4najXkHZp4KMscKyu8Xs462o7Qq761akRk8QcKJB/5O3BBB7
0YSpvRylCI4pjkBxFsJ6NPjyjxaKAJve9Y/hZqtZTr8ofrROskyL2Bs1zNpzieAe
Ju7hF2YUwL8eAinRq7yKl0lJj0HqpOkpFd0ul09BFcykAQOCphjG6qim67V7xPT0
5fJLuvIhMF2CmOKBLf+BsiSBUClGrrvPLYC8gAGSqLATxspNThbbJfelWezkTvwM
5A75OCizLWrCcKd65lFgNhGz6KaqpGABaOR620KzLTNFcWRCjlAc5eeplhfPFC8G
PnCZgaN1hqBjb+KwqwefT+bdaEEq9E0VUXxJWSDs4Ijye9r477hXhGadXzPLtj1r
OkbnIqFBHXlAzABM8cwKlqlyBEBOrcS3NB7oVSTIBbZnCZz6ei3dxy5tgLMl3l+5
jyaS/+7Z6lnDfG3X6AE4qpK91KO0p1ywhANbwLPLTiq9U8nWWJyIHtGyilRnJ4R7
U0mKGmHFVPuirmwGs2SZcfUHNVFfkdVPm2DqvYlTXT23G03Q4f0KqAv/27nqwINP
BA0rqQoDIqmlFiFfNk7q3xGLEVn5c004Ci0MG5I3JLxKOYsuHjnz0/hOZ8KIMyRg
fRfO5cGa2hClGviWXNrSMvM2UkCDlWTZm4rHcIIFbe7fU3iSj2iiTTbi97wsFGV1
aQWyCBvXK2qAfmxGzM1JTMliQBbXQ7rK0UOpx7wzwJzdUHTaytvoReZxNildFhyz
SXhFqb2AEBMCj3TcafSdIxHAhWhdCZt7cIl/t13Gwcjzfknj/RewcDNxk5lkbVYi
iPwF0adv7/it67o+hpOE0IIrBFOi+wU/EcwD6+wkBF7zSTSCG+7v1Q1TinDQwTJC
nrANUVlforsJqGX0tSLpJixh7L7Fj0Jq26i2w3O67YttzCDzW+BrcoXG9nmzzF97
GvhCPLTS/1RG+UVUNzi9jBGKCbQrXTLNGWfBdgK97CObyRYdRxqmwk4rUuBEyQ7Z
pmRb9FEwxm1gecWL58Atx9HMbpsOY8DYXhEmjMeiwsEWx9pOmFSnEc311ykJNsf+
HTPxDdf+piabUgpKwArdKnMEYazBQU0g455xdIVW+s5Rc0LZij2UzI+I3BWiqXgX
Eix/fBEHkZpVqbUvyZlD+1Xpgd8V0wiRe699zTXIv+zOpFhkIGaYxNBTeWlZL1OV
ENOidZtU4VFB6o+aL57o3kj3a+78dAtbJ8Kc1E1QrvACelkC1tTuhWTMYLiuNW0v
im939uQmni3vbDt7UcwYwvCxyjDTYC6NJ9ucM6V2KvElEFv9qhyMC1KZVJDmNbej
wTZt6EckORUdW6eNKmNvKiey5maEx29fa8LvXiajbV95e/nIIrt3akyWbAAH4PEa
3ZgSCE32C04BvEHDeA1PgMlgg6kgulBeGGguQr8V/Z2BuSLvfODgh18gZ63Yjjp4
tqPZsj5TL9eVju5Dwws/lucQgB4QkJ9usfCv852nT3RwFyPML08UP7L5BJ3U/wkD
ois34pCJF1Czu3xprUH0RL5wMdHLqCyQGNt4ynAtx8/zN1jT8T9S9kitFMLevB0+
HyQo1dqYQI4oUJ+6VOHo8i7FfhHHzkPnvljD+8+sbY0y0F1KJInrKGezDhtWzRFX
A/3roUr1M7ctO24xVG0QTj5miTBKH4I6WMTcCb9gTQ5Jls+xxgilQc5PH7lSFpT2
xbBkU6dR5J/QmGXqIFpuwRJejQeFDkPUrLLFjkPcibgFT0jGqgnJuJAVbQwsfx9h
eAlM/HVOrHskRyHYDTcwsjKM9m5qTAdSIckHn9PrlPoT8dVoFITWyd6KcuqT3Bpw
d9uMZkshJ2uxwN+LRzaYPRhmpeAf1J5pJS4IGh0paw52vJ1B0SYx6CMyQreCVYtO
EYpeDjkDBtFWjvwkdoN2Rpr8xAvMwuMUawgBYwUNugTSrPYbUuwt0FEMHOIjJPIX
kxYYxIjmggP17FaIETwfEp0g5dtUDKRtA6Iy37AwIxqjeBcRVIa9RDHt3FJVHSTf
FdLMZ4oJhpSuryUGTcvxw+xzhmVV+MiCPIgZDvroandtiAKY574EPTuKogIHykxK
F3QrBng9K+ob0YQuvPyJPCpdQMnjZb2vhd7IoV01AuSHM0caOwBK57BxqnHhMQHx
KzG1kZwPVZJiP/ymtdaxotysk0YSZgy5bQTceKSnvSkyhY3dO56F0gYZ2aGI2CZ6
98Tb5Rgk0EWevfAuc01fWD/58gg1FSgSg0Str2zkFmD30qvbfEAiplWzmhl8zBVq
AJSkYujmHzMFNKSD8j7fS384WqMAnSx4vnOB1/qRH8tJi4cRFVEr/kQeH10JRZjx
/K6Z1JsR7BCecENzlHQDt30+qa2pk5tjKiJ9rCmwcsCTt5zHuulBL98etbV6GaNe
+PQQsXNGQZOlq7r5afC/wZtU5+MnKbsIEl9v4CheOwq3AWLYKG4rNkMKsleizNaN
8F5oxFsNlzQTdVjKQ4zrxBExcMuh7SGKl3KZeGneMXcp6Us4AoyvkWX8qDQmG0il
4gQI2FBT52c5aGnCO9JreVssMos7U/RmMOjkKNQKXB3LbpiVL+ca8HQV6zcznOGN
6tgS8FlGGNPfJvkr6dF6pAI91CobWFtgVIao2qXnL72xnvZKpwdyXKtp3A8FRPWS
8cqoPDGliwfUXrakzFfzyZ0+aQdKqZfIAyPgAlK5HJyH44CNzKMIcRJViv1iWNur
DytVhNECCghqpObbsECDuR4Cr+kLJ+PsNHAjXxChjhu6BCFUsOPxBAO6vg7foyI5
ZohugsmdoXSR07itrKVtwAQEssuESXc4w/SvFq7/lGbi9PUMuutK6OUmEQ81PCzd
8QYcHhtbauTvs0zQwt3agEgX9sGWemjCG8Jrfs69AtwTpriKk8E6IaTcuOeoeqQp
ITxGkUjSVj5Z/FyT4/AFILlGD3hb7KwA89CgbfiQ7UZo+3g9JCSf41gW6ChODM0U
mURKGAamfXz0XbBanfiZcXsthlMGQdUv70JeLJJJ5sMMPahkU1zdTO1aDcYUjZpX
kSyZawx4Yaf4rCSgHUz1jOhaLCywrnPw1EQMWRUQlZpJx9zX+cKPCOL3+6NfRQVK
wuYfmBS+yPm1RGNKaHxQcqigGmMSjzn1TwLO/4srAdMt1kY2DV4xjqeGGxDmnE3k
5Tr02FTIGuOm+ng8jk9JtksotynM4q6HuNq7Dc343WkdLXbRHIlEblR0EMmy2HPM
RUNcFmixBzok9F+TRJbfrBulT5gGw4PZ40BaqwETpOly4i0P04Vzs/4fMJrEAIEF
9mQ/q6LeiMLBk1BHGBrJ2NsOuHBb/YWgIKmonFFrv2IkdBA6xjUg/wolIB8H/z9p
Gu6td6aEWYen3XM83z5ihFh8H1501Ah/KcEjw4ToHwyQsiTY3RDIOUBDSDD6P0By
VAQXAZhMJnwYHeC6qoUbHVIUhB5rO5efWrUxjTUacPJq11KI05w184IKiBXwrOZ8
xeqE6c9MBl8jmRVuSELhkNR41NRtT80xkN8ae+0pO88Rtgj49WdxCBLM0ftI7UO9
intGflbVXvCR1MeSfxo1rOPbbT/bMFjSTTFFfQefI6BZrTUlXFTjrB5JTxsGEhGl
tiXXT9A396oFTnmNjH/C3AM4bBNiR32aEJCce0N3WvEUPX0zkcPvixoVVbHpbf1k
+2MxZo7N6nvnPFR+B3M6k4a5QCsHOGBGKGwleq1VC3zKLmeAZYgDp0svEXiviZTq
7UatsoDmIejby0SpVzlVxZ7/h9VeOrXII0VcrXY4kzsyS4//8xXDIm0a/3pEA1Rw
udgyk8s9H8KarXGZ5J9eioq56+24T/Jhm83yZj7R+PPWJssG5KrCS/lg0giO4VFG
1cyp11k3mUxo7Hr6OF4708fs++L9UKJdEdfvjVfgaQoOKIAYewpm9t3/OGLtwgqm
5J5uMRFh8mjVAke97gxgOlCiC/6vGVFDsUoRvQThTtsyp9nyjiTTTyNQu9hRMRWc
EMhCHImm4e4/e9wLY+SLtE9M6BgzmGTTxAOtjnocID1A8SfwqXpA8nQS7MstgD/B
Ef5tiFm4R1lrGMp8GZVtoTFLSrINVhBg2XJdeFdoCI2TjJZx31+is9rMoYT34W7W
DhJEQSJfE0dnCtBID8TBFW07R/bGmUQzz8E7fyfSDxPhzsCYKE0nshUnaH3AVLxj
+WzhMJtezGAP+HrBCcyR/1qDY7oQtybLyo5iZ3FsWoBkypFOWrwADQdnfY7jkxed
rO/52BMqrGLyH2HUSDRGQNsMJL9Cb4hePgER0uXKIYhdGx3YWObCOP0iyDKCN5rr
INv2D6S8GvTV2wg3R9wtC060NfKMQ1fNENSPrIbzA1n6lEUeRbmZeGqGOXrMQ3og
L6IfAscZkjDhhDMwIdb3IArJhAtyaoNcPNRj2XOQ3bTGTo/UWyooQQp1N3OANSoi
cS2FevlYtBJFsLAnzxp+bIQPWD7gjQk/YHbCYMXDuZywCghk97PiZOTIhtp+WpqF
evY8fWpXITr3vBiCcnSHQbCej/YMNPn8c4Cfxnxbo8gcIQWCK/AZmDmn45wQu/nu
3VXKBYkKL2BssL08dS47+fVZsQoT/ouB1rSnL0ed2kh38NiDxxgrkalcF9kHEbi6
F8xMsBFlYVFqZyG79DbnOVDWT2MweQu8gWmWPEwxhcItbZ7YD0uhOS1wZxXSAfRa
L1UCV/mGLGmyDMp21LRo1qOSptRiyPIEfbwbg47LQmErF2lsXqa9OlBP/biMEiOH
llVRA0a1ixvc983Ooh8vaxbdefKJn+lqKbakfBTnQYmGj58PvdReGy8jFWGVvUJS
BWjGV3qA97LkyDZMxb7I4A+DttCLrEyb+YB8wIL8n9uq4rRn85j54ZeElz6n5GE/
bIWSEUSUrNT+SIbdXIoptE3JyKtmU1rufOLF6FVpfUIQFVT07wpM1mUNUk/REBWe
xdinYORDZhteAekcRh9ZRj2btrdCHasP+B8PLjI3HrwoZIEh+KDb65bKVHgoFV7X
4m/50er2cHa01c0VRFJuiVFzCdnAVChYD9wNpUTZ//gFxYUuxdyU7tKJUDGLHLIl
exWndfhPfWy++oRIAB4DwD/9QZGUuSKchBgD+yUscr3KWEeiFzHvsKffZcT5Xx5p
8gHGpbIi5bCUGby45dY2eO4UB0P6di9sHDIT9pFKhaf8J1Q+Z524Orvlg/fSptOj
gxLU1+1sw1GTfC9Irp5KAB1UtD559JDvbImLQ4reswhiiTsLs3qtCbN3expGoN17
EwmzRPSGY5ZIPV7Zjxe6BxpVOOtllmAg65DnVkYznaz9m4OE8svtJpvytsdhaRYh
3JxKlb/p96QnJ6s0BO/qGUlLOggUmZMcPZ8/hwcfUdXmfytUi4hFPHAOyIizz1GX
xVZtagxznSZJrWjAfrDfMzwPV8pcLp6PhFeCaCWKqE7GrgyqYdRc4zxkuhj8ayaS
1wDkdcjleuts4kBNwrnJRTqqHEh7UxX+N6D8B7OZKAm8OiK6vMf0/Ul8XFMGNAqe
mSseEE+T6RPIZafOath5XuIjcqKlfe/NDRmjpoXkns3Gt+wJ/MkcF9dW02+kl5CP
Tacu1H6cdkFuif/WwZ1w5cyQ73Ss5c6tspMQX7gPEdvnpo76/7xBjT5Bd2lekt/Y
lQLoWNxNTwQcwztho3IFES2VLqeyF1vR8NcBhjQzC7S5JO6RqqYnOaWfhEpNZd+L
L/UcWjO5LwYrzBVixrM8c6DxesEIWruX54W2L9EANgxzYKreM5uiyVrMJRlCDLCc
idRncueLOhWS3oLja4p5ZIA49d2YeQ1v2UkYIU3L49swYsm9dCVj0l4ZcwckgVZS
DtZKM9cpSEgw66Ds//tJUs64yJtVaxBaXIteGCTilkG3O//P4i5qgDbjk0DHZcCc
5XuuWVkKjuckVazELtwqhFOq4U75qRGPIEyGlgSIf5b4BoiwXum5rZBqpLiTNMZA
N2R3WexNNOYK528shjUIQLDiTv72emcaOazePuC3NhGhfpWtzyebnvDa/mBap4Vg
sUsNwsHmEPS01tbh45+NHATdVMokG8J3TcbsZz5hFdz2uRxVnDHzK4VlSkWPU/V6
i21NX0D++MbFievHk2tl7CPOE3umNe9pPplcmTI36wLz8ln68pZtphdy/x4jhDg+
kaWopChGalhipdiixWJJkOsBnWRTYuOCNjYPLSxtBgMV/iZb3To/co7LohZLT+s2
RxC+QDG7aP+QqJs4ZfxETLY3zY5upGx/SjW87hAZoUt8OKoK7D9mLTsUpjlqCZrm
+GM/K7wC3M9f5tczuW0WpKEMqnW/9CamBJ8ceP3vYoXjqzWvEirO1DuDITN5ehg1
0JFvM8q2XgdzTkzc0MmXc9Kv1mbY7EcRDv95+MIFEN6tCMGFatREaLSnlNcsmiyM
xMJX7PAYhR/LSYNO4DRuSr2XXdeLOg8Ed5nxzfNulGmSxiNPRH0rvKkDMP2ifcxe
tY6rI71ov93PEggB6GQSE2wPozQXdCAbFdb6dtEdRlQwJj0NvqluyuNXg3uuuE9Z
m+aeCbnlIqgbytqkOR3/20VVXhk2EsBcp3UiaYWOZEfqX+jcwcIEFJg6ngUEW0yv
bGfkSq3tISkqd7rOQcTCUrXjhiiXl91JCd3nW3/wbVm4M5FN2878dDjYr5XV3BbU
WxfNyR+WsRAL03z9l6wvOVKFy9MnfKVw3yHByEsIRDzy0L0p9uAGWUrkpL97pfny
7N+dV/AVREcmIQZG3dJci31Y4Ua8UNOr/Qdk2nOC+kqKpvStBdAWNAB41pMUH+c0
att58euD2iYi2P8M3RGK96LgvSoKOcSqwigvhd+St7jd/NIuaVVdySh2Wseec+AB
A5zPlt7zkNUwoh7xzTyjUg3mOabc+E3l8fl21+6uQfzTgl3bx3h5/Qz2GkF7rD5p
qs6KNbql5gBaOVSf6fIexoGoGFml+0/gmZ5jobrOSTgaw45TM+11z1bB1CgzD6gA
JLTOflUJDglsojRsbY+20xTQzwXSCSKLFW+e/m5gNeCwvu4hZOoPaEUcGV5p0Snw
pjLXUVoHE39e2EhoD5xZ/mtqzPXxq/ZQqsrI25GDH0Ay9rckbxVu/JtxwVQQ0/MK
7r3d5LxIHSj0aiBZNKecvCeBWypsIZSl0LPAE5dfvr7OLbTOARqPn/Ha+/aCuwFs
Hn/+jHt3L/JvC9UWIUZsLpKU9uG3s91mbibXr8lQl/ykTbfacUraha+0m81FotJe
JDJSmUi7gaR9OpE7+b7BrWw8tCXJWCtt+MwvBKVy1huuxMO8l/duTCtZNn8GnGOE
O3tgyVyNk0dQfDi2CriuQn3iweFydpWtYeUeYSuy8eBEuHHbqt8a4XGq70a4xUBh
GzI/XUY29QPTnPatL/QGvMjg+Mpgpqg8kXBSYxbAwBeL3RITeqE/iWeH8jiMkbsh
sEftF1ih6qVNaeI2fHc5ElmcLzvkTFEM7jsJD8a4t3hZpHpn89cHO2Vls12lyn8z
FhdWgALN1F2LKyN6KcRMAtCPiOXdrO/ik0PnnIXUBtVEL/h38imhBlSqcvV6iYsJ
0sSrj50jZmM2orbAzM9Cpz1odHcFj4ji27W7O4dSamEHy5rOruugM23QYWKGOYZV
hjPXuj6W/JELF4p+vo7+3gv456OiaUO5KEJW+l3T4lfWKwQ1uMK3T7h00RkIZADz
GVVtS2U6VX9AwXGfPYMB1mZSb70Z58v6E5Q45HPtQqn4kaDGOUmX3mNFf2D7jlLC
dVVTJ+1XWdCa9tsrP4BpyHzZd9eEoB6I+ahtEY9BQ83+Cfp0d2m2A9J0LJP3fKYQ
DoSYuAXcBZ23xM3h3OkPv1PZ++LMdLlHZP+GAnAEqc9mHGK1FA3CeoyDaYZnc+dM
A+gduTUdNhQuBV0Su1LZrhj5phf4OP1peTO+Kusdwj9/NkDauzkFCZ0Szc0F6p/t
McROnMAknjTmXzR26jFNvr6JVhP8QHoF1D5PLztB9ZkN81mdd1+TU2/HC8nnoKhA
TO9HT+R5V0+9WlQJUEwpm5OQWIqKR0cNlUKVJ1V0AMOLycIvY5lPET/2TyGzHGUm
yKao/NeKQj89et10Wbna0kpPOGkN++Ee4/UaWJX46ekQrpOwhn7CNfcNZY6N7vEH
HamqAf5XKxacS+b4dnbyVx4UNSppcXUk+UeQ+YdHiTIg/tNwEcpoF3mxGmZBh4rb
oTIthNZBidkHEwzxsh/GRIioVk8GwOFQ+ftr9wxFw9Ibf9N7EDKC3UoMEtlIaQjl
GZm8MATRt0/bz7LOogVESAZI7kHq99E4VARrf/oS2LMMOFItMYO7EbQ0xDDtWbMa
dvO66RcSDMAQSHRSXPz5Y6TilDRaJ1XRQfg0KfPRKa+7k0wMrTqWXuSpWCvr3wVa
7faXubPRBDt/eWNpgEP3a9F+Hzc1cp61RLQaq6aN0K+5r0zqS7nzBiHUTuEJePu5
YXFhmgczDf5/MYFcccahA+VVg9oHWkqVyWTDaoqqDfOWMlIET2XXtPxDGyyPY5Ov
dru1+LTw3R+qTYrOQ9IvxKJQO7XX0RzymPmySEzGT5UkXVAFSjO5y86ltuovLPP3
dVXyIMgR0xRJB1c8AegOIPuabdsAubdFVIEYUNMlExw9F0bG5W6Wr/K1KfYElST8
WEw+fOObBC/dPwjlYjiWRCKsoeL5VJcE0GbDbwbqGVOgufvhHdJl9KraeFWzoUKI
9m/Z0TWv73fXGmFiTV+E7HdHonVIMrpqf8FsMxyJvxm5yvs3BvuwMJ4D+eiirhQL
shnwpfsi4wEl1/36xZctSy7g713OOi7fvaFtvFDcdFg2XRmN6uQoToVbKgQBZV56
zwCBndDagxxuMQheUOyNJ0sOVmJJSTdlGEe70wuYRRZzSfnRpWCrRY1LfG+LNIdO
2RpQVFSiJoEXcTD0wHLMfFwjvZZCFx9E+iVQZcr7PTW8SKolX4VzW87HEtVQk5LM
rkxlxPkO5n3Y/0B7tZ+zdkKa9O/rrcTpAOhC1HQQbSUWhOD7ADJMih64sr1i5dYY
H/I4f9YH0UMihBGOA8+aByeUhAxOtfTNVvQBFX+9UeF6ZK+zCjQ3dohJyZWj7bjW
zLhAoP1lS/nrGHsFxsADUiy0w9BVuGY3jJgtnE+raAApHQIcUr8gWfwrqZVFvsOf
izbF4ltpPCUEWkShTzcmir1jKa7vK5eU5gSYMH/7hz2tQWyClKSTwDsrjFQbQBmh
VlFE7bSikzpSQCOX/0nfq7z2vexUPcHCIPbNQLclx4qP9rEYrzKUHmZIPKTBwpiF
ywysTS4oYKOMXn4jaznz4/DU+KhkHEyRj7ygBMLuvNGeRaQydigOhbrgVH4/6/Ny
BGvkXbHknErGV4I6XbsCeZm3ThjdiMKqCgj3XWAHQCAeDTKjd+gF8q/9n0N3Y7LH
YpATmgK0dVRPoDzOjWg6tqaC1KtL62ZyfT78oZ4/XJ6t9Y/SHxzp7x2iYX/p5E5T
fXZSnRyi74VfUSyCI0LnvJq145l6ammSravqzKuC1PG78qxi45NDFicIHm60IBJU
SNOT1fwTxM+8TUnXSCpvQdwVY3ohOIluuojWNjTP0LlY5uKJuZfuZW+HI4GRFM3U
c+qoD0CMCIr5QviYsDBqjzyCli9MSmdXCvsgaNWt0gGy9I/VVSJRa5gegMpw2gri
g2j2VSPsZco457m+KUXeKs35PIRL9+ElTOVPMJjyJ9mI91/MoRaQJEGIHoZn2FQR
0H0wCEXu0sJqdnQxQlULX+YC7K6YZiy7Y6HNf+8Sk+H0S8NeQv8HlOOCAeYQYBek
qHQbp9/o/keOKYDUmRZlW9nyxC68YEQTdNB7Nvh/bZO7y6PslLzUZrLWPl7HE2tk
0NPsUt89lZtpdCoqf6Q3TXG/fNPAEHI+BBnkGqgv13ZkIlLAM2vFTzIAYV5GplBB
EIJdvkpycgWhBHFTo55N8fW6nn0ZrvgIOCHzy9PPUipZ+01j924dUrgBmIFZxM4q
8fwkDxpVt0OVSv93PdJGr1tuEfE5tojihjdqBJcWo6mH+DFZeJpyrtQevLvHbtDt
02AdGXIz9dNLK1HgB00/Xz9O49q5ip1RFUGiVAdwXla+TH4ApxeZwtndSzADRtia
/2fXQKxUanURNK4b0mdmlONdHXU2ZkGaEHZ1tuvzJhdf2oyIyoLufDD2uxzTm2/U
Yi8q6aGy/8mlyPw0D+uMmkseSKoFGGHQQOaV8qb6tWWmx9RKFHJAw8i8zrb/oPXK
3g3/Jzvw4qjJlZfntqfgKbZODjxobY8CzMWaaeeZjY5V88VHjm/3hMN1lbYl+QcY
7Dj1n4RzGexShiIHsCPCoWeVVK9OAgP9oxKdcZQ5udD1zyumaElZYavUa7uxVfZR
l6RCm+qWyThtdxfG/Gnx+SfW3C/NXUEd8GufzDJJzoXrj1HClgELTktRya/kwwCO
nxkM9I0vo54Te2bOB07iCDNCAoBWib9NRvDjXKqAQ/AnTALJpaaUNZ8+pQU+R69B
PFSkQQsPhF9uoKLcCv4trRFW2P0z8jCixXHsCFmgNeylJb0ay6ts6rHf+SJ/HPR2
YB4CsSxgOaBXuc1Rek0zIV5/e6dlJPqU3/kTfemyoNVGnaIqkWsrcQnfhhwaq8V8
cSgLugvdaUUzd2/EaANWMv0zCg7CAi5gM/rNuoqmlzbKQOl/DdEa9FiByactTFyB
b2OJT6j3VyMrOGjDlcdtvxZ+hJLBrDkAA8ZazFeSjaUlksrg/nu2xHqdWyPH683K
/4HIPTD5d6+Oomcyz5sB1HgE+iyJ1LcbL/qtUHm8s95appwn/SBlmgnWK72z9kwA
bA3/quFMGHL7+H53YOW0DBiCSjJgESVE1n4oB8ATohQwTKPWSS9C76k2Q6izw97I
XAEbXKtJ/J5VUB/2SjAzZfNWzs1NWLTPglX5Wg0CEe75RRAlNpa/tmRObW9qCJ1t
dpoh42MSdhdWQitJPnDSjjMm1YT8AngATASLi3kk84ADugdjKx8kZaVP1l9R4oQo
fJVlRPrw9e+iwIJTYjWkqjOWIdE8ELakdvzzs2LiAXVHePMEBJvm3zcj0Q/8MBk0
VNn3+MEyCGSKh2IKZfJg5g==
`pragma protect end_protected
