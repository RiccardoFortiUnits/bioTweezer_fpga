`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sn+6ThuCzuC3A5y7+og6wva2+CkWPIqZSbQRVdHidTkqvkrVq8fjfzGeWumfG7pe
8vLBuGGODk0e04gFsuU3yIYX0wrTWHm9QcIQwoQqjCMpSGpeMJATF+f2O4Ax2J7u
ByugMOPnwKrx4yxKYQEy4jIWocPjq09QOQ9Ljsrf9NU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22368)
oqAqO50BTswNjNTl533uCaexp3F53R4XVrTWFHV/0tMon8hzxPXFYbpc4GwDQXuu
9G51MbSjnT4OkNFHZou7QOZFoTK938gqHdv4iHNbPvwpTMIPrqvrXewx4490j5FG
m9bkzI1+d+kvX0PFY1kSEP61pRlJwkxWYShSRZYacNtblARY5dOWzVWp5Cv/xrIE
LFtnk7HjQKe9qrpJC4yn1AVvCxs8mRYpQiZzntBIhsukIK/+/5Gj1zOrACK7bpBo
J23D0eskCR313Vudu3KdObBlypMjms8mVT9TDOIcRdqp76JoRvHOXeHh1aBBFOn3
lDdiZJugtFqb34ytva/No9niUDA+eI7gxt2/j/7gPMzwLHTRoTNQ+gywfQ4zqxs1
3rNBGdNuIYjG9mta/KSX7RGsAHvF9YhV0MK4Au5UQ0EKZZdJFQQ2kX9XbIiCopO0
veIetNgsnJu0Fa7pE1GwyiFweOn1Z+Jt95IWVCPjlwvkHkxTe/Wwh0ML3Bie6N8y
wWoYEOhgCyTA+RMhxWGIrjZm6TSu8LaPh/etMdMUUzwYzjpX8ZUZUReKfVvKeUli
+Pleiaks2eCzg1SZ6IR2Z559z1xHqifivy9yzrMvYHGF1wIET80sqQaSTHYZI4Fx
74X5/rs9A4F5uJmspuipkr52eBIzaMpieSlyjMUQ369RTeBO41KzfxaoS7s4Vpxy
6+cp6e0+hhVpzL0njHiy6+fbejyq90704bfvmrn3TLHr547a/BeBCDSVD50CzLOn
Lwfigg0d6/YkCG/A1b1Zg4JU6fpDUVPMLYViA1U3Ppow4MQHuy6MozDKkrlBC+6y
SadBe0O+frhoWH12kj2nxUgZj7iIgAT6SGEfEbC/jcW16AkdsDOcpxSodC8E6eM2
0AlGXWMoj90UDDNctV03a7T4u/s/zBBjltmYs5YnEBIQMaYVAobde5G9gI+e6xX8
NnCGs+NPFs0cufKIZwyXGemWZnypfeF6H/wUEh/cK8PlI//pw48kPBHQmGyvrjfu
JwgDXA9rVoENCTvL1I0eG6aZk8H1dux3qinuP4D9a/70RZASNfyfIH0Urg1kHLA2
BSmcP9DsdPZ0WJB+BPTQzAEK23stF3RMsow9tmhmXAGBxXU3dVB1IEUzPWSuubID
1MdeUvdrgAqymLzHhQBMAAcsWmDLqBNJtTem+x/+AYb8Lf+qoGp6iHO00ogqL6pf
8Z5a2UYmVuZ2ytDRVPkzEpWqg3ZpYVUqar75drLcNcWXPAWPf7lRYLJ7hCFSruKd
dCKsAhix/du5jzP8mqETtH90AabPsjbNmRKcF5OC2qZRgNK8L0tQtRvMJBRCwv4y
XE2lrcYSVgJGDGqgtpY7V4FmFXleCm9D7Y/L0I59Cx1nmAI9MPNHzavCCc+H3JFX
zItdrZVy+SVupAQaSE2ksWALKC+0t4Iptrrfrl9kuMT6fOccKRsiEq6Eu5wTbyZF
BOyuA22O7wYurGbx8+zDB7hvjdBoXa91EaL2Tr7pPk/DAQPVLuSRlcTHLcUvqfKw
p/QjhoeGpRfZ9n40LUOdA+BzYL4odhf7fAHvCV0hELYI/4oJ8bIVr97rF2s7Svp9
nOBN+Wq9JhRcyq48YPuvKZJOv1yrq9GvmAKSlNBwDEGXIuZ15wjNJG0UsgNyanfi
k1f7zbSEhfqnSMeGics3+iLXcyk7x/5Ej+emcAw7kdkLs6FAvKTW+EAZP9dCHuId
Ulz62oDxjLUyaWZ/3Pk9rEaEWdiwTSIHBG9/aia/78XIuPFeszfxxBfJp7g1ICPK
vYoDmalMR/rJ3impiYGLxBjkZEVD74aTECJSBq5WFsANNg6068pq/5cxP1bh7tr6
GjmZQquMGDGXj6v5OhMiDa7U0mpw1EbGs+6Bd9Ggzh0+UoMp2beHT2cprFLR+Ppq
wG+Ebrg39rMLq9DDX/nLI+buqvwNPRDDyHwwKH5LFyfCXZj/0AI7wmduZ+t6yqSb
DIAA7Fk9dmycdcHsDKs4LNdyCRxaMhjBRjPSX1iBJUmmXSiLffc3CliGoYhYAY8F
TZXQAJuKzkdWgt/8VDIMGbtGBkk2WLryGJedbozm7mOSz8JK5TvxK1WlZE2+OKGm
zZOIh2D8fkkC6OBHeySL5WmKCGNYvnv5YmVh3IKLVvutSfbZ+MM1xhAOmEFUaoOE
OiBER7twn5UwNLS2RnER2FZdD2eaIWLrEmdpaRUcS8jESkI0kvztjovscjJrmSu8
LFLWXnSC/+Qs0pivh9ggotvbCCE2FETZIabKtRTZTwAziQDEl/wrVatX/rHSPTkv
BJgYqpztR6Win29yFrCvTbkxX4QSdsDI5hBDv1B9Gec7kmdmAYzc9uLEAzmR7IoN
Zh8vu9sgHldPjMtPr7ntVMrfnT2iq0dhe2yMRbaXGHskVbQ1EBpPfAKIrm37Q80B
FqyxaF8RNcXGLIZnaQ0ENgprO0uAX6SKqScZHkZMHCJ1xurFVSt2jpLPfsvOI0lQ
RPyeRCKbqJWrU6cxD7C/SEkSFCo3CcNLEON1n0aQl+Qz1zLrqDgvHaQOYG22sVNC
HdOYPZzsGydp5dHFO2/GCDbASnKT3v8Hr1qbbTjPZ9GGzoe2YmXAj5hUKi5an1xB
+IU93E81naPxLJIQW5N4mWUzyiKOWDHFxkSpV3kZnRZTIq+rkLRdYCvBW4wlVu7F
MAw2h0MnUNxgmeRARUf7M3IPOjZo+SC9wgWQ5S1h/6bbGlxQFke23tuLyKG5Dg2O
HX9uen0cFnfm7W5syFYfbPe1JnBC5b4gQLQK6oFyZakewPXkh7IsritMGHNIFwRG
tUq2u52s+ZYGf/gydNDyESnEYqBZvSXfdHQULyA4qKNhZZ2BhZt9Um0kn4GJcR7W
msaJUKTZtrj89ohgH/yRyxpGU4WOz2C4xjwwed7h5/u/ckLZwiY2m8xOQ5NRwXCK
mabghtlIn/FFJgMnS8MlwYz52ODg8dQbBXisoJKjBVQ2iobv8YUCif5ox6L9l1KO
5UeiU+hxQ7PjtY1BruYZ7nMFgjcI0sDa56e0WmL68LU9C1cUaxux4TgYcby1Aw/8
rEtQc0CtXoYvj2jO4oLZo6FAz4OayUlbrhBKK66grYR3pie83J6ABfp1X0ToaPWj
3pd8L0jT10vJuGQo8E/8fi8p8a3tZfk6GmwmK1cqMGMapi6Gl3w1t9/Y2st0+mws
6QdJuAeK5CmAl+Ns7NFRihKAbLsiww9n+C+ceLP3EydHI8k3tfc+YnmmMMmLtEMy
fgFUTbkQCnCD4Sxw+BZ7Apl0WN7MRiASGP7etvCQ7RWEg7CL7wJM79Ik2BT80kbJ
c4P7k/HHDlYPTU+S2+EGf7HaO8ykXh6tyO8QU5TSUOWHD3CGS9F17KdJgZfIH7RK
PF57h3Glj1pfZ5dN7BJNey9wt0TKHv2Q5Ac52AQcdFkOrCq3aj7lveYgWQDU0yU/
EahkHpWJAxYncMHwK2HW/Hfb5I3YyuBRGoE3Aqljh0e64bsVyfClNjsVzqy18TKH
m+pXFC0CCCIn+HFWsVlefsfjZ49H8jE1jp7YsWbIJcjBUZF6T9nv0P3atHICkMuK
hO2jqGw5bOUDB8l34kG8G88sPfvJWW7469GVDNeWe4vyQabm+zxeZGg5O+L4sH5W
hCnMGVNkGQeUVogTPzIWhHHnjbGjYiFyOhN66Xbh5ZM8dJ+Oc5R3BGnOLCO/6kUf
rXgHu3wF8SEVgLWTBIvV9Z+fhbb4xCCWNSk+jkFdMVrXO5LZDFNM0qw/EuccobkG
dpPcAIuMJ/U16kKYDjh8fEVPRs5btQBXSiZlcYPrF+iSxXaDdZ4Dg3M9vmuX3J/F
9eQyURv/zxQkCY+HzgIzEhpRVgD4LWCJwiAEPy4fl6Cb4R7l8xkA/b8m33Rg/ki3
baQ5anTPI69reNGvMWkcji/lMlKk5/oXw41yt5OkxvmQI44Ofc1dNuyu+f353OS4
s/GSJ4VNa3TTmHgPSdYUfRyFOPB2CF57J5HSK2uJokc+h/GMbC5eGxxb3hoVENyd
bJMOk38x6Ja5AN1PlffHJWHCOaQzdHnvEzKI1ARHY2TPeGnyHlFrThRF2JY0DT1r
104E9C80lP2emxJ1Dt4gsNIZ6TNR6QwOEwl6QQCbs9hU/XFc2AelkOrNV+vS1YUf
sFvlsNToN9Z0lpZudnGv4+LekIHfOa8wdAhu7TfTF8uBS1yuGqs8hECj5kOqX5UE
RPuBXwK7w0LiuPYxd6yEd7qae0rwc4vZAyzbnE3sH+U8iXt54ZP9tJsDaJW8mvY3
w6TRJAsDfLkKrG21QDMRHSyZhDSkYUv58pe7oBnsBoAXTDYrkUwfP49hxye5bNpv
eRDnZUbznHEp63sdqe/K84EikC3YzSmhouXs8SBALT710TVkrOjAYvWk2vIAB4zV
+J+eDnV3iVY1a2l7p3trDmvSVJawCx0CwG9sNYHXXeW2VK55GTuoP5uKRs40PCrl
sSucdyD8ep3j5JwfuZ15bSkWJX4MHLiPXobNfxN9kQJAcJwb94Rsrs2F7XgaQQkf
Vz1qevdLYfehkMZOimgBIAYpPk6alWMmZ567kmTiMdTaEnr5PrYUjeaOvi/GABJD
fWDWrvGthcv0lcTAxeOIVj7BZHVx+30SUxWY2QYywdWm9X/U3pssdnzlFwDoJRC4
I/Q1zQWNirxXXI+HzdE4n59kEvmgv1/m7lBbQwfOXhMdAJZBS10MSYgJPEslwHQO
h3z/ih9aumlvnCmqBy3BN91+BXT12cVY0NDmXy6mcrxHe9XTDDbRdr3vjLtYByCA
aGh08gAHBl1DJCQ1zrggWJ9y4124IwxZbMLZQeot7LKVtxsuSf4ebMqBm1f1q5qV
HBHu1VHnx0PQLaXa8YN2G2x1pE9ZvN/Z4VFe5pli2rru7Jya6vYmi1sB6a7LTMtJ
ZnNU91XHzguSTUsC4k365dmEm0Rj6RFzMbfcgXAfGiY0eD8DTak9rA/IGI72lN7I
2tLgpcW78bvRNZreNzp7AmpTqKf9bZL14HgOncuRDG7uMk0sC9N0WJwcMNzTibUK
I2O3hKUxNsG1kDdmNuiHW5V2Klz7lBMrMmgv4NS/BywGEvJQoZ1kSM1rkgTUgGyD
sBxqHuiPeSuz1xgfu1zmRiRmBr7uM6EjyXpbmqbapQZi7tqEADSImtxT7+q+C4By
K+N8/sOqFAmrttxIaPNk9OkbsqOcqfk2lkm0RBNkCdVsziZ1iQNUZiR7kMT3COoU
0IixOW76kK1preDxRjjODdimD1ykFI2x9VY2QQb3RGCFW4bVCBY8d3Rcjp0FkIUl
V+qtsG6l8AyGYxVNIsk6v16sBegXOKF54RldpjRP1aSj6dECWucKDscE+Xa0UfhD
khVEIBKwcHwhn2Bn0C42ErEgIYBPi0tH7zsAtgFHoEFg6BLHVQZlYMYEy8ej5ti8
EUh/Lz9TfN1EujP2jsZJHN8bmQctwKfHMwnTUGbFkYmxyqCjz6m7bsM/ZRw+1Ywl
yOTTypIvCnMGYLDCYzzYCXO24YkoJWD4rnblPZzmPcW1ieK2XqrDPxaPM/GZj+OX
tiuZhO9gJ2DW6SJvB6bOQA1WQbth//TO7xTYpQYvxlAWPo2gozIEwLohmIRCVuId
6ISMppYFumLBw2oeG58SKbLTnWIPrs6I8r3qVAA9mf/A1mIS2H+hso5MfMavdsQ/
GiY23bZWd0AMVxxRKdnx/5tTDj8Z3679mnBUZRYpFKIk3ZUqXQb7AJXxWdVLMCI/
azBUSTaKW47+v8aYqSHw4cv89JL2CftxVCwZMF1GxtOAWoZ+1Qh/7GK9fjPTiGFx
AsDLwyJof48cWCh7grJ5tIABOQ6kWojXnAwgujT2mzZKCjZaQhhfdz/CejvnCpIp
nHBfIa70cCoKr+4kzAoNFgFy9YKN8Fcmn1OACTf07cIbGmV8v48yZJ24e54baL7w
MsredYU4EhgLAUZAfWeQZ8x5MV47Icmxpz9hb1GMMiRhixXesjEQae39c/vrA0pg
bo/Q08PJj+BeNgfIf/DPjmmON+P9ZjTnAO+bz0+OeEbiTzhEUhMJLqqMX90idg4e
BA/tAq2zrGwRAlDOlfudVQqn27jMGZ2Nv1qAAh5VT67hWA7G8+oC5M8Q+pTNSg+N
0kqE8JE26cITzuDTb7mzzGZa8HWdqouJqT+TMI6Ty6OgNLvc1J9OEoH5y+i6F7Zt
UnxckbNSE1sgkDpSl33O6ShgkWNMG7luly9x0SE/YMH59QghFm/vpDLty0V3jIfz
Md0hLgvdlxYVfRRZ93UkYriIQkktB7Xx+RAoZSA9hVeAYDaJVIJI6Y9XfRr3Nrs+
BoODPatRo2TJQHkblKkQqbhhmyYSdaLdJlzrAkYrGZ0+D04IQH4Mh0g3aAiN12xU
dLPq0kHsyneK5TAE3I9v7YlrWyF/1neLLWiD55nLseqw27p1Rx3/fST/9CN688x/
00/eHSwX9X+5e3uhR8q6yLiS7bHlZFQL4vHZ/NyKKfkHh7D7xSGpiBboinMdBm1u
E7Y0oAQCDpEHoL+Oz+geEmMLYOynQWnzZDW2qma++Y1IjEEhABNyPWQ4a3lJOd6d
w/SD+qqti45J9YXmta1oMtklxag7BuQRTQGW0jiMWc9ccB3/gNp6hIqSyONVL1ua
E8tV4WZrAOD2uNe1RgC5ACD7K/M+bOJhcBJiCsSX7hxjr9pIoHho10za0oZVMTR/
kh/KjqaLKuDuJvartUVVX84g+OvWziqGF7wkAXIDuIWiCq5rYXOWO1D2CgziLmHl
11ORt8wv6qykS1XsegXqzMJ2cPs/LEi7KL7G23QpZFXkhbmpRidavTNYy/TF1J9G
ytZY5+3ZRWQ8ALn5Z+6JGXbiQJbfmA+SU9mcXI+F83+a37kMhYTbV6PdgDZPtXyt
63u2LnjwvB/paeJ5bkDH5bfCYbixSPvShhUN2ncl5d4UzqxBKCgNBagCu2ZuN9ZM
l6UDWpXuzmXFS1SpRlt8avcxs7iebN754gCYS09EEXgK21/ALu0QM+pQs0zewJAD
V56WFg2hyNBNn1xx+wTwlKSdD9HqUNVT5QC5F5i6DI/x0l40kbWN6jVW2wOTr5Fd
/H0DOBn4co++ufhhpZHMUYImc1FZRWzpkEgbTX23mvstpRAKOReo1lk1h+IvjM5+
eR9cxfMBBWd8W2jGTTHO5QPmhWouysZhbArw66GXI34IEpTxuILWzYdUVOyYbWiG
tHo1hzYqij9v5dRcPTD1zBTb0O+Ltyf55xCXtCtkl9H3y+cyRXDd7hDukaYpRPTZ
ZNKLLVv6WpA4c4XiK9gWt7d1FFCoRHzSRsOK96GZRROtjZeAE4rSw7APy0Cmbt10
HYmm0LUtp/AsR0oeaPeSJwKG+/AGEPK6wKDGReO79N75P63kzhDwJWMurkA2laTX
zcQa9/7+2rfNlpTbfAVcJkGuol0YtsAvq067I26L87hvQ/FVLcLDRH9fEleuX1uf
uU8Cu5ZdzQ6E4QWtdUs4jW60UpuOLB/7A4v1ET43Q3Sk6Wae8I7kNFUU+PkrahaR
YaaA7p/5Z/yRNzekocyl+HVh2fvavmLKnXsWCrLilfw2wtNS+D6zZ7KMPUKe2QBa
tx4uwK+9BazsCx/W6uhxbVzOh75XNqPS55RIJMtdktEI+3eo6VhKCeYpiH2SB4Q7
1o7HUQoi9lAxdoKxdFCO23vFL8MSBXfnSCiJvhYCroIAxdw9Hg4++luOqlq1X2wH
nL2H/v5XNfPK9Xj2Bi0AOSt2BfRyUm0pQgRZ+CPvj1BcngHEyz+jZBZvKuXJn21I
3Ubm4AfhzUQB4kQvNrkmgZ7RRn6gqF+muYWX1HCBt0kIC3ZnZeHzLLezDEPK9Hye
0ELrCENELa4NY0d2bRLdQp/Udf4t2IP7YBAxtjgooSCivU84dgWD0/q9NLJgr2A3
Q559pJRCbiJodWSZg5URTv4hO3J5Fk9ISuGsKuotgMgviB/OMBsclf+pewvqp3ja
FvfkSqI4lKu8xAdVWkjQirZb94VMXMqRTZrtw5t16+jJJ83AyPGEHKvQy5XBZnZu
3RxZkTXYMdAznY9KCsBXWkPAm4wOcSyYHGOqZEMGQEIwG3Wk/T5gYqcskeFCFuwF
z0WrTRTD9BWcGVdsEZxvXl5P0WLMQPEBjFFx86O9v9Nyi3ygd9ONtQ4eKvx6pU9m
5fdFMcsEmEZtWXWq2Ni5/v0tiHqXYkz57HNPQ5IiU9r79ei2VqRH4O5kKkp++FIH
vowBRjtF3rQltIJj5ahWIUJrMXq9vYqEN06AabqV5IGNvECbF/1R7nzXeFU1qKlD
n3NCNhCE4TylyL1g4Wf0vbNwXyFc+zgOHuauQxuz9VTPzSY1erd9YmUbCQ3jzIvU
U0NUAxdXwojPb1Ok4vAeYaFRrhUnjZ6bQuEIeu78kizB8ZNqG3P3ejNSW670wEe3
+fs34HnOsd9z0mr0Sch34VqrxZIilMHxKzWlruK8EEJCe25p5ohM+Gd31obbYfbo
343G4pNP4jUy8mD7FbnaP1BgTvTAW28l6peS5kMA+qwfsPXCT5zFgQ/z+R553xe0
q0aRC1XhwYGw3uve6Pg3iXSfBrGl5vT3zGWOWmdMKokOcjPtdPC4xPTvmCg7xtXa
eymsJ7AMtZkUsiVanPeMf6RynxNrQdy6QgUmcUkMmT+ugipbdCttP9mJ/t9sUnsX
vpk7TnsgAACPXg9XxK+teTSryBwwQA1OZW97xchfVGuspVEwKPXmkGDKIGuGsJ+l
9o+RUo8EzM8E6MNuR/GTIxuhgChB6mcb5cXUetuWhwsGrzH3eqOjVidTjfv8SP0z
hJnP8eeZYVIcSPCVDklmuo7RS4BIJN1koeTAuJpvVKiMsyF5vjCAy48+k7NKpGEk
EmBND1KCk6t0ikSahT3DOcJvo1vXvzd7XSkgshGanSFg2MqANN5wATY/oatBZady
CRDv49OoP4oqIxkp5hKdpKjyGo6TOWMBZfMJ9A7oSxhsE7jSc2BeFTKUwf9yO7mH
QGgr2fOHBG8yRoQVpsFevioY9D+0A6OP27uwyD/3p3Cg1nj5PMd55E6tmuoYNomD
Dy8vU7/4nssDEszKvPK8cyzgFWdMOqfN00FblB8ZyrjfdkTBAtqdDSY0DAUjQU8A
2hNxLDh8xwjT8U/3hgKu/E+vDVrJxBWqg/OoT0zsq4BaOVmdyaH2jc85nhdmwR5r
8Gad7HSsSYP9KDDfFpMz/EebmMF9gdfq73ENGi/Ii6pS0HVBjIB66c/ucPniVlH0
8o5079zzQOXYi+qT7ymK5KFZER/e53mlqjDyf6ji8ZXtD8FONV9F1dIiJG6KSVXw
f+R/ttb9XGcRLhj6zvHRWC9NxvjP/ljz0mYTaaulZcnH8IpRAr9W/oQSHvermsmI
Zj6t6k9E7n9Q6VXKwJNaSkwMT0b4UpTJfp4h4FXBm0LFbPwFaXZenDBd6OR1sXL7
m8aRmFqqYDDZSVjcN2YxvgAjpOTTYo8MV4+wR5thZ38ZkhUF94wbI8ACrNxqCHtJ
sBUIJ9gbhnlx5+zRI8vC/K/MM+58haXbMtkQ6cDJxMTVVQF4S1yxwjALlL6LnksK
ISRiT7ijVAfgaFivscg65BoC6AD5NKfx9H1+w56qi2cw9Jp7DUKElldiNVdJ8SXI
OtRW4DC/EnFx6yAJxZFmhurkgUFJpOehRsWhkN2y1j3rR1k0T+pGMJtb5HAiywWN
5aXsFBvXwj7sJfs4Z8xyyYrVLJE1PkW55UblqvIvNUIhfKZUlmMtzUlBnjS0mGEv
3N/Xc7JaRtWqDkJJkR5e/WyL4aK9WUinfRuZuff5UtxHSMAdyhcARg2TZFOgaJHc
PyLCmtCQWPMCuFcUClE9RxItIwCvPaRQX/5F9a5R4vYo51gfngN/QbBiizhyaCaF
KWMP+hcPAMIZYJt7WP/3TZbkWdlsJtYEigiZGlbMvYv8Ga8gt31x8Q6t3FMdkbjq
QS/3tn16NI1AZdlsGn7PoxzVX6kxws9hgdbexlESUhBWqfFtLz1TpdigLJannxGq
p1sfiBiNo+s2lTtDNG9IgIwLlPasQq/gBHvNjwDnAZoJhQyIlOWdCup9Q4808IeA
iPzcPGI2XuUgGu/3pz53xuPmrIrkyILhMJhNTvZdiMHPuENONk2B235JMkNueQlp
pU221hPSlY59P8DqyLYR4yK0QEPDOQGPJXqKXTUHZkD+0FXSyNhv1ODEjK5EWOa7
9eNrdrSVwBwGzG5QsMV4dO9eM2q92Oajw/i686B1/theXzBxjP+4MyYJ70K1KR+7
lD3jjKHQLhtV3exX31zugxpNp3TF3jVug0aHf4ggpcg5H3cxpJGB6TdYsSyEQ5/+
wEx/vBjly0/NVuLdsHPCqfR9B8N3C26oe/J59LsYomXvG9x1CBq6WCDSFRdoxIXq
InMnaqPHliVzF/YicGIBMgCHJ2YTpYqvO/y1uz6Vp70+F4S8PzGyhBlGW5cxWc+e
als3L2zUuSG9pFcwUNrCO1Md/nHO5Zi/htfNr7bCzzuj8ttvUla1MsMPd15ql0M3
F4rZiY2xlqhAWwIKcXIJUhWxJ7kw6KJWFwUVorzu78RdE5N+HINRlgnYoU+LT7hH
Dj6WYr29SMLEjDzV526c99WFUSfhADrh59+jW5p8F2+Dp7zU9Lavl/41wfQsuECL
6A0S9qsVCxlH/BuobTJXKQooFZ16QqPIosacUMqTES1KFDPDRePufFV4efwikLUm
tgtMiMWhDurCQoU1M3lJY9ng9+o4uyf5u9aIFxPltE4G761wavIDtuyEL9WWKTl3
VmHM588RJ+sBafXI8LnTqetmvUYG5DD97Pcl6cVZDed0+C+JziYQjmss7w3lY17K
4zdIjfjWaQm89LpIr6J55L62wTMjcj8CcXul1U69aINe6SHQxXbHw4rxzBTiBgWA
rBsX61n5iQkaLQdNrEzDJT8IrTqHyI3MSa92beDdS10WYdFhoBQjcwR7mzgFFKZH
5cXxmP9jY/GXV5H0dRzkis1iofeb8PcEAktdU8aOoK46qsMDz3SlbN5+9zXmyHTI
MtqTWy/yQa45TOMNPb9C/tG2DRAQDzzDZwKo2WdTSXhJI4rz8rD8CQRyStBjulvx
gurNWWZYBttN3bSkI5dahpMQAWrH0l/qK/+0JyBQhch+aWxG0yZQGR6FcacIbCHf
ENvqPlN/jPmsOOd79HcxzGZ0QJMA3cZcMNoiGqKplh3fE6uLE1JS6rH3wvN61giX
WunJmeRKvTfJkgy6mFkMgX3XRz4HzJjA1/smBJlkCNjrmXhOHWrdIPuULTz1joqy
ybMRddvDkbwFsPfqx+7pqVNoUpdNhJ3nmeaP3vEA3AwLUgX+AWs01W8FjfISx6wc
UrFxdWic/fskMEOCLTtYyqxPIJJPGVVNf6Z8yX3bL/1pLSu9epXDzcst7pVEYOLp
v9MjgqkWKnHcZxtBNN91MdAizFDgGvKm4R9NLaAzXKp7tRud42qv+/Y7//WDwaEw
a0lKxdGnKYhtAyYVy0k4iysBBIi3YfYgXX0zdOOgbIK3QR66OE8uj12yRqGXg90X
yD1G3wMA4czTxKjnxQ/21bpOBU8SqYcp4Zl3+KqRuBgKR288oVpQMwHyDiAaV71S
7xx0lFyp4pAdGihbXYaWiKzfIayXmllbiSp3VHMculI5kH2hKGRP/Q7gzHppU+bx
bkR+s81i2qcmLwctElnQ6EuiHks7aKWkwEW72ly7Q+lkfBL/nXmQL1+Dl3xABCcY
EgTY+XYRDTJrW7SrUW5jEa3uI4XtBE5Y1VsBzKAKOd0d2k94sL2yhmx+IMX6s8vL
IcyrKXxH8eYXHsuXP8eIn+ad8NM3NC7+1PqHX3nx0vBwsFQL4m2BJRTQfi8RV8av
4kJvVPWLsgingInoAidqqmszG9O45TGiCqrb8tJxf6yF/cX5YklPc2pI8c0WGHyr
yV6KL3x81lC/8bw/As03rNdo44C5E1C0osnsz3PH+dXMDc8VkYlt/r7R9dGrA4lJ
lo9arsqCHgrAHYUxF/LSz8CoQx19662nq+RPBjiZfanPEQPNIwv/hnpikxoLUzOM
RV12DJwP4F1krPSGWPgZb8r/iortn8BqRXsTRQ8gSwxW4g6eSWUM+02jb1XW8XKE
iSX7qe5D6VoEJepmO3JVT/KjzHsJa6oj7/Ra2cyrP0HtvAsw0hAvFYPI7yzJYIXm
BxM4Xv4UNXKYB7HMSWGzPSq9CFue7dnQOaKdlZu5p8S43VOSuISaUzX2LIsboSt5
A+8YzLWXJiHCSuclocC0HFRCrphWSbC7QGny4+2ztHRdl1jwLFyx/DZiweA4/Peq
gXtoaEmcRw5ja+PfnHH3CLAnDWE/sv4jGei/q43e7u8HUZWmA39ujDb/q8YZy8HH
pNOSc68j4VrQUUkIj9qnOFx6kxYaWaZen6MH6gCo/G3v5k15KlWI10B0qpFT02Ze
c6F5mn0SlPAPsK/2cuaXEIB5DzRwk98ecDW7rppSZgn5HtPuhENvojtL/pbIS4ky
up7s5DdEJf+7Nl9U6rV7Z+PLVLof0jl0iGdO0Rjj2e1OzeCq6j4lYpAa9LNIFdV0
oaptedz1F3njkJv9lFHE4aR5sSRoMeKDI+XO43m8+tt4IncySSLItsVP8SqJOMX+
xOAdDd1S4/rczbUg4iYzgK9/n7fZzsnZQHhmBVWPDsI52uno2Qf1uhajO99Tn+BO
PVPim4lR7RqQPn/Rrmu75qk8cOBmGkle6tX/BjOV4PhcNMXZs0FSJ6pzCmeS/hkC
DMD+fWuKDBh9UY/cKTaYywfNORElhSmCMypa8z82XU2netngcRhswW96gIwEJMSv
bIDNsdt8KKoykSKdWJWjdhWbZg2ufjKsBflWayYoj/o8mIlIPEVA6chWYZ87bp/L
e0D3JP0ifnATpACQYloOuBe+uUHol5Qc8+j0O+M6nlIiFQBJY0z8cKxWvAfRWli5
j2U3pUgXWlpHMo4sC17UIV1xCC3RJoTag2s4XXttn0lDH7Fcu0KG90niOgHLLTYc
AIIbX4A0KU9OtkQ8l02uXPVLHJrjahp88Mm0uDLqGy/ZQQHUO62CgaTYZKW34rVq
yhnO7xECzFuxSUAHMx7AmsK9to8jKlx1GUO5rym8mWHdmehmCIT0AnQJwNvpV/WG
/VhsNrfc6UEu4WYsvaDiQOase/eWb68p8ypfQHeUTmYyi0Q00brxN7AI8zJ2fmHL
ENFP04dSQewOniqtS4bIpdKzJQ6ktAmi7077gmx7uJKkDs1a1xotV2Xjcfovg4c0
3V4gz6XU/9d9wr6kdSoVdmpqWlEN55xEvin4jJmxSQbTzLYRul30qPyZZ6dm/WdB
AsY1BD8igw6VcCSWW6USrti+42ow6IqhWeTv/PtzKHB6YR1Ex+xhHf1oESVusP1O
GcWm3sL/9woZxAKIPylNJ1i5hi3i6KAl8OIleLNOijzgJXUu4ycApjSt/W3FddPQ
8bclNtsrttC5vWdrgn1TKMFknri7RCpEtSqAjLz+4v++cPI/bHE5Ip7AcgexD1YE
w6vgdBoZUllcu7OQydGbdv8SJJriQWavMXZvWT5KpDGJzd5tAqYf6I24iV6/DPai
7xzyhMABexIMGKQGKQWiBkCA4HUr/+0vlzuVPMlydw0yiQz41ENht+Jee5WqElTX
B3rCzkHO+Ax5Ha/UIoMJ29WVRLQeca84fRyV3OBxZclKZNO6H/V17egz39zniV5B
E+bUCqzBEsM5N3OU+UxY+yZ6lnm1vIulFdSANxM6H9XC8AyFfxtloUJ4Ejahpjv3
AojH1Jjs6L422LNsAYcpwsO/BsJ1lZ7L0gjmtj8rGKmyFL5WVAjoQBFJfe70ohHu
5v5AU1Lcwk3Jq+WWu5cQdHGjcNyEfm5fvPOlmhRo0ycz0lzMA/K4h2m+9SU388OD
OMtlQyyhDcZZE6Jx7KeuWkhXlhX+iCo41l17s8rjBkrYYyFanr/s3Zq2VyUeiXOw
laP/MztSL7PRr+Idsy6NGeITwIfsUbqS7TRayC218Yo4XBCIqH51I8f3m9P9LqYy
FBjchQ7vld3lh6sn04j6QGQ15lqVeFGrXdHNZzerPHwIcYdR2+mLh60Mvzz0AivN
yLx83rqk86IaUVkB1IsKCT30y+9CwueX5a1LwtpFlVptOxbPgHXWbCO/ZCrjOTWe
YhgynQ9LAMG0EFMnw2oYshTMDxODExXaixxKdYCi1cbINVyz10+9+XLQdgrz0uzQ
4txDdsfwGdiy6TaypWCK9VDaeG+tvCrkzNBU7DLJAV8StqNvkLB1/C4eSl+2G9Eu
fyQqKPbi9B7esXZwHa5Z7HO3GJzFcj8wJ7HYwYzVA8/+HAoz1qxFsZPwekaZWlNM
Oet9OTR4TPw7PKtjCNJI2ytKvzgdszVFe0STvXpqjcHmSWLkcKDubML4jdy+B+lG
q/DnUij/smDh3HftakjVy0plPxjg1MIhsTMIqaHxcbpFf6hVhDfGF4L71l0hmMRN
BOQlY9AqEmCXb4Sm3aYUH17nPr7L99ISqqLM8eSEAJhgbqwj3g0S2I8Ul8LH3bnO
Lk3AjNqv2m0xeagcgv4V+h+t9FTSYTWJ3PgIW8q/FU00mkW8Z6of4Ueeiw4xWC1y
V5Y/OGJY9GuAEyGLeLB4vcYmIj9ihDcvA+5F6MKESZcU2ifZxT0VhqmL2ddrvOE4
jOvvxEK4f7NZjEnmES9ufFrhRVRVAw2F9ubMUrv3qk5N/eahY5axBv7LE0KKRslm
qb19WuX/6o3I838J+cWww+pEP/ek2HRKcwyDa0eYuGUMLNMPI9P1gne6/41Eh+Tu
sFB7kA+Hqc7TYC8Ro7Mo80spbrEBdgZRGKNq8OxL2UPscTz8v3pwJ8jpaS/JkXhG
sYAWmJ4cj8RaSBhERM809UGhpzLMFUaHxvlifIMgDT3QspQ/hH1I+yYVWl4zR3ZU
M+2UZaw0F2aG30uSyzihYO9OreRlGlC73JRn1KGfp706RtnN5YgGFkV2qcEFbxgk
k32sT9QqhlAN/aJzqdtTVckl26vxtQ/ciQVweO3M6Y1GFj2lZWB82T1B2dWoTi78
7BMcst3MDRHrnqTaq4V8ZaNXPUg1BHjQWK1jlk8Gaf/civbk2hla/U89FDrnzV1m
/RzzC2QDEe2YTyUpcoxDlmXOMS0D/+p98Y/mP1mot8VchBlV7sxcfFtj/a/q9Jft
3w1s0UGDmhkIdL8kYC1SeEUlJnbCWTDA5JIwOzGSyMrLqVBiB6rl29r5hl1kT95D
0il7EmHfUsy2087hhO1MUlWnpeeIiHhDj2JmnAmUq0qjCGCWGjT2AMdCGJ0WJjqL
nWI+bnW8H5+q1fDMmLDdAT97/8Lh+eOkgQcMkEeIcmlXEvgAQ9JIpjs4Qj0nBN19
IWrXD/GhzydWJr8rp5bQzM6rIb40+smw2GqtboqWDEuyLt/ePws+y5POPmyGlULQ
rzEDxWDfHBScR1gk8H23rxhsXFrEu3PaEm15xWfR6XYXcyYd6m2Rl2Zu3wpfiCXO
Mzl1ZSpQkhruzkYyJyzfY5jfQdVmAC3JMTbvxL7ET6HaLTxzN3dcfFyfB0OBmpca
pLJ64K9okqpu1rtnnTb3mvqN2+SAR6hXVs1s3bJgVOu34LkMaZ0rEPsgz/UpsqkE
N5QY57J1c1qY6ML9wzdQ2Yjmzyy6ZjKZibezdZG6ysrokSYIEw76vMaL97OlPOJr
revPDpXnzH0eOQCOXWkJ7/Syx+oDoYcJuLDwTru1m4gdbm8K4w896TPEyrEuNcPe
wHdYH9sMKvfNPvVoG9sxiExtcSbNaNNvb2kAQ5yxBK31+2NDsN9MyGrOlyIim8tX
ZdM9t2w1xT1DTSyNG6vtzkqrz2D7GsyR3de071mZgAgLuvWKLdi0lPMtM9hyuLYu
m91mql6XG1RDaVhuLnuCC2okIrod8GkAemHngMpycN7PzrbUjKJLOj9xAh0TaUSV
nvU+szVXV6s01BaP5Fr/XNKLyzOjPFVJJpoAH0z7f7/41i0CDyDrHe7NVxZDcwZK
bEa21jzA6wLzYXPIKpBnZbGawXZWaqNobR4ut7tFuMd9XzVOORBK814mO20xGRFQ
VawYhhFHrZ/qBRbKTvz40p3oJ8ilLvFbHA04DhRKhoRd6EnwTQxlPCGIJLrqr9jp
Cmie2ilVT2NRwo0wH7QFRtLh8yoqNxoV5BWLG6zrsXUbOVI7/Jq9xhd6Kxkc68gu
7VVc4tuu8A/8ri+3qqxbBPtJuJp9DGpD5jd8m2mA2UI97hsSN/uE5M338O9ZIzgI
rZbYACAR/HiDC6fa/dlvCyLYDbQnP9JyAewA/QeP9V5TRexLB/zF01JNyh96BFx1
D3UUq4q5+ByZ9Luc61A9rSwa2sC1X1XhdfS6utk/ThAeq3xzW0Vq8gNfTLGDELi5
gMy/J2bb87k738UmhsIw4NOBc0oV6uOjhgcu3oXePb0d75n3viR5M3YTJ194fpzw
0f9oTTkAkez3pRJPs3abdLRWgd0zSAfxSkCS5jvSX4wtHVHgVSSAOe0Ekux8UmWY
60CJfmU1yGGHuDywG+YB1qDZX7iA1nbioI40gtK92tXFFdBl+qc9IC44VjtnswB9
3J/6UBGFWG/jy6b09GJwn1TTbt5LzM4lwAbxgZzu+tJ8zlWppgXF53ts2AWrLqJR
GgZ0cCnOcSUtheOsuXSiP9QG7YG/6fptSe192bq0KyG+3Qwlk11SYnbsKosrrl67
ruoRsZyC/xTuuYTaURAbyELnOFe7b6cSV/QFxDwS2QqO3+g89ENG00tnYdGS6BVn
po2CJYJDmDRYLRYrj4IRxWer/2XmfHC8Ql5CNBg7aqtoeE//QYpMSwKxr0V1GZrs
Ig7nS+YsU+3LHSNsJLFSG18CNSYMHL4Noe3IXFEPdt5/BODfBbwRgATSBa21jDIX
LqjWFr/b92TKre/F3UmrC+V+HHx2sTR7ENaqgueC6RXP/h2UGfPvd5oNJrEHRCZK
WpycLEcuLLMNdPC28HDQFmW656/Tt6o5u5o3GbB98rLUlukEE78GSUQ39l77ZLSR
juH9pkziUxUkHRAlRChmHvdC+Y67Weg6ON3D9Q+8NGmQbVDYrx6gPK3EUo19MS6u
ce9j0mIOQNe0J/vwpho/lCcczWv1tn6Fl151iqtLhP3hVAcbTHvB4igQht/YJQZX
TeEh6wg0kTsnEGlvMIj5elRoDOW82RPsC7c7R804smZrTMlJh4SpTR24EbzOEfu1
1aEBcJc46qV7HrIzHGrYh7+cCMHWPefynE3leOH3uLVYnjsonaFvQ6kbBpYpeTPO
yOXnqS2J/ibRH802pWXm8ugGFi9heDViPbNUKfju6x5xJPb8gg8GCPLnRXDqO7RN
XziI9ltWbytrPToeigwb85OP5DCCuLRtS8PJuYvnVRtJ9KuNWgyucazJBjRAyTgv
dbHI+jA/pBr7qpomDrxDqKw6I0TePvJJvnj0YYXxuwexP4dbHPDu1jwPKLEiB4ts
Yn+Z7rQln4YT3NPiJLDeFDdyQeFGzp6TDe721CZv1wDVLJ5cppHwghFxstkmqmJW
uAackOMPkd992PPT2mQTVPHroGPgjrCHjTry70fa1Wmx+wLKJO3mlpb9PPIpclk7
H3l4nKPl/aC3vJ689L1plPRBFYy6uau/0Ba2L18L0LmiNhdLMILMcTarh2q2QUvV
3euUQeFULWL68HrVoBD7ecVzQhZCDupR5ioG+SOIC/0ub22aMslSYsvRnhnU8euA
oNsxNfGqHBBOad7Fhgc6I/AVLhWzIRSnpfb0WbA4eRj5cAkPkQ10YwATfnreKrax
5jylZQBvcCwXaDXgi/MepxupzQ5Ragb+TWrFn0BBcBajift9eRt7HOctbnFQaooM
ovtKPIxN1rBvEXdqL/jfRWa+sn8QpSfj34LBXgpyN3asGn0kbjWsH7uZNQDT1nYc
WhDmsH7GsaF07YcWfVKCtnZhKjhHdTnV1oCg57IwZtwWfzxan4n9ywR7Lce5C+wf
gChlRpItTzL6BFMMuFCL+1kDsg/vAXdBK2hLchHBx8UwGTACxJznjzc1fOCR2Qne
zwLQIiG3OZa20lZvJLb6c41cf4oaJBhy7KAo/G4gyJhomupjWsV3Vj6UbwJPYDfr
q9gyYTb9Zku6D5UnP5R3OMiCa4Qx7nPqvS7UDSXDYzWz1rORKpMzjfzDh/bUxz1u
9DJck/Jb7uUT4RyuOiXtBzccgad7vef/2Vp5rhsC7SWcRQ7JHz2/2iIREtMQiYa8
kdlQ9lFrwg8ShTGAeVOhI5wXkMQzulHsGpaE0KGFvOmmIj9RpiTD4q08y459wJvt
gA7Lnj6PmYcVLqC5kk1SxnIftaZLGMkoyANxWx1iqE5Ccv6HAoR9D2gxIesXMSKF
2FyhPDR1W5g/7QxTLCz7HN+8k/f/zvds0hlId81FSArtxV/+AdatyVJFN2nDoj5f
0bbvSjEtq6IZ1N/pF22LhcI1MsHUv7R06uC/c3BMLgykOrXxdS2dIE0Vz0jxqMkf
2Ag0RgswZR3xYCsUa6UZACyjzKtJBdO4CSAjPgTzTvy8j6LlWOZuDYvUpA5sGuN/
Gshd6T1j7ke109i7q7V+/KqmYxB+9Ww5ygTTeXRXgioI8UHd0CE6gU5F9Q2vrsSH
ZCybge9J8ZR8k668mf9tU1FB0YawSXa2tMEeWYkRLQ8441dHj/Q74lUhpp1im0Kw
PbnqWA/vMO5Qo4YS6DVbLlHX/MXlrWRitLjJS/9/gnudwwgld/brmSZksKL9XAKg
xHxrLhoKbWTm1YgzowkG5ioOMt8fX2ggx1zDizEafSwBhwjd+vYuneMlmATj5PKg
TVxNd9YsK88sMYpToKwLFTJYr5omJeEPswOBNs2/Xb156mzwQ4cok1JzVzNN+s6H
ihu1M07txzqaTft8EIlNtXBDGpc5Lhc7rk6TsXbOpFV6Fmt1mAVqxp+1hbMyJ/+v
6x3dkls1bosaxEDrNq2n21LGfdYq1mXI0SRsAdU+1z9V/dPOavQuDoLKkRktGmU7
KI1ZdoFk6SHG/IMAsrxWfDpd55fJnEh52vbpZLtwfA2OtwzuqhXPcJ9ZgUlB+O9B
Iyz+uWvsoHFSLizrD9l4O9Um6RT2nSFJjP/M6bDHh2pqZbrZdAFe4PiJOjZszAUC
aIgQM8fkuqmx07osMm22Zg2SdBiAEHhpz+jPOwQHHEFNW0o7wGPLALKWCuVCqp9O
FhAiADTrE1BTzwnLAvfU34OaJwVMqwZNbC5AKdkp/2M3KJn34LIGsQUMM+ZYDe4m
s/Kt9RcWvNcCM2bCIL48f5s6nB5mDEzfdfkmyPYj/Y4ppwvSFpZW2zqyHCokwJV+
CK/iJEt6zYWoa6GOMDOt1VYtSDtk3EZbk00asjdel4a1pgL8xdbDTnNU66GQNYPc
yNHX4jjBOmV7wWulv2uGVXORJYLxTFTvUk4Bf9qTehUN2wUnThCNw2tcG9m/YnKJ
SNoUz8pheGYZs3yL1e+Dlu1kU4VcpXzX5dClIxpCbXptiJ2Y0YqyRZf1Xa5UUFiz
SCFh5RTnwJ0ULdBjwZwglXrtVU0/N7OXrEstdp1BpHoTdk/fy116NypoTh//7DYx
WUcJydqi3ZBp93CwwUegiH5V+lxZNzjmSxhX66IryOe7VXXZeoOHww4IWqzxoal0
aHzViOkQ06WJzjtvL19SVPTwefj23ky4St5P1PE0cCXbSG+t1lQ2EotYJP6d391K
dyi8ApcTzVaTFMGxXSxUKD4TeQzFJdPT3kceAdvN6Z06rTp3lAjbp5ddGx9sDeqm
8EE6dDqn+9nyNDlOHt0NDZU0j1F3Y1BtJ+EnccZSvtQncZ4UZDpisdDhnbToL6n+
Y5hdKKWDjl/rg+voRXGG5Me9DDewUUvUCwdkvNFwDzxR16ouz1u7fAj1/zSSpfZK
AjXQXzu7ZbSmVTm5DR4Irq4AMQb9dWHHt/e+JSA1KO2GIyO1ICS2j4065u7/q7D/
FSxtV98LpLZfiMjfkrcmJNn05p6eYca7nUnjKMj2s2gWSATFrpdSJKdH1mEJXFah
GMRL2btpL4qBC0DoQ1fWl5zreB9tWoF4Savu7CR9a5TJBMzeSLbXOrEgWAE7+pI1
H+7quZSQODtX/mxkrEaZGUoX+UI9gw4ADY0SVxvSVr0FgE3lQsO+BNmJ9X5GrROv
S1eKyqXa5COynZiljjDt+Y54RMFY4jRAVERs7kmitFZeQho8ObBaYW7THvOperQj
2/SW+tLK/iotirmrdn7Xk1Hm7bye8myaCRckO8jx/5V3WKzJ7+mnTekMCUdc0Bib
vj8pR1UuBfy5CqJ0Ds3Xv6t+Ach6vV0Wk+1LhLabyicFV9dhs+3CTsza0m0C7/Tr
XNrVJgZpEQ6Nkjy8N9t3kQmvPAhQD+Agd/Mr7x8rGfvwyLyw1jS+6YZINhdh0haQ
RogrH4nE62yTMZftjfLHU7hWqsr5yyXnNstq7MH9MyEQ4xqvWRFUdcX4G96sKHOQ
wW4q9NSo3OG+KgtvGsZOHQGogVUHOwqFS8rcPUUf68BngSyp5zV0Ko7cUkJeSjAp
PKFwbScR8y7FzhinMTfeRwwoCa35FpbIEZa1apfoF/bPmn0T9CuFix3kWL76OQdU
cruxp1kAL4ZlYxaVp1TsObrxps0LPfAVPoPkq2VoVToFxCalJiOezF0e2TUGvkFW
7Yaj6+qre0eUOKcjZV1mtc3KeQeRFl/RpBaddnPn48H2tuUVjiP7FC3RQ8gNhU2H
6WoE+KSHzy1n1HberK+/3yEqWEmiAMQVZzImRO2mqGWL+TRJMh+NKqXMCGT16Sr+
SIMY11MFWDd0Q3YZBgL2zA9gCK4VLeNz48e6zKHPvSGcU5yMYpCoBjJv+CNiThjz
n98GWFB8+QdqGRr2VQL+bWwKDPG7hm7jMhSORP0HfSn1UZmK3VdMMNIUEdIeyQTi
PiVX5WyeNZkiBopWcqqRdclyzwmAWlDZGg1KPZjQycnjC/MZ5+hwIaKS5MRZXV9L
wXVhiztWwHiMwvTN1HojtHIEIIxbhXHzDE49QV/ZrS2yBguvWSAaPB6wkRKMOWiA
gZJBpnJUzh2WHsn5BlhL9QklTK53d4O+KDexhpDHXCKv3qIFRM3aC6B99qT2UJ4o
S58MLVszjMHW+HCRJT8kHEbflLYNG/waFd+KcG02rYesjhB6TwXGssf+BVmIsPfv
T5/Doqqj2z9/fevYs08MpdEwFjKebPmWfUhxORFbd7DzQw762xMK4UMFkEsYb7iP
/MGkEux0v5o+oNSo3CXjRaKpb9UCDYDvG68ANocYpIHlO+E+6jhEDL03NV7Lpg2h
obDNCcqRJdBeTVkZ0LuHxppTjvDCQj+Q//P8ivPgEdc9cibauNPhyRuYGV45USKY
qcO8qPJIzw7sS/Ej4+iAyakXjOQzgl48uN1NhbOehBIub0dWBPFWxwn/QwmbhIpr
7CAeAoexZm5WcuhLdmhqkREvgZLAAl6hay2mawdZglHDSkbALD/947zhfzLguevO
7EfP7cSjcc03SfsCvI7zHYLSjMg6ZCK3TxniRpjbyS8V389qPtbooe9PImHN7yC8
TRoLHvPZ8DbbDPajNKXpfSipb0IoqtyT8G2+UpZqeO0mzWB7HBhmJqbIDyYr6NTi
Tf5uPf7Dd0ErlyPMyV8iG/7fLdkIgPhYW78+eBG+aIJpxsx9w801f6KOTEs937nd
6z9vJD/HgWuUsfNQdH6dnc2UhwLqaPcRC74o4wKt5aP/BO5uPg4S7IG248REaiVv
yJNylOUjfnEbFxl5MI+icYrqMwKtij3iyGurw8w67rGlcOZJ7U7gQ2vI6a+yzvTk
W0AZ3ecmsTvt23XzZVnPcdApUZL3yRInVKw4w9QUUwB47ZwONmZlPGGGNlq3964W
8jqwqvA3Z3MtDbC8Kzg6dUQc98O5ED7dOudtcaux1HDHvacIHZ1zLetziDOWSOh5
02hGUsksOe2HXbaO/dCrD4XzkJwjyqXjUAXcP+cOVE1q6h5Ttz8jSQQE6DBMuOOR
j9KhY8Z3/5FkneATdeyct48cLbd67/44FdCWVw4NkaGaFeFQ0hWXd0OI3S9cGIGD
PSX6qo8xnoUEwlYXqJ4as/jk8OUKVK/rxEfiuJkFm4XnTvF5rDmmTWpiJZfqoopc
Caxi50I4Ro9CrcsSREp1kStsYRz1wP+A/VtbpYRRPR+vQIggxLhZ3Orm8GUP+JdL
P/gUfd6ob1cz+SgEk05lp7WuhCt1EYF432xDkRRo1G16uZrbvI2lTAAThWTxx9eQ
+X4X1T8W3emC8wwyT6RuI87heuLp72e+kJljfM8NxKjUZlD7j2aD66hDDA3Qhxe8
60knanSGY9hzxdim4EmKPLPewhGee13NjW/EJKZRnCOAunEaNaSklHbDFBhcQSXV
cBMwB/eGb0XZBD8sXuxN6l9IKidr9O8YTM3IcZ0JxtG1R9JhPfEVO2sA9LK7Tl4Q
OVj2j0Ns+s0sU8IPQfRdKzxqySFq7pdS7ru66OcjSW+eURnQKgPLt26WzXQP40BA
RFOhgFMY2hr91nS8aZMtPX4xung1rixNXMXB030ujV80DjrcUfnUscJm5koSYDfb
f0ZrHTBUbZ7MsewIlbJisaOFQQ/Hq4vH7VkEXwXzfpiv8/SwwqjZZrHoXUScsoAK
KkBSP7lH1jDydNwBDu3nMBSq+Y3TpQEfPx1yqD/ztP4rszgADoGqElofCk6plxZM
0+UfDinwW+InX0nEw5oRAtFALbbuEg3t7qO1fPIMqxOsvB11ePCMKQgJjQjuvDZ0
mNbmoIgs2lOP1UVy+yqvsacSXPgKGd4K0ZvsgAgoLPC2GOGoou+4woCSt8PeQJsJ
i7ZU19PUAkC+RkhUw5b7nP/mFbZw+T4WXbQSF5XGRyDcw5NI/Wtq1lD6RtWmU7px
n0cYIUa3HjhbVIRKW4203gh2gdXHhY+ZrzuYWIDqzC414Y6RTg3aTNFabu0q2s5C
Y94Y7UugorvGBSKpwdjun73UfajuwwhWN6Ps267bLdqVtrq7LIQ7T//wlXFq2WHb
0nNNGCse/us1k/gG7yjtuGXls09mtj2adem1BrqFufbEl5hrt+xQs7FanICwOQBr
383yfStdF3Y91i+940B1bLDpC2xgD8PHFAkB2yoq/v9WAW+eXPNnIfppSWp/hVNy
KeQpxo2j4UkkQDIYmODaOBUhQurbqlLG2NxjeymhoU2gXaaewzaCP8rNAaA2ak20
/BSuD0jdZgXNGWydQi9yvIrkv64xd3v2MMozTrEzzRd4bAdwnKJfY5BU6eJNeF3X
DlsoZ/gJmglPF/tUlz9CGIPph7m1ijxcTqNYEY5uF0a8v3KtvIzDmpdjFZAu6PmC
VqQqtZVgy4qvZUyhaTeBjtFL1aXRYh8tN2RqWqurZRU5xtly6pkyjF8TJB1NnJto
0z2sSz4EzpfgKCVmSpYYwrI9wumElIvsdtUL42ZXMc0YXiLj5wddwZkNdg9HbNSM
TfRg8Ab28djxXMWSXMyxr5q3qIdHuc/ssFDxo1RbhY2v4QSruSOqLwkJf+GS5D/L
GOvV6//Zc/kxv0uruJLvmj2ii99aD9Vo1c+Mnvv800hwjKPLuMpFZ6zwROM1ErvM
nt5gn1lrdqK7ql9BeTxE5Tbv0eFgRis2d5c8Xzz0ZQgtPv1sPwLPLt73jsPt6qZ0
EkcNTQv+Jt88ASvptuzUQKdYUb69RYj+fW7jDckMiOY60o4FDdNFt4ROyZoOUd6R
KCqpkTydcMWqjRH7eIZOs87ybPBbugi5f4P7eV46nIAWHpa+PxqH6thmwdvOC1E4
V26Vn1dCdUoj0eNQ0+jN5mPD6UwuiAtKre/OQmJT5lsFhL2b1NwXW0dBQVR+nhf1
z2jjOgMJTB9ayz8Ej5yVqDclQXSRxUsdHFlUfQ95gUDIN3mKgD/7iwmEJRk4Gf7N
DmK2kvvw4Q2HeTg4/8kHsphFq6xxnSEbSOVjjj/XVy6Nr3ABz2WVBsmvXrvKC2nY
HHWXyyFV8wXb/MWVWhB8Z8HipnblEfdNq4WckcNoNns8IdiLESQt21W3+BzquCHJ
P5j27aP3v91qgsdHTD/F4UmaMrVSdAd/zeMQflXX0xcfxqzWMqGOeLSb7DcHBQU+
newUgKWLWUfOzLwjx9l8qxE7aKkUdK8kbH795T1lG/y9/nvCDaQeGMzfwffgQ/V2
votrIaFf55jGbngCethVECwWhrRhUUvzUh7elXxv5qvvBDLZpzWNJmxFf70qt1is
8jkRBKr3Rb/rLsZRCrQrsO/6ucSOYCznFjMo/2hDaRi7Ile5/jvVecH2dRysAL7R
RZWuwPPDND3AEb2rAhGo9nfpy3qzqSI/99W2X8Bgyykr4G9YEsJsJsWCsGAuA+Wv
RvfVMu04ZucH5fuNqR+tpmAnbi2CzeffRZCj1wzm/mppQSTkQ3um++/3jZ91c/fN
Nefia0lqAhwKc1ijXCW1YJtlBL/5mYLHzoxy2gADVL43j0CY3ZLqo8pNx6shqsKS
fuh9RJ+YNfiEJpJS1ZkKE5enNGQU6aunpvFhIaaa4Y8NYlErk5xNCC7oAJrSwui9
k+o7M5nqV/8tHlg2xuXqQzgjddqsvV8qRV6rtmaUDQ91/8Xkg7NPjJ0UJNqcWx6U
VTH/+/PNcqV/87Sle8V5omzKioiGkF/sWR0YWqQ3uTDy4bXIJzbhj3AE423auyCj
0SNLmIHX7mZplx+YVZU2ybGxiu5QmWRke90xVHnshPjktB3jQ5l3vsbOnaRMwOfr
ntgrJfYW1DCrXVoM3WfjzxwyiYKeG8BeuU9o3y/fZa3g3NdKhli0gaaYVa+2m4yk
9/+EwUq4S7VHpKodxpck9Wx4kGCdgRm0QrOewqr2Hew/BvVxtP6jpENQ+DecdLV2
hEY8gL+YfA3+vrIo7OlEnD3snVQyYjFEKvU6vnfM4X0JnnenqWlT1po4Gj9ghGqX
YbB4WDCtHfk2iea1ruTPy0w9GnlvRkjIeDdQlmoTM+BBPp5s4jqKxpwpNnnzPw3c
/G/2oG1H+0sRTjEFKCJjLt3KiUGbVa6L+f1WK97itwQDRVEud2NZ2M+DeDkS5L+F
Zal8SjheqNfRdBW2obU5qjDZByQRiq9I3BoC62FkyEfXfGtbBYSZ95IfD9zqh0Br
kiZF6UEgH9BEHzQvl3OhSeXRCC7VOGkwm4oF4jJTNKva2y+jvywu0pAJ+iG6NMbA
mevYVHReJCFGyKZS4RNNQwDt3NmSShwSfYxNNwm6V0tqypsnBdES1evMSLWKtdlz
9WV5AHETTCzCBZa15YVi4LPREma3ijKKg8HFseaQSAT0w0Kp/W9CtHpaRcJn9Vrs
5l0U+21oG29DQ/aO7gAZk8DYZJH8iKRztzbG1SsucZSm/s33QGiZS8RAYe2RPsGr
gU7p6aJSox8HrQEGE0GSY/qOG7V23xZW4ma36NgYIny3kylFtE6llehop0IrKPZy
61ELcZd8bIuMid0WlN95QYo/wljaqTwwWEij00M53rqetX3G2dqenRVasvTYa09E
KTY/z6kee/AvHINLCQrQ7H4oQk/NODQ2wES+w+l6YvqNls9AIaragrz1plhIhXvT
5byfO4wVyOr/5bhQ+GtFIW2Yy3UtH3HYjvzXJXRYNP51IwQgTTXL49Yv9n1Rv3Zo
IV6p5nljeLe5wwwlkQgKpVGBBvq7o+/XZ04Zy5yy5bIHM/q+/Yz5tvFDYvukJ84e
6Mkdm7YT/mtXQu+d59CKkhylfT/2xIEaoyI7A6cPXtCtTvvvdYfVtcjZHy6hwq12
nP42/5XmhIvUxlLFaT/hvrUhDb8jkYY4macaM/ZyIBul5Sw+JVTNe65RMQJY+87u
vuQlP8Q3Nz28UkLlIUH34ZPgurb7bMe7vXkLCjGYq9Nsf32FuDE2dlcl4tYkf6Cp
JAKUrI0eO321PXYrXVrSnSk6JSdW7siO75U7RtCFa/FzgGJmbJTVVx3qusDjehZA
J6K2e/pC6VGIQDfjWwV4CQKONoj9y6S+LGnCFzOPi9DKryuG79PDecvMaOekLaoN
qIB5hl4MuzI6xrl4P2ukPpSKa6DcNDdvtnSURAmnt6t1TZ87MiAJVIK2i+4HVgLW
Ya9TFpEJROa1Hm+/qCbt9QR9VAQ+EJw3SKeSZy8G6ZugmgYtNQEK84+/980xaOFN
4pRNleNhTRo3nCVhv/dJDodufdAMnwT4WE95ngI5yS5JkjFaIlgI6v76gxoj8yGS
J8QEO+FdUPCvUDEQQzERSTSisR5p8scWpObhxbfSzX/x/sAmzh+W/3ODRQMVv//D
mzbNnPWegO8uybPs1ySjEa+zXLnZoI3hcEHwhkwFIGSpfd8gxFBB/TsYNDzyOwxt
ysyYr9ceMX5FR0aGwln9uChRbCRPEc/0jbhNVAu6bZ6Y4LtyX3lnHcglOeEQH3yJ
zTAxQFXWX1pWHp/mPPE90UKBtHEBZ/m630+tH0Zx8NPHVuS/ffZxrMqxf9SWMVXw
tchT0GGnh3qSVCtucyf3elmW2bfRMFdqkhQ5DW1SulT1Vkj1HyxTSGMKkSDunSm2
pwlvckSiOWha7sO3kIvHfj9PTrP0LxK++BJ4U/VIXOdgWYze2FRdDKs5kJh+DLzO
tO7wA0DIKoPFe8pYJoRilG1TFrpPYCBf29bV+6b01kHm0pRu/YcnMTBlZ7I+miLH
fBR3DyZw1lrERrpnZHHa9gNm4boLzk0BEL/qVM4ng8axreU5pxzNOPu/tQpj2oFp
PZenIc1LUvrnzFbOKt472/x5QERPMFoufEFTugJUofRYEgnFzOQPqfkuC3PgIEPX
sjZMSKqG3mX0QpqBg8qatMwc9hV3ib2Oxbp4VYuLDr7yP/pGWo0SKcI+NOIwNHwF
rh9J+r24ArbeWNsKg4gJCCxSMLLxFrhJe4d7VRZU0pC7NWhwEMa99QTuFzi2D2+C
OE9/8YObtajMnzSeSkJVoZGYVX7HSFBN/mBmyoDN+pMRMgUtFrWz94CA+mA8KmGk
lskRz48sF63WHUjYROab+LM7JZ/D0mM0GQ0h+LQrxQ1L8HxbGQ6WcyPTa7OyJ4xa
BOnne+wol5zpAzG+EiepnOjORBABU/2gyPtsovwx+i4DOTJLs0cxaWTVlu+eEsno
IQbF8rlWFLaHOpwCaYcyBA9hYCKom4qEmisfXap42lUNV/i4qV6CdZa46eencu2I
cy5e6pkVzFUmuKEYg8pbiWFfxHUvGe9JgZRaRuEuyT5oVcV3cweMyYVvnQdMKgSh
uGsnMEP/zRhB+XS5IS//IpNC6xj01sIWIaibMFL7Mld+qcnmGqA4dBU//zsGGtk5
PYICplQAuMGCZ6fHKTRwfFMV/3C9PssjEnZjLFxHNbc7X0tzB49Y3zARXe0McOxP
c0MTRyVPOzXMkMYMYLeRr1+DO7syVi7j1eGcX7mcU98Ws8RL1tpMHb53Vn8JxPpk
h8KCsj083jCNslIAm+1IbSuwSCB7kq9OwJCCqxtSlXZ6gJU90XLhFsXVK46xVk22
eB+88nWl7nBH1tQ9S5TJ5VvT9SvA4L/1eOyD/uvXE8Qe6Yc7Q0KGUIag6l+WZiYj
3Kwcr9rgArVpsa3pAzW6rogzZhsxP3/ExeGnyqSrsMxWPvKfCKSOFfMT13xLVzzN
jP+DuGE0JUDvnsQsidotp9ujmE/2YPEiTAYVmz3Nmxyo8cJbNK5Lp3V8biKZFZkB
LXflQ+Ifwd06kKZCA8OagdQ540dGdiLYxTg4T9+RAeasakRc4w2s2DXbYBVb4NXY
aXeaHwHc79h6NBtO1AfpjBw6tzizkrMI6+n+djHZHo1GeGgBCsg1foVGjDvQj9ck
v6SLtqgwDAiIWOTJEtTlnHv2SoY8Q2A43ZMxIKHRs+5hXeGS6yPatIZF8u2OtLxU
xHg0zrzB7QNIyNPwpkUHviZVCMXMG3sESdjscugB4+eLzQbA19byk1/dtq7Jumpw
PzN1dMugncy/hCsL0ZS9G1M7Tmuh11ruSqfFbgIg4XzeYuWt7JblBdpwRswISZTR
PZ6eRkiYkT9vx07L7h7X4mElRy/Rk5O2Nmps4BncQ99dsUENmRgiwEhjrt7aS7Oz
wed4ImtpFvZSTXlJZH41/kXPzhCk9HeQSI5y2HqmgOYBCKtvuDBDRyrwBbCNzed0
EHaN4+0fj8DhjOEQaA/jSUARFWWr55BlZzV+r0QAGvrM1iEceOgEYCW/J2icteeR
7jwjn5JM2/8jXcTHClgds28LBYOSI+P/d+Pj+A650YR9FnggKbD+xkT75SYsXI19
8v1dnExeiPwtUEP09cEQHfHERfuqR/7xS1Ns3XHKijeUnvKDVurTOtbme+JgK8Ps
ufmligMdJbIT9KJeeEkWHELAWepIGjJ5Xe20RTQl1uBONenkPvCM4EmPPz3VB2FI
8yMYcAO7KAKCzdF9wQCo/PbcWaCRKI/eLdDWN1iqFg74/PgXWr5Iza7xscU4oGsL
AHiDawtgq41U4LFtprTkdl39lwJ2k9xySJBGDmNWvzzemljgqlPHEf4DETGLygO0
Ao1q045teM5Oqbf5MbI8Tf7h1o07Ik4rSJNZ1OGZj1zHSqRBIYL9IfIRqC/yOxFA
0n67OElqmI7N3r9WYL8OrMYvuyEnthr+zASKjrSdwmpeH647hC+8Ban54hu3jYLy
9kGfnYgjbPYyJgR3Soe+GVyTo64og84BGPWtWDoBpnIWLpr1/WZi6y0mGHhgdvp0
uRLioT1uEbjH/trYLDb4rg86XLt4H56VQQhIxIThFWfrDO5H6V97L6P6hoFwGtma
otTJvQLXZKaUUjlFvMh9Ckb3OhVrZAKVI+cAE6TqKpQlhmVinx0LIrp8+0YulxLo
mCWa1tdeq2fzbbL7HEG/bWprk68Rzyw8sEsC27bNfslMxotabJglr0/iJiKPD+lj
3a14hM20+/lwLaDOgRlOGieb0lTBtjCStID3XcV7rQVdW6PYoO7bPsgNI6XOu2iE
qKzzGPtviTN3yaHbhIOK7RSW9PRauohTlivBxSDCNgQw7MyKOnt0a6HcnQqibtkO
+nLSuBqIhrtzTCotdDiOB2Zr2RB+4AJTrtVR3hKm9e6qwhCjY3t9Mn3JN1bsl87N
lWqdmn/Ioou3EhwNtPVs2ArhGDb0MFo3hBFIUjRjX2NFuLpao96TMokDCXs0hkpi
Cu+7cYL73tfhoDCZg1TywbacNemHLVgQz9sQfWUAaDvqPplAQhmgvXcg+NWTw5Bg
W2vXE/z0LJhfZRpUH28Cki7tgmU57ff4q9+fS7c30kTN/B/ZfeHUd7LRxks//USg
gP5Ow8UnxoFZ79G6zBpRQkI6yYX//QrNMyQ+6tR9Qh5fjFqNZKAnrvPHE28sbj1O
FlYRODPP2qyn/05hE0cbF1arTikZ2JxiaDuHtUIqUdwfXeKjdbzZpXbBrm6H+XE9
rwdupq3uWfAvP7LV8rcxC/+/0HR6ydh+38Sc89dsJLxu73gDhhQAlJ+bweQFnvIV
8OovTb3c53iQREBti6BuXCt7H1fm2iRN1rIkur60xs4Wl95QWEJDihUruSeAl8Dz
sPP9RcxZ+XJf3IcJtsFRdzwrnUssSEcno73cry4pi3HMNVM4BqO66dDzxZXe3qAp
jWjeXFGANIYe1GEopX6Ajz0atiXeQheZD/oH3EcuwUoHRzJm+PIwMuXw+FvW8mBF
rJAZif65FnKUpbR6uuJmRBBjO8Tg1k0dWe9PGaIDG9zgh9qarNkEf6Sbo8zTdkhr
`pragma protect end_protected
