`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Lod99HdY5KsERxXN+dTqzI2b1+lF4mrgJI/heeKnx0X1ckkLPaXexP2cfL0trElg
TcBqilM9yHE9LvvLi26CH8XmZW7NgzjeYLhr3brd+8D5iEt2hlDTR8PdOUhvmFtQ
bALSxk9jFNuNRRFueHq6AJBnsNSQZ4FvUmUADphlKrM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5344)
fA/v36VRXX6d5iynlrgHyXAgAKpbQYYF4HCcCHNPyGz/0kxcWyy65Wh8k20ptl1P
2cWFoekuHLTfaq6wDksL5e53n/1IrG+MZp8siE9rv63qiavLFgz4OhHiQNOEM9kQ
apS3SIvZyt2rSN9xfQzlIh4LBkaB2NVGCbTX88AZ/JtvQ4E2BbgTuNjREVhb+xsd
vl5QEbizQDhGibEcJuIFtOXf24Vp+Ppn+Dx9XCXIT8VzZgHT1RAaEi5bwV2qhWwe
PzrL4NAD/2/P3FN7mijPpuuy15mopF0Z0clab0TJkJxkMjicz8gbUIv4BsZiYApX
U++RgEBXKsozxhTDnFikLreypHrfZmExEbN69NY1F608qkG3X+ekAXvL/i56CXif
13B6HEYGW6yMi6cM+ThCtAxe2xbKTR3k/XY+MTqayWZjcOMt/uQ6r7a1nyGDfTjn
gVfpTtgi3FZZIi64buB3/M9QzgGei1rLPE+ABSFkYUuahFUWMceMEWOfklKLDIJ4
p/Wv9jrrPqmD3DaaZs+/W1Bzdp0wl6Pqq80eRPwD50DlHSb7D31DZRuUcgI6sw7M
mGhsdU/kxoUFjXpYrslSfXPg3K/UkhQg5K1EgOBziU3YYp2kkUPkKOsindC5CjZ3
kJWIcqp4qXkW7P7S3JDwukUUoLe/bAz1bQdXfo4MPFCeSxGDKRJ1cLiqy6XzyIDL
v66Yc7IAtBr1ev9B4tUHFlt8PG0SAtQt6rbNkZsioE4XGDOrxy2Cb+x8y/zs3+wO
S61tlkR5V4L2CH5qpzjCOCdr24O7tj8ySYHoiebsUBEMmy6/2p9XTGthNOPqPrQU
bdxN4WFbOL6LQdNOowV1QudqivZplW12sbSv0gtCAi7qQpjIfWsvwHhuO4BwLyL+
rlBHNwPCb/aA5WpFQ0JE0SiAwkPB+Lh/njRRszR9zKc7TOnN1/1ZdtlfwuROlBQF
G/A54BNep8J+q/Nu0TNSCmUAg1935kqx97POBraNtzTup50bfVSItfg6di/RXMJz
ybwNUV8JgxiUqzQHlyLiwJnjeiYNp84Fq7XVq6upy+u33nr5IcpadywyZ5UW01XB
hwvvmqeKXmWW1MRF8psz5KtjfYpF+lT+/keYKTv0W5S4B4CSoP24lKq+AvXoW8aZ
vqk8YFGdGf48Kzqnziyc38O3TM+YXhk15bzAUMOcpEtWMebVqi+drUqz8cdlZfcw
nnOiS/NL5O+l/BnOABJe8h3K1iB4xZv15g6Rcx75LlxGfQiXPrSUWwRMnppbT9Ag
/GZZ0Cg9C68pohVFe3Knn71QbdZwtFkxoEkvshaiQHTvgHBmF8yn77NnNUxKiTgY
zlVdbVnZHEQUpEH432RcP9YWC1ehe79uPF+1zHsEH0Lht98FkB7zSo2I5rN81CUH
+3X5vpmRHmLlCcxFHSdmecTtMLh8Vo8TEI/aejUWFd06kqexENPff5G9xnIb6CtL
7dPZC0qZ49H2JF2+J4OW5ECfMLZb6GXrrCDpPUvP5S2fYPJDbrvnsjBLSkFvASjU
72pt48jMUwvQI8Ajr+Tuh3UgxJ2QmWWi5csfVC2kMFxZOkX0HTKr/T9nOh2I8jCE
nx8mX8gzp5l/TW3ZHSZAooMV9C6umXos6iMHcBga84CpBnnMxhs3IA2QD/sVjb5M
fvc9QY+i+SilFHP7GAkFZEcnEPdrm9nGlbKeMeFdwEYTioSJe/yzQHYljgV+v0F7
slqPXq46bepew9VOxaqfdFfNymJ7Q/OVkk0P1ARwL1z/CQB1bjWYT4qjSzz8IC8n
Nor8AsPI9V53N4InuVAccIDTNEOWgwSi8kHUMlAdcjGH0s0i0VlKukrI4xXSikOm
i/lJmI/cNVZjrhzwVLLBYw4mZ2b/cASEwBX1AKEACDpi/PZGLwrWP8+Ifd1DPqts
j+ofRMZ0/euqbY3fdYo4WbGB8CAUJ188dNnEsm2iQwjA8UQ1QVA/iPb/kkj8MBvu
o/vw8st/5XE3jzCjulnTq2DKBs42Cj+K+y+bIzSB8FU2dAZ5JXSMYCFnCxhkOrJ7
r9nVH4Wq6to4eKwlHkQpiC2puLWJMO4MCrRlsQE2ZFe8qJGhxUJcD0pO14gMXMce
qQQYZ6suEqc+D01b+tDWEjIY6kAzhCSFUsrNqELN5AibZl6lcwEYcf4EJh2D6zDM
4TgHjaHIQtUgN3yHqxQiUAA2ZqZGLeKdKXJ/bbOU9zDqtvcQuQFxVdsmEU/fA3VY
yj8JqJJ7aXtzrtcr/HxvF3MQzl6ud0+68hDikpWgaV/6SmBK5dqZyIKabQcg2t5q
q9d6pHgrT0Cs2UVF0SnZNsdXKtKWgRpNANV5zSkhNtkDLa9z1x+1an289FAFz7be
bKQTG+NalL0/diSAJlR9rEv09oXBIvw5Wpggcz/Mn1JOz8Q/Jx2whwwwhNs6S3H0
DR9psbqOVhP0IX0MHaPgljBJIpuRopmFFh5vhG84jSmxAW0XZpU2b4KLa/C7MMxA
EqKQ0bbh8FZEiPKldbcjZfz6sXMPG7l0DBe4RvYNO8p0nfKt0GDTPFPfNgkByYqV
hWkPQg9l6IrwcSZ3PhKRP4+y8NERM07ID2ZBV+yVWiMUVT9w/8EBdC7oeDblQ0Al
iKbWpDCF6kQDU/8bis76/80G15HFZlrszCNraPJ9ojodyUkE/kzxsWxeO2Xj2oRd
LpseOu2wSntfF+/UAu9n5QKldbkaNV1sTSKKlFHjLxrjQVmA/14ymtUfBlc9dcep
pMcYZlYe8lZo7XKD0xY5IM8rvD6zIVIzdYcLI4DIjP7io43CEksS5j/LbzwECVJ+
smjeMDcH1bUmgV5kxbZxaGHvSmTmvz0Z+WNcW2+6kLPvyB+n1W5fbHLvGoq7Y+M+
CED9xhQd3urENrAMaw/D7UnmkfJ8pWr7LFxigIpP043SRhgJOnLx5l20TkHBVGCx
vq0sf2BhdaUyw9r1xZWonH+ggAOilHP3XqSAqllMiEMfOohB0HQCz3uITrIBiRl/
cJKpdAaJb2kxu9ChKDWAfOIkCTnlbqjHTJI2vIumAxfIp0kO4T6Iu7Ma/b4IvmNh
fbun68YiVwzUUhz0rj4jDXRjwLJsLec/m9rJmoCbKFXeNgkkwBuADMI00tw6+5cd
0llIR02psue2nIdusRIjM463UcVBk15lnQC7E3H6f7ka59MemadHldnmHLmWPwZW
5sVAvNG3k4z0cCoHwFPYEkjgBw+SvI5SPD1qEWmE/yyY9hSdagBmOvtvJtnE4ZeU
xJkHuwA0GkW4rZ57ATG8l7fwNUlSZbqhD/3RS8tKFyl9TVab4pPEl6gQ/W6q7Tha
jQ0QyeHOR5VGRx6PX6tI6ZD+CWc1gnEok+EA3nFFBNEtVZCvtANtc+IKaZxI0H5Y
Ildj0rkqSPyLhOsU47sUOMRmxRdieFwtWLk3vXsVNZglR+uLIr8axQjASe0KuVqM
AgaM1PwM0F4ZtAX5E56hu11ZJP/AEv1GU0Z4V6+ZZi9HW+Ob1wP65iCWehNMmmWn
O+t8rXkyXdV48eCOz2E0dFg/g+8+b4hxwxukV77g7b1HQQsAJo5eDJ0zNA9yUHIv
IVDE+hhVc76nM85iFcbmHpMS6rhgLm1yPj6SW4k5rCAhY09DY/ZnqDPFF97sMBWo
vLMLaiIfcw935kM7iF6fWRKsKDT37bkfVKc4NmXWdcL5YSvY0Y0jWacoAGLqzjOy
JVNx6hSmQBQcmwFRhX3KJYOpRb0jViE2CpNORgd4uWnmxDz3zCG4/7Ox8z/L5emZ
Z0CRTWj4y8bJCLhsVN/daDwwKWbNeJGW6nMyNa/9xVBG18KUK7d7+EPHY9l2W7TP
VOb9t3w4vkvF72wsIA8K3O10xsEevIbup1rJGBL20WCwQLI9LgwvM2s+fGg0vF6g
vb7DD4yKVIrGyK7nlLlVI3ygCehaS0r+pestRXHBqXzrNDxtuaghauhrLaPJpYoE
gGlKEeBWlelJEg94zXlTIa0Xvaq1YZC2ptan/LjGqjaHSn1s7peUco9UVG6mcHtV
JfKW2Bt4Jydyp74qw+zlor6KyTlPpUyPjFSlf4IPiK3uzjpgfxQ1BtBXPVeXNJLS
s3pYHCqpGclzM46U5+0PnKNGTkl+3NN1VUhmVpA5jeZFQBclteRBp8brzmtg8IUX
/vIOCCV60MCHV/hd52NJNc+IFNL2gj7Zzd8s3bCBpdlzqzhu5XIGDVlL1z6dQEeN
i1id6DnccV2uYCWDmmF0xfByaTuj6hPVQs5SLJwn1ysJT0tGE8uiSbtnJYRHcZuZ
IQVyHSoF3Fiz7WGWpCMhFIf1tKM6pc25Co3DrrdPc7iz7gPnYPRABTV5i71cvfko
jn3/fgTQrc3ClZetfpjz1iIDzSA+wfcf8NnMlgEarb9OV9fp40FGGp97k5pz1ViC
EKnygHsiLrAPpsPcC3ITDO3zsrKB1Gu9LDr5x8gWJTYFImITWU4yb45S9sj0Iorw
3ftjs5IAa8SDp+G8CNYZvCLVkwFLCinCSV7XJhCiS0WPISbTaPbB4LRyLVYwOSNo
HcD2oeO/njv201xPuYjPTIoKGcjCLCZViYrYYIsg4f/ukewXhxABFR3qXnFywWJy
V+zpmMwDlF6gDyKnhq0IYzSkpRIz0Ku0U5N6nLdPw49rB7GFQxKTmJzu3srbx1r+
o+003E3JEV9IET2CXLFvaI2Ir+WkRBsaYR3olWQHNjTgKbELz3tTQf+shrL03aWk
fhz+EQkLqT/N15halpkRxBnHB+U9Wp95j6WmA8u/CAW3WdwFxFLtpgVU3AkFpPuk
XwM+ZRkU0+Ovk8rRpLXfvZAehEV8z5L7yFR1LXZJOBrNxJXuZsB41UQXF7a/e3MO
izUGy+fAOHkJ+rQyUipeJ2zie1zr6r9AUho5x0lSXCgl+4Sfw3JEUV5THEPdDQGO
Fl1amjwYLPsqqwY/1p5tnSOBgFiouL5RkDdi0SS3yu0Ow7uu14uIWiMC3lVA7rtA
G2l2sktVndYVZJ0OhSzTnJYlBZ88G7N+nMOCEHAqyBpBGm3mgOdAvd4mNHtDVKUG
rhZ4I8OUEso175Mu3y2+16x5AlnLt4MQBECCMr4hD3oyghZOWbLMzDXUZd/vAvve
EBzNfVvgll1yG+ZGnio/v7FERvD35mC3GHaJzeZqFpiytaUDwe5FzAE0TSZMqAWb
W4OynKYB4sR7lhM7PoMZQt32Gonl8847he0zZZt6KcdJmV/OvPNOLfgu7csBSqUc
hgQ0tooZRCMrB36HW7h7QrB0CztruwcNkqpU7BLjYsRcrhL+aJ4dTYx1QEzUyh/N
0iKmNMVN0CBKf/vcfK210bG7TQGnYEsiWPs8T0omqohd6D5a5QpoxfSD3mZbSa3t
BetTmk2UreWBuzo6QEYFJiRagPxKzr26gSjjcZDZg3lesg2IFE8n/8Ofc5DMLHSf
Yp/I0SVh9/XB3v632kEfeBEwC2aHNPNiGVH3aaWKX4lKIaHhDQ/ehaw8SFucnCml
VhKWdFkY3tNX4REiqd+3OYKk86v4P2RZxct34rilxHGzVJqMPJHLvi4t8NpqbUf3
+Q1Rhmhuwk5ZHyuRaYBNJj4/psagAHeYaVBt3INzjqz8XQg9K5HvtnGaSptYTIOt
mT4Nc3N7dfv+aKj3u4BYSws0+Fh2/jdMptPM3K+dZ/+8hjfNR6Ril6sVG6jfk0xk
DNdD/+wpXcRrHaKob33sraO1y9xcCmpE3mrGQMlj2CjuerE62XJZtxaBNIvvVbiw
Yr1ctaoDC8WXfv4jg2yvC/2D3XFW9yPHpAC04i76E1M1ai4pznRjbXWeKPThr4Y/
XJg3+bbAGsMav9icxzbL+VQAOtZ9ewRGiWJDjt6+pkJQO643JRB2gPPSuWPiPysZ
JUi13223c1UfAiXw054086yZDn0DaXis03gitbl9WzmDrUp53+X/t4v6AlqYx2hJ
oI6gHHJQz9ZkhaNwLAdnj5dUsUQrJ5AWV36p3+dlbw4YNq7OAuzCTBeactopLyrq
ljez/3gYmWCdn1LXuZD0L5ZtglLUZtEWmEq3RF9mxZbhfn/mPecYvXH/UzbEzEfE
ClTYL/gGxfH3yj/NEK41Z0Snl2O5bgaPde9s6IljaNaS/cAMj1yrGUsfpRj8+mhP
bB9x35HSoX94LBZqhpGY2DOS+Q8jU0wT0k9YDpJ1Qj+kzSpVjh63t+k0sVfp8RZA
A3XKTmQh7zJb0OSvho0sTlFsuUU8oWeuX1uVcH2e6q4UM384GdSUGJY9hmwAuHXC
q41gKoVDCJtN0ZSKO8au7hK7jofLBcpsaJnIkFntnoJsW1pk77xP1j598TxWpfdG
u+salNcCutnWQ3vwjJRrDV/LzTVC9OzLzf2m6C5o5iBJx4+8HKBbJLHp1sfktrUJ
RpUChfpIgwHHqKYQWhjCjylFEK8318lKLuKcY6xhZgJvd3SlY8oOfqTugLOFLApb
NEvEouX29+dqxmT285UX1rWGPsrwPblGZUoqUQEaZYn5gcg0j7cKy0XydH8D15HP
MAm8L+ZfTfaBBT1e3BFDlud/wsNrsyfaa0PENimZ+8fcBwz2vs8xGNJECGDBW5ni
wxjVd78teLWaRF+8atJFDqWcymiRdWqGcm7QI6apmDhzH8x6nFav628V4qJH9pWF
L+3Ojg6VB6lXHE3Cm8hvjzTx7Z4InsOKdiKc2rH/K3grtQ7Ed/cbjNPICdjdxhaz
xfhpFzExM3dIyRbo0xl2NYIzxPyXVLIlcjcHaaT5ExARkNFHCtYOBdNrjwQ/FKZ+
PSVbUinGScjc8ACoRRbi5I2p3o3v553EFzgbfCs4AY03w3OnucIwl2f4C6IbgV3X
aJzWybK+j6+ykgc4rSNFebBqATx3mGEDayqfhtuILVhMigRT64Co89IVpDaiYSns
mAQSFCss9Ov0cQtlh+go5cOIQ26thZqxNFF4PyfHVKveNVtTcgfrbTsS7GLSNGUK
TarUvomK3lukMFoLD/w2q0T6D7mW/kvU5IzeRGvRRbP5+qqvUibeI1NqBBDQNy7q
ZicZMVqZmhWPpVYW0+Fc9vBEPAaIYtGz5Mkdp2YhuQxaFU8T1GhPKIUFfpjbugeb
esBmTDw07PKURJsA/pFAcg==
`pragma protect end_protected
