`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ps4UE0OpFN1CGlOeP7IkVCjPPtQ8+Bb+Z+16xFu0K+U/zaBXfVM7V3zaGmvU1n1J
xAeK1cQ2hki4dZI79SYyR/AgAqRuRNOMPxIx7MptXNo1inqTrIGF+W1zWfygIv8x
LKCsg0eLPLGG/Ua4oaZOWWlc12RiGuhsdBY+gDli0C4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11312)
z3Es2Ur9HeX39v6bxunIXi3OtFqpvde4nKvQLQYsZAdoZV0bZ7UOhiGT61CO0XyD
VIiA5UHVuCEQxegPKFBlCqQcBsOvrOVh4A8Aq8jtBsVskV9FFShfxhNLt+tHDb1i
AAYvySnn/vMHpSLwwWEpKiPslV9cWaecO08QU4S7dZvSFODmI3iVRq7HbAN1Jyp9
1jy2H+34OPWhrgfwCD6jNyMyJbVN1IgoHvrpcXyd+/JUGEMwTdpqpIxO1UAgk6/h
KS/anpknD9hBxF/LzrW6XX3wz/ZD/gN8EDNGJfsRKGWk/cT/K5Tz6f+hCgtHsqxt
10Qdz//X91phipG1jypHfFUhxlQtv4bMR/EIMk4v5AD2dtOuMlOBv1aC9XgJO0mC
zGSUsz4YFVWdxMwGJl5loDvzXwdkznsJKhZWyVH+80vkJgNb/epPdyeEZosJ6M5a
DtLTMUqQrI0ZxCItuZ+0B84zRoh2m54KPgXcRo3/Qsfc+oFhquacPSkKUirzjdbi
xAt0wtJxHnH67hfPtpBU8XTsHR+iSrch71GNKzx78Kd0euLh2vi27cNFcw4Xsyys
4g13ZH02Ft/FY+KWn8dGvAEm9n3iaXoupCWADu/QGhDWk/QxdwSP40biwqrrm/u2
z0kAjaQZ+gtNH2U+BgglwogwQQxPfoDh29q5VTvAQJH/kN4QY6GeYZ0jAhQfvH1k
R0TORI0ZxOFH8TwnGty42gmBIRoEPD+B5MG3IrZ4yv+W3IvGkAkt9QWMqW4ayTNd
HrvkojIeRT9Qzc5EnRZHqgvuGfXROcvLN74zhUFB5K6bixtsBp14mJmG6E92eXnD
IN3mPfmNcZpoJdkibtIfJse4yUrFFxaAN45gk0LwulTQ4Uyj5qtPvQMDOr/hGVaS
T5/4iN4T/XIoNjnYIXYiaxPzywdqWoRrd9aZm3Y4CvUZ+uqXH0LuzZR+kNnsvQ+P
9DPOs17CqHLyqUVaKARcYCoEBCa3X+qsVh9obcZ0++IDOjTRlvxRQMnNHDKW4N4k
3dJPw0O0CUjDmA3g7GcCQLYVwVs7Ccj86c1j7HOievt9lA86kwtVZ7Vj9ix5wUEn
giNcyrvdrBMLkPCQ2mPm7ZTpPdAa+zdQE/5fyJYedreAfC8jx6Nqiu40ojqxbcGs
BFgYsxzdrB2YDrJDGqB7k6W79XWBx4LI0PJ3ungl1wHbvjF/M++7y7PEaC4D1NCy
7aYCiM9xTelhYtFpc6tyifyufvLKWiQ4Fcy3GSdDx38g5er6xll537skK/bBNKbl
RO/SqNjT5Rd8WNpnk3UmoANMhHdD4uZSIWdYnmcRQhYPrPbLfaOVmfrJH+kfip63
/GKtO1lB/d5yCDwTINsBbIvcufzEkq+TAII/iCn7OYLOTxiw5zIqNE26KUjeP+ud
4lQZ7oiUFPRuduBJ4D+TJuCPoex6ZmSUhUmi6j6xHLTLpYu+urAczdcGTQV7gKkU
1m6Zhw/q0zuNQx2vDvQPx0iCa68Sv1Jv/tRy1b25DiksFTMsUtWezyhUZl4rTzCo
bhFyaSGsLnIIq8UNnAbkuGnI84sWFHU38MbYxBYmXeBdGe4m+q5Z5Z/MMbuvWNkD
+gjc3coeT0+f6X9/2DBr2tEWvk12jRauk/8BqHwPhZXeUJ3WshpiRXIQQBiQpPDI
tLBuytF35sYYw47kQZt5eE8U4V+Mx9w2A2KE8Gy+Q0gjF7DzECn2aHWtkplVHA5M
ygQGW3HLeoyZIPLAzU5Uu8w8IwSi+fdpUnbU0SBtaRdJRC9IrlVYoqznbBBhBoTF
OdsVi5QI8dQyjkmpMQ3yoCYjjvyGk5dGCTifhGaFG0BySqIJqeAi+OOiSYAYjv8b
CHBY7UGH2ZMrc9zjMNHOUFEO67/5sWj1abqMKQz8dAgI16NLa48oRS58715cHNNf
GoQTBAC1+4xezUXr0fB1+tdDdeyYp54nMu2XHKS2JbrFMFhqdojhwyx+nYjQRqkK
Fqkr9eG1w0qgQmEKRsdFzmnxwz36DsEqI+CFf8dAKZ0F5CEkrQwRW1sUhpIA/wz/
oacrgvJxtT2c3dKTmjmMwi9qrNaMczqVAgUPdOSKiCqNy4T4DR6o/eQ9e7y+U2AE
7JKfG15Q6+ZNbJqPxYoREVQq8Pq4EQU8AYsFKnFlY3sEwhFNelL3Yu8evdUbEUmg
B7XYYfQI9X7gbx7i/AsAwlYhZ5pXjzW/zqHs0dvcTL5YzwxnVhGdmteCwNe8t0JX
f3qKKHDmRJUjYF/qnM2rCo/myYhZdKHTUpixr9/seCzjJksUS6S6tc8HR2zpVd7c
47A07fXGXtE3H5gLmpaOTME53M+ZBmHu8OAYevNe7WxAU9pAWoc5t1k2cUu/+Jy1
WDdVXO6qx8GCaNsDupeviINjzgzDBBdkR/dmFmPt/VBO9uO5wT4ugtB2AwEDFVba
Wp7sr48hwTFE/iTKlsCMrNUna9pkF2EG6XUcBu0OmsiCAt381mhwg6RubQANkL37
db4VrZkCT2uUhDUj6K290oghd+Ww11G/6qG1az4fA0mUA7brTpvcIOLlj1WfSzRn
2PKqGwv2a1JtEs2Zb1V5+rBi70vUDC92GiUuQ7gSd79yyCekJrB9g6ZkiUQNXL+C
U5kmCg+HuDywT/4F9vqrnIba1PCpphLB+8YFNHI3HnMbe1ScWczFSuyHoT7uaYei
qdVJKWnBLtFvdS5/WhcVu6V+aVWwEna9fAwJblXr0aEDcucwCfLTmOux8NaV9ojz
8XYWdNFuwpvUaWu/HLFgn19ZomocaGaSLoSjTlwFdr/A5nnxJeqka3Bea7DL2Wb+
9ipqiDfOJ3PYDSH4Eq8q9zeK5fo0qCysHMvL2Ei5G+T/+jQsA748l5Nl/knK9Mlk
PF6ca8xuTBFOAD5m/5bQQcxlE4M+jwfpT67glJ+3f9/1IzbDixRlm6hJem2+I35z
GyHudc70QEgUZDBlquyz1/Sk4loTTkfy/DCfb1037LGxK7vj6DiQ736i74yu6ecp
EH0gt/JTbT2CQLaOTxLJoi2LwW79ihoEcbPm2e1HjtCXmOuFPjt7Ep5W9i/2WmBM
S2KigblQGbhHuwu8S4EIjDr620VrlnBU7yO8kaoj1OWq6EcSbAPN4w690941a4ZU
SuMoaPR0UB0vVAAPSSW0evesJfaSDGOkY6Pr06JtDG/ukBlk48d18IeB0vAIq/Rw
hQcSFTPEKQ9e/Lq9qwW6VUPF8FYmw+aJoMFCFbFCXfmhRez80jCeZCAHsoTAs7WG
EJEoqVlYdu58R60uy5JFrczZxCiQvFwcNHsPlyQ76gSH820kZIgLUbVxuaU0IxCA
G4EyI/S9iiPFI97WEgRC5FEwiaJWVKQu2fwq0Mybbf3nSbzqQy4P9/p5Q5aDm6AA
ZUU/F5S4+hycZoNxJcJQ8+P7PeLMfG+ooVpnJ50WmxYxmPJF/cm3ByVIXBmB993l
Op96Y3vAFd7RM/5AyHbPC8cd0nE8GzIMfQmiWIvDC66MkG2RIPoYvDoOTwGUPOFT
obihJaXc3WajhDKFVOIKan68ez9FOSCh5xALRkmVE6GFwtgyW7GPcaUie7nsqNvc
p4m89m0fJtOlklLVzfW1nVSXW4WYQFilx60tazaFpXs6L1oMoyR/rlTwRp4mBkB9
Sx4w2h2XmAXHyXUdZjsalS1cobKs7D5Umh8gQrmTK+zauIgabN9a+PqECrRhEmFG
pC8sfl7fbjAcuxqwC9tU4/IkiFBw1p2pQ6pz8aGhqwhkZHmFgFv/aXzA8BoirZio
e+HQNZorYw97phgnNutMelY2/DJzS69Zg8KVmTzDSE32WE8KZHUvgRvTQlXVZm4v
RP3X54fqBMrFeCH8wSaHtRqzNs/fJHsLXQRCan5Dooo//VMI2nA62loISqlE9K1j
C3kZp2MSPW5qPyeMZ6zI3Z/L0xR+oZSAsw4Lf97/cTPLnEx65NeoTFZ6Drdk63X2
O4Sc+Hrmin2L+ZUIyYtSEhYKYbNi6MNVl0b2R2iB0SdkOzYkhSwZ2ityjimXurLr
34U61twMYtPaHTgT4Q4wvYgviweOOS4KRgA4nv6/+hPvPRRz5piuOsEa8YckNfyu
Smp+kkRDoGov+R/1k4FktA8FvNDPe1fCWw8DYfcUOgEc/4DAZvEbTUIzkCL7WwjA
iZfzDm+e0oRtThGuBhg4OQXWIZXKXVbLHgg/CT2+/yCDs0DIziHnsmzc91prmmY6
v2yTWj/y2eCwy18dAVaNAAIJ9c5HetvE/P7l53a9tDvdtCu4JzsCtPVpiofs+iq2
6fPfo9rWVKpBdaMV05LdSusZGVOCB1CRsa3vmGNBUHIEaE+8Zw1dz/aF6ASrDNI+
dfU87Do4J50FUM3uCBf+D/FMrsfdsjJ6nY75U8ARSPAmbs7C/6p9xVLAsIg9UKaz
WBZR2EroPREm2OqLlb5QsSmPMXy73nkUeCCL9w7+YH5uGmWiqN22SSoX9B7TC9ju
8XnHKULWa+M4mD1VErYJJuoTEUtW1Jj8R7lpST4/hFG3yLirPXhERK+Qr3AI6j6x
mVBSmiqFulbKBz+S009PYk2IhPOBoWtqS35H9rEGMjmTYtqF0HAW9x2PV9ezDcYB
YGyV3t6Jnh2+qN7zUlFWotLcANNwYh+qwc8fiT8KHyaLvwPBY5Qt5Y2fgbrq8Dzy
hbdn6rnUYB8zxB5E+1uhiKxds9mhs3uZJsDh4gtQLGcOkoej8d9/f/m9Sh3uuF3a
k32xzLgx+g+Tnhc4M/ZXllGdndcU8q4LfDewExylcs5eb6bTNaifDOefKTIeVj45
Z8/uLzejqkwmsU4Yme2jNMsoW+6RuFXR2QdEW7ACcQPeML1uhM4BQ8ElSKOyjqiT
OJjWAWLPFdlJDnonf7jI1Z6dQlpM4lc7Ujy8qJAU2hKXuSwuh2E/IRmltTvaGIeo
yeK3Ets6DdOQswLEIhJTCQlrXVo80uDiT2g6ysHa2esKxeeThveZPugimsa9Mgbj
axIjRaH3QZnLR9IagOYEPrZDL+ypz6HPJWqXyfM9WkGlEDk9xqVGzXLozh7iZ5uX
jlzqON3fgybruPnT0T84JVeBKU1QyUE/Dac9YOX0nsDmA50uxgXkJ0dhtvAqmfhJ
U4IUYtPLMWPhKY9A0bqmKOpx3sfePRjj3m0rHGlEOddjY22mAzABds2mecdhWa1x
CMa0YPgpt1/2MgWnrn9wwV0g59n4AatWOADf98IdbfE9kTs9fGm84o7kKvTDQZ/7
emuE4fakY3hmA30dT1uOBUSd/A5rLyfyA1m3XIbkeme+3K60CeCT0hQxhradutbX
XVHe9JuY7nV/dN6SMx2L1iZygZLRBZGnWZ+1sDHCMMSY0KxqToDQnzlH1w2viXsu
BS1VqvBJ6UaLQMOJYvGpI6LbUG6Fr0LD6IqHQmZUUarucnGuoPixw3hBDM9W77tx
Ro5gmCeu+rKOaCapyIp75gVg5l8YFdhqtf7B4qvK8gtJmK3GdEVDDyJw/smS4Q5t
VFtL7iGARUUuARRAyTcptvJ0AEVMaKLQJb2rTVVhR2dAxUplBZHElwtlKmhAP10V
e4vDip3wwdfBciicpWuhekM+Dg8YMuI8BSrKYPna7B+Ei0yq9cZECfn+tMFunIsS
O5QPAtlv/HwhPR4YUddPYTPMy0tD8PuOjJfdM7vl6LG1AAPFtw1QEsppIrTMOA4I
Yrmn2d5SWcCp6M/xlxNjKPraeYKJTk6hLUtLoePofo2ZQtxI0QZh8SwN0RzuCSDE
vxkdpCswcDNUXdtnGNAqqxeFLGP+iVbN87S+d5OW4uqGR3SdAqOC8TImLMNtB7bn
TcTIZGGzLTkMlL6+mA7oVI97qbfeVcRnRBPX2LJmRYelvK/WJLL7GpWalVojgTH0
Xwyp89whbZyJA2OidbhvrHh3jbgpmiCbtEnFnehfQjtZh2rpo1q4cpNAEcfV2OFb
p39wVwrcgv/r8+VuFoj5qjrUDRnOgxKb6NjzV1z9Wm9HIEdbVKaqLGe9WTZJHqBW
IuXk00MlNuj33KTNwD7EC6OdZ/rfyjK6uiPvc3UwXa/gKZMNjeKGwigkKHoWRCA2
DGN9XEfu4sWYVOH7ayItRsTVf/SOyCiF1ZEqkNlfk1brgfBiZ9HJjO0sAe9gemXL
uBtGbAuUBkt3nlvPA0axkBYFeGB45zVpgw0x1NSkHKX3lPZKdPLbfF60lTyS/dxD
eAsjIA7HhorwCdG/jkOahHTdkGJhSZfVAxa2VbEcKSc6Cj99kBxTJj0FoxFNMUM5
PdVQ7pJTHFIFfJ8026x+9DhFKtf92lMdmu2JpQhPgWRgPKJyHfcQP3vHzyU5DL63
HqdK2tfWxwKW2BFIaYT85kaAAcYjlVilkw2TAy4LmS3YYo/Rsk0E4+6vjxHHj8aQ
YLagCzof9U3gCKLSn+EVQGuILOrQIktSoBlEGUg7ZI6drfcBcsr4mA3Q3Y7rLQUW
frPt75se7C9fhbj2oiIfOGr5aiI2X8b5vTNw5GJBHnK/U7eeAJMTHy8kz+C51LsK
/eqErEAZnV+Ci5wnCYr5ghl1p8oTIfGXHtuMmJ/KUWn4mKteZwl5k9tKghJyS1Zo
PjuaaLikMO6RHQAQwoFEst9hTDhlmFpokI5MD6CtZ4PogdCxDgLZdLrFxX0shbDM
3mV2MPbC8WpzFJ4x62hTmOuFufQPAS8jiOTfFIMKDZ4PEV5DYs8zQKxtiKc3AAyL
D1958yD6mJMxEvHbc292Rd7D18FPLXgJ9vsu5LRUbnJpma5jpNYyjjs1Vyy/7UCM
2h4vsSZ/7KOf7TdGyo4lYt0B0W2OVG0bv8MufkYD80lzWHzjtx8skRl8ex56FjD3
I9jf6ihDpxUwpWUdQqXNrc1Vc1NrrmqUtVQoBXL7CtOeieH6Vr6OEEgbjH6OaMtI
Y2oIUbvwq633RjzkRkn2dQC9fS8BTn6mNFXEhLienyhOD9xHvJkmlZW3wMzuElCo
hqp9xYj0bYilwZiFOPnFBO7Sd+OQLS/AlORrc+TzDZdRClDQv+73+fuZ8eB1A5pL
t5V+qljNeZd9bwibCRIiT6w7fGxQAvZs4gggRxuqg+Mc6kLsAi+3dKT2w9QKM/8S
FYUGrBVJiD48QBFUcoqScI59OwShlhiB71v3SKpJA/PaD4vIpOZ9hbr32KhG0owT
I08lVTp2TGDIkvs2xNREIkWM0fFtOWDND2Wz75dgadSWeSE0hRQF7GJo3zzIZ4Ve
w6we1gJv6g/NKXlDQ4MYBhUO99O1KxWe06rddE8G+UCCJ0iytyStcl6vmbs7nqSc
tNlYWmppNcjqoQ8zcofV9hKQygWUF6ZujafRGuQw9czjTfv0tdNfreRMn1LXBNP7
8LCP04cOEdP4bgT5UpSGLSYZ/NjDKb4U1Iuc6d5K8oNyZKzHHGOdTkc2C2RmKFGF
TE06OYmhq/mh7x9gtLhyoVoGx1hhUfFHkHRJ4t/W1PWRsdHeSeLEQdzgPu5gml1D
RtguvwjddDYNNI2drrz5g/Cv8/A2XpjMY5DmZ2myBtYmzb+hWgHowmdLylTKVKWe
HwrZEd3hD31FkZCeQcRhuY5Bt0prsNubt+gTbG5CW9VwiLp/vR/iuEh0trnjCJuS
3BtW3Tu1IJPCLV+pZdZ+h1gqleS7pZmcGLkQ85k37xHGIB1OMtoWGBEFQ9fWYfTj
nC36sHD8ICM7R24u+ON44KQPbmk5wtS9jIajO/sVupOnWu/AgGFiQpItEtAq540p
MspPUpI0GMhXuf00ITLUcLH2O7hOV6foGnD3uVRu/ZJiUvq1Uk279TgrAyDP2GZE
6Oq4Wyb7J5OFyCxDCF7lcaShfbxGOGiaHJgVneUkjYl4+8MwxNKmx/QalJC4MViQ
/ojgHNqDgMwrpmLSIjDfPAKeLfVG8Pnv0920sR/17FgB35mUY1YQHPJv0WczLos8
e/g4d9xuoo73ScsfNeko5zBtq8FFe+pnOPVKwj6HTp6ZJaHJR837sAXrB4h/gSsA
wSJyaS/Yjm1tb+T5T/nYNYHCyHSyM8UBrCGu5KwveG+v6CZ9cWf/i2E2cHKmM5Oc
hGRut0ThshlocGg03eGqfXvY5FIfwSFGUYv183avUjlamc0Fl2UKXcL3+/R95FRy
eXhHGw/QzDYyrIBsF3VmWpyRxFbQkS5RboIxs7UctZ78CWipHPAuZSOBXdoTVCFW
aetu4MzFXAyhpSou+x2gDbj5E4FdBSY0Lo0/ZYqQXkVZK9f0lJ4uP7KWRIRcUYQi
WsR2ybv1rcGvU7cTd7qFkYwHIUz4LT8pNMU+Ggu1bDXt/RR1tZgVU5c64leL2O1p
2SeR+kryw2+QyGzNHdW2Ha/Twfi7SngtMMTCAZQ+zZxT9mjXKJQVcZGsJdl0TvHW
DNybSbypX017Nwr16BlDSDUQN5wiNEfNPaXMiiSXjm82D7bd6KBx8SPIzqgQhQAW
W4gtEag+PnpAc61F6noUYFD0Wdljw8iIE73ozgi15Jcg5p2h68g7uA2U1chUfjAR
SsnHyy9a1kIlILHeuS3tuzJw29cE9HQfmSmSq7BagDQSn9OlmIxQ0nolapeg32L5
L/AN5Rj0XXvGoALRrmI83Sl1rnYtIuCTJQKbjWKvJW83xKqh7HyH5b+nxH9Mhi2u
Cd09qZSY8Os3fqoL0VzJnVh5c4ylNFUR9P7avZvHECIpJzQM6C0+Cm6LTmw5ydZJ
0lfFInxu9vEUETZ8Fz4Xw1olEddj3Pynng+LGSVji0EEyTV+gpaSC69noeMtwrJy
bzOERmJQlk3uTH98RgumNPP/JxLTGyq9pQOu27JXyTENPyMZm/h4V8OWdv3PYYpj
Jmrqq+PK7jt+B7FosS42zc6OlbPVYnYwkrCVOr6eQhQsa8gD0Ck1W9+5icaGz+qQ
VVAVHRyzijOjJfAZqeBAvRf9bLhIt8R2jE1lVLo4CUbsBA/CJelkL2jbHoMKymv7
+x9hlz+76FiSo8iOdOFTgfBwjlo43bjDraMwoFvwQgSwP6Wyq9TA7rFM/lVTLsEj
P/UURB8yFvYHV9ZpS9FZKtamI7ttGkCWRGNYAwY8lBwUWGHW6QGSSxo81taKfHhL
Oah7rrUeuoWokGP+cUTtLtITnDUW7IXeybLuBjigkwx24VUd7ZzkrjCKWNGYyB86
ZcgtifytwQUx+Kg46d6CX8lKYNCtG7fukHGRMOQtS+gPt4epvHg90BFp6/hgBcln
G6Y3/7uV81gZvAiBNdU0AKGo+cGPKUsAPhbzFNw8rWT4NZUB7tx0wDlwjJC7lNtv
wzzQ9VweN34H5O4HOoSwKTrhtyu4APHFb6AfxA+vYHkNXmkNc4e2xwEGrP4ekJcg
YBz6aTwRstR1gushlnvDiLAHvrvxJG+pizJFpChiKwfI+FsvfkdjNK2AWyDtoYUJ
90rrXDOWci6BgxoQ6snBayt5qDLeg5mXL+ZsCD3bXoRHUHIfValBZAIXLE66NdBq
zVUXXIf6ZTRrZBqhb0DZJ1IlirTftc77kFT21DG89f5n/m+QHeuzxzAJNwIRvafl
kJZl/eYbU5lht8I6dxqalR3RzcgRZuW1oQmHDI6jPNv9+ST+Pk8lm5E+8DpNmYm/
Ua+LMaWp24UsbEVhH+tkdIE9EgQt8hVaeUZCIOC5FG0NSgHfWnXSGkFTEU7bz0Yg
oCx4XQNEtW/COey7Zxyb64kmfH3tlpzUxh/WpkEZPCM0VTJg9ZQZAD0W4dAKvEed
icuTIjqfyGCYvI6k/PnVRslHUkneLL7EqwelkqNA8emM6Z5VSblSsKJcL2lGjCWX
mTjgguio9tLRAVRykxlgO5/AVqBEDbSCo9/DUzLCgOfB51+BmZoxWf0OZNYoZMM+
f+YID3fENpg/Lrnj1Y1Lp36q2YNJ3mE1ogGuIDWr4NVXG2exYx1pAI9ed6qGKCKv
yrUFMJGrPJytfr5NoZsfEiWFOFxR+OUcSsblwnaVhvZ1xXj82VIjHxLUPb30IlOr
eM/52BHoTlKbAAuhV97fHxCUuUfZXrvmyktgiOhokPAVC37uBPzeWpq+3zAXivN2
a64ta6dCC4tlO/iQBxX06RcnQTp2/64TwU6WkjDB1wu9wtlLz0pjaSZlM/dNSR3d
Swq/adgsbIx0GzAXDNIhZrWth5RNrC+fVVtX4CDf5bFJ1Ql2EDZNzWsm2MvoWsSI
IeBb8X2Aeu7+LkRpYRcWpzCmk6oiy8mPFAjdc14b3l3LcZTP5g+plPeqjRjyt3TX
DOz+Ou/CD0SkAKEAcCt6JgpZTVomT2fj909moheqqFA1zyWvhp/ApwuCAw4Jx5Xo
GaEHm9gkBVyp3R3gcEgBxHzew0eyJLC4o/HjtJaJq3h4rOTweqq8ILbhbz5qV3ZS
J2BQOtQug5yyG7P2jzxaXyyvQdSg/nSrl6oO7EuykhO4l0Dq0HImCoUHYXl99Bbe
2SZDfW+YwIKvo6PLcX4LBpI+A0opUKdIQJaOs5e7/Qv8CJa94qRBMUBg+yHBAmEp
D+0yw8WkkZeMA5Jb1EhnaCtrfJD4bANvs8cW0YgcfFbeZvnZ7QmPHXmWf2/QBjM+
sdsw9dmcFfeaqlBup7aNEIHI7ft3G96I1eyMHWejHMrFgvDyttFROmBSUG/TyFVw
wh9B1+HjbTU9FAu5lHh55YZ2IEfZU8n3/n5kS+H3DSqejrYeWxX6VjmX6Qexl8IX
Jx5U5LJM5kdf5GIdJLMU0C/wqtypQnkO5WR9R6ZaKSQco3AG0JEM0B40iDWalS6M
zrCFSgwDu7ZzUA7oCad44K7gGwHVJyHKh+yB3i3IBenOjouwX+XB6CQ7bTATYSfv
XiAQcDDXsrJPw2cgzu4VfIMNX4EwxyczxSD6u9TduK+jbe4y10anibEVQ7BhIF8R
F1REWCRLMEnSfru+evFhBQqiuODLTez+PukaCcL7VF+wbunyxGB8xusLwBse7IjH
RgLIRoB8iK3MpA1hDUIcG9iPQjWUa7dSYGPl7E0JfY6Ww2pUqWjUhniQfl0TtX/a
kE5l/ROinVHGuHF4AhdC7YqVes59mgbpK9dhRCKJQd2dFKBPWGFOElFuR41ELZLw
ZuhhziCpfiyH7Ah6OccxnWHKqBxDIsk44Zvx/DelFq8sISX5S/I0i7E1jFDkG9dE
kAvcitKQT7LkdUgWl1Vt6oyjCtga9oo9oNrPgCC1qZ6RbTXZkUsWoRdePUPLxERQ
n8o28mYW3uA7f0PVUs+zvrmoOV8bUmw3rvj24Lvk+0CzYbIHsdJJiYIhyvp42qQf
SeO+G0rqIGHKR/w/GRguL0H8/VyeswJiJDVwuPY+ozbet9hlckUUkk5TPRsUJLfo
tUOwuuiW5FZ+DZVdSuXiWGnUB2F5INKlIeJrFOSUwJ7UqY119UVwn9tQnmP10QL0
nY/RKYd1IE3WebA84U5sOE3BqnubiymGdKX/boRfy479JgLDJ7+pUw/rEBNUvjEo
e5QqETH2toswJUvSBx9FrAqtUkLj4JIKSgq+EODSVkJUDmwxepj5nwJBsYQbhiRs
Z9/3XTd0J6Vh5p0PUdVTd5qJD7u2s4lMRMWrStVWgQvnHYRNNP+HLJvhA5ZWkcPj
lk3f7crAWJiiiXOuReVSWpnE1maCT7LyIAcNKCmkxwde/k2B+IMNgBm2SFBsfHz9
f0Ul3Ga3Hhuv5OhzSkPKdg6stVqMAVlBkeafH+R6QULnkp4ffgT0U69CSGwbJCnL
2PYciGSPPzDeNgSJJpcDFbriB6f1Z0MlMqES7BI7UH6nvHXXBUpAZuhctYgUVJkX
Q33TuojuONCqTLBL9WPrmMB2i7kZVS67S1CCvhtSCrTX+EUaca1UOfxYTE7OTQfW
jzMSNyN4obMzaYBriYdLn5Rdru993L1+ZuGB3PthC2UctV8JGLzN9zqE6r1UacTw
cfrcgBQsLxBOXkJM6V8axsIJlVyCEcUorSUlzx8idIzH/u6TDe1gxUl9pTr9FS2b
4J5WJgk+mf/sxXb8RTEqiLw8U/+QjTEiisvDrXs8CyBIDNMRvcGou3fXjHg6n4Jw
0qT1oDfXn4JOThJL4EtugsCXJyNGMmkuENq2luFTMwTCQhjW2OxrtluB0oYKa7x3
ppeD/glkVZjWegB0mDHrK80rSQhFY6dE4yno22xZv6teaHvI90lxiPHQhCGLakpF
YPuD6616099tgHkchYY4YORjVWxR8L3iM+SpMtreQ7gU9RpvvhIfGVjAOpnNInvT
Wvp6NKYEbnlXa9ZUMyr4rb1wAkMYQ3oFsacal15jgytrBLRBpsSMtny3tOzT2Ymb
8IH3H5WgSwlGiam6eeL1rKXV1NL+rqeHM0msPJxGbSYAhSoHEZzDyjHhNZp0bCys
PqtDeNAnTYEcn7lguUW/MPBzbzhzhjHW+QZlFXFIgxd0ZOcGGm7Ip48w7kePk+5n
k7Rw2Eo6xkoDYpJVN/0i7iLUhej32ysa6sZvaL1nFyXrkiRUEfemnjXclKnBNHV5
m+BSC1Qb8J8qJrR8wnb3oDX5t0W/9flnuGvBV2n3CFFQH0f+VftSQ6Dzprs3e+Bf
pwhW3HQ0DoBzEZr3jJsvXo8rMjo+H/MgkiOwq3E8rVN+HkcaCODR2F2fGD7XLPvQ
SCwhAUo+pEf5P0JXIBoDz5jiJ8OdhXgNeVvzAYxKHwzskLFOzoeukI23932As+6q
boU2jQtTP2eDuhlufhIqLdYp21GT/5MycfodyvHehqK3jOO1XSQg1Rq7Gp3QKQhI
73akaxlXaycbdlRt1+Qi6V3A090Vsp8UlhdGYHkQDRJmboTAkYN+MaAAEgxA0N7k
dVZ1E6D6v8OusI4Sl4Mhff1brNSMJBPTTUgGt8d9Y0pc/eRdAZ89mwu2ZD1xVtlD
LpXMzvS63yw4QaDtnAoZ5jycITQFgnX0pa8qUvUbfapg/5N6HVQiHriyEc2LQEzI
p0tUk1LlNvbfK2w/AfdzRSiHWj3pZI/38ZTpXZCuibwEM/7pCF5FipB3+WqFNYy4
QJpEi7Kyo9EyDtzKq7OYxTrbTWo1WG8CyDU8EJ4uUMZZAWrzAS7KZmp+rMuU2EfR
h1+1Oss6T71eCmMN/LQ4+hf2eC2wtGsUYuH+zpKR3hLCJ8+deMBZinkeFtAR6odv
/NV+TR349O/0E9NYhAKVK3XFQz6j1BgSM+WMizvzINK5wPY7y8yE4aMFHzYlla08
bkz4wHhjoWT/toT2glySscRKy4zKH8BKLERV2LbyY1lFOvJB+ydHZdTW+/s5Io/o
GIpZz6YN/4yCh8IZtWwkUGkGbq98U8F1Z7qzMbF1qqzIFrtKJvcABf6X5knrmE44
G+WXwEay/93iOeF5kZnzUerMz3d20/gHBXM9PT8igNIAdKQx5B2yJ0VoLfAQgRcl
/PAYQBkpLnsHl+PDxa2Y5tigfVdbdaIk46nAUwZKr+S101ne7zv73mmhay3z+3tg
JqW53mkq9FS0rmCGd2epPLgFYSszgKSyZqEQVvmSkdrBxM7LfInNzW7Fhaw3JL+I
NWqYEbb3orh9uPr0RtXRnupdz+gddkG9v18mP1U9Vz6XxMYb+Xc9TXt9QmafVUGQ
cggRiQ2eKAnr84iyDbHLVud+Dx4gw+gAGUmOK4jgNqXEvOqeNcEyOxGebns2V9XK
PUPT/WhGC3cmV1DScuTYyhSnlwC7RkhMsKpxr1GU7m3IinLRxVb/T1y8w3krXE6A
MriR784VWPT5aGCTazjceB5EE0RSvC5GUOZ9mA/YeNtXgMYJpi9EL5ysWL0VowxJ
ipexaNbzjMmjrMdQejt8YIz2xrRl8dTBIqoWE/nbOw+iH2IBsDICjHC2hcAitaJI
zuqx3hSX+WEnjbftmAskmf3cezkSjkQ/u/WO7+ql0hu8BBXmLUhGIXz5rXfEdXW5
2NkGuQXJCvtJWZvG610bk2M3nEX6f3nkjqP0qDN51t0tF1K/tV1krnltLYT0LPgv
THmXmFlqjxqZugEJXKeyerSuxHyfjg8v1sOI20Rl+4ToWNYRKbxV8rMc4WpVft7a
NLoqXn3lexzV6YwxjNCcfPiOIJF5o2xUQdmegMQ/HbRImqMZbhSHL71FeDAiP9uj
GyJqO5Bs/4rmWiWeNK3olcGdqGNXZQEcPUEw5nrexiyta0ckOFy3yd/PCn+/RLdf
FmXEK+MW2Vw5196Hf0wS8Mcfh1DIk0XwgKkjEdjoRGdeV8vIk7OsQrzOrE6VoNOm
Z8Cd0XhqWomPlN61yEPaZqDQJyDzj4PuFMfTpL0m5JGAcTVMZjpr759kpXW+c/dx
nLEkrVv39AmrSC6Vr+5/4lkU7b/Zl053CzkXYZ9WvRcLNSTJdkLcCusE0yra5IQL
RrpFAP8oohz5pjZDXPRQwnxzuk+lt26afFHRSxW8nlwtYev3F166IEZyb7XxG+G0
2vwpYpmzbSzI0kQOL5PBfZpK7HE3BPshSqCr1glXVTjVZZT7mTn19WENLWOmLne4
OnvDBVC4xYrCGn/Wi/WXDndhZBb1ZjqobMXcv2edIhVz4CbsPYgpshla1X+Pu6vv
Q+JPNtoIFVHRsDHPrzKEFUX33VNaP3KWs8xAAx8W2vjEA9I84zht30lx/2aulUAW
6+ZrRY/bLn9wPlEtS/ciqQgQOM2mPkvI0SCxk8bUebx8EfAyjnAxHoZGxgPfevqO
naiwHg8/VCVSb3M7a81akZE3LvorKCQK42bJ2uaKo1QX5STRcIR8DrwVxwRQy4NG
UFxBP+pypZOeHHhwrVKLN+d6WQoaUGg0oWy5X/QlH1JfJyrjUnAz4iyKmGIRGPO9
LmCnKRX3aGAJXTfjJzCNvJrm5qp7sBPaBcZisCW/Ssi4nivWTyesw4WGeq7CXgT7
E2o/EQPcJO2e0GUTsKmOgSuYKiHNkhTEwXr3KQYxQ5+6bHRKrg5ykt10pHV7/tJo
u3gqF8nsHIPajTCImdpum7uTpngyaUIwwsAzje1PQNbbigW8ZyhKwQ+Lmh0yfrEJ
ddNYfROxM7RbCmWWNLRE6qe2TeNb1sDcK37eeF9ZuIe8MzE0XoMz/AmNDMDTXbie
woahhc8CrxT9Xi9PWsrfvg2PrRpPzxXZIaIk1HtcEp0=
`pragma protect end_protected
