`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MAsv+C8BRcU/6wRVZfCeCoVQiNxlp972HGpIlmLEIK0ksgvuKTekRjs8Z/rkJBK1
DHvixn7quVqE5YcNrKAzdklZ5rr2B0uAt9E3JYJu3R8j1vmRjZ0JhZ7xaoc+o7Zd
NJD5jZhGCI9lH6Wmg4aPET4sjzM7NAO3gk2fA4oyv3M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18352)
AMdcjMwMiAOSYw0C3xR0ONrZc77aZ/jwPoluRJDAa52IlmllMygUNvcMyB9ap1yB
jZSc37HXt6rqRSjhyOY3SpAUzPIq/lOiWQorKvx/ALQEpYybQNN/uZ7uMMkABXYb
n9Cd9C/1h4pKNA+k0i8SvWUrIYrmf71mE+H1ENLqpmJnPZMcQAlUnfdl0bLO3dvG
PiVqLSHeF+1l8quKbf3NiAO098m1qDeOEDab+NMVHIHzuh+sNqyKnCB2EzW75Gy0
KFYRcbj4hQnj7ft6/INwqCQpCzMT2dVwICcdIRlSDqmdBKx3GpVLAFNo2NZjSMjS
j8nAPy4auExEp3klJgDaWSUuDSt0pvBg4CygT34/CNfPuRtKCgebIdW+wZ2OVmsy
pPC3/yjtyVtE2l4P7FX/nLQAKNHzy3WRL3GQs/G9/21SC1WZG04n4iZwqanb1dzT
ZO3rvleI+NYc0rHDxHOwoe+D4YjseZ+JmTOJ3ye1xfOj/wSd4jZ2Q6dlXVIFQTHE
M1WTRNkTsJtGsSDPLsn0Zd6SuRPzrW8RGGtgkx1Agp9Bx43ivnRm68+amwaCHuLu
IpLr9/jcN2CIQYo2DXsYDNq6L19XftBGjpQ1X3nZdmvbzz9EOdwafuEqFVf7i/fP
LajxShCgWOKqTJEfmAeyq5JOI35Z8RP04tXjdtuADor+4H2Uysv3AGjCOORj8nLR
GkVhnEeqsriTLGPrF8ulRwvy/jnAHd7VRmVecLZEf32L8FXTGqxyz6jd217l1QJA
2ItF5T5eutt3+p4JIjqyHd/qEaHcQFoqbW94powXmR4D/sAbEJSKDoVnJs/VR8D6
xWTyAe2mGwe4kb9CCY60d3jNIZNQR1AzZVJ+Iiza2Nsd+fPQ+6/3LT2X9HIqhR3B
2qOKfZsw8aMW5+7ofygkT4KGoYlZLP1TqIZqUJJDwjN49ZUpcmWZ+Tq9D3UKKI6M
2QdbnKjzf3qn39UDGvj1EjwGt35OPOoZzQI6966vVBrhWpdCwZ9c4LW0G5pqFZTH
/aMKt7JZso5fePiyGMQqfFuG3A0Ro9bOclbKK7zTDRMCt3XI7R57njWsUK6cSRDz
w8mNgmhXklEyKrAU7HIa6E2KOJrbIVqSLGjE8Bh8X7WiwG26rJqNrIKhN5OEZfqE
UwdRI7qac3Z5JxhmsBHQZbFAEHYi5Kqx4OAVuVtnMPym9yMwLEBkjKs6QOw4FgD0
Cx9xct2mV0b2yORl6UI52yMRC8hL2ErJ1juec3FAi52zVy2EBlpEM5mu0SUim04+
o1DmPB5Dsnsi+vU1x+I3HEmcijBtDPlUspJkFxo3jyHDRxGhxG2dXmlBvabOQDbx
8RnLJyTKdZiSKKFo+Vu7PsobKCxArv3GAaWqe+vItG1+e+54YNzXFQCyhinOh0gv
Y7uEyIr9N1CXWOALIkxB/5eLkiVXnereJwsnlDOSXH9MVI4Po/TsbHmvSNzeW6EB
W/MuBPNJKtmWrogznl6hFVs0wvIK1kWraaZmq76hCSU+SS7qe8iJt83zz2d7VAli
IXfAUE+jDTxK859Hz6U/V/bM3bjujQTuaM7qpN6/ojKceVrONOqLlC3+0hXIEgOQ
YvCVIsA97M5U+z/J2On6Q6R1LafhI6DSGJmuqtkabIASPHdSBqlpmycJfkVI/JON
/EP+P2nbor8tzX8+z4serokElCCrJEc2j+DwP6zPV0MOPp/6I16u1cwgHOAQMJcD
aPjbzhgn+kuM7LzikNP+iFPVAqoOt+nlKRR442/dUKpz2aUrd3EJyD8I0BYD+mBa
IzAkPQr5GdhvoiqHHdt72z4b6nBOMAFRmuXnlvUEJWsaHkjBHss21SlGkdZB/n8e
OEb35nQGv1Ll3hwHa9tKwqhpo8NEpcUWjA8RK7TUdvoWfY3XovPste4hhmCJPPKR
d+qg6wxHWwF17vmfuu6XNxPPTF8mty0XqKxnrDA+NCL77HQrjPxb3BrxhvSn57zD
8GyunGJzgw3skA0uKKQMtDQ60UU5ZAOD4981FuuQlW2CKUjpEchLc3j2+mlE+jfA
iX2WyCYwZfSDLWtW+dY8DJ1so3vL/iGioDTgH3ft9rGNe0otC+ZECNXl0OFHg6Db
/2zOW7umGgP13qHNdhIJCJ+RbaMNNLmrsMBHraAlcNilfXwbolTdU8Ty1il8Jlq7
g1mlHahBvpk7pilgPExAtnJHjZ6wIXBBJi/Q3V55UJPW/sXKvDDSScYV+FBO+uLf
zxukMbOWdOYXqe+Rgv/i9ONUEVXXYfasna2+0WnHtnhKSlFM2JSRttcIjWuD0LmH
lNDQ0k2jPMD/WIr/inVoVVKS6NCpS5zZJzOmEHBVt9GxtFxzCmy68gFThYdvvVjc
BbHlSoDQlCC6LeM91PxawlJHGvvN7fOI6OMR4SH+ICWgxkQrvRDTm3whh0pu4b5d
IdK3Zo9mb1my2jWQWZya8l+Qe5PWo8J9F2INDQCKNooZwqHDRgbRyK2+ZkC479+6
mjmtNaeJODVJ4ZfAdSbNzThSHZC/1W4zfMAnTWmkwEQSZgIlq8g2Tc18U3Q0gHOk
IL38SMWmJyQw5PcwzsJhmwumyrsjGs46OlSmd3Zr0eL6ruE2jcFK6GUwoXozNAZa
yM84q52uwBmDo0oaU1L+RlYXfDaWqu/dnbuTPSS5rh3FonQRKcnIEHTVpvWLIWA0
yex8Pt3GJabKXR42duCC9GNv5slWz3hUbTxnDSEe/DhW0P1ywra1U292MhpqOVPq
+yc5C/HPz3THElvD0oAK/VYKYODqNF5TSKt3A7AN4QQD92IdnnUUl8d8mfXz04N3
jSjHZea9SvmJNTuWXPIHoQj0iHzrBuADazUhcxMf6+FMUzsR7/6uHrM8NzYDJcjg
4DjHkCTs8KAhka+IGMZSM1nvCQy5Vs8MgI/jsh1WKZ24oo72m8bMGMZrzi/vbD5/
Bpsa+TrIVF+HiiDWBWG/u1wdMiH2l/rKYskbTBnhrutLzIgZ/76OHzfifUAljo5S
+sJgFqflfyE7T+h+ohS68tcSEFDnlKk+rt8CNKkkTQ/3t+G7Q/hpPsnlxk5Natz1
2lRUZ7DNK7unW45LGt4r3Inx8PSwswZ64xCpAjItZv9Qr5yAuSRefpapWTVLp/jv
ZUos370GtaZNrEaa/0ucF/oanH+WmEuLI+hIXdHH7X8bUkUcEokM7yDdSycjZjwI
DyD2B1jSckiz6TrDZRKn5fvMm9m4ME2/oxv7Ap7iQnUh5R55/zeWdDahwqGO49dQ
Vtvw5Rg1aE6AoYEuzr1pnFf5MspxmpVcV9wJdr93gb2bPLxfj1WHR9BFLdDbAiNm
ivoaN9pz5e6lQ7L9Wqb5SJWGmeXe9Lo17uGYYPcGKtuqfpNPSh7vcOzydcC5lwF3
5nLBbGkdyRJQIGiw1CK4W2KflFoNxMzvnRUydV9zuXRdHszr9es9KwxH58BVESQ6
6uGvhPRPl1TEQf6dd5PFowR4WAkWXRtjD3HnwXqdDNuJc3rsDM8QgNJUKyao9z0E
49c4X58OIDef8+za9GmW8F7h7A8ZS1YVEOyF+aRIOWprb8AymWocgb7vRKP6GQem
D+ho7+O81ujkTgtK5ECGuOd9ogM+pg4AtKMGvMvJhvEwuw0WYZxMIqvJf7AMFDkI
Cx/M/C1l9iV7aEGObujAXHQWTps48Q0ticiLCh8V4y+BzxPO0cVBS4aluH32otA6
ArYBSfO4TJBF2hwUAOe+vDdw1mvoAEztUHYBlMg+J5UaqrewM1zDPSXyYLIwbHiH
Pgrz/j6QtDIQENbjcauwRUiN4978jXJ3K78asoiAVVGogvnOYeMOgwUG37tAn154
bngcZG9KsKlFTtMUt4Ng8znQqU2lHVl316DOq2Gp4YU5doi41wr4Ukhvhvbbe9qP
UwGN/V2htApQb1e+nNLGBzP0U2sQHkU/z8+w4CemG3WeIacwukNwH1GcpiDefI8i
76qqZvGfq9gTBRX56K2F8hnCAeqZLN+eTyiWdWIfV4Mqnr6xDzynb0l2Qdwlzjz9
Cgcw3pnC1BE0cLoolvorhENMfqLDX9ElmFRZUX7qAf8ikw1qoLqPh5XrK2gfWxQT
ZpxGqvcZJ3POuVrJi9/eoMcZHg8atUM4hXpdXQPZ+4GBKSaFjaHH64Nr8WsxoG1k
HNXpg0CYWzFCi9iwNOlivYeuA3Y2Wg62jatCKobK4JISHU1c8JFfkkSSmHE/zXJZ
ux9BeVmNWIyc7E0++4tZY1svCzDBV+v6nPpvFbqz98zWn9m0HxlsuJdK+dRR+Fa+
ZQVxuLZ8WkDODuW6bEKlauHQRRlIaGPPFyTjWV/4QV/WYEiryySZ4PJt+FdBDnyy
bika4t/gk6OabfEXfPZ/2+hsysLfF74IXVGuir/tmg6xG11ahS1QeVRkIxLnyiNt
ERGqcDfSUGXGySQjqW1VSLwseCGT1SZfv2vUmbmHtD3kK8X532eAT20LPl1uCT8R
wFCo+cyyAGExCjZVJ9Xr77ueEngP08k7j4Vnv34YjnP23nD3PDHOz+3LLQRltIhr
zQ6NhBZUMZPz/2plEh8fx/UYGtlKpYgfQ9gpTc8Hc7o05XZygOF6DrqJRg9pFv43
QdyWi+i4CJ5VHrheQOCI4Rw3LPYmCzEBrC7JFMI7VM4m0woAxLMs16HihT5iqs2O
K461ab2OeI35cfynBOxOf8qufqHGj/wkFrrSCEkM6sLRek8MMlMqnfCY567OxyVt
I0qGBD207cShDPbapPj8SV0Gs7q/nTj5QB2YLaydMTeZgKecJZjXlXUqICVHCYHD
+0yJFBo+AOvKuRjJbkG83tm9nzBBFqLd9X0M3C4zXvrATwzHFB9SpJYVg6ZTuxmM
rvOxEkzawPNz911m7wN99PJv1Kth80+li4r7z5Vsh+gmDQg5fNuZ+ScwYcPPzCIG
LaLnA0DVQYRMWdVuI/Xd0Sx5h/JSAx16Xd+gZia8leorYnWHuoXi9k8wjNxTzHpN
HP8Ct6jWB7gKUBG5YKO1x2FUO2qdxt2uXMteRYbnae3JGj9KdBJsnPx+JBUtgIL2
Uc3bF0Hhl0Y8r3pRb6ZnLmFoZMlJcrAcB6l7KsryePilZI3jA97ODf8Y60JbG6Q8
JR5R9TejS7c4CEkawDZmMSLgPEXZei7KFj+lfzCO6VHF7FDtQq9V4aizYV9SVMDC
+S5H/Z/AyASMqXbA+XD1CoV9IeBaLYzuhP2uA9XdOquo8cpVI1WiCOl8kYRObLwO
Ukl0GE0XV6QecXkaZbe5yJJyWCj2t1neTH+H6gqSvxacCZfOfzssXMFbLIOGL/uT
7X6247QHMtYD5uiKO8hqxO0ORZN/OvhlrCiCMUXYjQ98TEi2yvtcl+WyEksoS+sO
OFzbN2DpFjACGhc45aLrbuOAniEmiWoLJeaxVRm5T4gdBXvo4C1DJL+LX0focxWm
HmikGRJznXZkykFSwcd8DwOr8DKjQ9mBxnBJVVc+u1M103X9ycCqm6h/iq886amD
ZdX8HWGK/a7CzJscHSo2mcvASxwm8Ani5y1IN0lGeekLMJ3ZGWI6X+KZt/S9Fxsr
1Py8jf2r9biix5+iONzr14afHXFcxRXeiHMTTzfwVbX1iSOk4wowdbIXupyIr0/y
fpsF/XxG1AGc1+M5v8d+yFsV9jaizxBUeRiS1hXvvg9fv3iElWQ+gX63/xTSHkSe
mso0qxX+yFOKERP/6vr1btWub5qsKXGHFiPbWc1I79wu0C8+cgVdKgSU9NBXiIAy
N+GB7x2uSlYprW8vF3q2huD86ShBRm/XG+ZK2Va4Y+dpMlyePnD/uNrTLO0U5bB/
h3wuRVwgyQxBbOUMMDCqGuJSmJYE7+Kc1aCsJQ43klYKK72GqUmKBwWqK2vsjss7
q+xzvcZmpno8UxC6YyzKaOMDMwsjrEmuNTqghP98MJMTnDpB6SM9onOKyILRo3Mf
BkmuL8+2tCT6lF/Jyw4dxE34JKfeb99UBa9+f2aaz/IBifWe0iDQxelHyX2sDEi/
AxLNusyxQrJ8uOeK1ruhlB5QRaww7YUYs8Akz/SFI1ydZmnmVO/UTDhFFPHGbEfw
5q8DP3jXoooLyUVAZa8RwgSYF+pk3ePYAmPam10iF8zUzf/wHZSsqgVowSxfxTOG
w+NWp5hmJLTkij31z+LW3BhwD3/kdsI6bkjOo9IwhOuAFS7CvrIFdEQ8U6p269Lo
aEMgrVp7NYfuCxhBDeDvQME3njHW7HYYUPMUunAR4FPnZrnNoXPKFK5dUWvFWAmQ
VoxZc17kJXzaSx+G6ILIUYq78ko6u1Y3q1vtOdwiFAggm5dEtU24s/TAJnq7QSpq
qKeq3v4anH9pOIHflUoZc/1FYRHs5YK5kKux6lFginJcUIx0pHrW8R6CVcKqzG2a
8nyZzFLHF7xTkQvghhr94KXKgRh2G9/k5JoNQchU6t+CyK99zslvKu9MZIEBZlta
ApP58sqrMM1I1WYj8SXlvbMbh4TPQi0Hjav8qhmcNA3AoZj1UpDi/apU+Dl1r1lU
uUlR/+DohxBwMzVNbfQG0n3FcsROIqizvJHNkKmaCeOfp8DViyrYWOKkWe3FR313
XLBC6rQJOYTDGQDDarZEoL2J7LaYaSUKtAzihWHVG3577FmqLvyhZyVZhHrcDjVd
2eVla8bRy6Xb0rvSGkGo5yNWL24JsxAJjwoRMEneqTdGMNQRVgqe1ymBlNiYBM+7
i7cJBG+9pACUGzdQCF86jmvF0hnA+qWEgxbzDlDozvGeXr7vKePpNJAdXljKGTQN
gft1c6SFuu9JGBB5D8BwX7lYpk2NWUoFvRMbKuXpOS5hrhkV+EkNT4VO4mXPPsbd
EkxRJGnEI0xqDNdukbqZkuU+mJ+qNDy3/eq7xp59agcLeG+lY1HPnL8aNk4+SUbq
7oo1/Sbt2MRwIbdpitcRYLNeuKb/N1rP5EisFIKLSDTpGjxuCm5r/QYylzSG7dCx
y9MHAnJvZEe2Ccsn8M2/0XswLUHkp+Z94mnLhP/Vln6u0JeY2si431egu7m1z+C4
gzrQ7IbhbJL0BdL3jKpWIGwwL/Fir//2JXEMyaGL/RHz3PhNGOWpyYWcByBJJJXc
MNAMcXkZg4iNyuAAeT1d626g3kFxWFOvaYWGGo2kkD6a50TsCMLdlxNcbSnKUUmr
3CMs8PPZCGOmnGed4RkxhW/KLB6ilNxCZyf3rS1IGs6m7OM2o8b5qeDmzVMl0G+n
4SxVAEWEKeOh4UxiqGEDpknXK8ix85MZkUpiX+RSdHGTghxndM+8ihC1ezCbmU6g
p7YSYi3iwdjBztbQsdYw/hRrvEg+4spQylqS0FXjzqPU6bbcqHkaMr3b0S3aU94C
OVKpTGP6sHj5LwZctAQ/AMwWSEDBgLQhlT6N+J74ha9tM6nneqWf1mgRsOJe2k6L
6Dh44yD8x7dkD70rIMlgnmAL+3AgU+lGVEjmW/7qqWG9tolKDyT/4eymFCyWwwiu
rzLqiFDSI0IHv7pha7R4lew1W3hUDAF3iREX9GN9bonpV1LLqgYFnx0J8//CBVDr
3kA1NFyc9ryZ4KKzK1Q9td7zdM6/LVL64+kOthXWr4SsQhxOQgpI8MCaKkSJlyoT
n0v1GIoE26MhlJWuqLLgnyPAXhzRGkGvjZ+fQxaTLtDKdObB9KYxgWkYzWj3u+2O
dS03gTwTKpr2K2TPBX1e/wEFZf+QNgeYfZK9hDmrtnwyR4hRYUt9psFfaAAv6nJn
4Lxglmbh4foF36alwJFDHOAKUk0lQebBS0ZmBZ+FvpHXVU4L7r8iJTYZmbXYYbEo
qqBrktFmLs4At4X5TBh5cVShotamBkuaimmDVZclvrgfm4Hwykc47CV2Drm8X4rI
JjZY2DitowjnDqW3CRPG2C17Q3B3nqOuBGjDIrp3uXlHrVNpzfzMjB3gu5yhoihG
A2OLUtPg4ggmaaXz1fCH28OuhMIBv+agk54e3/06uZ5bBRrHYDSzGWb+Gh8gs8O/
FxtqUBmkVIu2Qhpsej+zSqwabBfRX12UjYgOvDkplP+NgopQui1MgZp7OzYKvwKg
BMGPewUkCBOJ0ZbfMhSokKHSbJsNxoKkLzUmvWclYjABfAR67jESpTnr92psAfOj
jwj723DPV6UTPZdFjwCGt/TDcjwVvTMkO0pv4W5NwTUMgZ+HojVhwpC5Ebav+mQP
gHinNWzfAFqbVh3pFFiELmiGTOh87xlZFNs3/m1HpignrHdkVu/+FnDjdcAPcMS+
DmLzrCudYdPwUUHUrpdPrac1YfAtL1G+3xVQtiweLhWNnhc8sBTQuZ+hUMT68fBg
4qiEDh6J9oDOPZjIt0j8lQFcgtKHh/lnVKGgIs9jo0770wYR3o5c496WbEP764Gu
L5iiG6sRYbWYyKY/2/JSvinkQIAVauMkoiL4pcBs/wNU+Z42OJbPRljwkd41vvW6
6Wrvy1DrgRBzgrnYhixQ5OPFBPaazebXkB28eXQOOBvh2t0R13mOd6JPwpZRG1Bn
7X0us1KSUcGMGx+iknXIkcxshq0c/BTMxAbjIIzFUejhMmV9b8IpK9rHZbp9aoCC
5xYcYfrqz9wbJhoBOjksw60T3B3yR/liYt5tT/A4C9svq5YxBIMVdM50IQrQrYAQ
cCHWFsur//jUos/dRZchO5Km0u99cEjKPA4XpMw48n+NXPnE8cGwyTNFCuUlCWcr
tHIo9m7lmw8orUp7OuzHxO3bPlIDSI6yTvSJVKYjy5IG6vlOFHRT3M1oCTPn73LV
PS1/fY0AVmq3Hy9ls4a1rtLaDuAc8l9Ag7kOprB6Y+oUShWctSVEMz+/K3krMkf+
eQPCuzpwg06vEGPdIBn/lsY55pQHfCQa/0a2Ku0OBMPSS2NFRFkcyEwmhKYzz/FZ
NM7CjhTYPgmgSr7Hpd2FaGywP9zjzhVLaL46E2wdDxfSqEsWaRcggZeXIdK3Wy/D
2d9vI62Rue/nFbHNRPPPVFLw4e5dQZLxyuCVXZ0Pnz3ZqcY/ETD0wkm7IutLcy2t
job+3GTNuhKIBlg9KcgMUIojCL9yU738N/gFItOwVEu6TXBmGqXct56iOBbmW43z
+6YJXArq1TorAMaxWNgz38pM6i961ESI22mWz3YZ6ZpEEFZTdQ1cpU+G/iKt4jRy
MZnYbxntQRHp7Ft49bzZV1b4f/QwuSBo2NswegvHz2vqt7IXr8jWm05z3cZugCVn
ayOKOTjrnMXlz9Ygaro4+WWnh52rtdIg4DuN/dRteqQeMLh7S27Nchh5GQY5NCy8
0OKyR6QzUtiWE+Szcp49VVWMpO3TxYBLHABRBhfi+d6r4Yn29xVuMU3Unb6zGKo5
ltyHwplrIXMwhdwX7gEaTzX9VzQ6uvOf91TyhjYGJltRAfpds4ZRZv6M9WnYeyGo
2OLdnwk9gHOiCJBSiZuVont8pfPRpcDSA8kA0tYIgvVUgqfpAcQXkX7m6W/swJdO
insdra92k2URwhktFR3iNprz3J6IHQpf5xI9K4m7YVndo3V4oeZJsgSbvVkwPEca
ZM7ynf0/wTFxbTiZZ3zpRImCAzbOI4jvfOhN/30sXv9imQia6Xx8DMVARqTa8cec
zXe5/DZdmuONnq7XtmwnZzRsIW/tS8xOjv0rCemxuP683BAnum1ZtIX9VbLvlsKP
TSoCP4lIUzRTmu1vyqDwRw31J1Ifa22kGVtfWp8N3RYUzEsMpv/Fte/FXp+ei/oY
x/QtcxkDGkP5MOzvQZcAuR6XdiY/vR9/3g9XwrXoB66hhKmcH4ExxWIJ0SIr/enX
O/xvkh6rZPBCTwztGeRl1h6CMdRvrGvpbqnrqGQssTYzKg2FwsL1o9be3Ch8cHsk
WWX5tCO6gIQZGU9QHXk6mjrVH9Jyfd61e34qCEZ4cvwKUsArFXkIRVPT3YmJ1bh6
m9cdjazFeIqcRGjJ0S6jwZDeYCKjfNStKVSaY+a3KeYmYtgg7+MP1CvBZfaPcLci
UtxNDO4B4xnlJ1OSHU8/ZtaeTiazos24tXHl+V9uqaycYq16uhWCXmhbPX4Kxks2
vq2T/XCcLVICTOC7ZBkws1Ji8S73CRFY/6++Y0BRFO9LRRUQ2y7v61IaEho6mR0I
ZHCFWhWeM9QeC6rkN4bNCQ6iDyJHHBGdY4rHSMaikXNbDmlhzxk7l6bEjVScDnbO
60iR/5D4yQ4FCa7aOcn1BMHrBk8qm0Lvy08MwbcBgK/IhaO6jiHp4to9HzR41bEm
v4+aG9wV9g2GftoL9qwTkV0hvEbPNHVPmCLYosTTJ2B1lqldaJVCdg5tcBu0ENoN
b+bTgndNUBeF1VAOgGLtKCQ2zlp6wryRSoryoM5RQ6cU1TikFhf9iOH9PJ08/hjw
/gnuSGGPWN2cVFMl1ZSUBsr8wRnaMNsVlDDRvlzmo9g4d5OyjEVRvmsGBFR7qe2K
Pg2dIq/Bbwj4TMSxTRyYBSlgbSA2c0pm7DYNFC+DKmVUAlumeJBm4EehINBVmd89
lFLvL+i5NYgFDEK4PFpzl5fm7lsBeKLu7OtgZAcTjzuVHJPHXhzXGV85ABaFOMcs
+xfbhATbKGjntYzH+09V0jpzsslfRmEeW5wpMBRerzLLrgQZDnEViUFOchCZXc65
dfJPFr7NC9xp/pcZLnpH5J1VjuChGEotbYPNNXfCYsK3URNK/4Cvga4B8DHkeVZc
f/DuYjUZk5dp5i9gIRCT4zWESRlnqWI6CDXCHf6U6ise7z0Yr+gZySFtC2OYMyB7
bXvKNZVZOjhi9SW6cbNiHIlvmpdRylQy9EGs5TxiAL7KWGPPOgI48b3DfsZh06RJ
8eWfNvqDQhH6jhHXCky76IqCKR61rmaVCa7XyUgSq8DvL8nuM3pg1evmuk4pZbvI
uwtxPB4oB0pFUtPWClzGqWxIwV06/+AuWcY2j+GC7oGw6V21gVsj98UkdmiPCCNS
b0MSxRtG+PHMV59AXfK0YoL49opn1o6Auuhc/XaVoZKhMxthwvu8ccTgWgZclvNI
zWYeaFsFhupeQIEvZAXxCSRPTsEdA+1Hc/lGUsu0H7qu3dNYEzh14wtGLKQ8zpqb
/3VE/woGyzo+QRISPbA8Ctd8raHIt/KDYZr6jmkciUsL4Y4Mk4sQ+/vVFAA+huVh
kvCxWb+UK0Oi/Idiyj8rV895zf39WgJa9bSM0UGFuPM6/PtdXSgD3uDpjIkEVk3w
2ZUxnkeBBdD/T58kvvBlKApJuqQob5Pfls7ekNfQpHEM/jjVEaftbpdsQgMoc1zY
RrFXQIJEgw90B+YqU8wWCsBE20S4OHd6L/7zW19tst/81MWF0Zv75buUYlKeuS1L
RQ+n0AAocloTsk4BMLPfy9T5xaCC6J+5/ekj3yUepWxcVUq0qJwZiLMfX6WXOBMv
N4KxoZ+ds+PLED/Lh88k3a1XNMBAez2WfGpFmnBM/RUIBVBtbkKBqozOpE4qB9x9
FsTgqCGakXgzysq47x3GxuyQltlqNg9X+zb0ySS+BymGG0fA91olNVKGPzTRbCfS
XvsrS0MT6gse6hPuAmta+AW0jwpOEas+RbUjfDsmwyZC+fdu76hdgOmbYXvGdjoL
NWkC6NsROcEc++P0AeK5EtFtHKgDJEpPPQ3RBPlyiNjZe9nuDSyeFXMHuZ7/s76o
l+RdPBbI31EevMjOPySLVTzWI1TE8SwyOJ+URFsoyP1ftA6i61pBRq4Dv15GqbfU
vEZDCzlGWVeXTktc+LGZ86kGKmMelno+7BUp5vBmx9rHijacF6wbCQjYVjVy4Imr
21KDIfaEOrDzCiQpKn2Dtdk76wvfjeEVm/gH140lxCssRN2gfgSMw47IFgkB+9YI
t8itJOfTKC+1HYfhPm+PLlm2ktVzCHNGWlVMt8KyZ+Iua4Y2np9xvlc3OtDY4rKK
UftK//dB7ml3NCnCudKEBj9oB2Oy/tPucc9OnZC/imF0d2MxHr/6Tynesjxn310r
8IualzvIrFYvB6x+7eD2G0KpFzaXTqD8ZprrplHq7PKbr0iBzNDPvO2y5kmCEcs5
AK5mCUd42Wq3ljzXowSeUx9vo9TkWf+TE/3fY8Yi84JwtzWkfY28wkGMu+81LfTl
W0tIHVLfgN0jY4ElyXXXXGDjWGzd6aelrftFwaXA/482ETiaWenJDZJ18AZBu4PS
e1LSKsGBequsebWMZ68vaC7GZgSvsxld7r3v6wgEdBEw96RuZJDDboCwpigN5eWO
2BVHI27ZxHbuqC0Ac79HH+TvwBObaQu2mVhQTxhoiwJurm/GpZle/y68j4Y8xGEB
NuW8qnCoAGNnQoVrBSgiVS1Oqp0cOBpT+d9c02vmPysJmQmLGvwt/T2ho57EEV2H
3CFA3W8dBNsg52E3g2032Ma4MA6ojtLuMkiHlAyy0D2bymiI62U7V3igkja0e6mu
x8CdoVtRKF5bQLCaLcsOALBJTFjQmEZs1mHPd9Bqpaio9fNGD0iIVj/mJ76nNCqi
3ne95+rxrML5IuT5WC/uJYdbfp2NNILHrqtmBfAtEmgCD62p1jm9d/CgesU94lW7
dkTVexkcDs7lqgolEPfVfjsVyC8GTXL1gVAY5o1Vxdfbtq/zX7sINKthKbq3UWGe
qAAP6ddQdbBmr+4EJX5Gf322Wv9V4c6vnENicSJP0P7vW9A94SUoK/QA8r65b/68
7Y6dgX1bTfrKEAaK8h19jsrvCqYycpkELtczuLNus5b2PvE6bon6IN9cor8f6lIF
gIU3ztnWRW58Y5heNRbl9FJ/STM6Y12olfuhIxDdsNZkD/mZJA9hwnK6FtU9uzQo
IdY7amC3FazAtY2D7JwAOIjj/y8zFItEMQGbBobrtUc2CH5CA/zzMTomCGtemX5I
POZyjRSBqqXNGEPBAFfeUSAozW8nV9siFEeIYryCqriS/o4qQ8LVZWV4/Axb69f8
2M4EId/1qEtcgB4ljywPN6jz1W38Ngv8dunYSoWLlrVZ6IRP2jzpjY7VHddhB16Q
VZ11ku6t88Xn8GuhONKa2yD4Mnh7hyejc4isBvaBiNdC37OfB4O6hxjl0x2G9Fsr
7ihQePgdU0W+9dVvdbj5PRvON7gEq9bRhqXCQx4gaIxpoUSMoEW3rfbA2cqakSyY
AwqM9e5EmiUX5GEq7rxZG2CH8k4x5BeIYJ7RwvKQFFvdWWWeVSkO7kUZuFqwbTNA
FXhzcgZiAuCxz6zxQOv/y2nSuIRQ15GkXwqlixLrWRjjrgUNBeXUj6ijKf5jJEQk
hgOnpHvX9cxP0Nj7QRCCIrDmN3exvWhA/VbHw4K0YTwl2LiBxuFvQvTFbIHV6BOi
JftmZXLWNtdn578TWnTQPdBb+/nK9qona4EMg1EiL+oWoAcNU3yBYT/SN8LM8RCe
qrpEE9flnNp2BcEIgogt4y3/zQP7RPTK9Tkvg3C1/RGsAwSkWF+ZE3GoIfvr2CQx
W/7nfw02QLvDGUwmpNs+/m/NtjUACjMrjgZf8R1pXmMG+sZTedP4o/bglZHX6jXA
0LoVHzrtFG6TQ9dr9n15xwEJXF74T/AzmC/UKBe0m4rE6KcWXmQZkgKhqfjqcGiK
zs+fYBAQfs1LCyHtsSgBHfEHZtW1UiAM6gRUQEuUHrXpwzrnbdpBYASjHSZIaDW7
xP82jJ+xuJ7jQCpGsckNQfC+P6cLXaFxajNJRpEEHtYiJI3q4TTEIOWyxo+LOHGb
zRusP/iBnKLwwukvz2n2ag+P9zDRMZ1qULcmZpCjYu2fOhy3+iZDr4yc+qFiMKfN
2gmEwCLanFcGlhOI+x4r/YymVOfEtT3kipIBoQDUYCB7YzMkEoyCevYGkdpXkm8j
5EonVLzdTgDS/wlkF1UlK7RBu9MtYP+gaJVAdbRtKim+5qAuOE9oXqIJ27UQd5Us
ttd7liEHposFpAksmfccUKzjN78i5WHwjpjZ29/bnj1ORaUVa5c0tgIYUmIjaO/w
TXlqlodiomjM94PJM1162dDdm4x1/vao229RXWYHrKtusteHgGTCilNXzGOtGiF+
SrpCASP9WjkI305QEXHSkkcsdWlGzkvL5ZtjEQHOSSY5tHIPEQS9Ksyqi6rvD64D
pw9peJQKlqq59aoMSu3phov+TdIFpnoeJZtCLrsXqrz5isUeZ+yrFz+/5wkprkoo
710FrwS2znzI0UBGF1oY2JkQ+35497J7mzaqvcuwM4ebuLcStH4HSv6Trxt4ocy+
jHflZTuudemDa7FgbnIpP7as5icu2Vc8CYz/Vnpa49AazXjvtGBVW4+TezFk8/Qp
Bz/IcErkNC4b/f4iTp+jWlEDPTV77T8bIw95QkymAncs8adM0Gx3s3El1xbkWnwz
MCm142FbBy8FDqsD2AGrHIuzSuiXXOmebViYz66gtmY7PbSGx1QCyCeOCYiZ6fYm
7h6mpmgxTZkZLnIETTs++s2XVfoMyFDS63XkmYZJoJyMpMBEO1HJxAUUQbAxrigN
RFZXUmyHVsdTcSv7IzDjD6QXzaaCMMrl/bQx+gHACr4CrESpFatXw0Qln6uoQ72T
1qRXaJN/AbEPpO/HrgQqreuZHb8taHfmCb0/6qxfFl/Kwk9S7aEkRGLs7L0H08AC
RLoCawaMCUBySPyKlSHugrtZxp0ZVFR1jrXLYq9+B9ZaLOQR9VI+UCMTQnPJkjJS
v7aAy4u5AZ86owmF+CS9sLwKG7uMxpe8WoHiv7X2Q9YDAnrTqzTQUp/C9fe6cCB4
MYqQUId2DszEhu3kjlGnaKRzglifff7UKkfoEizlCcGY9oooxQ9+nQ6sJRqMjjZn
MizSR4FFb1kv2gs2TXu2vbXlTYv+H1qx6HeZ0ZN7M8bEGFLo5/l83qv+qXK0J2j9
XXsklixMyUAUX1EmGH0V4/JHmUaDEpET86iuQT/bHRibk0JY76LDCSuMEPlBH5KI
zfTTK3pjw8bVryEYM6h0OVj/4sEvdwGlWPUEJad+JiOM3dB/bsC9aFufBomjGrGZ
OPxbW0Mp8KxkJgUNeTs/cO4iD9w6UalWmsbJ9Hx243wTDH9ZzEk5xuvQPerVxS9t
iUBah8XIodjumfysR+mCOmq0mbf7r8emfkDIHpZEepWXoc1pNa26VhyYPpWT3KcX
RC2xltaEPgmn21bChPV0UgVa1k2TYW4LdHWZZO6gz4WpggT/tW0rssCvkQcUXYji
ITgYHwPO/h9p4c2K427rz2La8MhasovSwUfeB1sNJeWhvzINmgfpLCg9ZFB/nbr/
eJE7hOSwzx8gcBc1F4hvuilv9+YVnKn5ZW9Zgeydn5LwX2qPlc4fUy5F6Wy+Auid
2eJkUGf1XjnYMDPZbCKdqyM3mjQtoD6UGCsOnJLNYj3zX2Tm3U+zNj2Pa+EEU0Ju
5PPGwtUF4R72b3zXSHIUP1b4AkOLfG+2aSHFwOk7q1I9h4DlfCRY2M6Mi0qdxdtX
05+j399Txh/FNmCtCPTWS7zuro5VtovaEPLuc7GBJC3teoV4hpEyqa7tb1NNao+q
/HETgKCOloGAwswhrqXMPxkfjS5RYXDHc42cdVeOJn8E3EPaRk4In7p69GiO3HhQ
dO+JgkGTNPPizNk/gjqEIumNcVwZysLhwNP9HlpPWLDQ5rhEDekBU0I3PqgAsJmF
d4vf2Rz8dpm5iB2CktuQtDgWDr4DalWLmzAXvQ4C0pDLe6iG2StuFZb6vy/EzFKD
tE3cwvfOg4zQ426Fw1O8HzGpmC2Nb0a9OLR/AVGvmRKkaX2JCjMYvd4GJScRmzCx
yrRPoNNveaemVeY0xuB9c645uRNfeo4rh4OfAb5OmFecu3/wzekNXjRleqGW4XwU
9rRVLsIQri0SnhUDzE/uxKKB+qq0+3aoxbBszoAximDsJcOBbiZAvkpE9Wa1adaV
XjTLNTPrOFXCy7bw2Jk6G9AWr8S4xKxtFSEKny2eQez79xmJwyCFfn1k776pQp5c
8cZYHD/b0JDjHraarSN67rvpuAmpTG1TeDdoNp6WrCyYObN8Zh0u+sqdextw7T65
/qZLC0X+4IWVSYjMEnPkH56yDxPXLXERJctK0hp19OGKzehrQRtwSB/zqI0a9YeY
D+DgT7u4HzHauNss7ERKgUkvkbNKTmW8Jiy8GPite3Eyb2OtViy4/TynyUeO4hQp
7eGbelqan1MgLD4IFooD9KQxNFSHVRir+DTMHlS4IZAtWwF43m7GwFxujblterxl
F8yfhmH3LFpol+XLVFMdb6wRTuu1+1pncrTOE4NcDdEXEcd5X/jdaf6iwO3cGrSy
WG1Hiz12hhOf2H/P6iFTBkrkBpYtHXBh9fNRxhABDB7UGOd83c3xAqNJ/p9mn9fh
yVwYtnq6EbNfamshwt2fcYDTZTW+ao/pMGKoGx7HWMh4EcHwBisABo51/TLHlHgN
0p3Mj+npke10hMtH7O39wjmm2Iun7GJbxyBmpFrMhdEGPVE3N/Xh/Oj8KX6Ton3/
EZuEpnBKGrf9mUGwprMHo12Cg+5NEMK3RI7AjXn2IrfbXpyaP24Eq9O5rRVGzsgM
nbZl6Z6Zaqe6JuKNiGU7u4Wp26fMSJh9M5j/AdPyvCIu5mdkUlMQsxeH3yqim/gR
tK29jG4Sw/XKlBGrEMbGV/8MhJtzbRPSsR/5ZOcx5wUiJBBNrSYFmnFqpu4Njqlx
0lBV7ij5jl25yXD4e3PyzI/b4oAZBI/4PFvn0Oo7ch1bEyvqrUT6CHSI0AEq0UuZ
XWohvmWH0swSIPbYV8c1XhO6lg/xKeYdUYo2XnA2rROL5E7UPgWXp3bhVxHlWANw
HkG9gYBH+H3to6zy2gHY4fAkwKJI1+g99yzhxFog+TgRoVDe9BlnRMBGQZzkj71i
JKLjgPuVjmu7p7CGbKGNmN+FxT6jRNm/uHLf283SYcmx5qDPj1Zyc+KwTk6aTbWe
2hWPbwYYdAzQw8ucUlKE6JxPNKEJmgY6SB94ZJ+h+rnLWTW2FtcSGSgJDYaPNMC3
aZnmNc01k7pdLpVZX8H3goy+SxWGMEVqqKF87TOCGvf1QS6BnwVSm3L9cumFvGtn
tk+loPN0iAzkyldGyLTIiGTvoyoqdkTYamGOh9QdAqa7ToghzO3Uc94uplqW8FVB
UTFcHCQlpxiZWwCMNdCW+3bhontmdBjDI5GRuskTPtqX1f2JRUqyBJrX3Fx0n+3t
kEqQZrFq1v2ltoLd493jzeP2bUYCsuPBC8frzOEh9srY6dW48ZDckePDNHktAqPn
phwj88otRe2kB0z56ZSTtGYuDDLIVHlTPEZfxB3yFEtJH4fhtq0Q3zwq8filPtPt
ccrDemmenCsu7rcrvbKThUiGgMSnl/ou5Kksrm0E4wsnYqhcz1VNp777dr9D0zo2
lgNoI6vTRnPCUYhSVEbUrHbT+4RbJvmypBzZSf0EaMv6El2Ar/ivp3yLpNP2i0eL
H5/ckvPiqiyFXicwYHfNwqUcv/gv3hs2JKmoGnAV6I32rbabStBxCL2jRL/0Zupr
dukoWO8CiHmWoXdasgLYhrrANLu3chudxhFuYQvzfK7HAMRf6ePqEGV999G1gsYD
PVAnSmUW19xzah5WjtgdzCV8KoOwyaedlVJMUCDP/cuvwcdKAMfQdMkL6CTHf+cz
edOt7+LySDhL7CWHQMb1zZ5blD7m4nYmYFH2bAvLbqlO5/TjYEpBRVz/qlB4nCDV
aSrAD7qY/KT6Xp72cQsBz+lwH1Tyi/jNhZqGbac5KmtjQx2vMkdIVQyHKlVSL5at
CN09G643Ee8cA2e0IFNME9iLFNJuORIjzw+vjWkkpxCIEtfjgr/Tcg/HAWWmhB/A
pObI4nUAImLQ4Zd9WJhQDFLnujhorbzC9UD7ZKF5yKUrnqOreNKzGgzad7Z+1sw/
ChPBfT5wgOLiuYV2rDTWtLOrP7GG9E74mXzqK4o+xm3lMihra0Z09BQO+Nb4tvGv
adugv9cLxy0GC97+L5rc3DXFOAGIk2TsWu9CGLgL0JlNsoUVqZsZbOILvUX4MWYe
BjuVvUZ8cLGETP3hdfCNr075pPw50VmMG2krUBn4Wx6FfiwubQNbN5vFB2XVsxX2
iIJT3wJ13CjI0a312TvEwxV/Omm1IbD8UabMWzvkGEnfdvAHaJK5GSm6ELt/V9Gi
k87CQ2DqEOHZmXjn/9y8JUFruDFH40pp2lWOqL0+qjXeXlV1zvdnVuqMZ0j0gVlz
XKteXE+0QfvaaDNGFh6OlEzPJGVRIJrV+ney4qOusn3ZYqBKzpbkDkA/8CgMN1EO
bt0Z681owSBqY1fWfqYmdxZA1o2m3dk+CPdtbRrZ+Yy6eWdhpwPxyUsgWotfUiDN
HcoxhvhcqUOY4gjcDfpHTFfBjsui3++L7trgF9K5VRWVH03HoA+nBQUKAw8+hnIg
Q6pT8QYYWvP1LkomTzsAYlX6Hm/yx365SIdwwWpmmZjZaZup3NpEPQZ13L0RbMdg
qlfdcc9lW8cxqufWT/CWTSQtLdRzBo9EewWJi6iMk3BHLaKbWWkw5mepMoWlwMhk
Et5FMEjfahosaKZMo0hHAWDmCLsWpxTOCLNMuDzjHvXV3EMdw/eAVYwMnq0gW/us
CeE9Z/1RC2pv6sBnVefoKWyIZY0turhk/QtSPlVmlbuszeosbmrovJBoEN6npWWN
ru01frXnEWdcWe5a/A4fRyislkPkNDKaGvFutV6BmvZWkiUPrAz2WinryeRNvyUN
UKtM3YnuPPf2fBg1B/7+F24hKFsipolRsDljz0wCRbKXEKZ3HwRief//Re7z+VXw
P7zWjtnSP9/KNCIJ5G/+S4b8gtp3RtjwAkSqckzSSPDOu0ay4lKyEYPucTcMCrMW
O81ak8KLcGI+DpOoa0sHAxiZSx10AJK6m3vCeyfE0T/eQl8tGwcLXnlenxrrqe1J
5f8M6lHgTdhSqPn869RZopxL1PPHQH3okabZchN1uSz/DDKb6hYGcZRwoJlxQMCl
nPfiUnTVAd+X7wznTCxs8QkTuiWbfpCvdUkUa79VTMndVRAqCXnRa12AYjFQXOPL
iQ/YPjv6ydXp+fv+npRuJouV8jmDiF/l2UBuqjzh/93qRa9zdqARSfJQuB16hbJz
0EyXZU+LLktKeVSL0X/IIe19VYdcitYP7g8GWcf7aVFFjnSbJ4ziWe6vOxi156Zz
TNEN12iSO0oLQK9TRhvWlSRaZtZo+r5LOS+HFbA9hjgFEAkTh/6SnFtIYcYJVP+1
71SWf38/UKA6wZnaiXTSRQD5yRJHsuOGnK06WmfruCnNIn13rrAItszgGzBD3zjm
kCfh0hbmBram6pdL4Qrx5LO+F/OWxvE/VrwD5dWe/2gBhJRqc3uxyW0/rFequSwW
F1ZPSLbBkNI7EXpboxI7nScvczIK7P8lWDLnwSYkTFTClqn7/9xGQdUkk2h0bVfY
68taoQuLQ1pfLoH9qD8EOfK9L/1rf7njlOBjLwmBMdoTzyKG/9HP62WXnIJhBBrT
X1QgYz53jiJ2+8cCUiTKfvVh+ZaO/Qm8lmSnf0KQMjQPVHpIcqsHX0cH/QDcipv0
RVl9Ls2RRq0BmDz1l6AfeJhgXDhdqjssIQwxDksbw9y1nOTA/iEu5bu+ykTpxYbQ
9PxrQ9JFdgIHsd7J07h80VhcZ0LofR8ASEnO2Ue/rVqa2HUpH7NoxIIV8dj16iO5
LxkMkL+uq/rQanLpYdp1qlpBYMfEomKEiL3XlC2R3hLqbBI+z0IofXiMEifaltpp
4AjmfCofs4lAT09iFIRVgGomK9VQcimUwmKUwR9iNUNROkGxUa7i116pa7V4du0/
ak7YL8Cu5mW/MmXSlE1TBWTkVwOX4NOKIKqUs5iwW6ZyHj/Rkrnbn7kpUZlA8jr0
msyE7JigPefDidfAZrCRrqnf+XFQ+zcQsW1lEqPYyeaoJdh6GJJD7fWXpDITVb8j
2U8At/YgcRB3WC2U121J3VnB7Xd9wjskR6D+AMqqGYKwvZVYGQZdaQJW5Ylzzjjz
Vu0THvZA9sz5EXUDE6muGjPDqqb+L1Tg1/OxCJ1pHLYclfI4Y885zw4S/xR0RQBx
ETBYRBbvskh6lXNplaBF+H9KKuFDeQUCcMHM1kTtgrBTNa5wKmhiX8H7omtGwFcQ
j7gYxQhb0ZTNfXisZA6Q9+ooXoxcz2ugpZtLhAcxKj3CVzrauZNvS8PIsYAJbcgS
QVLqjYGIztQxX/23QwDjvuidmVvOaif8M2ALQb13LnTYpLSb+2S/mneUJ1OkIbww
ev0QSKX2HIu3DQzgQXbZDkkkm2w46jDmt7d0+8ceXpuEckyZdeSHkAuRSLTIy4ox
lX4nntOD0W0+jn3FTYDPeUhNCksIPG+ddZNAy7fB4/+DcJnpYiMg6TbJptWlIgIs
UirdqowQMoxgfwfN0ebnBLseor5EIWyPG+lpwUO4qmFU9YoMpzKip/LHqTquRTXJ
dDTvyrW0XkbgWZUCYgOeKMd4WIP8VGEwAd7roh/Ij85MiewFLoV/MlRuXH6awLV7
RJamDGJ7GOZRibGjNidH1YU6bL68Deq42qyDz/YTATtxkjwDwGk5YXtPW9ia9don
8YJQa2lq/NLWPKhDoixFyX5UiUI1pabdz9ZCBYA6KFtnq8EZvrdB51INnPMLmphk
nKtk/oQ1ZQt3nQq9N32i1COisVVFVDKVB3rjgxqCPOAXsvOVndaJ4IjoZM8VqruL
cQInmYEluGcT2BAWKT4fRiOvmv4E/vnB2V9qIez4TXV6vGIDYmQfUzZH6h4fJWky
ivLVz8k1DgXqhAY0o0v+v5iq5z+PRcmRley5WWyAjBcnJ9Cz+K0xgFfgVMD5Jb8A
BA11+0rf+a+v1FobeeSIFGmjMCHZYQNBk27vsr8YFZhAxO9EHFyZhRBGNoOmpupk
hH/vQrg+qLPduk2D17Dt+cFkApXyXaWYpW3/8unywfVWB3yo/+/zHIPYLBYhl8bQ
8CKXSpHeLhqud6lVKD4FI+o0r/pgk/ApVru4r8MdzzdTBlXXVrvaO0SlZbd9XcMH
45tEhcwSfzafrodgSWwdhgEez62INl7TNBnnpc6ftYJuU6PsA6Cfj4dh+H0LGj+K
JhWbO/g7ziLgdDtWfrR2gcjJPo2Uq95CSMMv2NLY+7MJnuTlYWOzEdhmWWHunhOf
nZkCktHkBiJUMcQv9Td76U/2hZe0GbGX5WMs2lLw+YUm23w+2Qhs2OkY1/tHkASx
w7S4iXMEITXR+D415qWYxb9xcrT0ZItYPrgshboAQggb9f+wq2aoU4MaT7k30I8a
Z6bz7t/vOqQkFXLBZK/mq/oAu87en4oX/AOO7qJnPnWG8HAm6Jd/H0f64qN5w5O5
6jLWVd92QHgjMgD02/zTqW+CjonqnCmpG//NQ7DY/9HPr5vmk6ZejdX5w9wOAsb2
c0tEi75/SDh/huUdrIc4kl9TKyF+ELUBQyfABQjfVGbZ6Fp4TyeiaSniAkFK40c+
UVlj+s48PaJXgQylPmFY4H6D2FuwlXbFLp7/GkGOBhIW0dr8Snwrjytr/LiIJp6E
g1MDZEWSjwC84od0wsnN9i6of/QpuW4T9QNpcZ+kn/Fsz1jicjKuZLjQ7GNEjUXD
VUa9SigAh6egBP4r9j6Lj6xwHxlrhk8ca78I7KG+UDES3cyW4e/UM4TZj9sNSWj/
a1ZVQ7fXIGuGb60L13cLhQDIlFRitFwa1WJdgW4ZMRstO9q8OfhUZ4id7C4A56Z+
YgU5Pu9Ucwig7kOU/MA82y++n+eJj3+3tZSkMTqxEF8NbuXkwhXxq/hc73RJFxhU
ZRYxXKoitO9VKve90EhKyv0hOF0bAkp7DB/SfvGbBicfs4wl7KMlBidIZriSq2ed
lIriGDcjJ7uZdKpeE2VcycXWoPcAEv8FHcXGrjFMjKcNQkdxiscQGsW4mEOimYsi
rKz6nb5dD7Y1Y9nI0pfxOG72sZQEsfURXkWs4yX0+oJjSoWT7tgUmkuZoYst00CE
SrtTptXOMUroy1Mr8P6kAGVqU74VxSXPHWhOWgxlC/HPv/z2wI60ZPZxVflAy0C7
kd7nSWv37wxXEhTjtN5g6uOg8g/ELxxFdHfP9ZzcQGEUzWf56lbSyzOiv/K+gcke
vW08+aF7KaBbcOIL8iSiN2EZJPVRJjhKuodnUYI6XEMqy7RoSYDynBBZEESnsoq3
YakOEHe0YSyj55gVlLn3s7JgFkpaEYNgX1SKyRQ8/Rd9IZL8J/N5ZLb37Fuxn9yl
TvxT+GwiwFVwdTl9mGofsfs6XAsbxPxMWlPa5ERLYm0KkCeRwThm71GJt+0WG0Dq
8Rq+uX7oCltKWaXwdizQ1v2/LxF/1UNullSm6TVsff4Uu/geQndyr3T6oc3P8djK
WFranxkaEyRSTGPEkIpQlP8dCggCAgRA8sdHMI/SNZDj3Eqs/U3fNd7ZWMb9p6k+
5lZOPXtnI+tYA2k9vtbJ5CKHG9pDQrxxNDNkzx7roOavqGesSM9V+3Kx2oj5bP+6
UnxSvLxxqdXLm9zMoep85iI1MWPKvk9Mp2pLPas8f655hXJAy0kfBbb2icFsK54n
8mBgQb0Me6TvqtpjQZtgEWCExvdTX52hmxIaxzQfsGtkQc4NGeyKUyKrWImoCa17
dZYBtozR5UFFr62oLUPQ6ClhZpfQeGMj6CeSzMO8X+ihtXyuty5cMUmbj/D8MTv4
VxrRXS22OfioSQPpcRZSzXYLJ5UmQFgH0ksNskpP0BtLhNO3yHPlVRUTsfX2TqES
bogr7+GBqjotoQXP4ftZqCu4m93oNrEUEHS/ik/0ikljXBIrI8GmUbnD+4rfgbBJ
8Eo240Rf5zTQip6X7txH+GwnUcwFw0ZgYwqRH/Ydh5rNLX1nJ+QO75ZEyW5mkC6a
Xvom8GUcAYvFpDBu7bB8IQ1D04aY2jTZ1wYhW4yZDCpgl3REueCLth5YESZzaGpm
0jBz8psD7UY++d3wGb5oRb/KWImWJAvfeHEGS3gDNTiEEi1CExKR88v8ZLpqNwhy
9dffYDGXbZl/ha6JsMQkiD6k8lhW0Vo8PoGD0qCmErD8IV+8PM5rf6JJ9wuTAT2S
3ZKu6IJctBmU+a6d3+x68/klRfSMWJc5DzDLOKJYzeQhmtD3WFDgOb7xtevheYlp
JhEKA4Un/39KwnNMIE3osqjrRBuqU2BC3b/DjPmIQc4JQVUb+NvW8ig+wacs0mPp
nDIq+OFP6nJPHHJPUkghHT8BRRto6PuuNMr+KkLm4CpPAzMrDdBYFTLWoZqYuMS5
F2EKDIAQmHdO4C8/E2dWWbGPDNI1+E5JUv5uFQhvXkR4vBz/I+zK0mLgIGW7LJHq
uDEnV0qI1c8OQ6I2hjeEvNk+hT/+++avZZySmyyPh/gEifie4ynxqrCdbHdLfdKy
Lqk/qjzneG0Ajo9jVLmwT4gLqTCnlVJbWvpaDsPs4lOEnR3qT6kqcq0Y/r0qC/fy
rh68dLboGXH6xSruUSJl+CyxTns+VsK16wf4qYJBiINUcpP6r2VE4bKwtfwgKcNS
wsH7EViGy8tSjhkDQXz9Rmy5gSd/dNf48STEEFkGAi4zbI+WHTspTiKUaPS7qaaM
k2VsEK3Hq1IolP0hW31JfUoY6d2jhnqDib0nu3SRdfzM34mjbH/fVuG6/TVRwwEe
dpewgM4e/OQz2OFK8u11Roc+BXtmOkDXneZSTxML2jiotfUjOXGvbXh+TFQnuFnv
BUN+zVSom8Da7ieZEieVaZTa21tpDqBswoCPMpqrFqv7KmLKlAZHc46+Ikh8Byc3
WX4vpAgVIVQW06Oh2GH92EQ9IPhCvdIQmtcPyQ2/HSTRWOSSu7WtEgen32A63rN4
QavMG1ZL2RhRJETM1Y32gSvIup4D/pSrS6QPFvn/9u4P0DiVYt5Z5ndK3Ic6ctXA
bnBDVmCeCKT1W7F1IO9ygcwISZH6CtygKIEgA0U9cVa5c5jkhRB7G6QwWmEHsA3Q
95clWzoAinx1Kov8kvPfJjCzFYhZC4IGf4QFKIULsabaabBLgPyD/GtdRWnV2jD9
RCYBEwRzXnmuQek5Dw0UL6UhemeTWyPx2TjBDJaZBJH8K/2FPdkwoWGWKpOpPMHj
ptSQkWcFVw/3tTBOH6QjqvM3kUFUkX9PPa1NvSFuVP5kZWcHfskQ+fq3hng+epH0
decFf+wE9x+1iw7SOH6Dy+lJno6vOMBRo7bNP6QKToriYRTxzTPyfe0dBD1YK7E3
n4QTBjKjbtIfyvJwf/mpzgB8gFGjPcqVKrSBXeLeAA71O5lnPK4pLiJrDX7USXzd
2DStitz0s5DuY56qMHUAcRD7bUEg8MYFkAbmtS5YPgYmSSHvR4K85nvl1/yIGJ20
kRbj58kld1tKqnVlFjaFKJwsyUEDduuSmjg+D8Epuwrds+YGP3LRQmGHzNHCq3qH
3ihH+nh++z2fLgq0TpuB3uwQzuOnzqzh8agEDE5Ufb9OVpExwmN/42oWpUSVjsOd
1hDf9nmpZ6pW1pF1wMg+fQ==
`pragma protect end_protected
