`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pwQvZugJxJdPT6jWbln41o318m2Mf9RJs/mUclcHXqjMPNoGLPXEr6QM3JMoihHr
ZRzUjN/xPuuGSKTFAhOkBN9uWZM5eUDAjaIGCj8zONssAYIjidXMpk1Ix0jyN3fp
6NV4W0bLskcMXrJ+C6wZH5tJ/eBFoqIvF0fc+R/wVZs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
9J7tvczN+BiOMX8XbYq0QYO4KXP5Ryo3Xpb07VYB7lqf2MCtqCQTpp3X/zhIvEn7
33et+BYiY+rBzvdmvSYZS7iWM4Dslw6BZjO13P2Ev9rOgklY7RUS3cditg1mVchG
+nJWa7O814s1BtJXTXFIijbgUvoGdiPW7GUePPpZDPLwuZQUkVWNtyeeKR44LAXh
gVmBX1Ywn4IdlHy0U3t65kcGHQMNTFo/tg3N4sdUnXL5qgwTZfy7pgtvgQqxUBe9
hlJVOdq5vr/i1oDolilDVY4pXCvtA7ybu49aB496/6tcBidKGoLnvy9nWM0pJxdi
pkW/YM/j+v9NVoTPU3tQHnC+G95s6eoLs5FZQ0SMv1oApuOQqz1537uXTHxuXKDA
alMY3B2ah1K/+m3fjrumWu1/e3YETthC8r8lAqofgj8fkhGxICFYCMhJa4zX3cWG
0eqBXv3WItNfgHfY5xChELRiVUfT25DLzquvP2PnVRk3saHL8LfyGa3+hcT4pOT3
4+Gpzy2ApbSBVycy16OdJD1ea8+uvni3Agn3iNdWR9fXPio8RonX+tvxOrwJerZV
KeMUr3ycBCqafKUXjOTEt+wImVmtN3jsBfIg3gM6KFZbBO+fyeR/zhV98DyV3fvQ
k6RQQOdpNXiAXinBfADkkpp3HdIUHp+XSY8mhnoGvuo7datk29NZremmIdoQVfV1
8eYeuYLVM5YXIN93WGsW/89SgtMHqTaHWkD6w8KwV8ZnEtN+TdrvEM8JC3iYwUbY
vi3DuEp6kfiCyK2n5ZM6trDgsm0sf9V2BdATkGayTCMHE6GBRcqchNuOK1wsHJzI
qiEnp39IwEPIXkLFPKT1oG1jQhWJjzG/K3rVE6i3VnoroqrStwcr998jIpSW4K7Y
1m0jEnPYyhEPtqwjGntf5laxeZFJMR2qT+NOyZ8smhk5UqnNArwr1mFlYWn77S4d
Db/wICGh8tiZIDovx12tZB+i7hQkJS7YK5wWCUtxlCO/IE6r1yLyHtptGCzRtZk9
TaRMD6Sm8KTnSrW9qEHLD01dE1XElfVi6Gr0c/sFkQXXpYU6s+LzUfLcEVhNStMm
cDzzt6fnsdtX/+Xcxl59Hl1qtFMaKltM5JFx/oOPVVKzvnZRmgLscyY+pURnYQDp
F6FyEYfo/1oDLUo8t1edX/oVgS5uGpCrqrwEsXbPuntkl+vNxzu4z/oKFI9qACkL
hm73TVRkf7gG5ZLPB9gKglFZxAvALFHLD4vy4nZy34FiFJsLUvOqblZZqZW3IQG/
jeGmZ6cY6PbpEM24ErE5xVCo0rZ5VQF/HFm9CbTckDisfmw87/TBoVO3qYTffNxg
RO+knaoac1eddZuVIuTfX8Mzbifojht+40bsiy5BOG0OLbnXBkKyjo9lz31V3G5+
NxFir4B3260oE0LWTkJ7bxHJqc92EhGDgrDsvO3l4+zQxy6IPZg6SCURUbVWpWhv
7WAwilY/wuS95HyWWxZkUAnvssZ16/xmtCg5xOWmjILLR3Nt9ibnAAMmq2Wf4gRO
ncwryklY8+GjIEsQdUMZnK5JxMDhbfN4f0mo5mT1R8MZ+sGl8rnW21D7vDW5visA
NuTmAQhM4t1Xt+Ke0jZLpL+TMJr0jzwrwsSFWUC3HsRkeWqNHPOB2vy8UFhqTJqP
8oC5MDgB3KnVE30QFKpD2+hKF+vWskTVYLIybmXzS9C43WW/jz54jbVMl+LmUwPV
CBrFpT6D1X2uNDAHTj1J9YXHWnK32tfwKk4jhqAFQiZlQtCkHZEcW3hlEdELBQdu
lTshBMz5GhXGH9PaqJSwKiKYQJ/hANfpY9Q/xoDHcUlmvqUfgkypu2S//GW06dYd
9shYV8W0ABmUV/qaxTnSNhLys4InpGIBZ+h4VRH5QZ1E1YiSlSyWB4k1PiOX9epv
jqFvIYiQmkx3HSl6zVvq5oBYbL4nmrXPa6u6P0B1sLiwYs2pMj2IaVHqxLqdwZqA
TK6NByIUX2QdlEeiPQIQw4TiwFerXPXcQ8WHFg4TUp5GMftScTYYREgvHIaXWog+
oj3fXU1b6v5woiUtYsFEv/MPlWNpd5eE9wBxz5GRLCZxXbfjadYbhN59rRBoixoh
lFMBRZzFsh5KtCCJfbAG+Io9pWlCsBw8jGVSAOiTaNN6Dv600KgKpSRYq17DfIPu
JbvtJwHTJ6S/AY5YBit6ktxMzcHwEpPjeOotgZIMGO9fjwmWyDGKZ6bOnCt+m5kt
3LhLDkbStDB/KiQ0ZeRm9O0q8thD7V/T1T50ARnGbyg/T2p5er0bNKylMIyeYDom
7r7M/nASRHW3Ft57dq0da/ucT/aP5F/hVvzmecnxKZbwtpRQiMbHfUH/BT8xCq+1
czLjWADnsdSlWbpo179qW5cpKobFsuptVd/UYKiP7Fy8z27IjG5CVDih5zdJK1rL
Bp4pLuZAlqcc6y/0aTUpxbYZpEp6C0lMSNKy6dIBFp0cOcI1WQuub5vOwqSqXIu3
po/AWeiwXCubf4g22iahEfgc9oNhjtLXH9Acvbmc11Yn/iDeQ4hUGXaR7JLnpApJ
exqH2Dcaq5XiVqF2ATZpiJEMgSnQt7CKSFvfkqMVXh1EJj/89QcbfZHjz2DR2qvb
ax8oEd93VJBTNlifmF0cynvcCyvs3byL2Sj2yZmUc8BADaZ7elWyXXWtKKWrQpuK
g8gIyXEKTTFcKI5+OV697XMLsNT0P/oNVKwlcDvKssxOzEcJkXC6RMKmcVAPEX0A
oFO3qLNRmb0za4b2ChQqlQHhoY22hbnM/s87XUm+pCN5BIcAlvnlq0PuNdHDIWpl
1WdYhTczpTo3HIbmMkYNVPH/Akgr1xwmnbou7AiwECs3uXl7MuiYE7YaBdtCwTTr
MExS4pT6erWGIefBLugldV9ocXdyeCPBlicxRj1+7I/bs6dvaibKG4VzAWvlJV5E
t3iODVZcSFbST38Bo4UQOHiO5lmCbshwrwrFyWKeRUx6pgtL6g8PVQ5GJe7MHyUl
6Hnb0NpovB6hGqrL+0GsZ4QKOs0fkdUo7vaa8h+XYXp+IWJAmTuK5w+pUKnhyCwM
rz38xQ6PYT5VRgkwMscOPZ5v1JZGHVxpZufNnkzwjDmgTXBXG95sC5hYlLqZau92
N7iFi8NVndOvg6V1RfWlyOVly2DEYCsQ624wbj43IlgVI4M+ATjO8NfpMWju48Eu
QZ9JUFoN5gL5NT0KMKZkhovMEe1XY272dH4kIWCpppJdReEMf2qezD9waON3rKWH
vMVk8pTTwtYuvvIOiskr2ZH5+htg0ZQopnHYiJwUbOd8wRycGGbOH5+VR0zfpWWd
3SAoEDm4HvlgbjqLtcVdtdY6TXBIMI9TKyVmREPNwbS5pyAQvxV+fabcGN4gkf3T
QQElbxdNluTQFVT4t7ICytkjolWPG7sKqtgHoWy3OpDj4wtpnhAef32Ln5CfWGLD
jXlIfdA5P1hAUAuA5T3VPNFPRcC1I4h5mOtNJTAjKWjZyzrQPKQR/AuqdSkfXELE
uxbWV+cnua5H4KvoloCHJLR0wVoA5nUzbDfyX1Dj0Zr1Xett3xVmCuKkbQCVDtOO
027QjuIHH7/S7VZFVo6GlZx0jnFxXZpfP6RTg0oajhUVQlodaF145PZBUJIEhSgF
Nzl6utwGrpwuLthD/a05+EA6N9IPQWrvdbWEE38NwVUIvRZlM3mQbVfmS9VrDRPs
+/GTFGUPvI8fpiNe+oxoToZq6hrPz+KW70zO7d/kfBU2EjbvJwwiL+kDr0bzJ1xi
NTVpyuIPxhwWyQ9CY7+FevBquQXqFtugAJTh39mFwhWb0OBd6UNLWnTwP6T4EEUC
WfIhtgXX0IRqgj7/t6MVVQMHzSS/YoV8H1i2+wJf/WXTG442hxFeVE3OMbYTNd82
7OpWSlwD/ZFlAH2K0QasyS0V6mAQ3ij+wy0jWj9Ymh/tCx88Gmi2bBH6z8DDBPIG
p2VSwDoUTKjpPx4UwzTxAwgRPx0vd6GqXLIDLpZ/Q124si+6loHUP+dMEzcAg2jm
W0pgj9ufJFu1LEQxuSseCoyxxLhbWjLICbvbojVF8hjMGLjYZlJREsqSObj7AIVG
FjFNZWTZlWm7yrKNgCQXHykGGu7n3Fh9gBuyI+QbD/vBpxZ63hf9p8XLrPKvl9xs
qsufuyotoH1fGwk1oW2AWhsKTnMjNCeCQlGkmn+cJ4K3B4fGfaLwrDpaVoeAW54k
nXsfTZg++M3rS6AUEJzFdJ+4zl7hZeDI2Baj7497oYTumLMf3iwai2njv7lMZf7E
gdjmG+gn8qPuM57MQiSVAirWLOpPgpRYhjDCNUPiUxdtooLw81R/Aiy7hP4Spbmm
zRT0liXcWkwW4LENphDdwA335/XbJrSotZiZq6sreN6nQ31iE5ZYCiMqMQSJ45qU
nowfeeGKf16KPIDDqG/dWopDwypjPdMHpSI4DLGD6J0BFiozONDbS1yo5GJMcoFe
/2OKAEogQnSHc+gbHEp0ycUPH3U/1EgSEG+GtL+5K8CrKX1A1S0o8GU6Hxlvq6Gt
3UIacSssH9m4L9EweO6elQRAEcgIsgZgwwAmRsId+APWMRzraT9q7xFTo0ooKa8V
a/WeSq47leOgi7QqE+PQe0yC6v2sgr85TIRGcpLmaecYG+oDqzHkPvDg/VhkRwSb
uKX7HqXe1CmeB/kmnlqtirkU3RUc5WAQu2utdRUBUxDziR3wABa1mAK866Yl3ozy
QsupDmihv3EOSMRQ6YcZqD6s1rfCjPzoPgSb1nqiNrjdwuERZCzu9paWmZwefbdD
SuXmWGS1vlxjlqJ8d6cPgc43vv+CkZg66BtpLQpxRZ0DmH2wa8PZjtg/mMo3YYA7
zMgeT0SgH3Ig+zYdojbIF+kJaUv9lLa8xUJjt5qst9LooKzS0DBG2e6Fxa303+Tj
8eOkiJPB3lAv0Dc6uSkaMVlWwfmzPzp8rRCJhP2JOiXoDBSzBRpJ3P5ImzLJUFle
h2JVQDusBIxtvMcn/8xWGq7QCzmP0LCjybeEW34E1eZcgfWoKllXv+aQRuM+kiqv
Z6qWaTmFbXkCgiP4+c2li3iBOswvQ78SKBd+P1ULKsPqi0/qdjfYl4AhgQYhW6YN
ewx/uhYpDa7/HI4H1OmbzRFpf2rxMzQAEzSFFx6pElBKiWMT5huhCcw8hE9BaPSx
tkeUfHkt9B474qXOhmUYx2/6Pag5EQArAi0KXH9vwx5Lheqw5HF+0zMF8mxGZFIp
YQjm3fqVq1YOrc4B5CEun6MM3SEYSrSZGonPuk8cYibKINkR8lMaFWMxVittu3w2
c1RhXlQ99crbfD8al40WV/+6n8xtBWcueShj+nedOTzM7bWi3Jiu5txWsDWGItO8
00Ww9gijBc6NLF2dHGbQaBVt1tHFxfrtehF5UXzOhyMvsdVv3yELDjj8zg1pcnEL
k3SEiZU6bD7bEmvkmfXjJbQWbEpvd1BM4bQAvfCvbPsloz8sV2bM7mWJRqNqKT+A
r2bcBvnTOOyltAc6hjSTwfpP74RPbUtXk9BLUW46KoOddSmaBdVbjo4rVePB1hCh
rq/GhwPnFKqS0/vB+KaE3zJCkGbLMAIIYHSDgikw6ci8SHBP+nDAfyDwrUZgcnjq
g5oEBCQPzUHS6jnmMjzLrpNpZ5efWWGXMqSP+J+I3h9irpGUll5aQL8T9O3OLDAm
bQ+vKaeZmhnQbQy7bWmrWMJIZQu2ItqAsfaZvt8uJPyn0kJaye9CLRmga2WZvxkr
NAiZ3btEglQKtjpYD2vflJrooovrwhQcSRHtuPTDGbdj88FGsw8T/gEU4KS0rvfC
Ygdpy963I9/IXeJIx0KvG/AOFfupZMyWpA/sj9zZdbP9DTNptu8ZABE6ajRD4YO7
ctEd+ekWak/fnhNxJI1rUP+wwrufM6Rk6Mmcy1cZ+oFFyugWWrINR3vXjvNrvBLh
EZp75B5QW0L6W1cw39siCgyQ6LUBsesK7ptNIaNl+GF29Iv1GgK2krNFPFSBqJ/d
X6PWTj7PugvdhViVVmYDsWvVwI4BwJwqz1udoKwd3oyUsFq2sblbDQ/xE8LmYy43
XuZHbJ37D4svQ19rr+uP4nvJDP+tIvM6GBiQpTAWt8iRX/4yyt+0byuNjvqkA3Fj
IIpoYpfMa86qk7LXOhCXCUHiTUSylM9K6Cz3p7wzRoldzXBTgzip0B6WwTKg+tQV
5mVSAigjzraCLBaCphtykaS983YSKoUa8v/R3XdzU9JKqSFW+kQpGBKTebKbhMrk
2hP0ifhHVSNwHMo6DPQ0kZwYGHZMqPP+EpHSs1MVeGWca700N1hNzq6hKyz1Ziiv
KGW37Zzn9p3MiEj/Ig5K2aN2HpAamxRqlLxVVerOMVg6JincKcMDxuL8L0aI6NpB
WIm3mnGjMu61nmo0jCxBCz9YcoG0UhmTq1rRckLKvBZ86J/mAYVkXBgT5/eV8WHf
86StE4XGMRfOWvNs6GKin8mtzmZ6sb6kQjqQu9pIBDEB2ZTgFyina2lv26p3Mxnc
Y/5QgeEKVaE9qzBZc65Zfxkz/+UgHeP3wKxL1HW7kz0WDP+dx2qBjQxYkNyBrnnt
lcOYT0OjwPYCuW/yUrfKOTWR8RniTVtdEiGqSVhK1V168GOX+B6SeHlnu0HA0XrI
YmdUerWxXkcUBB269/YBOOaTm3yTfGxnxeVmJ4qYScPyfzlA7qVIrs+yZ6d8xhjQ
UF5GsEQOPaEQ2X6JrEzfbr4Hd5fBR6qAsE3jJtXNktom285jle2lqKm1i+1lQcTl
o4B71kglV2Q0lRL28AU43P0y303hlH30f3X9fQzn18kncz6CIP8sYLeOHJrEFwk+
bVbNTTdkq0+ZnryZJd0mXRHA6/1KutBvhSPQHIPtRZ/0TGL7ASBOt/ocktXF8u5a
B7UA8BdHY4wQVgPYxbvzOUj5jMKrAv//fcFFAhjE2LB4cOYavhirkI2OeyKvR0ZD
VOgL5XytGuclm9M/JaeJssxDhUQlJ60v4YUnGtQWbccy2QWPeC0ADREjWT2jPRz/
y50k++B7SlmiMZERf/VxmrKXqdRkecMrw+evzc2NKoa8a6xSqTILUjo6KWNtT1/z
eVqulIOJYwc4aAXjDbUQcM/4h3wiwEzouMn67pb98EUWZWFlwuZYfInQNkbKn9Vj
vkjluHx7TcDc9Zo6bS2B0n7VcgsRTu12hHPSg03I2m8Ugfj4y2nkhfC0VsspdFNu
XLmEDtdIw6YycZVFXpHMYiPBmZVXtZ/hK2fNpSA5a9AU32RHJ/BQsMEPAMPASHU6
tb6N0D6HzGqLPxoI82CdC1X5/8mSdxHnhFe6G5SwGZmxctKZVYldtdjlvzOb4pvt
MYNET1X+BHZQHof05xxWo/+ZScchbBSXVPbCLzmvV+9r4ypT/Dpw+KZG5R0AK14U
M4FcofjCrSQxAv5DpZvvUvy7+DVtlvz7Idh56QC/kwJgBd6HVcfse34/RK+TIOdo
2M77dh5zzEZd1rMX7xGWKJCtkMfyFG9xVIITX8mXFDsZnIFBNFd0jOiuqOG8ULfq
7IhD27ChjnZeRIVq3etnux/kg+LaXmohaRWUeFWrz0q9PoyF2gSU8riG7tBg0fYc
vKF+pke1BAfITlOAjA+hWONDOAU9cc0rJTZUmcbIwsRntifOPJN2bM/r2DGvxiIw
9l7JpcLLgp9rGaQbrVG4fjIQmlB4Llvz1JCdxV9W552FQq0KGlgJL9eN+P60igR5
tFU9A7wwEmue32kNrgZbRZnnIeX5oxx1KJ6LVCsK6N3nhmXIf9p7e0pSKqxfui80
tygxUsSaTFD0wt4HYNjbceo9Eri1KGESAJchyIvita7/zMvflq3gs9lMRuMKKvP/
bY6CJ+3ZNrZKGFlzX28OkK3PO9WOX5h5Ftm3dJ7grq6zteANIsEqpq7T1S/xmLh+
Xjo1auotC75B+6nhutb2CRbQzhAHI4lr4qT5OJhUSsrXmiHw9JjZFvOaxEzffByf
mtmpqZm3un3GDw/KdoRip7PlHmzzFevu9LBCtcY1C82erLeJd+zJPN6Ep/c7Swy1
q4dt+rVWafmH1QMezK5Qgcq03fuSlNYfLIiMyiXJIv+F4Xwrf3T3z6dd2tS5knB3
lt6/OCDHV5o4z7pLX6y1Br5uJSFNNKQsZykbxTCK0wsyHQeqY1MjA+ui/DhCDfFy
y05LDdB2HlkBDMfkrgD8e8eNQncRU8/HY4iPKepWypqta3xMp94798hv1XEKq1fR
qUucrBx+spPS26jr+X6pexYa3tO0glIXv3kd1c3h9LZAwzlzIvpbJxMr4p+mRceA
YuNWl726bTuCy3cg2reIjjj8/Pb8IwAGhrAVi98JDBJ4NMkcb0sr/J22ABxjbEpU
aHmlx7DUMK9M+mqkenK6VfT7nab3Q8QcHmjV8wlcf5wKU0yCQ43GuUYPFFnAS/nk
sYVoEm+iqoaflhxYZjtSrA6h6kBszKxJBM2UWnpItjF+arzdykR/enFE/DRyVfoD
+jcObt0MTxkmrBtzbNHa5lg5fxhslUR1q0dKliH+dL863DyGL34mTihdaL7x7ttb
1oAuVK1g0Hab04/CQ5ggNMpIorbVeq+R0nRzGdOIQuajp+sm3WScmw0KCXvRV7au
Yt92mUIcONb1/RBn0wl2V/rAfuNRcvtT+GYHPVA+ogjQsxttq8b2GfaMEep672Hg
yzyZ6nP0szPMytYpfHZW1oq2umwPJJAZZdjjSHGhQgcxWVIdkjbKfSQlh2fj4be/
61DFWmkNyOqEwLgnuD82PU5wQMOhIBxbRSJOfxwfy4EAc2IyzwU4Zj2d9C6o+fwq
F5CnorKM3vKCKHTcpZWxtvx9cIFeAGT+ADkJqdFDnQq/FyzKjOPN/tP5nWPJ9jTz
uRBs8M1EPGlS8uI7h2WnIQoBkAeABBa+beYiHv8GB1C8NLPCYAZHiWs0cdWkVppg
m1EAuADvjNhCSdpORyFBBLQKgNXczH8kn+JkgVAS1tssCvu13KFehuNmhGsfmsQJ
E6HhJPu6xREv0TMcB43eJS+GmWRp4RJM3CVPlkNk0oRgYrt61gbhS2hkfStrNkFR
ucItqVIAgWhWNXTD9cktkqKMJOS2HK4rmusQ2q5IIIgLjn7poPtZOyZV38QAUGLJ
4YWoL0Y5uUZfoeU7SVGRWzSLPTG5eVE1oU2Ji2wL6jc3nSvtelFqoYd7ghmSMWgI
7AvTn/LzXGXcfLHVXP+f97QTC3wq5zNx4J6EhcHwNRqzxUAogF7In4RCXL8bha68
9Z9Y/gHqSgHIo4Nkjp7Kb6G5kRbKaB5ixAxXjY8fmsjsS7XcYDBubBHiJyY3lf1h
5BkVDI2ErChejrynTgEJ3vXgY0/F8gtDuiKV9Yui7O73DZYSpyhFOujegU96zYWD
2wW/jHIGW6lqLTSoaVzBMMhNQpq2M2F7zUx1L4wRLEc=
`pragma protect end_protected
