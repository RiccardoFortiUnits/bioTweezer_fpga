-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
snzUgFLTNObLuF2AmeaVMnw7VFAy9lZkBoALYNd4a1ghJ7KWqG93NjvqgaYyBZmeOXggnNDIiDmk
rp9XBGSEdI5gpkTxkZ6Ulpb8EpSGha1PcCIg/YKUUvu2fkY0e73M80kHWaayYXMxSdyaEdLhuZvN
QTpftUL67wpYZk3aE7K3Hv3xof1etPOxQPMI9e7kI0D2L0c25NN6cOKE9fXifruxsKOJPk9sQ/aB
5+LaqclNn2PaWVI1Nvc7252DohhDef+3FftbVnGHn+JF8delms+oLrsnKXIJXL8dFG4ScwJ+1ATR
5SXs3TDpW6FTfhs0ZTi3eMbor3qvtslfFBUITQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
+6VNaW3F1ZEiL8PZccNl4vYzHnL+1TwT4RW+J3XQ1rKMr34dj2Y7+pdQQiwG1ketVl0O3i8Eaeu5
MjYHaf/KBTizsQgMua7ElQcPac8c2uGjhGJ5x0ZKP+LsoP+c9I+V5V8Up5ypOLz0657Jf1zmQODI
2xBwHhl3i+jFK1LWo8Kai6LYOx2CWCSpPfVhEjke30Ghw2ptiL8QTX1Mi9vDYjcA07X9S+U5YeFy
z8GWRmIzf+FGIyGQzPVh/YVALJPdhsVMmsb+8/1+s9wejxFJ70G00jlzEGam8siIhASWi23svgXy
yKMcqAuypWlHuJcmU116RXSkYDChjzeIKLOKzdhyZWNlKscybbK6hOq5Hj1l4EHIZViowVpYvSnp
D66DMuks9bwWBdUgagcFvIU778zduIvQrMWGRxbPAl4RptX3s08DdamceSM3AQVr3eY0L93Yb+8O
iCByH8bOg/crWNCBGukJncHoy52kB5E86FHYIi2gQe3tqnLdIjbwnjH+0Zm2I9RnZ5k2LZKm5LrH
eRGbAIMIG0NWqFXt6Y2TTE8U/6a1HEpxwdQr7Pv/LU6qsgAho4HjT7B+me4UsdhCd6v2VT/56H2R
NKE0/2F1z9bqDhM/KlxunxDiblf8SM8dDx/L3CP/3uBiWdpe7XxwbPa/sDmGkjEASXLjZPw5HyIw
pNRLqj7J1qKOnSoe5/twPYgCfM83rkMrjyWI0a3gG0f17na7JQy0D7QEK5earN6IInHy66Lol6em
jWm0INyRjKgfG0FqakvbJpjRXqk1i4GhguX1PLD1Z1GccvBorVhF3wNUY6WRMrZlelMqMyln5QOK
pqk9DRXLQtEcOLqAeBxAVLbCdTfo2+2anGh1HrMJUuHH525mPQwZjGul3dRH7EFaPz0pO3/sMdVE
maqi/9TWaaoUDLZdpz7syu31P7LSJLeFJRTAggabYoXmjSBLpgqDAZDGQkMKkAEzVjdVznXX9e7s
S5xjYhBV7x2JV3+kulWwBzxWQRtHIBHW0gKDqOr8nVi2hMV1EUtVLAbNzMnIDtBVu00Uaf5oeCMX
TJxXLMvi2kmb4vBpuwI5MRlbNz6ph3O5F5lFnZZC7EoC9ovjHZB6+A0BOA6lPoiSfMEK8U0eZj63
sDCoBt6lqhAaE0kVnq0xHbSl5/xwjL5cicRNqoluwgjzOLgBvDaVrSA7IA+/hFRfhg06/WWZTORI
/+VFKe6AvvvNNf5ynZVsD/uOWlgcNbp3t8rWrGjfkRboUzIpof7A0COxBRwExfSaoKUttmYon/d8
g9uI9EQCNKsHH1uTCudVsy1CIX3w+5mFTLI3DuofmvxLJYcyuHcbGBtSnIcF7wkUxsaIXfeGsFFJ
k/ZZ5iTcNFG+3TSVtrI2QcUowcyBVoLSiypEi+7Na0FHVFI9iBz9+8TM2ODXJzHGB742ZhbZ7IEy
8yGywCPjz1VIH6v1ThdDGqyOsLvnbjqJWuhXPW0YFtRusP4oXv1333mR3xKR2LKWdU4publDOTJW
+K37CbHvhCzSpJZxp76u0aHjdKWgIqPAhcjIbx2Gm3NhZnk1huZxWM74Mgb6XCaOhL8LNLlRDipX
zYkwOmLQ2WZhO4+Ygwudp3yjVE2idIh4bRtW4TJGts/DPVsJHN0BdxK8DOfBJGngzLdSMRyYbVF7
+r6A8wiyFvdynbauqYaN8Pq5Ovtz8gC9Iv6oQcko2XOEGeA586lJoX+m7ZR32rsBq3IALySvlXKt
1Eq8tnLu6IW1kLjY2iFA7KwHb0Q0Mt+zFUxCe3V6iyTfIrtPvW6FSmNzbBvsfAY9LvsYb44HMGG6
ASbDpolpVUjpWfTStsn7iee8xMLPY1gbpC96qUIsN1OzYS5s0Qml3OjI/rKSxjhtAIyqbGxc/KPx
fo8RxCM18oqGd7tlnDlBQhjvgbdneBsGgK0/zJzjGnyDLrDAgrBSou81iP3RyX2uCtvht3rgmYyQ
cgBxlNrk/6uoJ7viHi45oICCYMfwFDR9u+/qWSK6oRMVSqCLGKw25GpUIBYoLoNUXTcX7gmLDWLd
wNR7DpSz9O4bqwbRbPYvPq2N7852AynT1jjC0LlmSSEGLiy6/BfWGiz15ORgY3E4ekikabYemG15
xb65o7jwTECn76g3XWqrEpqryBNDYFgSlbcxQph6jQrmffSSa4Gc/iJ+Nsm9pYryKg83VIe6JsmR
a5uCEd3PTVEAmZBSSMcU3CO2HCT0ny/jDiiDrBfoU1PvPFMWv+6htr4LZJu57txJyeMEplrY8Y9H
cCSXP8UsS9q7QzPdv4lndfDoqmxWfybVMWJ1KDKLco8CcpvgZhKJqfvv2pZzmFm0PEJI/48uEEXW
JkSTFAr4/35EFKw17w0vPemNSVdRuzNYf32JXKTD927Ubpw9kwQD6K3Oz4nkK9p90Z2R+aZlyY+O
R+yjSvZPNrWy9Xsko652WZCH3aDvi0QgMMKgsL2DmIbF8Jj78qFVU3fWc5TlT4pI4qFSAgdHCxiP
dRgZmZUCD/qhzRFo388iipflvwkgveESkKCII48POvCV1vYCmw8udBrurSKtuIQKWY5Hf6Z/stHg
Wmt7DyeTr9wGnRd27N8uUUhJt30fK3nLjKz0/sG5NCO6D7X/FYwQu2CCzjUPQKiFN7B4ivcfhpt9
qRhFq+uL+dgLLRPBgVb9SupzZxYfp7WlRHpeXUTlc1o55ssBHKux8IUqv8j70yo5sTls8bYfGVss
f/YKZSDp5x+QUPQHy0yS+UgEu0nu3G9PW/bKwVAouU/JvO+m5k4oy1rmcmhd43iSr8cMCBql5zd+
TzSbAmvCZ8DXj6ItnEyCU4CBodud1HF5x7z5JbVwZfJKmvUlVlzouCNRElhK69Dbo9McqhWX9Y3Y
RqsZ/ZSBWGx6CJ7W+mj2lOoqAPO1nrUgMo3KbvFAK2BJ2LrjFbo3sGYBRZDt9leAObBILuxvLMuT
t+5aFg2yq05qqR3/W3oKrbX0FN3WVK2gGOFqbMcjhWuirdNGXTjWtvkOrbJca9x1mnVfYDlMzXyv
HuiPPoLIzEAiXB70ipsSo94Z8xdnQvr3tmq3PiQjNR1WX3As+/ctzy1IqMqTKoDJezPWnJ5Y/f0c
NwT+cMIh05AnfolUaewGBDcLXzjsndzme6osfQhfS83YlEhBZQzhqVvWYrifn3mfN1t7N95tev6u
ewkckFoaW708l5tqpVMppI9UTG3d23GFhE33BOsLBo2Em4lrB33zx0WlfDgmIwM9v/Y/LgksWmnQ
D3ZnhOYhPcHO33hk4ArJa6q50eQ5DCfn83patjky6V8TJFH1KSrsGHugQ0CsManNlqsh5e6OZaQE
ZmFrp5X1205UzK2VpZUzYLRp11vANQY4gq9L1I5IgGpC5d3mZdOtbPra6mB8Qp7dSaQBt128ra5Y
8P05v1pKJtU8fwQdM88yidcy9N5BDrZ+HM1rNWv4tigoNshDgmifWhq6dxk+iCCZOKvDyjuZWbb5
Uh0vcO16PU1qVhWej29ptbl4buWlEPhnrMGPzvWgm+U0mg2xWta/liwkSl6+/Z4qfv0oceOAt2bs
noPM3Kvjbm3Sfx0RK1IY9039UbutQQM69UBvuwhZMlE7HxxbmWOPoYhlfHxRyWcgK7WLbwKOgKMD
A81vSNaAU42bVmNr8nJl1yfr2Z+dmhFF2lpE8NuaJMHY3FKEJS3irpf+90hMGxX/DjPa4THWmG5T
d4STbVuAzI0QYQ+AuhC5stFLGAqqUppzsVBQ5ijUA9YY5fzS321EDSdDbciV/D0SOJoSxcoI7evm
d/korKEgob2pz1L4A/0aK9zl8g9PDoAIOTCZ307tTaETOKlmZv4NIuBC582aeUBOPiZAnPb/CH3x
uuvnBLqrZ49zlkVY+D6tkdt9HQAx4KEBWLCUAOjUkhi6QqaLB43GZjWPlHfrAPABSPQOwynyn91Q
LtZriLPTM7I7Gwl9bLVJdia9hndwESd22I9Ctn39vQovFsIQpHX79XE1z/D/AvsCzRwuf7RH99XR
llEyb4WZlZo3u7MFbEb5gND8ZlTDjBaXK3l4O8echHqcoLbte8yoVBn5dgz3rND4fuVy/7bo11W0
JB6xTQb7yscggI7Wzsl5RcD7JP8e5RNLsrAB3qZDgAq9JYMTcMeAL6JvecFvf/lFDOwWLASNEANE
Isjs4RvKQ51Gc4ZuCaxioN5oLJXuboXe/d29yZKEEE3WjRRvF9zl7ELGRlLt4NZ6nBTOM5RAq9/F
ixVuUplAKzqb0ONluyW0F6vOJfpgm5kSQm5HbEoALP+QWIE1H12dR2oNZNAEW4audsxG2yUjmmeY
OWyZNWpkWICPDKnyRGsEDWUQIPaLxoQVv7Rbmw8lnhTRdO8ZuTcm3iGNBlE5dJ8AiAM9mpzthyAP
pel/7Lp0QpQVLY06A7e+U26JyxvSAwmJlFHXPn3bBYf/f17FvtZpnlOl4quVPWZGdsJeYb3SHx6Z
9SDkwDhkO6i62XwspW6FhM8ZLArvTl8U+CY39FPMLI/bcJ3+btYZAivOpHfjGwcasq7Xy3eHgxeV
moVgHfgloR1a8Y+1H9yG2mJDN0I5isBzCnVdyorccZegiTgIZ3onANq9SCiBn8k8x+KmoEMG+waD
bJzx2DJiwFhlDVhfm0ElgAoFzw1TWREl2lyF++ez/wbTNeJzWRLfgD1ywGAKg/Rhf+JN/T1GYhmZ
XCPmF0B1kIR+FzVk/HROL4IH1WCJ1MYwja79rl+1Z0/h4CtY/1cathRu3gyypVQnSyC5Xo7uatJQ
owIOzSbe3emwcYkLaFHgkGUdHuaj0U1FNA3v1HPFTUbjiwR7DD0pEkh9feES5dUipyv7XqS7SF3i
9M3OakEdvwX0Rlp2ENCokiteohik+/RKxM8KP0QFQRlmscnD7tqM6I84XkWKFBjcz4AoMNhK4o99
zJKSlDxIQsT88NpE1Qe3atiI6k8yHBjYSbMnHuZ0utgsw16jCT1eyVkVMZs/ZpHL8RZ7dnCTTKQW
Jfx0lzRZ1MpWCVLcJGeoGqWAQRUHUIx9yS1pOAxT2NLIErLjFnPKpioAexdLTlgAwA6BS2AtUPKu
PTNbPUL3YNkx+TorpYwJbF35jPn/4suUJ3uZL14n9clfP70tj99ovJGMjLQKspT8U3Tog8jWqBwF
bypslhZLE6koQ2tT3DnUZ5bu+NKngIlb/P+nAEk47fWkLOd/gmXkQeOrN1XVoAQwuVw2UTu4NICy
4rreS5/bqMLE4Jj/+jOUuSRC8NQ1EFHpsVCYlL8/zyU0UP9Q5/4NSw68eORMxDBFMajtIb9Om+/5
Ev7+APylHCcQmGmxZ7inscMrwnPBcBvxONFx9U1EemU77U5MMuoAipzxzIDwziVnAusdAZiJzV4R
1SZ3OpJizpsNBdabOSdDkzqORG7lgDsb2OPLFXaEpZ9NDNvday9jts6LOnUDA3fhKI86N5TjBfj6
18lbtbVWCMhIClIG7ZKJ3rosY9z2Y1zJcR4vjdNDO+6uY54etKKiSMaadvsS/cKfoI4DG72l0rio
qrEzc0zSE24qpj/Uqh18j7qZl/G7AhoUcnqwZEgRuK7LG1/bYcYMWnRxg5D3ipirad4g62Jvks5g
cQlhF/jjwWOloexlMkjQYQ+FDRW986RZ/0Z5dB0CDly/kXDQMB2mdOAcENcom8aMIzWBeY9vB+65
p0UZt92RAw2cydB/M93sKIZrm2U2NRciV6qyFwyDNbUs6FQKFirplRfsLrgGDdA4Kua+6U2OqAG9
CrF/upuU7vpgFC9b4vrphhXDXG7dTqDj5LQlDp8GIMaNttbU/CbWPrkYo2Iz6UGQW7hJrdxqpRGA
q/5b/j7sxLTIGwoN53HWdVouNGZyj1vDnPgy5AlKkeV7Cbx96IGZf3wyB09yvI8LeuWCvNpryxtx
flLsX1r1XOOeJnxVGk4pSBGbTcxFmfeazLeGaxqvAWAiXXqdVYU8W5xWqyEpCRljeBv0/tyQurVj
qo5p5FyAK6BEkhFZ1hPEwz728JpHwZ0keL1OADZOnLuyACFyQa823DXfP/E4rrYNB4SpM6OvcZLm
RRu8MQa5QE9CgTqvSc6zzgFvgppBHJtJPJ6k5Zchp9BfVA0aQDeXsfN7rU23DwsP9rSkqbcl6Wrk
PPJgV6uWG0Qm1uGQzQclMYfthJlpJzKffzJjM5Dc/3YjhRwUaOagD0oD3ueqD4qwulVJKHg4QeXB
aoVakRhDg+/kMz0Y3o9BHW1ZUMqPj5Nv3Sr1IuTJP1E0ZPlWeBZwgPtTlPx6zYPg/V9yozrnPv9M
dwukB6y2rsHP5dt1lTMm/GSMW9eKgt8ZoBf05XPdSakt2SoDTq/rfeOn/WL1+rgXzWPMBY+XZjfT
RoBF3O+KDZS+LpdQHopL9ZHivXmea0q6+tUT6oDtJfQFiE9zuPoQsqY1fFOoOowHd1atzQM9O2S0
fZGFYvyX4UX2ugYOCRGTT8AC0pJEYnDU42vmXy89BC5zZAqTOtLj7NBMwxmwv5Nc+Na98FpwdDom
oedSBXCB9ddIWNVTrvp30IYR2PslTu2inPklFh4OHAU+BVkt0Zq5QUf5Lb7i3Hq0j6VJG7zzNHsY
XudsN1/izRswYdnk5MLVs4cDVbccIGwZp2FZN5If46w2IOB9uiCPZ+boL8bEmrNXLg4rqdhzi6bH
q80LD+q7UejrH5l9UZgtCV4y9AVlyQ67KQNSpfxqNaA3ktDO8rnrAekdBrxjQEJ+Rj22WPWPLvVs
z2dj6GXTmVil+086HItiV6+L08/Oc3bhVgJD0W3oOzTtZpyA8WvR4aov7B0bGCyuAddUNQCgfAk3
GXQxo6YDN+Y8ZQ4OmV2eN6EvuFj2x1vZjWufWCdmSnCm5arcnoAGiRpgPR4LQLNFuVCC99Oif0Oz
ni2mWlnHu6X1sXKfkmegZ5Z1NXyQlTcmtnethOb5wBoAaniEQJQtwVQ2Zet25nf2cQG8I3LO9lWl
ASvJf5lPw59i7TZfnYlyfxrgprc+Kfon5R0lMFbW707YEaPmR/oiCWrfd6Ac2NMEAxyYRJ72k2kS
IGyJic460vfVG1g13zQQjgv2tz6XaVNxH2wepCA44rWHgMfIJsIfZncXHdgFt4XkDaXOqG6BzBQn
B58FzFCvKwF5BV9mDqdYNrHhDLwyzEZVjPMrVFG1/x2ZIccUYcrFrSMnQkBczHJ36ZQgBxG/qzDq
5l8K9Doi5Otl3+elXYLZ1KxrQQgY4kEuDQlzWaISQH3f7rJsI83skQ5bK69I02icT2YOwxmS+W1h
nD19/rWWPjAj7n/qq9sq/KBKmUqL0v0XC7+TrSJk0vAGK8Brnze2DJGq5hTQyEkHnIhBAYcecuFL
RwFvsBDPdg5ph/MI3c6or18IRATWG1Kr0zWykmockq/P0bC5GU/Y7OWNatrvkq33Vel7zIVeeHT/
q6BHgAyUn3xobh5GKeuTYoq5u4RIcvPEU5BHjTpPLGYSb3RR3c2Yb3KbiYTSV4as4o9pwlNYRtMP
YTwRLHncPCp3CvIYSC3tLyZ4Rd8vyvpcz7QcNOcoSB2JHyYCOfAF2m4pCIKZfaxGtVtFF4DqVBw/
aQMWgyVF3MLKZqQB56WDCI3PxCUoI4JJNN/Zbjmj3jWfms+y0S1w2iD1BfdoOy1UiyUfazsDCUbh
aX1qslzksTSzfzBzHAAxN/LpRm/o/nVV3DutL4AGoZkoDAvrSmOf1B8jcaKD2UfwnFwrZOF3AcQK
1KM27ZDUwhO1nHjq5D/SMbmxqZ2388WtvDGXFSn65nyLb8y7XkoeoDReWOXQUSZ8qHM4apI8C/ne
+59gr5lu2P8MfvFT8ovqws32gKYcx15M1PpwEvwOkMs4e+QIRurtvkxeoHYrFf0AaVNi9ijUSPe1
G/C//vdR4buCa4TZDNnWL7tYpui0N5Zs4Frng2GlrzjZarEVojZ71TwIeOHChRhsOY7Ex4PlpVry
h+3xMIVp5VvP3Kk0DOprUdXnEvZkLOvMsUc9rKYT/mpmYu65WjfC+Lb4Y2PzqXpJ4S/JiCkC8arw
n76HsVPY2xPGLaYZsWrnYpJmROHB+zZLGmlaR25psfDVGBmfnYc6jPqkTuFa4zYnM5AKgsyQS9sJ
2e9S2kmoZSyH4B7QYl/bDMPzeeuVKNIcoMp1S8bkkhTyYPA4CB7pDF30ui5ZnOZsUDhlngcqrtFG
Y4KqRLLzZ1doVBWYV/NKsLXBacsoWr8oS2UqpkKdWJ2Niq59yYw/VjgM7mU/LvcF6wJBbnVMbvPs
QmI2tJoWHsIa1T+pDDUdjauuy1j4MzndWPZn5znJOrCj80WPOkvaz67Ptr+ko5uSKMOQFnqZUKU6
Fnjk8DqF++g0ErJ3t95xsiomBMVuKg29a3WQnpfuDyEn0jV9+zG4D7ZjcjrQ9MgnO7IWk4wmVZ1A
5OKIp5eN0CyGKw9RrDX2AVDVk3VdFtHNXZpT+4E7kJYKrzJ1HZ2rWp+/gfexPxiM4WluoQYkOUPa
1ickdGRQsmXt6aYXDW00GCxvWxoHvZXM/ZJbBIYchKMAMLfeGQA90PUsNxQ3oEQYBBQgHXf/3myJ
29uLTD7+l9dGX58Oij36IihPRASM6tbFGLrkUo9p7Bt9K3tIepyTSMsriApfG+XBcFKmiM4ymCnS
QdBFE03AJcJik0oz37CAY4nb3vc/S4QmaAqkPAfIyX1Jwag21vlgHC7NxBEZV7+HJJeXM06JwJOY
3Pb9X83F2jixqt9OWGfQocR91QipO/ocY5C+bRKHkDY2qRsGN0N020SrCDkFp/Q7vissAOmQd/ku
6l5rz4cvNAeT/GRyoaJNqrcBlsh5XO4AVwwq67Syd/G2ScO4nfI07VNoWGsJ9liYL9/fB+Y45Iau
tw/QUvBSAMg4zBbtWn54LYIL3yJNKZ3r4CMxzuU9T3pQkdkJeBali4H77p6g4BWh37XqVvxvCbv2
R0FrOQzI1tNWhYZghOVG7IyqjYYaZ1fL55/u2YdhYAlqxmka0svkQFuPVPlTEW3F9uklQ936eJYH
Jp1xffSn30SfKl3UCcBEszgdPqa64YKCZ9+rjG3g0Ewr5VGRpA/LH1scvnwoeqk9rY5tEtqsAkEE
WAGlyjeU8BQTxMHIq+5FIoD/rvk0hLiDp416ZEsmJ4DmSk1xJPyzS2So35XYHswD/wj0ZMF33nlP
MiT/w88f+NhAYhdFaxCPQZkvBNdMLtEIRgQ+Iz6W+po+aLCIz4TT/zVRVbqJXv24TvGVHfBq4B6Q
MIi851M+99gl333Xyedhcw9KtsZtJ2xsZclVxDpdaPEf4BAN2mUjcesopubfHF6Ipk0gSgf3XSfr
yKJA281KkmbzfeV1w7US+Jldl+Xw+SQiZkOnXhPzUmvTvvF6VoitXIMjXKWSC3dRJCV+B2zNKCDo
R3UcE9v9bAfv6BcaC7bcecQVVPR+XahCCaJKWIf7p+FkpFxOnZ22YN4YmmFfQUnfsDDxG7YoFp74
cdYzhyYZ39bURR0cu4lVL8AVdqk4uBgy7dDkocfgOlEUUQtRJNJfqRfEpwNOT/e2me1LKvn4UrE5
0EfCYXL/zYY1jCm6Frld5CIGFLSjQit3O9hNdXjhQDDNKrgL7qOdHxN5p9rAf/Mmw0arHH8mMXB/
HQOS0NOiZ0MuwjW/paJvIO38S5mZG+ayfVlwYVFIno0lMTxTQBQZbp7koe04KttvrnuQ+ee8KRWh
E8fdSRoybTQyrUuH3FYQpzg9pmBtKTfiw6TIC+Np4Ex+nDvGCLof5UVY+b4hc82x3HWOu0Z7dpbU
9D4UsAEzPUSZFV8bSyglMZqduXjNqItsOgVqR0Oa2Yqvd4TMj+4aq4aaF6A9D8NtgytQRmSP/pbN
NNQBuwTyyWH+0yX0LrJXJc0OSIz/CnY+Q1Lx1o48Lu50hUaBh/0SobKxAAPIQ8HCjsTyNwrdy78/
B5141ACOqJvpBlw53VSGpZ/R+O1OSrPOdZRopwRtvZOCD109N5KzGO+jiAPhWQmd5CerlCx3KKqC
SfINzTqYUFJILhryCeJzyApJpVFM20gDI0gXcpAvMw16FNeVEW8xYD/rtX4p8nZEnLzSrS13uWkn
K3ydBTQG5pI1TgX2H6BbQKBJZvfCDO6hUKu6ttMD9sxln8d//upe3NXNCxcyJX6xTj0hzXFpCMAZ
nDFdINxZR96ebyh4tplCbpgYZzJQsZ9p1VxqcJY2lD7/oOQ42HXxKv3kdgwe1VEMX476MnInjmOq
g24CbFKmgEG5Pj1yPUPGiCl3uI7X45juQeg1guoiJQrScRQFyr7cTZrlfdJYdmnxFkjRQ8laXMgO
KvDFI99eFJHtdRuGaCwi8EwaCBEhLIW/VilxnMgQx4Vt7x1cSDXThyAP5aI+c9N2FBBgG+eNQG0p
F0l3K5fBhE7sjhbTTUM5qmTd662grVmm3zNLR3POFekJaT3Z87MYAX1BsJ2LJCoFG/QnZuWKPkkj
rM1gIye91VmJWN/DUpn1d+vUL5q3sZ+z0y0qm7/NTXDCa7kkPSPTVxyHAXbkWaldFnHvKIbd2VMT
0dUHD/pO6d5YKd9kTvuGqWo7WOb7onKOqT7uZuPU1lcVizt1ylSbTOEZtTqLbq2+olNJTJRmP/6i
W/xUn113S+gmVqSxBT0wbutSkvUvWRsH3Idb+Fhx3VzszmUIv6opZGj/1RhpIFz8F94SAy0ZUbyf
+SNVR3BOSkg3g2H8+plcvGYOkr4CjVsYla93AGNyxIeK5v7A0wNCT3tkQ8Vg59uUSJzd/BySL8mP
s0OhCHc5wPiNRldV4EM9wYq86LuJk+dYMEgdK6jAp58TDnAEPgvTx8GKBAfOD5pPU88vb4EC1DmF
A6O1XO2hrDTgFbjK5OBOSQcevmMZFOu2wA1M4h8TctsPlKkpbxIjmJlSkfUxBlCX0HNrIBS4y4Cb
`protect end_protected
