`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qf9zELYJOX2pF2q2av9fbiQw+YV0TEpx91qkT2/2zZyVHzAvT+ECkP+iWYh8geuU
NuqB+rB4kGpoIDrX8ZTbhoZhmiw/ihsy+4bWbkCnx7fQ63YwxjenC5TLYJphwnBN
gMF1MoBI0H9Bl79SJy+l/Aux7E99vlGtATuXDbWNbJw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
54wmRrXj18+5FRkvuGdZKUOQD+gonsHffW8VF/++RkGCBmCmvDp8pKIw5b88GFBX
7MdyvazwM1CAFgXWMhK5MbAz7uXBhP85Ok32fDIPwcJTbeAwLvmUCrm5/YA+5Aot
pVF80VGhBWlbaYUNZPvFppl0CUKCivmmNkzkRadMlXx9Za7Hm88Icy2JCxnHKn0Y
1rjbuAfFuGRfhpN6ezKWTobQnNEdTQqvWKXBDRL4AgrI4xD5rH1wvpTFUzL8S4LU
9Mg6jzv0eWrLFKRUVKIDFkFAjTCk4SwUlVMivJ8q9SakwofZTskoeeki0CO2qDQ/
/gU/5SfygPWRkLMLs4nO76BRzBC9EZOyjJZmlTln7PohBAS0iYgSaSSvLHdpwjvc
tdnv0Gqc/qE1wUs6Bg9YGvi07WwWCeAPG9byEDgZ59L3B2XNuHY+sElvc0aqwEvG
/zEGqWKgkDrhumgTpNcoVVccJ/KKb6HgH3RF69UsLXrW/UcbZmQGSnOcjMR+kqY1
H1GgsO8c1H9v7Q7KK8Ltegmf/oRez53d3ysM43HUD8ouf2vTiREu8NLBsRA5EkdC
i5nYdnkIUSDgjt9u217j4gjbb3lyFDuOzP2LSDu42tc7iDXFtZwQiN4l+W7avUk8
9prmZG28oyx2VH8xHe0gtQUtUQaPhk9XsDgzrXoJ7zmjZ42Cw9CnO5KiGaqDBC86
GIxHNDfDMVe5uRi9h+420qNzD1t2L70F4or/ZMvRgJkhhtB24hlBPNijQWo9ZnX+
eyjG8UxTHiImNlUJksMZPpcrD5urTt4jT8Eci3beqjRAHPyaraHyQy6UeoNwN8Z1
cNg2OXaLUaI/OUusOL1Dw4s2asHWgJmLK0vaHIwvLQVKLRd1cfVJ+kzpkTxpH63l
7gmZzww69CFfZTh1e9CIPYykKnypE36lmFI6Mj4umHwqb3Wytl7p2McT3JCxQ0+q
I6gQOIr/j9ykxfZaq5j+6sht8eIsucswOkXG4y9EoIac66TIsYT5eKORawGiREJo
D7sc73TMOXe+F85b1uuRcNmlZ/at2qD5bw+POuHIp/swUiLuBJE+xaM19AcbcPNx
d8nFWJlZ5RTRJ1wvekIId6TqtqVburphVqgXIdEyn5twYeBUGGV9dDzCa83VG0ot
3gBvPjVlyStV3vQQp5pobD6FLCgdTFb0vDTt49cGF1uoleD3Ao7yNNu/jX4hkNPu
2Y67OEpkLTmCvXbeiYrQrVDnYyUisTHZG3zhQQNwBoyj8pIwut0TMX1ZHG1KuSzt
ZcZdsqHNZIXXgnJC9YbOpt72k3y7umZWZ+UM1v3GC9QZfQjU60Kh0tSlJE0YuW+4
lRJJMWHncKI1c5guIrDXEGgHsCx8u48BwPYd/Zt7Dc+tmknd0E7CE/tzx85XWH9y
cGAZRphypFb3eitTpP9RS62qoFAyfbfg+8xgGykzFodGEFupjlIsZp6IuZcC3tkE
/lO9Da04E43dmxcxXHSScPP3tA5QO+LPRqKvUc2Pxsml10xPnVsPNeYGma6Z6r+O
fEwI2CxTxbSby05GFSNBqBNwy5TFeCZt1jrncSIvImI8Y+T6lIUMTVqjEA7ehJmz
WEpuluozYsrj/3j3zRpQYFzuujmps12dRlbkQUM0rt098X/Sfd3QqUFCz5pImgtU
ycGkfkQ5Ud4S8EwXwP/Y9mMOKTa3FKRzdiM/YkLffdElGxrH4KHzZBmLkPTDldmo
qADn/7Oedn61JlWwhdk3lR/4GJRjBzuOeDlMrLkohKIDYMp2BcbQdZSeM5hhX2Z3
6IzVVZ9UCQJPmlUB4AMKkDavkvCgl6gqT819QX2YOUS0+WBXPC+NNZoBtCLLdq1B
0tePalxJ2maZaX+J27bArY/OGlcLuXfmOcPYSO1TVnZFHLwcPG4vmw55s0wHBnmA
L/IQCE6cwHBHqu632RFqdEiv7OyerrhosxuPfW1tw7uBDbL/0BHArRo3i8jz/tpq
kHSmwtKo0ygzjNiGDcWrprtps/hBiwD2SQ+SoiBNahjFFY63lV1O6E7im7jZdeEC
Ntnv2WnJXec70ixf8x38brqB8sTBMm9K4pEUa1TEF/j3gu8XwGY/Yop0Bojw6V8w
GcabiXB1FCYu1kdpIKmbCczH0jof86DVKMENZAhUakGcfI0O8z45WUQzzmULLs6i
0T/Zus5buKR/7DeH6sxC0PmRsaMf0xRD6N3TNIxNJ4GLPTTe4TmSxhJ1xhhwF7dE
f6Bmwitzfb9JUv/N9VRODQGgQ5ACU77ZSmR5EWgEfNSuLFkL80P1lNdb9Y/lAM/Y
qr55gpIJnSJnYVIk5fz5JYiYfBGRmapWXhuR7VLMZS02genaBQEtgO5aIQrM7J5k
bWmFEI0RvZ5W8eBFfLHwV8YAi8CQ92xS9xjZyhMV4lH3fV3oCkRMuoww0/1Bygao
7eiHDlBK/WMZQ5/j4DLjrkO9ChjSwiqejP9FlcZzy2wDEYPJFLFh4VzgUNP0jrgl
rluvHDUN1Z1lzXJszpR0AgTWQhVl3eBAUgBTACY6nIh1fTH2xz6yRxm+a4LLsZAA
6VxpYnBfK6n6xjDyBikotBtc5rZLhcHBhgoclyYPAZQcVr0LRkvfb1rCw26WI3sQ
9huUuenLc18XQuIUrnmKq6uG6Q7qDE0vKVBhmromK0fhejFVGRT6RK/VNG3zRmjQ
BiDzNLmZLXYLRbumRmSKylUuedhNaEYm5iwa6bUYsDP7KOqib5/GlcPBG9vnNSJN
KkpjGmBwH5MDEYMSBtdsQV/PEIeIBfYXIPyCuA33l2HH5w1NH+xMqcT2xDE666ox
GyAgYO7u2MwUBLHQLi5PErD0OlM/tpgNU2ytUdl/2xbCrUzg8684STHyalKCxiqi
k/KxyBXLJR8yZd4vudYM40RxMyh3A9zJIg5JBCC1VpUHp5S/GP3tvHo3XCz3L5mV
PhfMhowS2xnlgvt7SgGkXZERW1cJKjbacI1O81th0dtUSZl3LBHhBWdrAbkWvUbp
QCke4qRp7MtvJnxzgzY+YiTlXXCogX8ZZV2zpFZFJ9tHUwZ7/NsCeDeg5T89H8vY
Zu51IbBo3udljQvddMgd1Y3/TX3R7o6XtuTyXcQJIhFEETO6vaxdmIXLTUEWB8ar
NdBvWe+BxTiFJk+j+MAs6yVm07mGksgV9AGeGuE9DuQKyPxuOAJzrAPtB/AImw9p
Getonn5UdaaEq1xCX9GZaPdfs1issX6mE95J2vKHz7RY6hM/Bsg1vWiZHYIwTKZU
ziRxr/MVodkguG19j10MogfRjovC7gYIbMCIyP9ZWEV0P0W2RjoHxa7H/LFmGLuU
9kE69Ohjpajot4XZqbSSSesHih2kjudyCso6NdB441TbcuntHhAnxlXIBwUQllZF
5dxO+jEUN5VAp7T+kqpsaJAlO5T+6NuxVU0VIZoCaLSVBekS5QLnV5eERAeSEDXA
hM0uffKzJoY89wHC96smSUsUJWcwh3vB+bYmkJAujEdurUALJCH95ZS/KFsD+mw2
eymXc5518QrU+v9zUR85Ykuc4sIHrWRzC0hEMGW+E8j7Jni4NRxpmbAWq+sH8Nl5
cvpnthPx22VBzeoG6gEJYvj8cLN9GPWjq+6VOO0eL0EDE9LSKDGRRqaq9OTNil7g
T5DVEeiwNgEB2OEWOAirWERGj85uw7eig9CdUJFR9KKSIaqt/19m1MgnQBsIWqnw
qvWpAl2i9XOWGf66Xtw0A1P8JzgWeTRtE2QRFdZMO73VBN+mnKblvTJ2cDO8uSBv
MS0yXdp9n478RldxLv3zyqIhy/rT4z4O3kNJrSFN1zNmcgvJQbuGel/4VDEJiHz1
NEr/vzF0oROk2hUtPNvK65rBemWUPidaESx+RG2fv6C6pRiFPglv8+uqCcRRcUqH
tiS4nGwzn4J8DtQ7FL61viM9+iI59DgcquX5WuW9V2aXUVhOzxqxW4+U7hJf9x/p
ybTTJAgwLZEfQsyQS+F8lyp1bfHnETWXQgNdfuf4TgkRmI0AmhvURN1Buhu1viw2
yY2xd5lwHjXYw3pqSoUupVBKxvQnaBecmsH+OaYy0fKcyInCUSEF5UlMyYh8quyq
TJvOpYR8tRb/Be+A81sNkoy3RIbDsnV0myt9OP87r0e+RGOGLvlKu6gCSL2F7boY
7Yp0b578bc085dm0UJP3k3j4xWJWxyfTr3E0yhpFXBgXhGGbn4kiBsUqJyEMh9Na
Q5szmCNPXgcNnF3ANmvPpoN39qo8s2XDlN1LTwITQGOV74M7mxYG/Co4MS7/Mr6c
lfT8w7rR0XFb6YyT+6TDfLdYduve5J7SE2MTA+LwkY0/1fQRLX9tmXE7YC2dnk1n
+nFZq3EFErZRsH6g28WgY6H+srEN1D+eJIY1nxPMOy/Rgv3wx/ZoFMpvpVjgTB5w
KocpBBPi6296/LmM903ucIUjpqvw47S4+90sKolfmuAsEmF61Zgydt+hReVGcC3l
sBJ/r1uTTNHSZbW1VVRUIau76qUpgF7THDfD31/82Tfji2HHKFVIzvdpLIVhRQSe
t0o7nl0DkofFcEr2zi0sIcD83BAXQWb/voYuA/a85nv9lGUNfc8hdtP2w/n6ZXLu
mTaKimW7lioj6lYWYgbyscDhnSrXhdah73YBy+N/N+ZuRz4JDo0VMnE8Zi8f5PAh
0w2+lxdUvli/R48IhD0AwCm/FMCKUOfJFZhE41ChIA81yQ6+7Aby2CrGJoSSfFfF
R+CCEI/JtHhgOcZMMBPQOmaZ5x+qBC+8vBNQnVMlTFgOQZHDqhNmxKUDy1lQ+TxI
Ljiynat8NyZhAhG3ZzKi/X5ED+QbvNkeTWdB499AWB9KNUFsDm0vIUEQZgXn6xf/
3bu76upaIwT69VPEI2DcSnh9tEkvY7d1HZUvlyg0RMd42uVt+MiX1uX+Y/zITWps
8nF9drMtaIUX4SZYxFoZekSKHB071pS7xJKvhPd7DqUnQLe9daHbCK2BLCsHSOHw
Raggf6xoNzLZXWp+tE/j+aaAZk5ccwebIlE7bGZMKT44JI46XO2S5PTa4Sigga34
ipoH36HwurJsZsi5OFhQJg4IPJa2TSFWp0yD3gradNM36X8Uc6Wc76qCeY8tk5ER
RImpfJYqzzQuLeqcgo1cyd5WIHZxzn3mfdMHQ+i3Frf0RPYsFllEN0dTF8UOQbOz
jORTIRkdH0MYvI7iJzKkqlTlGQbvGQEv91XiVRFmUhQ0uJA2zV1IKs7xDzYX9uTZ
IY/wy2CRkjEv+6SKopm3Mf8Kfc0qMkUV1fnqwgbeamRzeLmDddpv0xCgVFx/S4xO
BjjD7sAFhulT8cA6Jo5w0Tw0htDppcKJFF9uyIRHlNZuw7masUqaYlkoXsk18cEz
ECYt74GM+e99lLFMI851koZbnm5vEaM8VUEhQKvYEYvApcnZjag/fyEQoVTS70eQ
MBxT76iwgCu7BQs/IJ4C37T0th+wE9U2wvu2dLDZBZ45Q1gJIL+Y5JDA9BOyLSMs
xufyeZQsirfb/5RZA8HYPvCbczB/R7KjtWMlw7Miv+IpycNU0aImCPzXQThf5bLq
TwlkaOZklMajFW8gAVjTig8MjDU7OYQucsV/izJFm41ZIDgFZ1gScH7kFFTK0RSb
h2l5fi1C3NkjyKkCALVjEnAge50rkA8mp57BgwTHp13Wj148aMpCduIy9sa5Bw/S
ZIY4EHDyHADjAns/FS63SrgpO4DHYsTSJ8IXMBMD/aUVho8NJ0WPejvGFWhurtbY
KodHgY/mjUYV1DupWlJ6vcJoFflJGfmvBXWSe377kY2PUE+eQoF1/2dv3+Ylh1oc
kc7Y/G6tUC/aTNwBSPGXmI/qHHpDozi0T/BjXhbb/qfYx/LT6mF24ULmMhd83HDo
GhBPwIawpGBKXgLC3frqwUCck1XFfh9pLGQo/HlFQ2+7zacGDcV/ONbYCulenP8u
JoBGoWVWEt9biZKlYVGREOuR3L/6BOlA7f0Px5xUNyHpdJSTIf4og2kusFfl7XQD
vABFJmBVeMUvQ5YlGJiV+ENPxMeW3aBHDPfiZ5ybVZC5zl6yKZCeV1Gy6zgrc6b7
MgrnQ2O7iiVdiofzRPR9+G/r2Mn2VAPZr4nexNvfE9UCKkXa09WIr+rYd4aSfotU
zR7PDFkTjm2s8lovI1E+YyZ8pIL+dJ5L6QUkF6rt7LB+mUjHE1giFnLKRlf3m6wH
j7TWOJwbNiOR7Wgclo40CJiPyhvr3tcD+rM7NNlY22IKR8ibalT1Zmf4Zx+zgQyH
5ydpj6HO8z7pOHy41rvP1oQoaQRDCcSJhW4rz0D3+QQ4LVXF6xUytar5vbrQG1wF
H//DBB6sYp1ljzMIDXddiIqnUt2L6FM20Dpvvcrefu2yJmyd1sRT8MNTN2WAEJiF
34ZtGD5XjiOXTUHJXQKCSvmNxfnH8OyOICLmafm8ItdvpvyK3mNahEr2rmJVic0m
vP3iKTcBnUo238a0mS1vTFlV9v/0bjUu8aBvmTV0Bg32iw67+6JTLSlO6+apo+5/
LJKHqwdEfAK65D7QTP9k/z0fay/BbtvhxIwOAN+yVG4a8FMLu/l/e7SOW8DH9TQb
CQxtwDaWJZLM2BGjxGEHaApLy8n4MAvYeYY0M5OH694mFdqjc8i5XTZqOKvfcgF9
rCq8Vi3rPUAfsnGhDyNlUdbQ/7JMldtpNv5NSecLPwTQNshsu+h8uQcHNu3G24fe
Flmx8myFxw8jI0s3DHAqJ1iPbF0dY0P6zeTZhr6tsmdQVW5OC66QCjo/1vlbuoP4
j1doYl7A+shhluS4swgc7XWfyPw2pkrdtkBX6ZKbczmWrMtf76p/vfY7P3l775rz
NJ5J1z/0E7qq0v5kZAx/YJfB8brXEJ5RmGlsKZM7jJTgbdTMIx55bYNjrzCVbqhR
KKJEKPJcaW9k3lxkA4uqjWSAxqoIorWvr7kTLiGWiWKeSTyq73ZErVA4ITlhvsOO
B8zrogfscJ2tTtEM52lkikRu4SXsxLsjOhE0bM9xxOF/3e43u8omdTgpA0Ek+7gb
xL838HajLolzL+v5RQaugeMqMHxabvbE7vzjpmPjuPVLxB7aKQi0VpwM6SyhZOx1
gtU5K7PsPmRhQdNtb+wUkxBfZHnHapn2fGKCudAhJi2YKQ/kKdGsK7CN/8jilCpS
hwdvGhzihZXxMSfIlHP4pC/5zUVZdbP4FeVb2FoaucjJiCXruc5D40kSNHCwYVvC
puld+3YmEuXD1FNqT9J1efaIdTAjk6ykKKQC9Qug+si0/yLt0qZbcXSf/AbBvtCN
JX3FvnLJhQUzW1DQihSfcPrc8REi2kkZiuR6RSKKBd2PaHKpLNPe5uosnbreEBz6
aE/4JjBMdz93TwvGW+dmSfVOtE/VkCzNc2++Vk9yZiTjL9xqxYlCFiLSHKOmkRS7
kOKS3drZp1+euFnYNAqOuSlXJiHJ9zF8qXO+AbNKGHWO1HkRqK3axDh/nbuhtLLx
VW0/kuVo4P/4uHEnvGU2PHPj+ft56p90yI/LLjuuGq8OEzOSEK4B+YSeTsF6kIAm
8Oox/xjDOzpQ7Pz45b8JGw1qL00iNgEyXuDktEQQxUCDCz3OxhNtN+apNxPR8QIV
mzt62qFs63jGjDyJQyYa13UHqlJb4OImiaAmMnD3pxAaX8huF0k9yfELFp8lzBJY
6/mpydZQUjad8Oty53f8/bpFPghP8ufNu4p/WzWDvulDSRtkyifZhfzY6DirqnIa
MstCpEFX7TLHwgwaVWnIELQ0EjwZuQ1yV/GawUnAZRI=
`pragma protect end_protected
