-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YaYQl06MoRJqf4rL/ngYmb/fuwT8Wo8B7IenbEMR3GZ4OK8he/eigUb36fGIlQrFCmutOlTRth8W
VEgIFZXfqwyK7eBNa+iJgmLRQjm0hLB8HC74qTkwnQeCZdQL5Aq5tb2GQ9wcU8Ued/Kx/wvppm6t
E1Fvwp2eMxvVFFTlY9YIPWXZ7MNoJ8RyQok5odZ5SpHNR+NMOgmQl2Uyc2H5GdxPqCXBdVdKSry/
dWIp5umh/BquPiLRsqnKnmVUqwH81VTLQ1+LFYmhUfpfqlScq59/FFOhc7ybVD0GenU60t501w/B
VZKii+2k5cCpIOG+5K3y0EqAXUQGCQWRiJmwsA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6672)
`protect data_block
FvIxztO63dvTdjuolJzwR20P/cp2FTR1A0FAkzQQUfS5zRww+psXPuyUwTm4lGXwVyAySbhRv25Z
sJ95xl2hbgO7M0wN6RLfmAgtcdrbTeX40WT1XPRfEWJMzWcmOH1auC7823rKIAOuDvEIoGJy+q6O
D9u3klwZKCZ/bLXVE25eTkREFuY2uDxsRUj7Oc+2+jEHL1XrsNg0MFEDNB+wcPMrp0DOqST1l7gx
ctUo49bo2UkG/JR+oCv976FgET4yXMHlfHaE/FhjGBAGW7b6c0SqasjLdAEpETSGQyo+DV41XfDn
qcujVdl0b893kDmSEQv8ruoH9c7ahi4twplTfa1h/mFTzoaTaviLAdBqn1wWsXrs9fTd8U0P2stY
GoHGuIxW/gWQhflw+wcfU4lytZQZafp2cMJzBNPfq3Fwk3DdsCvlds94CuEmtEKvsxUH4+PU2c9a
i6eEWmK9mzGpjC4cMO8IZCljDYNz4UxAJCX1Bi2yduU49Pwb4ya1Mpp1ebSFcumXCBo6yvDwVsGu
6jAHhiQ+xytzlfyQXDXCiUTo8B+EnNv52g6ltRQhX0ZYPqMeWSqwVwIK7AdhgeMVfdbLNOIRfjmx
xTzIFsKIWY3Rq5rXnx9U5u9/FpAHthQOT5uiSpCs2ZEav+KQ2RESdYA8FJji5mqpYEtLWmURJ9zW
Qgma3l/LQZhqtPzySPYKcNwl/of34KEDDQyXClwj7nMweaQ7KloxiQ4Za8xY8s9XZyvYkRQMc5od
vI/esAYYK8x3Yh5HU17phEyrT5LUIT7NS/F8cGgXRR67X+sraThhxtAyfyaD3dBRjiEL+yASwfYb
4Mc14bOgq3ZGSMXoPkKtg5u/w/matHuk5DyXLCrV935i+6VcTVpFRR3XgQaW73LxfrahD/A+jWB9
eUy9+B0JPMI4LmV6wvpuVpWmzFxRNTNG1fkTXyJjb4PWBqk70IxBWZfrYbdBrVNnjuThco6A0mVO
/kwBegu1Zhh44XD2m3bv3eSIjBI3o2bqT3lU3a//F1UhwR/tJMdX2UiRApvGojeiV+uBI7paegy9
Ud/ZWfETjWv5N8YA4hNEGtWByMgQOifWoX12LnzK8VeXqbAwfm7OWeYo20fxCgL738k1nnqdzZ5q
tr0zAbKRbLQV/f6a/UbWjGJhV9L6/VjeJ5BHGJzoKEtwJQL7TNoeS/g0nfIqnfpjgiZHB0DfuOJf
s7CgrW5h0AMr+ZPocGYIlUDWwU1DaB9jBEOFA1A6HYljMqx5lwUVTRdr3LIgNa1Y54kcTd1Ghl+A
7N2En/TBZgIGO+c1UucOz5GCKd/DXZ7WPLqfGq5LUHAaHAjnZnuSuBmjiAh7TUeF9q7PQNxamGjm
WD+3ovPb3BKdcHfNXDQuZ0gkRZRAFzlKR5O2ChOddgGJSTZUJn3hbxg9YFxDjPlBFF6K0aI8kdQz
S8q1CK6re9XKqwKqD4Q2SacvCyILGV3CR+oJSUHv6jPfIffqszAPQQ2wmydWyNiMEbCMO3RU61WI
EnVQI+TfaEwok+nfSB228SlLGmIf6+oPDAu4Jvl3a0mfbhLdZQSK3Cqv2v1Gk3KJp9wyweUuceck
sLWKE8Co8lRbYO8Q+uVciQEScTyLbK954rUsBKHlz6ij0+IHE4m7EVTkDJMWAeXKJ7GBkzglq9Ov
/T6EMMrEzBc9fSmTGVQA1d7e2qlHs/gOVKMSkb2OhrLyWJ/xgL7Rv+HjDQvZgAUwL9e7rpo/aFqm
e+2jszTUcFHlwyDn1Q1YTkfga2mmI52sIZi7mDJ8Qz3pDiml9vZ/CZVL660cGgBonN5DSPsSNJNJ
wOYaDk4uTSwUtklR9ElWtxP7+kIkb4M3YYzpmfheZMC8l9DaCnDuRPlQ1G+wdeCG3c2aYKVkIezL
FqQ/aAO9U7YjeBMuSDsBTEm+5ReRPseelgk3FlD7ObhR9DuNng1FQz3XEZFI3T9pSGheJa8c+rmD
hVCprJ6747sPB+A9vbIG26v1DkeOKSYPQsZLNBf4bw7fhluB2Gsn7FDN1caPAcI8Q5fovRiMIeAL
9u3A/WSl14hmbVk0TfZLsn2BC02KZREANxATvY/gfrjPeZzoI//LdilVw23nCmyPzWf6pIS8TwAR
eI3KOZyUkgKNbs6pKWN0Uv5f74Zcs0/IraiOo+J9stvFxynHlUS1kcxCSEj4aLHmGsAoyMqPMB6C
lX1XI5/br1NCGSxcACimgfKFkZ+dNvotocKXDEM0m0sY9SHxrIf5qtf2Vh9b0q3pGFZPjM8gEVZ6
1Cp2HN5o9Flnpvk3CBqiNuUBh+q6dXSVjapb4p7B6jCXh8aTpsGl+rcp3vZqYWXus9l7kWlZSnr9
qHbvOvcuLq28i4Q/L+dCb0p8WZrdlJvdlqLa5uKLVVz/8aVh/0UAB5yQ/m4InWSsuzzKyA4D9E68
nFOeG6fXepYKv08eGYHcSkikd3NIGOjHfXdkIq64oh9zWyB+yMCaSk2b/Ou93ZTUB9ep98EiYWzQ
FZ4TLtUTtfwibvjqDZkJyug8dgQyL1mr2neSsLP/yNValqs/nLPZhdRqG4DBBh0YT9L0SL05PKW7
Fac0XxGAjv/rx+D9HcrCPBe64ncIGsyfWkhgBiYBkyLX8xSslyoOKgrjZ9VwMmkyhUwDsfKrEBWc
TBAjBhblR9i2tEffRbFs3PTRGK+pqIIgW9NlbkC3IU9g71PvnnfeELZ90G0TQ92RggysTbEpi5md
ZOW1bxuhxdq55eI9fvgDVf9YzfDInR3ylJ/XHujkfB0ZasU4qfPCdXuCBnEJFGYevJG1WjEqaDsb
VtFm8ffndRGqDcreYezS8Iua4/KbVT4bWSAqkUrvZUavCrcfEqjnTG/fMTYwVnrymgqfs799goOz
H4QbIGEB9t/j2Q4iPh3mSFYY9go4zMos00BhcHA6UYX1z9LnvByHXdWFUqSpa0dMUKK0+9jZ7n8f
4AsR7Rc0kF77EVS48KuPAu4N384IaQGLevoXtI1btw/9ALDg7wpu55UUxvcrnLYSQqbPXudwPIJ/
ZyjKU8rY64WipUqbXNoc91JJGD2eLS7Fy9Hf/7187IsL4HoCwMiFkLdVCdynSRTsEPbcwE551BlV
EDWd7Yzo9wdfC2DBOcQ2G3bpElN093gzUpom2SxqRu2c5LBSOT74XAaHDfAOb2pZUVVZs/erZzQV
Fgrxbue4yv305oCTYlaLzQ3FeGwbylrkl7e+JcDVyrK+c5iuoNRyVu5UuzZMXzHDh96gkq/901hN
55qdLheZ1U3tmO+NghjkF/9O5RuvN8PYSqM2KsxvBtnkItb4z+UNPAwfi4e6L95fMa3Jp7d4LTcP
zFhU1UvK4Ni9uvcZeYkn3VRjgLb/v2aOdBM31rOPgDXL1xTE+9KO7MDNDZ+Gv2Gz4swEQ/t9Ux/A
qvcY+U6nInwRY+RveO0yIw07xFLLc0Ur4nGeFJbETw+1NwE2KGEbT0QLLeiBsk51jecduGl97W+j
Mi6HXCkn5Q3ojr5cHCd62HmCXctWSnBhnVrKDSu1dIDZb14Lb1Z5Y3qqtb1wGdijyZh6PZfp6X3Z
RMmdEYvDY2sLIMcZNXODVMF3cEfZkGmAd319ra+YxTccjvRqBjTIqV7Fj+ZTsweU8eRdH9sJs0Ym
wfu6Yve6QkflhlWZydnLswuB/mOJBDeTO9lbL4JCXwxVzl2sY4cwZVSo1kH3ajaMJS9brZpeu39l
aCXlkHK5LPA10TYJJyKepBxqxl50bRcetNW8pcQxnQDlhApSZhDaL4xQN+A6lQ+XZiTW2qaQZMLQ
vnu+cFFDbxVHqqqPhcHUZtCmSFWYo3cmYAwlI0cnB28O+/0ToW5hxvp8Nad6bVyaw9/8TIR3smGF
NoVpx4ZI+onPKJqmnXKJhptnouYliyR9U6brgf7U69DSzQehFf8+IIX72NHCVnF54V+CM296+MfK
6wsNHjXNkOIexc3mrPLIJ2IlH+NsDnMBuoldBYYg9TTgBRTTc3ILcDMKXPGaQhcAnMCH19h76RM8
PlK+bdz3SJTeDxokikXzaEACiIVdYksJhZ94KPRAF7LRjWSMx8AItzP3P4fQY6SpINhZjY2un84m
Yqzd7sFxd7SK5ztsYy3qvuJ5WHLKExfc3D1IWUqRrwo4IfQ9rRm0j/0d0WxDXQ4oHArivmWn76pu
n4tPT/wW2+JmPB7WuX+D1xVNNr98/rrPRRK30U0262D1YnU89s+l0khXUES8l7LJo59J8NPRV+oJ
OVB91a48pm+3pQkJbVcUmlaW2Kf1PbJoBoiWuZhsa1gFL2ijNH6JXv0dmdJ/uZq4mk0z928HDZ7T
ajZm6bKhASrULokhkw8Cf77nBNtLLDU642KR2ib1XSoi1nfE4DDrIpTsTURR7YJduaBio1A+xNlP
K1+YUzBBU66j61c9uc2mWOLmh0sx1XbC0R9GVkYZMa+ylvlTfvmCYjCJrfBU9oqbE1abFVQTh5lL
vsNW6GWVDkgERpaANI6UocHIfoa+3atZ0Uj5bcY/XkeKgiZ1NpQlu2BWzT/2DduSlCYpVbhK5TVe
YccI7/tujymigLWCg15vGZEJNb1bGW5JMtejeZh2/HhjzkRZUCTsPdJPYATsEYaFSRF67bUSol4P
Koe+4P0H+hcxkL5nP9X9+F3Ualx7aZF+arC/u4Z0NL/Uvm5RHQaF0a3URvNskBjG28P1SldXwTx+
yZzl1LmZ0wOMwedtOaK3MJR6ZvMn8et5jA9J6BIXgrjxPdMxdRWaGmeY5w/Vj1YATmI64PvdKJPO
TN8FpLq2iqqsh3uoTo83Pb5kyOZtDuidpwLHeQZ445ApYyoy1ynSc36HaIYGa2kzHzGn6U/Y3hZg
NDApbHJSFGkCubz8Chz4HnPZ+RbmwX/TEJxYIVIdpDlZB1ypWGiIn2XiitflTewdjobb1ZbOP82e
4YQTqZk/6S3i2IM4khNNKLPk6/jzOtYs0qJyb07JY40WB+NREtywuVD60BCmC4ojM8qMcx+GVF4x
HN8m5K8dTG6iGks/UtLIvMz/d9aT7mqmr0GzaePcZidqUQFn4rK4rViRm9UstmHZqCq5evypiJo3
B9Ocj3tnA0Kd1GzSg1kVXUrJ/Rx2mQOp3cA4o/3RVMWzbTgE051RF2Ydea3s+sqvTf6oSITmWa4P
KnmgDtSDQM1wAQgHMy1liI4cFLvkHKOL7GbSqNhMFzc9HU8MNop2M5FsNQCHdBKONJoY5GpfkCwD
tSzGJJn+qt/R8cWj2QksgobycvAvlbn5OAVPIbIdLe+bA3yzuZEDyZW/4pjltXAzW+MyNRUT26Q2
9jB9nrcG7zUlvl/5jJY6DkKkO5J7LYcH9rgDegGdxxqiK+C973qd8eBcuid/hSCJ9RgRnfGs4HAM
sVVo7z/FmDki/snDC0vDFA+q3gEuXaRWjvlpoMNu8BL6wdW81TsS/ZHsvZu1hF5dvdjk9g5Y2JYb
h38e8C03lWcdiGLzuA8l3tIvzvqeuerub1DiGkatUmVDFEszsywYC+9Cnez/+OXBIbUGmAvH/NZX
DXqLz/c5TCY5fipjLLV8poXuNTFwMQHhZ2wp0WXW4hRVoD0il3v+YEu8yM6FFh7levopzPQcbG4R
YT76XYXG8jhFPuabNpXP4jcttf8b9l1PL1jS95Dt7PCbAGwLRqHr1IArdL6MUHdILflOtlMYTlkA
KjCNREZqOASbYVc4hLIV3SLgQtKZ+YH/6M/H2JLfCDjzT9WW8HPXCBzjH0i9qcfe+d9cNIlg8sC9
nu7Ga+cFvEM1xmOZjl3Rs3sViGiQj4vb6RvOe2Kb6BU8+0ACWMpsBaUimhSGhtANwfXXxLxaAC5H
s0BhJGXMZLA2AHbs30VNW8wDHuI2SgLEgTe0FroJ82j11WweA5tDmvQJVKMB2n8C9ab1xN8BxC/5
Ce42QhBOgM6IsD9n2uDz7FfU2rNIR8JZb8NzI0usLWztLc72nJ3eJ8MWHmU+MkZEvjL3swEEPprG
b+FoHiVyhzq9A98Y9WylUyAQfTthRdFR8Oh25UXnaUrvV9DJkoamp1Tz11QJNnqO19nDvkyN1tuA
PWfmzCRkHaFbyU4UhvD+f0bbhjTQwMx4KUtVibNwhwR6U2ho7On6xHc+CrxzPmr/FchVWukTyH+V
gZtUojV5f768oQ5rMj6ZaI8nvEhQ8elcAGcKn1cZLIgqWWH8QQv+/uJuLzvIq6QObCP4VcWjuYVm
/ujYCMfeZvU8+43Syre1gVN4f0EjN0aMY2j5EBMMYZ3yuXmJHAw9MJbpuDiBJFbRdMUNrLTTfw+q
uRqA+GXXTngbipvVwMAEZA5m3VtJZqdFuWXvdddK9QT2dlVWS6dp+AormnOy1/ibYCHzwE4a+5Oe
U7OsHsJ6kMzSHRs7XqkSlRyANHHvhj5dovmE4jNHdjcwuW71CJQvihTpO/lGTM7LSvW2Zcmlx/G5
MhaW6EmvNTQXxCCoQOkVDpRp8JYSvS9AYLcWEqrU/IOHmofGBLHUiC9RFfhwPa6J4pCoGIGDOrDx
w1ZiquCVCuZpFhiHCU/hSv49yv6lZXpLyY/Moi333pf/OjT81t752QT98miUONXcJF6oOJ1J82mA
LOvDpUQI7+v2TShBQmuzJw2hTHDzYygNM3Cj8EXzW1jKgwMuLIM2+z48KIXeK4vsu7zxCVcJckwi
SNZWl9XsrylyetL3djl3Yo05D95e3rrLcWXFk8kNAHyy9jrhgt63y4GvTq9k+0w931EkJhxUsyoC
hT5fJJkVi/GXKDfJi3iSa1UiF3/XvK/Zjm6brli/yzLkcr3tJI7cqvncdJlF1HGc0rbM7Vo9rMBm
RKbq1QpLyOYQGAsi+XQ/4AKYHQ2JCP/Zf4EJ69eLcVqc9TlZK8QiCbtB5CYZ6oj5rimCn+yrsgrd
ygdzcxYnfVgR2LxYOh6tqhvTEjzL3FgVwGb1Ks59NKfDuCQr4qjqgxCB5YtqnoINSTi3nPkR3Lvz
fVNNyXnci+nC7fLxmaF9x4eRPtIwgxjqK/ZCGqugFNBkiJKUxVMhJ632d23HS8yYSNIodahoo16S
BG71g1gu2Qs7CY/VUpOrtxs0TN230jHq71g7unqx/cz2w2muXQu//pLlyHM9ukCeC36cxvQR+V24
ivcze8GXr3Vd6iw5gtRC8EQ//nb8HrO3XMB8zC/gGdzbFx2cN1Mn2jwltaLgLkvPcbxiUqi5fWg4
G5ewB/aRkg+eeGehod34n2i/jMQnDjEIed4XbksaNxBEChblrEgGEmZwP9VpTUjMJvI9SwQj8YVQ
VHRUYYi6Wqg9zUod4Q1GjHbaTWPBPqEXk1f5mhNEnrcp6UqupTvFL21UB6lG0+dGukPWdwfw03dk
N/BfJJVqrRAEhFLCjcQP68ByRoVCDLRFiICE7MlGfAwW9NAhEfTez/huxPcvSrccUurtQLirrk4H
ryWXj57u5cZBLmGA0AmIwn6ctbxMqfJoonZK0G9YUCbEyNyxjYmJwvOdog8m7AvdLfXTiP7WOpE8
pWnhGJealPFnNENu7zhtC6e1tD43Rdqalu2YSXqUu9WitCxEDeV24F72WXBzfn0zan7pdiizYtfb
ZFx5PfKTF66ju95VE30EUoT1anByNxO6avYEaO7a+uurtxAA/CK8QEGa17s3qt08dr4lr2JWVpGQ
7nCGFOgM/10D7Muog7hzWySx2MjviD7HhfWxqMm81bQj/Tu4wz0g3GLmPgm0UR00q3CuQ5dkEG7Y
40fZjQk3ZX3rxDO66NDYLdmuybHz5ONxGoWIkZSrzvB1RqTzK8YBTYtDh5YCN75GKlClI88jQ/TQ
JldFEzvSGB0GKdS0G4tZzxp6BnkkWTMoVXyQZ44FVFpS+8d9uXUlJZgKBx/ZvuSp50ZOHjAFvsOI
mNg4tN5m75pwhmdMortmeSmPZdK2ni0VQUZp4pm+bqlslSXvBaxoUcrfylusz5u/rHJaJJXWihFA
Advs6pjNajvMk5r3aIYBmG5trdSZdeA4vyhhBxI2osqWlarVbdWD1iqI16/vI5taXwa1szphjUxT
HJcA9Aqz3Dd5XZP5jt6WL1e1wHVSRm8w6cn3Qn0V5roNT9t1EXatFSLiRpfPv50FTiwadYc3LFvz
0kEsNN0baFSPL2LXNSXxOCbb62sy7yV8LShCrUnBx78BO580OPGyfekX7EgiLX0IgWltvNd1WcJ2
MPyAMv3Tzc6HZC+0aAQCUDNFSa/G3yHdU78gUqp/PoQP5ZOWrv3oO0MbYzGXuCbULgFysGGhvqxg
q6SFuNgB6dNnrZzzv6YPFDeLVOAsJUxf0Bxy7ba0siRddvPPNqG3H9TQhxsc1Gp8er47+xanQ3Q/
NiuJlVzhcFROcPkbjFdmSKaZeP2DFSzM5sTcUw3tyyitsCjZ3HWPxzV+CS83Ucq5Me02fD/y9xCW
3fRrQDw94lT2Cb035qdcX7yykh36jUOAZqkBN1t7nA+lhxRaZzFmwOtpSbf3p8vnK9he5Y7lRAAT
+AvYgpQm9mROmR9dlYSlXwJF+6gPP/jCsb/Zv7FrSIa4ILKznQT8jHDkcreNrQ/EksuroAmWWFju
uaEw6G98C73lhuWk6MOp64Ixjn7B1N21S2XTVLvV06A6v2O1WDf2iKCJqDqC4W3t3+/Dc78/8y0b
OoYOFAOpdGN1ywksjnXeWpcAV/OUhWoPHRChggqq5iLwQvMP4TFzwVHPWfS7LizjswCcE9lF/p7S
U5H0+8L1UgLpqDUezLFMrx4j2SNJU82YfjGjtg0gEFIqEJsVYZZj7jQzNLloK5Aef1sRFD20dCBZ
xc/yWUvzO4OMFA1PKNJmrFLCmVJa+Xj5VRdh1M/sEjKQ85bo4+Vp4AAkAyx4NbKxyXSXRoI+Tt0h
szMF
`protect end_protected
