-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YfvCyXpUbamzrSrt1bn3S78QRTWSgR153W+6e7cjEgXivdqlCUwQBjebGEurSF+ZYbsa4c7tYO2/
fGw+KgsB3RYuBxby9Ep1p5i41U3bGWmllHi8Ky1CXO/nVU9/mPcOUrjUJcUwpnjuyJ2bql/WaWot
OGcDbc6YnTXkEXNIkKLiGQJem8Q6rU808O6VpvP0SPd5cIQ4LS6TqItyJntJVmq3NtC46SfmdWcR
LjwwzT6i7CJ6iof/3yJYW7l6lPb6iGX22G1zoV3/xMa2NbDmIIYATsWxfRhVJSXrE9xTOpf82K7b
E+XXjnDLS0QST7nrh1ij/2tAh4DtNIL0QNkGzg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4816)
`protect data_block
pDi/xx7Kj4XoTzAxjQDlbsn0ua57f7fx75596z/Riyeq07sOqvCS07Un5MqnUtAm4J/4t/ASM780
iSEJ+5bY4IoPqGVzGZJ2cZxuyUhUVD+bhZUmGrag2RbMzYHT/wa1cXhSBwGmktnNHu9oi0zhMlob
BBjooppDRLcgXrlTEqWvzeE9Xftsup09t6OJweCKTJATYWpt9eZw5JyucL1SptrJJHWABz83zoko
GS63V6Y2mDw0ePalbCSD6tDTDKZyIkgYgoPFDtU1ETXXEDY5n0lnhHQVwdIAHyJoC67co5/zvl8a
ueopObr9lssB4OekJCG9zFIfrZfBaLMDlmNgkDovO5p8xK+i7TYPSul12OQjt3w14Vu2T7B5PzMn
lIjm2fmQ8hAqMUJmb/aEBmBQ+DhEGE6UbaJHUd7bC/shb1TDpV3vlG3O8CTEvshtmSF6+mQdXV8x
3H6b1x0xgl6z9oEM1QgMM5QteUzJ1X+WZWm9FuTbbK9kUQND4dk6EFV2iGJthtEy8b9nvHs8+VFh
H4OQ/rEbwmyosDZYn8g7Ie8KMDj1oKEgJE4tT9EqKp9KcHdOEzUS8H74kCMjENtRUqNMdWJYMzIy
l5kHIas5KewvUdRdeKYmsyg4Wd/3IaXdYt2hbv3FuDugG9uigU+4phM1gvM9kD1MLMEIZAPsFKG+
qZKNqbr4eoz9eJXoCDM08snYG5/zVEi/ZgEP+fQ2auxFZh28EeEwtijJB/mLsvRaJ0evrYTtiG5y
CkdOS+SbLGXdadj14+PR7Rcln5HbIHHOWae2rf/9TYacr3Y4mSOKIyvrbCeVDgxXS0w3ck50V6Kh
79TGWDZTxh0CXjYhsLpI3jTvLegQG9/kLGd9eFJ+uHRhM4rDhZV7IYmzBfVjTS4JXD/CN6gWUtCa
gmgxOsb6+oTMY/Xl86ck7gXudrr13uHW9W2PTpcJjCwgfEhIPkO4nIXHbOamNJ3kIX9g8m/0AGCs
xRub8PMWLUFegtCKjm5qbbNxHTzssAmXXJITyxalkdmbIkWf1Kh0HJXGpTF+878Sv24fuFu71HB3
6e5TccPfwI0GEnDLTG2FveyiOlB2ElwrNdqrzQgvyRqxr28t5aoT8CRSUwSD0a/23P/TbYPqgIZ2
EGMq6ALB2f+KngmiQynOlFIBfPTmOwdKVCgRoDrnwcKBoRdffvuLfBlOUGTpUMpIonCfM+wAv4fC
BgcEEOmtH7iqO/FVrez66XIvh5f2W1+o22u0UdbVRdlQIogM62TE0/NjJRYxCWhjjBO92MpsdqOc
gh5a0vnhh/oMNTtgl9iBweDE/wOw4VgliZ9UikOhiR+Yac6wKn9M4Kikl7orJkVLwCrejW5uFqh8
53QJrXhl0eniOapPsSdAWz5vPl0Erv9zuWowX9Ecz2ZZDoiQZ9Dy8BMUg+uSQFHQ9tdnq7FtjjWt
CzoXAS19PzKdmedMtnyCdkUBzvboqW0a47Buv9w4yOU4SJP9z/o/6fkKBShuVjMXAEorl8dJMsXY
lEwdMXbdeb3VngvZClrDKcUgHcZnZMhAajK4OfHz7IsYzPnAILOnMuXtzLQBUUbvN1ACPJr1GKpd
SxBK/AfO+DBAOd6f0VpxFsAqeH08D5xhNwUAwXccqVKd8g02P6tdF3x+p0koKhivaIUNJ3hPRFrI
YvY417LSbuOeMMrk4gaqCbzJDNiQiX4q1h3vCYqtEg3zqy2rD8jndVYcQIcJ2NA9wJ8bZHxqrgXz
MXN5V4stRVxeMx9UOCYRhd/qgllMYSZl3pWh7ykOmq8roj+4uR8tlnSbj3EBswGhn9yQ+jgq6OSF
v1zw3XnBdCRsf5VdaxEO+gVn8aZup1IKH98i2xeyXzo2zv22lWxVouSc+QWtNzq3GmszcgNVXqgf
p+doxrKE1AHHrY2xYVbdx25sc3kFpSUSVPEkXYOSRkmvz3UGG7/BjYBv+7nRDy6QJxfpj1Rq/y1i
Ecw3I1+0S1Byfvv5A5+dZLfhf4w+EbTtfJ8CiLE059Gui2K4BU7+FQz6IinzxHHuLWA2OksQSOTw
/sA7akme8mr2m4c9s+BC2xh/ecfopTXiz4O7gZd3IG8eovRiNg2x8s48GuIOpp4KyWxRrNF4qPyY
FyWxqQ9nNg4RIc9XeYihDdWc4uGhR1N335Llh9XvxhZ0Lc0RE+/2pDu0zkyzuVgXdQ41gsi34HtT
Ed2DjQ9WSQ7vsE/CnVEtyOmMDPK3AHw9h7tslZTAFJQwrN3Fkk+49KgttpORu4TT/usbfvRyVGHd
4vPhoUUxVmkxIYpxg5pG6Ww7L3rxBOxTFZCx+/d6/pGE9UhAxcsdBIAd+38jBai95eMbFlw9FiEy
T0m62EUVh1ge42O8dnAX38RKp+ZPZcbW706+es6aKYZ6canAj9Ps1hCZfYJh23b6jBZTJt+7QcPS
3+BjtgLiwLGUIVjCNQdv2sXZE6yIo9H2wQfcNqIV+kMWBPgJ5c3pp05K3S6xkzGeR0JsKqBTyBp8
ezWH5LqVdyKS2PzmTJDxJAipYB7GB0Dx044j0d5Z3mqwqqRcICvB6BOHT6tpyPdhUgJF1Zxed4j0
rSsKCwdbCr3ek6dgoQJu6inWzRNoGdMARGrqayEnLSBcmsWu9TQeZ47Ms/RWflVKvmxEZnwr4G1V
089s9eRCRHX80/TKpe5ZQsFzFI+3x3V0jYF25jlk3BnL3n9EJ0DYndOqdSiebN+4CWYFQh6Vy93Q
5ui7SHhzkVDbGqVhFoe7tJOEGKBcOmIwVmFn0mSbJEYVVfdMM/xThSlcP2TGYCXfPSpC+kyrnO01
ns2U0Lp72i4dUKZ+WErq56k45KnniTALw0paQ5soFIif39c7hjnUW6xJVWDn9zRjWv16tM29t0qf
Pdxf9MncjJc3wd0s6clJYFLVXARUTcmongdrUs1yycDOCGU/ho4hhbP85OAcsdrXloygy6+QnLml
IjSyFYueEmlej47kOPAIwdljc/yjkQOFxb0eq8W0BqL2plhfMyvYn2ne3FNzA6XK6VkWh3St04g+
G+l7LKVgw7UfmzRQQEI01BWPtaVjEUJ3S6LYd2QiNUPCacwEd04DS29riSIO6CBwSYxWJKIopITP
r1x5DyD10mg08gaLx2PI1FSj1bB9vgLf8kocu4tZP0Rrtl7QTCklZWEqjB60Gc07uDihA6+rHNl5
Dgm+OfnrWCAkxWGXs+6i0xQvFxXAT2P8ZKQqeB9UPfFCicLh5pXvXqKwxhVFCQ6XJ+BXPLOfAIII
/uIqngtbbrNzmKqPHDuZxQwRyxOO2kNKomUu8LQeEY4/L5q2LPpoqng6K3U33b/elnRQNt4mXNHH
/4kQusYbP4r76FxEATC+AA8zODxq0bl85aSHmpCPLjDW0RtKgd0Fp0fOVUevDsyDKqYQlUWYC1OJ
0bjs6hu2G/9yWq3Pj/LdMUXlHlAPdT0n1GMiHvwa2sddkFTU6KhdwaJwG12UXOauoBuaqPKfAy36
2wz9J2c602t2fKBccM+oux9rK+RFrHClQM3Twrq//tWaa+8422GAsqSSTJ8UerJNUHvGEK4ZoXtl
oACBylYBo6eozUn16+kpiav4KG6mKO2plpfr14BfEI5SYMVUk/wayjDTP/uUp9Sgw0n6l+o+bL43
K77Hlnw+Xkmq0sMtjI9gSltxawaR1BXyeT8ZeDtWH03bZpWVdNiJQblOnFeNXJc7tWz5o/QJJI8c
w4dFHQWGZXmh8xYGQF9EWSkaPqYszVMvN/Uvx442NftAUy8LHQnxC6jMHQ5rJYbUphc04A+dyB3X
vReoaiNUq+Quk/UT4gN6zpvl/k66179IPoXrmzOYtTnJpjrl9e4u4+d8e+acAKJpkBSU9nQqJiBq
gviikXIHVn+Rk5+qOXCnz3Pwb6DXBaHzpM2t8yBg/wBUH2whjrtVE6JKplcShhi+9GvZbPO6luaZ
ewYVkxvY2408w7xXpwoVBk1UgVgyFf1cOFba7vk6Y1+Ti98J1ioLPRf5zjuziCUARYrDrwayox3i
UnztJWCr9q8kQv9+nDcx4ehqqJTQRdnFS2r5wjdvqAp5krxUz5ttgVqNfJawh22fhDoH8GMdKsyK
HjW5AtJnJkYWBdAlz2oLRqISFBZ+ucG2jT9L3ROVh2yfbIRB2vM71cW7jqoFCbD2TtYKCeT0/2dW
z4l+TiWDA8jVLT4nEo2rEWC7+CEM9oe3n8iBN/08arj0+KRL+T/t7qIlDnYeTowz35+V7UpgDmDh
tPh4WKdqyGRnV/BpRRn//GJzPYayCfuQ/lGVMX0P+q01P8xsEhGh37fCWetW0CuHaVBGvGiDE1j7
QGSyefuY8ECpFodyIxHNpNyMcwc2bjCuwj/t7Cy6yOk+IHDLkRwodwKNwRXOfiiadL1269Hgt+Jc
r7hRCtOwEzXLYQKc6jcen3wqwUSUx3hWaQ8SvtfMhapyi2vY4zt2G7TZ4TSPSc1xmka86/O+Dr0o
PS9ZCzmny4iQb4M6N6x2bStfk6e5X4uFvvD0CPqNzcC3P6sDXdrWQAJ4su9tY0B1EoPhGAo074MS
fw+u/HJOHo4Kr90nT393Nu2BZl0EPpN0j9UKQXTPoJu+JU5sIofmPG93j8acOOj66ioPnA79fY13
CFXZQJvhv72v52VGtiLhWEivPxxjrcmRm9Fbh34IamWYsPTcFyQAqxxvvRM/m9a5ghCe1Xu0jcdo
stH2w8d51B23fU6BvGSfkUmujKYZM1F1Q++15uUya/P9eD/3VHYc2VciNYNo1c+ybfE/G2k0YE0N
fnjwlxFHfN+wkpo3bBr1RIXAcqiuetHREASqiwG8K8UNfRZIbZf3wJ2tIx9xuozogNzkRB/4BqVj
wrm15KEckv2cDTourYK015yuCpw4xDNRmmOVG95niQo2FIXieD0c8vyYyF+1DwE72n/8cu1iJtZE
23bM4wJW6U69VOPS9gsQLBDP1xcd1dUnOB3myTGDBvALySPoUPEmuivq2yCjb2JfcRBxnM/FYTHT
3jFbPNO2CopN6SEdqAdlI618hxshaOpJ2UrMk+j7D6rjqLClWvhWBe7DylHzw3MbPqoykyEGdGUl
5W9vOeNTHpjgMIekzcudxJjg/7fXoave6jMvPk1RdDWFC/VZdmPYI8EQHgQvbE/CnsWADXu4ZiIJ
PsSjwFrYDInn/ASEl8cTJD3Rh87D01P4S44zz0Y3ZPK/wQOLIxS7ZNZUT5TwGusN77wyOmpvRBT4
F29gnEMaJ9NiIZc45tkzMbmuI/M/iIXxRuhXJA/XQuohkHapM6I9ZtQ21djaS3Whku3YL+THhseU
41xDqzhmHPFlTUqNk0iV8IMFv7xJXDSps0KD3qus64pNv2iGHTczuh30DEAd9vKQqvUGa+VaPOke
X65A0xY0I4TFM9OOOd7XzbXZZEJobzKAAcqf9wsWRT2qS0AjC6dIoTPrM42Ixu80YqeR6kncRppW
nOf0oh+nAitbcuKWgHcf9kuE3DqRPsMruZ/Lq3nBcCh/bJTyD1OHWhx0VMX4UFhY7umx8WMlAwTi
79kD4BiuRRjaZElXOYTSHlyeW3ePoM7C8rmxO+2k11sfcWZFI7X6INgMoExWb8ODwpF1chL+JgAu
O3S1D7wZNEmVT0Thlpkuav5PnarvQeFUtE62MAWTqP/AfwDog27Q5j8939q/iYOqwgaMYCkRmqYW
0WWHB0lZFjlwiW3FaXtEuJ8FEpp3PhIxdo/eL8U0uqs0737lgWyXfh3Y4tapZFLvtuDhhq+A7EjO
8tY16uwRC3wLGajLDjuuI64HEyt0+brbvXEoFwO33pyOX0lyyE6CSTm3BJAI57IafBNJBPRQjMJ5
20ycsUzDVoEeP+6dimMu4yarqQuXYDKe876DFhQPuYOQot4cY8yEeYW6Gf3CvXIUkQXaspokdMDS
1I16ON6rMeFZsbifyIVg2WbZ5yoF8p92gKtYH6n3gRxFEKLtJVGuJHkM86hwvHxe+lIWjQZN44sm
WKnjmnKZMvpfETpOoWWHAHxfa7SGi61rSdtX8Mk7HIsJsFBNdLETFjJV+OBpJMDv4wed9q9Tf9ZF
WxYgS8hQHgRQQg/+F5GjnNskrd721AgnmdVBa33RVxGB7tR2FNzrtAjLa/CpcJ6zrQ4FCy3HYrm2
yTDLmlXWx0LJ/a/A8gBke05njf/sIjKiFMdQc7dfS198LSx+qDdLBZGfD6cpYQO12kkSoLavOK/V
/4haexjcbn86tS62w+lq1pYYdS0o5fNCtJOr10UDZl0YvV2EGYTEUcI+XiIZ63Zy0TyITxZeSLlE
kLSwrDfBvqr8QqpX/EzXz7LJVxGGMapA5d7R7IB2oDuBYIHBwLEs82CJv1yV4BJ/7gJRwbhv76hi
8hHv/W8mfJJmU438rPMzDNIdiEirQ1Iyjlcjjw==
`protect end_protected
