`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JkF9iExS/PCmaAcSNRTtUXX8huDGrRXpVKN9Ulj/0cAE0o8q7+V9xlaBnTd7OHwT
i4pGpbfwYSJ0sU/yLsVP+gOaiZtFjV/8YHnRbaezujLEtes0esiwWjTxlGB6qSYo
xZUdb27EaLwNnStRK+f0LuC9Ig6mJ0S+MpHu0nfcpH4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
ZeKbZ08fkkJEnp2QZTkjvVvuESyoRKsUaR5pEZ5iD8/Hc5970WZAO+1hDiWDiNbJ
xv2ra1r4DzUoN7hR1iloYqa7wUSV5Nl6IcjjHJnu8um03+ojOyz6Vc3N1cKL0Sbf
BXwF4WLUFuqKYkfMjt7gHbvth2XnGtuPwzOUs4wahxw3ft8b1ePeT/z5DIdX9XBP
Wysxu4lKT0JktP+FGhFVjhMaA+AuUFbSCGivxGzeYXnERVdWA7f9JnNSkCcHm5Ha
1E3/sNhALTt/cD4P+fNIqPkxklwv7uJstw/1DBsXWqpy7spze8gcomrPeOEt8WjZ
t+Pgsw9xzk3hJVcjrlhL0QtJ/wBorkLav2ssqO5/rTdlbKKS6V5qYwxrGeuiaHD6
kc8Io5KkryuuiYFXoUlc+EBHvEmMhzKNjyWF0wBeit7cV9B3l/5cPzfpjMzFAplU
cOAOUB6o7CdmsDk5H1MMc1XJGBrPqHDd0tQs2u1/OYajwd0oDOMKught+PmBKrq+
BMC/Yz99NiYOlEEI/36ZoNIuvePtoeWZL5zD/9QCop8uF3XhPdQW4iE5stwVu9xm
DaYFfBHCu8k2MwPwSHF80sqV1OwGf9J5h0o27FzMtguFTZJpq9E5m0tSwlcVuTJC
JuKNLNU2pXifJ04wouTJO9NeNccUwkAaEolxjmwthFuSXoD7kERVmONmTwflCREW
TtUb5MNtrNTPuTUTQuI4v7RaNPl+rk+Uqxrphn43SsMEOZnEglURIyWWaSthWbpc
ZbSXyS/6zVoax7iExr344Wckmt/1y6823md+2gN3UVhV5P37Bjy6bO99uPY0tUZP
PNI9/GqhwS+4o4kVUKoxxVt1Qysi0SxSr8qwCkzXKMAylPudcrOortVlL30LxBSq
OF33jGZEsAxTkS5EmvAMK7tSCHR5ghQAqxuLx1fM8LdycS1W0rmuE+SKuLLUuGpV
IBHkuIUR0syCGyiJ/GiW1Ai+kOgds3wXBduQ0JvFhcM7ucqPUhWlEXPtANxome24
dE1Asj5Ix3/811hGRFMHRXSgTXVApEjiPNA3Sq51Z/Yj4dBoc/yEKXp2qMMnmA8h
1oKtQ857h7J1TMk/cPlwyy6AAkGIpcTas0GSFhW0PImqS7bc512LmqOAvWpKvIN0
SONsgJ6+7023oTWykkbbdQo4KwN3o5T2yRMMZJt+DSvsf4+6gT3HiAx+L9vEsAQT
MvDcTYavrc40HVKrNyRdYSgWrBOdTkGiTWpJsRHrWy41JI0qBB6nmW31dOkeJjTZ
8dmeIzagTDNfXN+4QrGFOWZ6+29IcQhGM5pg6/vk3bY8kqzVjkC3ftvZZfPIkHg3
qK01lHvNaKRtbD0hzCQPHwq6CWXse4HW4ylGjpNRXlMhA4kWjt5LNu6XCMGjumF5
MyWO3VHhNXKcgaNjVMPUfXA8GZemUYMPPriHJUpNMrpeGFvNMUVQ4K07Vigqk89N
VJ5F3eQS8eS+m2JPRbLqm3Zzb/feLHM/yKspbvYpkE1b76758R1tLGTPUaTgb9Nl
vKx2J4IlHf/Ggeb9upGF9sSgRMcIbYgHtVGkbMw+yjXWfMFAhdEvFspqq9llLCjZ
FbEU+BlO4WZoa0YP8tqfLaW5zB6LcJN6F8opdIzNbvJjC1uE5EKiXrdY46UhP6EW
7dyOkQ8teSC0bpAL27oz7gaaJxKiQgd2+ZlkNSKjb3kI5tXWCDQnOk9lJ/3Akm8N
8gZQyqxpzEh8q3K9DN4ltixoqO6t7+LZeQyIWxUej86BoC8XBkmbqa+uANFd+pBH
RKuZsj5ryRK1PLO2U8Bf3rJjGoJ7lYQwCfWf4iP5F4/Mwr2Bwr8XrU4YpkmGtBdm
6SZDBt69Im7KvjI0heRlUpqKEdhyiA+3lN3gYuB/ZEvLj1q0YJMmt4OkV8eWCkce
4nMvvA+6Y/SCleNiTeFU7uniHEVML2AUmSUPb3Iey6/gdhGsArhs/lsjGJlwTyo6
GiG1hb54zF/wT63CpWsIKz9QSq90ea5gJbbZR374t7X3jbOb6v71mPGxeFIgpROC
Tm8eEa1GuMF2cKdrXIsmfHGhsnTXjYqukgvKi+AsOvWEK2LW6tNa9Fx1ROaPdeFf
5UM8UPbNfYZD3Ajjcc4iORv1niDKumNp0UliQHEuSceyvw19aD74WPR+brKfsvfw
7CYpybu2nLW5MFdskxzBxlN0BJwMXvtzfwkwnHOpwZnl+aMAs6XBBHITHCyFjvOP
KPJrA45eg1dFmY+AxhDUnEfSwOAiKktx20tRZ4SY5JGieMTa93FhwFsYLq3Mkuaj
Yrv+2WTccFUBjirPQGA9IRhVB0z0x3n6EWqJbxq3ycKyfkvHyfWpZYztHf5Ag65b
pJZvl9T04cwD+wBwizI1CH+f/+eGz8ZVPHXA1dvB8L+dNP3DGwB5yJD1937NIlGB
60a/FExXk5agEagWZQVQJfrHw7pfsbkMmDenMKf38x7vzHLZUVvM0JzbG4RTgDQQ
KUt2ase4ceqL8RSUPIPi0B0QbyxU5mJILF9CKd3brvVt0Twxlap3yN/TKVEMlo7k
Ys/yKypAQSBTpUyAZkf64l4wBpW2pxI2yd3tXY9v6GcheQe4IyPdGsW8X6EpeLp7
IZ2ap1OPPhk3bakRT5EIdQMyO9gqBoyPi0r3CHZ9m9qIZTsfrcsxORDLdMv8eNGP
x9g013tAHtX0kb8hcur4KwHzZoyueuqOfwmVRla9O0ovWj/nSNshGaZ8axfqapVJ
KApXOmNpsAtlTlwC+Z0mro1gicYeSyIL95XXXmmEZlN3ujzcBphjTeKEdA1mUXRl
dTXD0MXbYKI0RWd8k8QpFeJYOCMj+AmKEixhbT+C+9GSJ2JGFgnjNowRymL5owjq
Y8Lq0hyDQBcRyfFYupYBFKoLJUfG4B6Odc0TcNoK8AwfKS3av3z9Zh67CewHygrF
f0mS7h1Lt6Hl/BsjhNLFM+e4Z3d4Y1LNgkY0XFo9dRHHNG+F2VIE4n+oRUjLZgIA
U+vG2NQ9TjZtkH53tBrM6FDeIIk7+tq2RhnBzecHf4Qfw2OJ8L3siicrLi8uuqZX
vc2aFxxKVpYN0/lOsZaXppkK/xIqW98VEOCgF+DBNFVMhngF777gQKxsa5I8PCy7
gieTUojDPy06ch/kNnuMAP7qUbq+ydSeFylzl59NMNwc9rzeP2h4y0W2fZQLSh8d
qb89zomukvaxfp2S4z1EUkJ3EYIrfdzvLc09E+/TXGmg1RT2C4rt5slrUiZlLj0F
dLZwbLJ/8MfIbF2S8c3nd2Z9CGC6x92EMuG6zvgx92VhV04F6fLawI2Rq0q8qpEZ
LTSU9nICPltM0Cgfpq9iaSXQMoPkr3QQzFD7SuiPgB3nktv1STh2wgtNVoJfTjyb
MIfiZU+qrho6Z8defxkC+5r64w2Yr6l1c5Gie8cwJ8Z7xdI+socss19FPDWHOGF3
hL/ew+ytF1fhzO9uUFeTryZM+HG/yGxHRkDrp9yJ60wFL2wU4Kmd1WMc1EznSB5F
GMHKEibDiyh0pmAGFnlGNCWec4ozFb9W31+oPrhYMXjRhEcj0Azteukjl4Wg7onb
0MuILfkl8NmQhV25Oolb6tneS1gfCkidIEd09jf2VYf5up2qGDMqJ418Wh8JamLB
E5zMuQSbKZ9XB+Fn60Bd2EX+fbYRkU4P6A61OQg9+eIiIGV+XtI8Vc04wGMp7WqY
I78vwiFyiEHw1hBEApWNpM/zp1v2XIGqJT/2s2vLLbMgeO8CKEFKQpdL8Qvc3faE
r/B1eMt8PqQIzbwV4S27abv1tQo3Z5StCnQE2/qC9L3SYEww5xTbUNTxSDBCugoQ
Izyz+hF57VYg/NAaNnP6Klip0uVxz52x9ujM2+OISHktN7a/paK6E5FKjUaJ7JUE
PHP/MZPd5H0z55lOx/v2q54s1H/oCetN70K62U1Jpmc2vieK9MyLbTCqja/Tx89U
gNLSYd/haqEiuPVCuRAbnp8Ihpt8hq2q4KltJ2P3f8pOIuHbGPbkeqj6wST0iJHg
uPdcr1Og0/w4C2tHwKMzZrx5BCYFzqeHbkeO7J9O1g/qLqtlpidqEBcPNxYgSyiJ
FAX5HQvVZcCooPBhjfNwUoVsfaoty2qRjjps/gWj8nAjaeb38StPg9OP7qHSSAZI
Vv9h4563ckjd1nYQROSXjonptJkHE8d+C5dYM+PmwTwNhV2zxQUH7XAP8VLaAEuh
ABrz+fPrqp0wSYQSG4eR1EsNRXnLSLFTg9b9uJ0BUmEWghDuZGedpZ2TkD2/7Gtz
puG//CdEXRGjO1HGYmNV4PP80H+YeGDi/dzumra4AlXxrdGTu1g8tHrHjvo6fOED
j42c80K1zyw3XDmukqtqB1sdWVRqtj/dlsn1QsSjIrCwMYta+AKVSQPcvfhUN5qf
cJ7ZUw5G+e8sf9Et7xxrdoEoh+bg3FStJmikZhT8tXB+XAdMD2vELi9fWOAvh5du
vkVREHMwSK1atRENRp9Z6cZO1UyrOQQgR8nxIM2Di2GWocLA2O1uKrqrT17BmvNE
HZOfSsDZR75Kp+PU5Z7F9Z2YthroR2At2K/CL9iDYUIpZjwyJMCoD/93GuYdZH1u
6G1sBsYrHPcdsLIkbzkpm4RMA0AZQZr+jOKoAw6vC1175DwGTBqkK6IONt1Lo2NK
18gVGGr2mABALyyJiOCndEnkdHBA0nERG7zF0kZmeAaF+QmJxggP6S8luknXix/k
mVlxIgkD/49EQKf4bEJsA3TJfxT6DcB3fw56+doQerPwhXd0rEleHu/yhs/OysnR
rppqWJAPmEcqD5gwasLx7Uv1kWjcpXM6FSOhr2IeRJtuKcSPiGiZBWXfuzaQe8U6
li1FEb30RSe1QweQORzCReYieVmp8MbSZyF+siEu1/kSg5JJNO7BKQLIK2TA8Lug
q2BPzzNf/MxQd3WNE0ZbVKXtse+WUM7e0nm6p4PCAOvowbU7LiUo3dodMC6dvBGZ
8eMRUvHDNTHVWfgIXurY5sSHubuPzcV1wltRWYeaf3PA4cEQlLjygLsp/PcLTJPF
D0zf2x/+05GvZGu7SnB6Bl0uXzXb9nOsiV2imX515gzMeKOx2RvdKN53gTuJndGr
ACRfZkTdFQC9E4tB9Y4xP8MUmmi74hoqfk3rsMFkgbjmVi1QhyvjYlc6OYx4d+UL
+EJznQaJ7TQWhmDJLPMVmRtuOQNxU5eNmZp1ucbllZGN3fV9zDY5d1y8W3Y0ZgyB
YyAZRiLwsypjssD+xV48qUXqFQRskhEg/tNTjdgOytpHoTyDOpUTKD+CXQvpegtr
MeA1WGUZQusHtohWIQuYgobbrZ85LUEmUHS+Rrhlbs0m6/c8KGPoChRCXX9uf5em
TKlixxV8XyfH4HfawYgHZF9OW721bXK8pAexbssVx3Vlopzj1RadRbbJRStUXkml
4k5zoEfLkPVA+L2nyjgSy/KO85W1JM1aN1meXvSW5L0dlTF8GUveshUYf73AwqjJ
VlLnOyayZ07vlBgvQ9h5E5RJQA4TmC1INDCo8QXcynB0kx0+/lzKRbURGmMoVJl5
r1rNiHff4C88nY+zn+GEQbzl8br0XhUVXS+C79sADfE2UFnQ0Tn6INb9DM/WdwMN
0QeI+RWqZiHwkPec8zeCo6SAIgeNKqlAIZ518cR8V5Jr5wrLcIMSgqG4XgjI/QOV
JeC7Y73OShb9NuIrYDwrL3CkJcZlr/mBY8CAzBQW9PRKOtoC4V8kSRXBbQIrHjtv
3fEmn57kp9FrY9TGd5L1/zI1fAbbd3TiVcuZSDeR0NkKS2YGcpOuCM9TjbwkjGtt
pbd2IZmz07hQs62cy65jmfxz1D1OF+rD3aZvCrPdzvDL15vJjDYxa5Gu9MGHeICi
8AefBruZW5UMnhGwR2n8X7QGi7Ytyx0HxWMT9WN2OLQ+IuclzJNXLuTPQLwLOB7t
E5VrHcOKEmuS4ys9k/rm5WUiFbPZuBfl6SCOHIJ+GtfnkhozmmJgJ7ogWNYvjWjd
L4lUUdBQAh2Xp/J0G6/Y1TDTRJW1MHffJUTznAMoPBp1PPaNdCuNXqrT7v3Ggyk3
ZJB15JGmasYrKeAZXhxI+QjLkc1UnWBpl1mqyPpWSW+KGaomitqzLk1Rd8MI5y07
oDOKq7LL3z69w4UhQ3ap8dTxfkT+QZRhhZYPW75d/zLnfhvhfbh7GLg2bhCYl9hk
7CLBMaWfSiuJy7k2cMZhNfInLtZJr2+8mbNv7vkzrAUfhGITNsc39VBOXyaN+/5f
4om3HUxYGMI+JnITpeqPffrzzbxFnW7NksgyDK1Ost7ukvq5EirNMgIE8NWB5CrR
4BJjCD1JQLWy/twS9+ywoAU8zxvEVCveoidqE3Ix6fHYQHdDERt2nwq2IZxewJxk
7ssZmOYPunPH1UlgfvnPx2i8bFOT+GiL557lzu+58BSqVxr2gsyaIrKfnfpY/IB7
e1JCABFy2KWd4ZTf3PqTJZE08dZlCCpS+zblGsOM4zhIR6XFC628RzLC+ROOqV3E
Oa9l0V9SaOpCUhgmySJ6dbPivO5EFKUAG68zffP0Mw1X/DFfvWNN1q0pdRQs6zdS
tAj2U6T79QmE18dzHCqs+6DcQSssL1YhZqLnGj57JnHacuZOO1rIw/WhW8rtul2m
Hf8eWfAV3KAZZK2/8IzBgOgrroudKaKEMFnHyOskW2M4kgyuWdU1itrVqIy8EKH3
9rVaab+6G1Oy2EMqcfoRzT8yUtf1jHf2l0d03Nn9+DabNyQ1a9lTsjCG/ZtHqi5n
mcAFdvKFcUHDV9cs+IZ75ndKeI69Ope3ifYObVF5nTJdocZWK85L5fwM2UctcX2t
43j2vc4Nhp1KKojAyBZOtfr91h8zRofXNTO5gdOrWBhYJmQ7CozKETVed5vyGs1k
tOnClm4vAqD7r0E6Wrq2ws9w0Jw/Q/0c3Iy40d9JAMFjikP1HHAdPY2kV2uoH0Sm
Ef3Bt4DtxYD5A76ex4Lmy4YLw3OOxEoYremowj3KxSdPI9+UUZi54REgv05Xa1rO
1biPS7DF3FsV0HxDNPgjAPoprBgyo/0l2HBu+YwH7U6qAEiPfBnbQtYitljVdfSY
p5d1jo5JwZqJIU3WjAcLLo2JwDkoyyCGjMB6zYGrMjmJrZ5gwCIyrc/RiodLzpkC
pTnGIaqzpqULS50+HK9VXLWkG2e1ao1kyIqAxvT8IaqVXkOP4EUq37rY3NoZPnyS
X9t5MNqLVyxd4xKCCzThHybvojjR9GtEOc60OzaT3svPiaDW6wORZms2N+WtTVEI
/vQUvakO86cT44yAnE78OalzZ1GqubUcxhaRa4n67iwjMhjCUwI81xiyFDl36i+v
RTiQjQ9T+/dOm7ZHRerU72ZJ/O8vU15IVwCG80ui/+fyhsJG8fQcJ9nA6S6/FUsS
TwceIfUV5G8JzWxe4E9KCQ==
`pragma protect end_protected
