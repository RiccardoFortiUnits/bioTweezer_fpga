`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
owp0jlBR760NxhBFeRgBx4i6+R6gyBwSOt058VQLwfez+CsxtK0bOucSeW6EuNmI
4Luz1SOZtNcrSnsbFWYImfUg7VSOJJuaYPjgJmyFh6eI+h/7jmH64TYr6ppoQTla
/ehiVKgALLZRkOScA4j6ABMDXGBwb93UiC6hs2ja8TI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7920)
NNwTST7K4WcD0rUR+OefUuXJ4UnakKnIgFTDrqQKu2EP01VdNaFbKhMieZ82yu50
sWRJ2NBLwwWTJ/tUxd89Bm2xh1WpU2pXm2MGN1Fv7P6UwNJyalwi+ajJOa8rL29g
g+dwc8KlzltwNFKBgYWgnXbR4hVitLJRWEKBoz+JxYNSHaJOjBFE+VWmFrmTC+g6
surxK0VYWNFjNRuQvd7ELWi/8UyFOJblvRLszliUAF05s6Os7IchvlxOuXauXGAF
m+qAZhnYl36gULA+bgPrDcnKUltLhEshvgmvFoQUjaviYe49u2I8Q6/RxuRVl1Nq
UF0Ev4L9WWln6fgjq23eTuhgjG5rMcMQQFiAqIl/pQgMoLADOUzi5S/jJW422WLv
xFIOJdbDGDxj2vBG7vJwrPaOVoiSSxzNi2lpbiragJ3qsd1LIfhYIoehhlqhtKkd
659cUpAB+L3Cg7LnQdBnHLdB73jTWxXrXSpjcZnpAdybgPRD0CuWOh0VkxeJYoQ6
AHiYiFXsoZOWU4eKkDsMYrn13Li2wlT/XMaGf1TUx83XzucE+LRCm7iYtI/Eutix
hTxpQmyZLO0AwnFqgKnk87ZUMxoNI/v1kwHMtUkY6cXQ3NDUszmHFEsrGW5TKbNr
2gc7xC94RkFQ2Ufg6q3xNhMfH9i2VRktvUGOO0m1TXhCup8YPnIDygaowhsiIyst
DVYArtDnv3U2q9EeKqgx5NSnFAdepiKbhUsiIsuIJDCzh9WGAQOpHJSEbF1G9WOB
PG0mNPnIW5WbQrFkzBHahoAmoFfRSUaSHj3RrRAHlMw+J0oopr9fDeNQgbCYmjqK
pDzzJCnaI2ONfOq5xplAs6/qjRpjFSNI2IxkPRJwWhdMOFVBALxgnXv777ep6xRq
FzXQNkQr6Nm0r59ePk787DxipHVkwoIAqomLFXKKhbKHhL+JF/XhCZlKfSBumMME
Ub8HOBVWfQj3PTnBgFY+HGWJY2hYBn34BO7eSePzMxNCgaw65wGZ1I58P+OccuUw
3xygeWnJmMwyeDlLzFpeLX8Ni1qrPsu8ocEmLgK7FKMLlj9zMFsLaj0wL6dzU4mi
H9Setv/Rcdqx0wFMSTnlZ6D39z36xknYIX4M2UuiQfbdVA9AoNJFes6nnGnz5fi8
os5HWqu8Ut3g2fnx5x0svfVWBCqLxPNbT2iC+yPI5GBe4DfoE+zTfg5N10pZwfBX
gvy9F2fte++QHsRtKnDqhNz0Xp3N2SH7OV5hQjV/XEArQC7iEOZ3sjSOmvk6OyBp
WlIjji/+sb5Sx0J24a4PomBIvZKp/C94NTSAoSqeBRgvro7zGUqMwqhDyaLLsDtz
HyM/5R+sAWMyEwfUWP9H5rRLEaOAB9HpOG2/hjAuW7DET48krF1Mnua+YinpuubF
tjj6v1EDrdAdst4h9/W0Ujidku59rEvD10zYP7thrYANvECtQEswUAg6tRZu+MkX
8YA3xv+wWbjfy3n5smsYQ/NuK8IqmiAW72Hpe6vP7e+LUhqM3e/OarguqT2YpF4R
HigGgKa2ghaJ8DRkhwub+5prNn7c0DCPPYcjg40naRFFMd4wshv4lKrgQjQG1DI0
5deevLCl2n2lZ1AKg1FQtiRVd7TtC/JUAuKjYi7XbyfuqsiDHPOQ8m04ZiP99b/r
Rs54vEYFxIp9zN0yA87RVcYfCZoB7VUYGMVAu3K9SVJM+RjU57sf+vhC4kb6MrUI
bOZ+dY9sYyeiBL4QhGjlBTS7ua40qYPIbgMTQtg/yaR3ni4NFbgL12xrBWll9VHU
IsPtVv4ZoXyykJTNjzx8rdUBQOPRk7JtnfbE4SgWQ3PETp1v6PVhdgsXarmjMr7W
McE59ydfM9N8Y6Zs1mPGdbuN9yuHlDUHgQSUWpr/ouFD15CysA2ItGj/F7TnGXkd
V6RZYP8P2irOR2T+Tak4fzueozJ7APzSt8tEsf1hHCSn00SH09mUiFZk05UJvNzB
NUVsjVmM3WPjETM3dOBGA/U4fjFDwhC+Vfe98hw2xhI8LieAjjYGz6sRVLN4faWN
LkroupK2iopTCICrnsW26x8PUuZkE6Q6xzdfZNKnHKtgf16/JLFcCLCkiVHt0Bvn
d28vMOiEupd1UuuVecqCqECMCwpacpwAVcaN94guc7HjhJS3K0bbjyvi05tL/BUi
zBnqpLhmdcT5HKQImUThO7IsOV9YKtUg4t3lO8iHGnQMPdL1osUvWdbZsIJ1Pxnb
HNEM7w5+YoQO8ZMWpVfKtz9w/CKj0hO85Oh+Ss1DcgD6tHpwrJT8rk5rLhy2Orh7
WmhVv45E8H5n45wIluY0hPLYB4CfaPLf3RGrQrd/GpmsIYhND9BJ14r4POUCsMSY
VOOL4jobkXIEGXnzrmF3aBGo/Xe/RtzZu4tKJSnjGPmJM03BYRWPafKkcnFS7o5y
QbJZyHc5Jmg2WAfjJIHeDej/CTc8EihAsOcqPJEVwoeVRF4bD748XP0Ku0TPwAfa
4nkB8E2FkLdXtGwDxqACLudgzDkp50Y1d+nRBoCflXu1Cszzf6g39+6fyVn32IRd
LGWGk6N21l24hrZ7dIb6r6tiEhRoG9PEnNi1TnQmyKuOCjZYf+khb1KD8YIP+QOX
6KQBSAGK8Me3WzAiaj/lQ4K67exuVX/KA75BceydrQHTHWYCuTlKXbAWTDk2KS3h
JzU6WtngdySkULj4+The3Wh0JO+hfIDiKgcrGIOy7BYfxJJXvW6PizDymJW6wAau
6lK7DXtXjbTJUgV5rps9EADlPi5TNdUQE6KfOxpHHNoCX5JpExKoxHLO0z7P07cp
8DEqWo9Z7p0+sJupLNrjm7gABSA1/nf/zAQt4486g5mId+qnYGwqOIGwmMcziP9z
2dHo2hcxhg9XYJuCC6rWfUkn18WbnFLpB7fMLnQE2F3kqbiJd1El6HzW5uZH4bIK
eSjaHRUJfOxA9KKvFlzP256ogOTk2ducqVoMkGKF4pW8o8DpmRP5ZEwuMpJVh0fB
WPRDJfEgZBiLW/6U3WMOZgIM7GZ+Pp15+bXJ1lqjYBg5XoZA2LPUyhdSVyXgviix
hf9Px4cL7bHMNCt1KCfwNO8f3pBGaJKXAPgFuSFAdyE0TBm9+1RfzVzfsdCWH8CU
zKahcbMXBZy0wnYExFz0B/w4sGEg8gh6CidNPJwy/WdNS7OFlmKadilhAfvtgLoB
OF3+y8nzjfdfww0zlB6szUWaiXRyVJLgc/SoNpa1i8VoH664+IZ2d3f0J5tjcwcr
BoDnPZ/o4L3fdO5E9GY62QIqSEEdgUXN4J2m2+Zpwzm9GmASqr9fwDuIQVXumzAw
foJ3meqSF4Rfs9m5JQTyiWlsyvnv01m4yucqekil5R63SlEe0AmQm3BsKiVDeWrY
IRkS6LbmSxf9OvGlRIbvEFpsbEMPVdp7I4wChChMVWLi+Z0VScDjESJy9qPZ7WDa
HChvFl2PDkc4FwSfBcNK+kORY8NGbzHApl+v52mXEwv2BNpu6I0NqWSjRHOXnqNC
oM2LqRovn9s5mV10mD4JO7NBrJL4mwueL5DN6OOzOjVUrgbSW6iO6Wd7FeMQ7PAI
U6+5fCadTnI1Skr0cCwoLpJueEDGRWYlg67qHaNkdjg40ywm3FnPaeHpIdRRBteB
cD+4SgVko21XbPqadHnLirRhWAIjo3CQgbhpBxvNe1DAD8fxgPrWgkapyehh/aZq
DZ+d/BaGMZHZjvQNOtdBfrkmDEiR1/vMa/+zyK77ZZGpuIuS5JcnpP+C1+RsHxzL
L797v3olj1s5aEpgysHvmrrRm/wSGTy8EAOgXbfWg0CTFHjexr7zKnUkK4cKa2t7
gg0dZjWmOcJvn3NCvEouX853zWwcLYP8dlOrdziV+YfOy37fE2X+37NAxDWHh3Mu
apyk+WXV0v3fu42P1p6Ujmirc8aS6E5CDJU0wQ3joP4pBL3f12WFYvI3MHfK83HN
X97nuOFk6S8KSZZVJIB51flN4aD6NZ4yjqqc4dSTyxDczE8HHXjQMuuuHUcEfNS2
IDaIWjoyepuHYeYUsCr04rpcIW/eA0CIyKIbWZI8SqG6fPlRAv6OvYVx4Cw6sk7G
Vc3mtjnmfZbd0R+CuntaL8hurzCMYQr3Q0YUvR7AMVSKNtCaepl25z+5DxeL6XJi
7g8dn3tMQUiTNgrwrAugvBVBwljv+t+yPlGC2nCq57z5ZN2jXB5EblOAGtx6T13q
lJUqyERgxTaM2YpdY+ZefNuSwvMJ1gOHops56LNF16j7FOWb6TOXnohBK7lJFIVi
s0BEGjZWn5TI/Zg3S5gBliH4TjsxotFMoIceH5JkP+2rvFFLQmvPLIk1Apxaq41E
sJ9Ksfuah+fmRjP6/1Si+/6GC03T8PWM8cWXSJGRL/4Q5fftY/2IXhJe24YLj/s/
ahiVJ39TsNSSDWEOFVK8l4NnlP+vZxGHI+1rD8GPOeymUQybGNpql9F2xPsZF8pk
0INq4y7ZUSWwHSAkFhYJj+RuSuhYn8aNphoPj1ilBle5zeihsU1PTHC86jJ1zsBP
sx2gvbkRzv6zxrvxaQiNtTO31PcxmPmlV2S82Sw4GgHyadbwrXCiUILsmqINdPy0
sTOItA/Wbt+jFjDNkd7O5C1Sj6ot3tdFn2FpMtbjiRnKO8oOC+djK3qf8H4/Yzx/
u7bAmMpl3+00RuKG3ZOyeaRQTAFKUVsyEmUJ3SoOVd5oXUHFXUN9Knd8mwA689Ig
+nX3Y097foIQKZZO73e0gb52CohKMVUJz+5XjgF/ydZtNtOHhKRalkshllewGYhb
DZ0ZDz/+2gv84XjkskrybX9ov6ZnIV+xpEBE/FG8jLjoSZ1xWT1hxh1QD5VC6EHf
D0mYe/t1d2J/AHhWFrb1vTd2lSOxyVrDyFbbk3/4j7Emzl7kBvuygXgE6GJh2iEt
8Q/ETxXOI/5l46lN6VPyPEYEcHNfUZNYkYFOMEfoYXdEfPLIWkP+dCg2JfWfYPFe
oHXmF0v9ZGBbMeJGW0vt1+DoOATOboRtC+dE3uxuZHxAEr6g4DURv7C/ulbOch1w
lIYmkCsEyjZYzyXyqN6wU77czgI/E2LhulBW6uXedbuRzxPLzKiJANElKgpP5A8b
OtxOYoBn8/Cz8Cuf9aPasQS/Ih9ivHdlZ373Mlfc/zTOFneJybuOTT5GAYYZilYG
9Wuc8jh7+1KFyg2xsCnVWmWEyT17AEA4E3rCfBc7HmB5ZcPU6QRnKCCCqTYoaSKo
hOkO2S2C7ckjgwGzrlJtC7icHdm9ATGM/tbLAvWWiMtFRJ+aqPOtvOwxctP7bSYU
62DhZpI8OhG1czjl2Q8m6kHowK4AI3piroguJRU57/MweMSVwrTWvo+snj4Qbd4d
+aQOmALuIjbn/Nx2XH/CJLtv0WpFsrPwv+UuAM50myPDcFtarXkyZiZ03G3GPAv0
+ojkES0z4+v7x1nb9CRVOsyPI2utxynBA4+oa7N01lhALtabiAlI+/g8gI5b/LcL
ID1X7egRgQR1VtyX0iXTGGxgB/v7ICSwjHWAxK3Rl6GQhlbL2CnwrGRqdTQCwWdw
ywVyCBpT9kw9xQjyQe0tUKp8Vw3gCmefD/w2ZfR+G3trEJe+ChXpRXhCtHxxOWPV
jU2jkIUcwOEpvxe3mTbmMv70aKYXKsawvKgxf/VXmjtQ4FBUhmd6gxWKGlh9rnwT
tP2FpCuaN4Xkr5QZ4KgtTvXbBbLQFaql4K2cNjNBqu9mgYKOvS9sh0AiiIfRyrCB
HahZx2yh3hkMWs5MtPK0QCXIW0rFxqlyg8r9+cB0QMbExXugvVwdfzyN4EX+0/bu
h6H3oNByMVi2gxb/es44KaBQsK2UgHRU3Wt8TuzIp1HhKfD9qHnqNsq4DWANrCNx
uUd0lu0wZ4YAIhrE6V9ceL7By0kV2NPe0Qg4+8Pif4QsyArK76ZuH+BjSO/XM2pX
wu+EU6ciZldveb0gfrpVWHux4FLorNKuO1OEDLHk45Dmeo6uqxLG5OLzGXND7ibd
LHlhr9fz9XkBChkQOOQb+j/A8PcSNbGI0Eg5yeMNVNrO+u1wEuuoRX7Q3gy/Hu+1
hz0ksczKtNSsXRlGdlxqP+HA368K3DtIVU5pPxqrSZcTYcZDcP8Sjci127jw7Q+q
Q9zI5HRSWEuXHCkjK0Ark2AqUiau5CrmKTbUeYh9kje3JgyeBUVv3lkG2zOc7Z7W
hz0UnLE1TBBLPd6yobCSAFy6jK5puiGLPl2c1Gcl8GtXzE0jsMBbvs/Ud6+DxYiP
I8mzIK7A4zCpM5yiMlyPCauRfkD40mt1rVnMg+Gfe4YvjxgXiKqWkNRFUrUvcZJb
yKd1V3l1/dQEfx5sSq15Ww28oZnKsu7G9LwQV9Fc5bFOG72kNuWANpwWFMNAt3uZ
vKngl4VHIxH36YmqpdSPsBAWRnVot0JLpelVNNvOoFMWdwvkwnTm2xoefXmKKvXa
w7jOyAAqcL2rnwfBx1qEjJZxPfulFuoKDXNsB4WEfSRYUEk9kh4YWywrZClyurdv
8tGeeHTjI6g9otgHS4rddC68/J33OQrWdISifHtXDInmW4skxSQcxCLhWWA6Msk4
6SW6JONuKvZowI2vLfkm4In4jWbpclErJiqV3UfbzCcRY0jURcqy2fT/Ky1QQYnJ
1x37vdliE4S3iWbqcwjc02FgGt5t8edEHoM0Fsnmy4OdKY+4ntr7qc1Jykl7iL2/
Ky96g2h7yVFjjAOBv+08vVAxYtR6dPBkBnkqcQ2edQg2eKeRtiJc4APkW51HVSL3
fjAQlQ6HZjUdhg3Z24D3Eu+E0pTVPX4Ict/kvjqWXTGwj8bpRW9zMwcurHfT73DG
ShFusifra4+HUZc2jcq1pgSDQbbUKcFDNzuRX8/iSraBuEGu3eoppzNUXWlZOpnL
8QuQkOuCYxgrOMtSZCDtV4uhmUQy0dtDc52KnAvR0yKQ437FggOdemiqbgEDmQ9a
4kXl5Q3e3i5VoSvXHsbJUUsWFo6qZewQODfXkR2gJxNI3IdsVWJlGfKXoPHWwfx5
KNMy4WNYvs+2w/PKuKKSYPAwHzImlj9bVr/Cd59dDcVPyonMZC4Vt+BaQywUpri1
W/nNt5lSiG2k1Pcclu5le2ONZr0SyeYxEcu1La2vijuruG0JvNkoXKWQ/Ga66cTr
jV7vSce7CrzpLIh/APCaNxRddQBSfGk/rKnZtjof2HDbzXKH02iPWhz7olZW/R7C
QC7tUF2wrbgLF0j3dpnM9i6h3QOInPA9sBKTZH5nA4VNmPBkls/wwY0RDujPYRNy
CPHzx2BD2IJB071+dkT0FgQVR7tvseQQrYmrBuCYn/DBFWq4goQxRjMRa5mN8Dr0
yn5b3RRx8HXgvcW5xZHZre6ndXelEfbsIBGEQkIERH2l6GsigGdFzSv3f0cvM9fA
xrtuYy8Ukt7MPY/IuLBiL3sjk830fz645cZzEshj2xuaSJuM77UQMxoKuxT4BNRj
0ZegKhpoFaV0LzHQWVItJ3cf7Um+eKXOL2gWMnf+Hl6Kxm2Nkq4feqj/uaG1co5O
hrUO/oeH9PN+dI69BbYz20BXohymOOI7j1hR3nLjmTcXUx4UJCcUzx1KK4lho8Oj
1vFUjCBAisO8kItMnqm1mfZ/s+CcrWZvPUatKgZoHncr8PeX+3O6px0HVjeVRKA8
wezb0GwkQpMO2/g14kLxMRNgaDFMvCbrGyOAt3s6AmH7bCSets17OV/h2cRN7Nkm
L9rE8TaJd6RZYL5drnO3b3Bmlt8qX8iLt0uX1SSaTXB4VnGAJAvkGQiEZ/xXFGfy
b65OvAOlEyt7p5UCDkHDuZ/e5KI6/UP4+P9XfcWt/p7tOHE6bso750++cgDl2vH9
2RPed3Z1fvVDTyzby6aIHQHllKYmjBKmk7DDFRCtFcBcuXSvQN52x98WSXCegdH+
H2Xcx27ErzTD9uioYqEJzqchO5/SNBVHDMHHiud2s09vjYoBvHFWnFgKrm4j4pT4
Y8w4Gql93DREPnSoDw05gBc5IxbuWBW5J9ycCquUdQRIF2AhealUaz190j/HX75Q
dL1jcHSwtWBnXcPg5V63gywQtIqfSiAHpuA86QW/mLEOShbVRDHPcdLJ22M3cdTg
rckYywWlQaMYsSAb4ZbzfCdVTzLwX+3ZdRfGCgVySm+rggob3q9jSZqmQWPwm+hV
LDtffycXTqVTbk1E8Qoyr50RjQHDAH98rwjtqIYebpKVmgl+kiEkxzOj15f+ixIq
LnCEdaU7R2e/GJLlyeNJW9Dwbe1sDSwglON7nrswRkV27f0yKcj7OYHs/d0INAcy
dvRli/j4k/j5zY6g+U7+kNLQrBWxfWHSq2QTiNxCKZitAvi3ra8CSRtYWlTOkN47
DE9P5E0cO0CMnj5Iyi/hzjDhyOhxQtOPQJ2QTbHsITbcXqICkjsBpEFawVvJ5Q7x
0ErrBqpRUmPK0v7NwWEQ8Kh6kS6AuYVoGyQIRJMgJyyBeg7J/rcNfDXQXwyP6lI4
N1nH6t8pvIhaXHYxawy7/zzijs2SWl96ywxafqdM3nixsibimsnr1/S8Fwx8/LcN
w+wL1Ji1E+Ow+EgqYP5WphJZ6UetObxWhWCLN5v6qtjfwnUhoYIXF8/iw4oghcTh
zQ+0KlQWF8Ig5FjA8ZTZeScOwHIDF8AqjuKlkojEWxNyOQdSQMg6ZBhW8Ez9EYSq
lzP+Tu4yQs9Zgfodm2jRQf01VdD/8oXeydFmQViKrTbpZib8c3kW1QSFl7mRcl1Q
tvxwFXV+CPvOAQTCU9H0wJKeY/rqevn/OV33ptZEajHyhQ1vkx8+OK719b5Grzgq
UwKQu77WKfKr+VbwYrE63Mrflfdb2AGkLQl3n+8m868g4hFNUIiqqQAFmmavGypP
qAr4MaYp2Dh7pFnylDRpJ6dC6oSnbsOzV47C1+btu+opNnH1yegEfutHChM4hSCf
sDUBWFeU3Atn58xlk7i8y1/Q3NPgAv12TUsUtPLeKYHAvX4BuQGjXndj1PrX24Ko
1oHoQxTz5pZI+xDJ5b6aLxva6H+G+XEGCLNUqXck+KwhUwnWeiNKwHqpI5P5rkht
Dgf4yOTM50r1Z1iFfzSFn5UXwSM0wjomCkeFKqAdOFhpyIWU1QrUo70qDn1g+p0C
6c/0Lar4fSvBeTae1uM95t+WdNfVaYd2SCEQXX1agiNhIfhyCxFEQZ6QF0KGW+eT
1ERekr7DfewmSULA638WNb87/KGMpVkYkJx9jtxxLnv2TZbs0cjB7Jd4ajcj2w5y
CwjVBzA4xQuLJocaE+3uExvEXySyvpGKGMIr0c/pLzaVLcgY8E+3TwVCv7+D5TGV
mhlCK0j8GlnVqu3lK0qbPZa6bH0rJMWClC9S5jWzly3vWuy/q9u5th7xv8L/2j/Q
OXpavEm4EYHMsR8UPJ0WaFXX94cY+1wRqMxQ3DSZ/0T/JkIH9wR69vwjF9vcyHeg
/gK6HFBANVH2f66KdneBLY4TnNQrgMBagbikaRzu+n8yt82H4lrT5/divfib6fOI
IYQvdFjh5kj5SftGuxxtAPkq73zMzl/bKTXhw+uETjZMXUhdl3HoSNwk3RtRSAwE
ummYbX717KkjAxLDh3ilz14Mjem+/gny3p5PmbZ0RxbQfYhy4hlV13ny41H3dtw9
pQbp6CYvAtXSLJw9jh0pduuq35LfZM4SzRbHNKQEN2HCJDHn6ZDHJ/NgtWbYbrOH
EGPVIugd40KC/MMuf6mArB/ad4kEcN+dgCdQWp50XM+J9lvA5QhyHnRT3hUm0VDS
sX+q8dDIVqQROemGvjZ6+882U0LPwkFyHIEr5TRVKy5ZV77ftwZl8yT6Wj+NeCzQ
AmEN3CPFwV7evZK7mICRn80pFxg3dK8CnRZRO6atNS9ZkCSRp0lWlMjECyGTtLhs
HBo3ONt4VjKg1HRQUYOSP1dpqX+fpXGWOMo4O4sKBmgyY67kYm6zpqvugBjbxyaz
o9VgOru0pBRwtlX17SJevLCYfy53g/f3kE6oRFfwkbQqe0PBw5YM4zBPysDfF8V1
5sRaYW+xE2G/LiTK6YyzwCnaHbkgEtgw0RUBUIG4dnatqUXVW9k0hTTFcZnoSZiI
SsfZVtbPpWEeBX4PNPGqq2lzPik0EMM1KJ6pOknUZQworNYLjr+cRWUwdN4UBjN7
3beKRWoYsEKjg1GPytXCmvGGyD+jXlA5Oug29GvxEph6D0GPY6wjLI3aF2iT6biX
Z+tGFbWr5KKZOkZ1SjEszRAI4bNKr5cOildgxpZ8BHb4PBq2EWKsdS381rQ+zBWZ
NJLttj80xXSwUWVH892HowfiDynvjhCtFjX9Maw7nL10b111CRM9CIRSnp7ZbSZG
G2IA2CvJYgQ1uah1u1jaEFhSstn9yYvuZh4eWfAK7Tb2o0aVaeyzV52ILim2omq3
0yEZ9P0YP/Chnccu3DTmRUAJN99FsJ+24zmm8NRUVui9H1itiHiol5WNpp6VdITg
SHo/T0a4n2Mb3XHm53fl2CchJzT4ekGpXzpTk9VocrfWEBrvqeoG7tplC1TGUA82
`pragma protect end_protected
