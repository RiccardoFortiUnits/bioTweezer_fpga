`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R0trRluKycudZmKe/58oHlyMzWrB/tQnPiyr7I7LPyjJOlkCnpmFaNpC0iGik033
/9bR5Bi6R58YAMeOi2COPBd6B87lmvLsUbV8ywEJTjB78s3lYSFr7TIbpVsI5R/q
4mX1tW9ley2+J/u9xMacrWXln0NwiOhlF0TC4lo8PaQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
dqDK5cExTI84mnMHO9KIqpEh8ANteT+p6iEb7Al7f+A9IcE6V4XYsBL5EjAKuOim
xWwyk4Iu16ybeQIPf4slJmD3tTmSop/bypKjk+ufRwbOQYjtjBYgDR3WH3XVqTpH
1oL9ZyVX2kz1pHye45Rk5VQOxTzDjWMIEkEjVL1h2cU6QRIljpMRfvBCDBkTaxOd
wfDG+4Cora87U7lt7UHz+UlCol7AiiRSEpozaLl4uRnnsMUxpFcHKAYKfrN2Sz0P
/FqRc5rjP6fXQukI1ZcHdwHMrKrzNkkd1543rxCCWfVtSDmQL/wc7AHHfWckIzwr
YPriIv6686H6LqADHhvhj5VtBTa9smO6HsYvXEZavBJuxm6mt9onkprrQwgYuoor
vsTcEjef7WBxtiln6OeYSZOZW/Ymq1D1O2Barkck0OkwtKlS2RzgBBr/jKccWo5o
HFR332TD8yveWBKG5pbIZ1Q4DeX2vMfeFwL7XicypJXcG0B6qvznUjkA4tj3Mu7R
0dOxBkXE6eT3VkixyMC2TjZbZR1F4VaWH8+V/EIPsDEtFQ5MaJdJ3qws8cf83Znb
tZK2XDad5dmTb+4BqwEeTlMh7WiOUSZAAxjPxnD9AI1Te3KufYOwMqMBJbZfCD/W
uVSCcQNB9yEzrRf/7wa+RtJan1zSU9YII5+K5Ov/+VlcmkIOXcU6MT9nEaQD2+Aw
Dg2U1FlmtWSSOCSCY9Pz+507A+kU9izyc3f2eIh1NSOyApnlUUf/rCDTc7Wwx9kr
T7F11qlbx+a7jhcdhSK6oNH5Fv+n8vDyjphRoU0PBjJwE+v1Pdwh2jZi/fnmY6r1
C6wg0PfGB1NG6OjPD8aL9zpV+ncXloS7iQv44/G+wyxGDPwgUmOGXtxZmpIUMe3D
d99tgkAAHxofvxM8N+Y8EsH9DphcfZGzsT3ptrUJh6+WI3MCI6H6LlzxPe79cIaR
IzD2AEh+AaAat6pHLTXzRR+c+Y6uFdO/n7jzj2lruSwfsOv5d1HNZUbDwxd9acmy
fHL0f/VlJ4MvMUkE+7V4PQuNrz6i1St2zilIRwLeVBjQi8NZEb+DeVAu5h1S3l7H
dr7XOqMzspB8KTGp5cDNi9zScMkMkaRU1kn7ubpVxBdGramKwwwSSIaDZctqEJ9N
/ZNr54YyrQrjRImQLVSZrVGFR7Sd8bHtUZsaL91LQqQAjNh0X1YuH+ucp5m+TEqH
/s80OORA270sReCkJX9sH3Ljj9nVcsGgBHPiR82ZMaEOmuUOy5w4GU6+/jA+HY9O
BN/OFL0r7S2isk4FdKtOBzY9vPFjZxWS/NY4H1KlqvfcDuKBCWPPfO0x3HT0I4b0
Omcq0Z52/WfFp3InSDjOnyy63RMcrXkDPvNlj+yb1HScv/OoOzKlTiMrwC1DaJ9y
OLL9edazCqHIqy/HBRzXZouYnexuOoSRHQiuCrhUVP2B3hLws3qUXKPPMWzKBGh/
foPl+Ufaxsw6HIDMszrrcayjoC1frRwlcVh6CVasDw9IEZV6LAZfQ8WEhroCk7fO
rYSNmy0/xJqmJZ40I3uIraa7DQBvVQ2hMhb4nPHSMHUdNsseY/j++Jk4eW+x8olX
a7bBMu8CQ9Kt2rV6SajRb2f+5PFiy2pZR+hhnYmXVQjlgdVKnc5Lmd+pDeDGAPpX
OODkHhmKSy7vKJPnlNBAHBU3slA3KceQxlVcBt/Wr3bkBSqskUKU0zkjyD82k+PL
zSY0Lb4zc9q7E4kKj3GbGycbSJjClyMDzqbGM99Pr5gI9sa/Sf5Mh32NWepMXjrn
+HPlgI8Hd9Aq7E0/oIRXjMVEUnC3eYDb+vtkYorUuvO3UEkTPJV54kRmggjS+Y7i
AIqXC1+0C0DLRDb9Qhy7zI+6rJSgAr8DX4rDoLVFXrhG8QjkcSeZOBREZEPgx+6G
lVF+HseH6wm21Q5THy4503if9sdnrPDCVfpwO3U+UVb90zTzn5yeKkYUm7HOvxNd
xixGMc7he6dqr6DVESDZNObQKInSGUrL8aylIF1OGQVEkx9Q3Zcf7EF7UFmxqKeQ
ps0QJct0Pv/zVDSAyRR1qJOx1CInri5sSTBWtC+gMaFK9nlIUuMsXKwxOQhihTm9
MgkR+9PqpG+GiNJesbpBt5MnoA/abaZ3eVqfo5GGk/nXOgh/eXnf+IP9idcOye9L
oJSz9xZ2fjd99PKiV1as2bzya3Hb410T56Bkz+WppfAW4xbiXfCqK4X9WheHCiEd
nQkZeVHiscKRcISr8Rh/Sw95zGEPmEhopUDLCq1DerfXlqajwGF/MROZAwujt1Gc
hKavYlzRXS2bS8xoJSrvB+4plhxqbmS9fobLvsL3oi309nZgvxppw2k/dqTLVbph
vaerUB3gfo2QIfuvYLuS+DJaneA1C61Vm9dufGBiny/OIhPtTwMnlvTGh3u+tm41
EquxIlmBJr+25CPnZmNUEOIefb/RxaVuvaRa5ci1PKPcDAP+d3FwhLY8myieXF/p
AVYVl7gCldFSVFClia+yUmt9l9ev7TpzHX49kQPyjjkzEZknoGsv627Bdr407qjD
F8GtTHtcB+2h3URwkm0YLLKVp/Ue5FeckVFmjdhjdfylDr09kbbiF5FBQ2BVjJ0T
6ow3EK6fqtQEGkbpMTHg2FCuv2iw+2DwmEp0Q0ypB9f1ydUW7nxZmzlHhDdf5IBg
wn3k0Dpb9+NC6djhAEuu/kvm+b3A2qJPhqINIliadA/4u65xXLvbRrf5uSrdP8h7
QCicXFLDYOX0TVwK8862iQJYaGlgxFHAo6jnf3QYMlNMheZd0pL62MXQJ7UEvrko
AFi2VE97mrYvNbdxMJbnmBWXUKjxeTkePUKjCsMkIBnOSp6NGbBgrIzDc0pbfQSq
BJLccKJPvcbGZQ9Go0CDkUk4Z0LBTPWw2Wn4Gi9IBSTp9S/Bt2yapaoa2y0yb2ie
UCaK6wqVPAINMRTY9EQZK039Bq8T0anqVNsP35G9zp32hL5dMVcV/PX2VR52FIAn
H/BgF1dYtgpumND8VnwZm6EFR08nSgwmvfjKC4UPfE1LG2MSZclCyHiPZ2e+UR03
AJJBfFUYkEe5jSBwaYqqQJT+Vz/1WvtC7QZhYkBBD8ONLOAp3cxp/XbGE0A5lATe
ZnFZ5LYPgbhaJapiwy+bokoR2x37ZGYfkLF+TLLfZ0SNsruOyCryCrnFjkX4fDJo
xaafKFcmmjIQTzA5nrXvOoGWnCU5qPUpiGAobyGXwkb8POZ4rIHJXUHKV3xsZNWE
tVuQhmqB2IpFBvjS24n+pA6YJ8WWMPkBewLBasWfVkj3rMgNfAr2NDeNDwPTDIpp
hgDxJXZ29InfNhAb2S2BEFHajz53DaY0trlsedQF+WVuQd4ILqKnHGjAyA9LV6d/
g5xTd0nT8yacQR4jTF70Za4/oBLcu+C9DLsgq4igIMZjjzJy8dpL4EfU1w5Q8UFd
vtt2rvEW6TwjV4TZjnteI5YLI/9J7rPkoq6CHTe3O2UgSZJxbg6iXnzDiBsiXPd4
S8qAaN9RPbEyJlg0gTfhZ/qprKrsuvUvUWc6RSAVIORDbjeTTNb+O2VK3kJs42yi
zOjd0s4MhIuvIEKQRl04QMEoUtSgcICD1a2GiBwtwLlMfyCVCmRptbjTUOKqnnpD
VP13cKT5Kgm4B7AolcpajyHVVqefcRY0qP2NqyJX3PfB7Hgk2m1d9BC28+VX5/mH
hNlM8ijvadwH5XrLMSUPEcNrNEf0FGQVFl2PFkg895KNe6intC4Id3+1dxv6TEAq
eZvJvxnCZE+kSQvun9JuLYtyh+Oc4lDejBVzjX0LZlumvc2waPBrvzcpdZar+0R/
XCPuwKkx+P/zS8O8e1cT/RouLCuFDtR7w7IPn5o9Fu12jkIIdETouK9FKZUOVJC+
Ytnv4Kd2ocnJIeYv2d9NrpDSu34m2YCAP3/dYKEB5Zyn25GAXsJeU6gmRpJhOnAF
9zl7JrQaQ/8JHKeDnDjQLnTyllVge37AU3IFil/lm7qhiBqMLCu6pBfAYxt6km0C
UoYZLLs2uebPWL5UkTTfAu9WxHzlkDvT8oocKjOeGxaU26fjWWhbps3eQF7zy5P4
u445LyB7WD54RuejG7gtal9/ccpE7pI5xGXYopjPwWNBakkHLaJkPyu9eP2w9sGr
LjsRXHFuyB+fKrSKE/ao01lTjf+jSV2DOOOZcGFLONAFl7osPamSEjZNrFQvnCGm
rg3t4gdL/nPjw2m8Q+ih3HWVTzaXwIxbYgX8jihgsC7HlLYMfKtTfmrclLuYFoji
qUaidSOWqspcxgRCVXkMu3JV4+2xU7kKpgaZ1QeMYOUJQeGJnyiykarh7e3V1TP2
foNbIDDxQ2KZOWquegqdQ4IixL4bksSeDFBiVNZDitFez5IUP2iI85sV+E5p1qtM
x8DPQU4r2qgmtfWWuiU9GxxIZghTbnIT/1u1rcUNlWgTSw74EBbv2APMlcvVVs6C
Jie+Koux6HS1FQeyFcYnS9ZYPzFbZg0DKYrvTFcO9dhR03/bxdTBvuSHN+Txl7mI
YZ2OZ4TzXf3LWZTHt9AgmrLv/o+MUXcFyfDeem6a+DpGuQ0j2xDmlbNbJpoWCyZk
S1bXOhOGDSNWYTOZPB3fUiGamndayixCC/55iQzF957D/FQWZiKIvsI5Ui2rXutC
SHOfv+AhZi5n+GcFnv3nwyQtyCZ3oMAqqxNPv9G60JXJmmSn6vXKM4XCpoZl//Bw
TDNemss8U978P/+UBXOdmwPsZbruzM8CrFm6DkJb7rMfvglaSi8enTj8CE9wMhD5
SC+iiDSwaQkhpSJbdWuY5yN0zG9FR41wnUP8WMtSqT6ptx/19u+CRfcoXX3bK+B8
CWTYoeQhUC63nj4GAKuQSn0BOP1VgJARvURy8EKLq4/TKhqM0BTaHOciwJ4460nT
FNk0kcSw0T9DPoRxjevxlQ2ui4X4t6rRJjsiLQYD6D4D1bRFNrmTz9CzJJwF5MfY
Afieh9LD6UoSSs/M0nGUDvA7Dvii/xpQPJfMugw7AGJnymCcSsnRJgrVYjYTTckQ
321jTc7WH6LFuylHAscaOezI3QO7Sda4wX+bG+C1jJwp1hLhpRMTXkGfetO434Au
1xCK0FQjSB/arpWF9lU6n1+3XPHrymDJdSisb/U1KQd3dyjleNHI2zz3gOGGQ2KI
lRbEqSlWZ9XI4m+LohFXhAqwzvyAZLZRiRi9Q2eEs0sbK0jl69CXgmYHu/YLBgU6
ZxZNbeNB0ahoBZeadSvmFj90VXJsa2Q8nbvBw2m+aIiYrp2z+56fiH6CSJYdnB+T
OV9yrNk477xVdX079qLhM6vOFm5wUU/HREfi48yMlmhWKyYGRdcgyDebGQL0qVpH
cfcXkCbPtjq7pLdciT79l1HJvhjZqXNzEuKq8EecokUIvt6NBccPVOSzgJcpheQy
RIgGg2RAkl1PB8UclVLwcKnmMYBKuvbBdXScs4Uzc95yh9r5zJzb4IhOlhJo3jgM
0KLLdNOSvhPBl/F7MTl/1ggPNHZGVa7U2c/KRSY7G04zcZvkX4DLJ/2Ia0nEdQNW
MeAESjW2qoELol64PxtgK9S31+lKesH9HCq8jRUJQkjKASH4aIgn8461HAItPsb+
T9CGaRxNcZE+Gco739H7nKWDBqZB20tqbWO27RATmDOUtGggFRkBUCkz/gBtGP6S
LHu2UaHU/XMJ8OPCu4EoFxX++LwWoKdlc7HLGuVOfpvtyDEy1ZZiRYI2XFTsXpem
bNDJ5CrTEJiPnUtlaUYUTdkpRP5++/WGlJDHPyJqBmUanFh6tsnU5JtTQxy+GA94
T9O4LkItpxMtHpPzZOU1NzcPkVyxmhoyE6lzMCYqUjYagZo4y21VZsDmAkdzwyQn
dysY/cL9X2dR2UbPPFDQDBnaCzw1kDfRAvvhzI/YWtj7vflzLS2BM5zfc/EDL1CA
LWL+0Na//iJaIKZuavutvU0NhXBqVeA5IZGTAvDml46wuW4b1f/HMINw/932bavK
WYB4/rmELvoQuv7J8aoRqCaVaje9y0tLhyw82vU79QAk3gnN3e2dnSKN7IzQ4TW0
0n6qNnYSZwsp0cpoUizAPHN2ReLRnVsysMTVCzL+5qVDf8XhhnAEmghEeQxc8Kie
jpKI8l/jiYqyXQr06iVXrJlTxEpC3iAa+JldVe3QV2gac2QsuRHVF2LpS1zYLpzJ
RuNCc5hg8Ivi3JKuTc27S/fgjtSA3iX+9avAeKUMCGjjc/WO7MuXE2t8fHV5MjT7
sVin6dKDcZs0c/13VUuNQM45kfSlZoMvOiAG1Bh7M6SIQNGBrQH6L7k40h+T4u0R
nVjCwGwl2QODui96Ls4cRDVxYN6I0P0eSQXVKeRcFot3fevCnBjyqNutPWpB234W
s5eyrOT+sXLmlDF0YUw2fKI8iogUreiIZqZ47mfB0N3mTI5v5cNoWrjyukUUrBt7
5H3TFH7aezIIwWicdGubd6t49bQaWbtTf8I1CqOUXXsqJyk0+wzWfLMGEcLT2mAj
HeWKkLeOXPaKDf8eznXOBkyYi86GU/AQx4pT6Qs4XGDtmaHVj/MrSa8pblPPZ9pa
3mBvsL195mX6qZI8+iK9xJyJo77rIwDQopzjg1pV38N2azAHOQszCUSQM0448sDS
mgVLTUg71rqbbeGWC2pC1GRUKS589CEsGllzhiI2dzHCnhhxamYYX0swJrg2489z
yN8fjX+ZLcFXkimEf/1YhHUgMTmt9qIjHV/GJhE4NTVQcW9gcQFMBYnT2kk5vJUW
zaaLYnrpg0lF28To3/zeIqE0TNRz1lkNN50U/uCVRZcoCHHVvGEsyuLSGjXnkv3E
eRUFUpbPKnyJFbLOTUuF8xdKFpNrqn9wEaIZBFff3Pvh6S3pITD30nckmEg+2D1Z
yn20Jw0UIX1BegZ1lClCmdE7a7aJxkkQoC7EzpZLNbDn+XSXWZ8ZggLLJnkk4lHd
LkiQLiOQHal/Gh5uhikjxlZ4YztgnuofQCDWmPFLBR9lUFCjbqBhZLA+XWuUY6kn
xm4wcx9eyhE7/OqjHw/lVAQvbt4aypbJugGA221m9I3cz2jCaztKXOu6B2jlaN9K
y2aQJ6u1+OlqdvnPEdQIPLe7u83ue+EWkORdTFdvn4AOoz3WDiWHvNX+FCQTYbya
DwWwtfQV/sGOLuT4/pcinF0XAwt/DQ7WoUQKL+SUQg1yRvJtuyu2pHZEoIiP+6rf
LjkZ9mxad14nqiFisHVWnPfETXjC8NMK/PS1EJLaCnSJihC8d63+lzDhlwIVUvJM
PstK4shkDjQu3Wb/kwqjVW2SS5rvZjKYdmhLZqXH/110ho4izH/unxENefe0vzhq
ZsmvHGRxYrldZCGJaUvJp3AskYKr8OeJaye1aMgSJ1HcwgptyGcffA/DkKLxpXkO
Eurk9zZdCcl1ARt8dh5iexncMR6xBtYPAh1BKwquk2VvtTfv/G6CXrzm0OB5CsGQ
4OUlmRMnnvMebVCz2f1lNt6Qj3Biwkel2Yr/sF90HiLStjhq3wbzDRIDDfnD6EuG
lCr3+wUKhXqVsvvVn6yKQNBUZ3yLhYIGEPQY3PlYDxufZvItz8n6lhXCo6Ap89RM
Uyh4FWxwy3ydfByRpmYfiw==
`pragma protect end_protected
