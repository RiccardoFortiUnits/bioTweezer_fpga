`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gYMm144QaJVuM3obcbmNtFwY84BIzbjYbLO0BcDdHSkn6PAJb+c3qiZqRKNXlmQK
o67EMhNAUKMjXN+bEPR+XGvRJhcuimtAxWg8I6kCMIR/f/mP/mCFZ/gbTefsDFmf
hGy7+cQH3N9RP5kw6MHOxdbiGOxFDFa9LwmqcMwrfs0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28160)
WYT82TpCE+egmLnIjR2SV/jwt1yMr8YgOX93D0+yTedsetmI+oNKW6fT6vCKV/4O
rUrnvuoV2mO4raw9Gnl/6a7uzQGH1mDuzxJPm90OqrCa0lfNWLhlTn9Y7cRBu3a1
GN588nBANEhMWYGDQsblpbLK7WRPrNzBsPRhCf4fvX+YEvFefpZunpf6a9aghfIx
AWXcpqMZs+pHMTw0qsdRHnq7FEpLnmM4Q+Ds9c6xief+o1o38DXRKV16g6wY41j0
QxOQJwBWQZG0x5B/KZiEieNRTHieaOM++rC902wqWz2ERz1zaltOvTY9DyjYoFhQ
CD0AGYv+MqlbBzS0xtttmBDiB9Hyd5RTvbPjTYTrphSfWPKfri69aTlnPzc/G/I2
xSR/G2rc11LqEpp3wjxVlo67qsrK81mh4kh3iH2VbJ0SzhmZA0N8BQaYeIK1sJ1V
yTpa4cjhSOHi/2MiLFxVVjHb5K4+dkj/7uPJhIzIFmKYvM5X7dftCdRruPJdmfhb
VjeGrOu0jFOv/CwOVjjlQLBGD7TJ4HngD3zdBLXUBQu17qBa5w6mxgETgnCNQI6o
mp7WOSC8DQPpsB4N01BKXKcShP/jKAD2kdEfAs28KrJ1l+nyUFz7pzZ5n+uH+q6G
bTU3DKep6eZnRIcGJo7uUsCVG5d03pm8Ugl71+LwGFEVxBbYiMeB4H54ImhBSbEy
phxoMvtqfrTJYWWKUyjnDU69u9TLUVKLLolY/x1ONPq7zqTKaYu1sTjjr2maLxBF
Lbn1IeuRFBhFeX+zFLWbaiviWRj0XagC58u7EjBWymsl1RCWOhUgutUVYB6xX7tt
eWPcoP9SiSmPBlb5ebNrZGU3O0H2aJtoXrYUXYIQnBCj94kQya8c3pcpjwe3CNzW
hHd8GRfyYTs7mGnw82dgVPK92CBrWCr6uZ+diLveg/9W8aP+074WgQzeUCYCymA5
jXEeHGito6LT97PtWI8IKdc5wdHe3LJOR3SQpCu4FtxlOj1TZhMhgfIA1zfQOUyx
/WvwWgRSO3qmIyEyHg6GLi8z13I8pAqnfUd3XFQQhahE8wAHoAcJM2kHrmuwu+iO
fTMfI/T350sZulebIQhiK6ROTG+A+PYMuq2SctRojkWiXroReV5IuIshseOBSAS5
6lrf1COMQ3VkVU+xIYoNJoFpziwiy5XuQhbAlZmg6zJt6MgLLLtmT18o+BqUiAbb
b1GANChf29fPBUwpOkJx3Vl4NB1DlwTRgn5BbXNjkq2cwQefJ6Z/nNuhsxqJyfD3
hgxYQCL/czVvnjntZU56VZGYXKvhVzP/pb/QgG1bRGrpJzIwQCAXFMuvTYmf7uoe
HzUfZckuXWtk4+E1W73Q2yofDmG3sw4w/q9Iw/mPcKoO+TX2wy8VNSQafE6hFtU5
b9gvUuxdoGBZt+JrqFE/0KJPTLRcC4Ds+hZsdQxmCUX/EjUh00yBfYEjBX/9+uUg
XRjyBh6z5ND68yQtybEdg58NceeWQRjViH9pHwMhrAHnjnKE1ms4Qxb9RGIUAKE/
Bt+ukXB3f0frCHNX5o0DEaht0x2vKdGFJYrcyPztvm2FlPwFafO0aWVk9W2mQwVu
dTfPYc5Za0pfVBeuCuyZkGMmYfPQWhFNP74i+lWz9TIrNP5/Xaz78mAu2pcDyfFU
HRGywWRRovbZlKpb+lIkfOu+qk+hvDqx7ZK7mPuxiQcycSTnScfy8hrfjjYw2eil
Kx2KYAL55n4s860r26btkKPHv69c6MgDkBog37HJGXjFrJruZXKsO6AYjuQKRxj8
EKwmErOroVjt15x9r1sRMI7cJkc6ovhlqSRmy07CRL4DxB1Q7icrBPn5yDYybtf2
PKdPGgCnQ1mOOkmWaYmz03Qimg8VUyeRqa9FRFcmBowd7jKtOySRZez0OWyWC1Ib
ozUpc/itbVg9SRMHGO07Y5LF5vERwfXwU08Bq/ZtQdo7YS2fWn9LPuN+9WD3A8T7
rgTXswotXR09IPTvqBt9bRYnqoHzZKua32eOA/sv7uAKYoVlEuvDOcXryup3DpNL
UhTJ9GIVR/tXF4CHGeSvRJR21BSm+hcxwnnlwl355NCNfudlsyPioFxCn+ePrRJM
7sIEDbAdVv/unmlscjzCyesR4m8peMFF30dR3MUuq/2Ty1w9YeA+MBte0h6WKkVI
3RrH5PDsvTNgK+MublUFqqWsAYGAPV54czVdlzW8UAgGT1cgNdPzjhYW8HSqpY43
9paOsWXJGnEmopPnornvh26p287IY0NgfU3dmFmyYnqQzYjO9khXolv8kU/ympoj
s1z4zMn0EQ8SL83uUCloClNqXCOMcg/f6238+6pJ7gb2onQngc8JEWk9HMWNcu2+
+bSvq5c5dHdmwekXPukTKrZ91ZucIeytJVl7pJQ2/rG6ahx8TMVi7PmNEh+Zv4wW
JfsGFVTI6ThBUlJEl5owNbE+FHlxOmE7DXeHeABw9FPe9UXMxnStls9TbA8S4dUx
QkRQY/Mfj/IHlDQzxLRtnABRwyUICUj7SkFlOmSEloJ50QPJ23fimcUN5VRF76M4
5uia6qNKZCryPhsjormGv+MGjYnfk4D9w5UeSOWqHpZ/Yra6z6cI43JvUYgHv1dx
MPshy0aB35IPusw+9qLbgxzplh/msvIybAJyeIrMgGyQU50MRAyetOLOIVE8GYth
BhdXkc5/ZjQDGgboc+Vt+z4w+md+w8Bd0l0n5aj5zlPEAY1OaO+JuxvhV0jrHJ1K
kNDRMGhfFTPyfFVz60z2/tPFFDbn8EmKXrJ2D8N5z2inEWvNIYZcvO6w2hiQznta
RMb85mEW2+5+1u9ml5zN1094Sk3g5gJgWGNGTPMHb9MaNVi9cQEreXEJMl7Lctl7
7yzHmV7D9xY+5u3UG1ex1QOyc6yf0BCwIrSOxDuSffwVY8qzD3dyq0+9WzwuT/jL
EUatGrIhL69pL9oLsq/1HfHBFIO7XRtKIxdS28GmZm6dPWnclf7KUlA8Pr8yKwzf
+64aX+QXmb47cz4eJXNy7Ts60HfmWhLMXCiC/aYfepdIKdE3VHhOB6vaV9ZUtsNj
/hso4OVUQN9R/yqkoSwc/4v1KSGApIMlQaWWmMn3XSfuoH4eUH6B+s73qOZu1iFV
JS7LgJMJub/0eTq0+xzdd3I6BJJcLrNmfqjmixL/kUiI0T0I85700NBsXaLW2t5y
0uI6sW+j4PjkvCQ8pxsubPjfe9AAgxRjLv158JiEAnqw/yAWZrGlO9bOk/0Ndxyq
CNSNrrHJSqcl7jUWpjz2ZQjdNpmFGQkXYPBMH5XEpd577z73Lkb6OiEP5vy1LviD
D3P6zNRphSnGL/ad8Ht5bzJpSDoc+AbuZHYWDPptDMMBLoZ4b/Ih32u1Y03W+6wT
hvY8i4l96Wi5g5dgAk+mAuzUx62OBfqbyuU+YBRBrSQYGxhp/RRl2RMIVLTht45n
n+VBVrq0yK3W4rK7kclYJ2h7xAoa0ndkFaaWFDpZuXAPvClVgS5PuM01gB99GxDN
/4pe9rNhcbkrb00t/YKoHPfam5iTXWPzh0m7Azr80e1uCR3niczEwGrL2vj8hOwd
T8UZyINaeup9Cse6tyd21WoBF8WDw4iQfEcKF+NtUewr9OjzoBymzQCNrstus0Aj
rsGHgp9K4/qt8DmodXJDrI/KEGJhIHh611A+c0tzeAlOmiJCfoRUOMpFM4GKdirj
YRHwrigiRZmX90Mia2zALLvrJ7zFJ2Kzl2rg20JSa5s7NK6Lgz6SPTY7tlK+A7MV
8bYPQNrIkFv31CSnJ07GWHUqpMIsoAYbd2Pjq2N1QqaFXgW8jpK5NHAq50wwTYYt
rrNcSxnl6zPJ9Fy/QKaxeQ6z74azIQ/wGtX6c4zg9FyD4AyAYJd8RfapPAKY0nH3
0wMaQn3pG5ccVrF95y22+cTYhzzCQicW9zCqCow+a+OAxZuOckOxTeOqHsnhQOpj
nmxL1XIMtjXN3AEjPjils/YPL16jsW3tJRgJowlCowYqmH+eEDOnZLNeg6SRucqI
khcW9xTa+l0odyeKeBsRVEyiahr+Ibw0cHnxQR1rm7ZAe65xUcciz2pkG242R565
coVwzB3+0v8+N8PUxxO36TEJhN55BZi5yBZdd2J+KTngznBH1ZWY63UOW9LY8fgJ
qi4+wmQ8IDDH9pLFdPgC2/7o6inCywYZFoUvqdpsdRNLM+4FtIWoSLUb33kaElhA
3GMiVQt2ox0jtmTtBFJOZdV1wjdj9mwbysPpX3nOG/X0W4exeQy2q7QyhJdf/ruJ
JK2bFlxevM3SulQGrBcqU7k5Oi7nqOpLoLPb4FvqCUKaajo0eHOQ5Uq8XhO4NttK
+T2H/26JYn5e4xZk0bpJT1XcWWwhbMgI4ZAdES8nN+pxY2shwVyXSAxcINThkftx
MKzro2Nt2cdCP3+64Nzt7feHOIzfTTKzKXhzlTbz+XEhKUOkwcceTqgj5JWoZSYR
osUHvONjWlmzZ+hT43XhE2UbG6qyJdTvHtxl2weNiOxBnYz/iQWKUIAvhJNolUs7
rD495ggQuk43zDYRSEMgE5154NfTLkPpnceU4BAz45ahv0GMRj4LZe9p2klG4gcI
XR/4W4VmX4kxroI+Rg+OrONoQMIT5hLEylY8Oh9ODS6siKcMWQt2z6uQJ6gfr8/v
jUT1pFDCdAHaiusOUdrxN0+2rw6zUsJO6aCfO0zMLg3WtP+xNq5xmn0iQbqXkKke
KkE1xP13psjb9wy4VNHU2FH8JFEDeowamO9M2LwKcNGIQzX/I2h8b4GlZTbeebS7
Z6Hi+MDX36j6an0H7F7q6eOILGVgL+XPid1b4YMgMSDio8AokDJnswzRC0KiYlmd
Pn2iFxv5fU9zfIWU0AbskafPX9fffpq6FzTyKCjFueqfg5Ez57U4zrPeYbv0ulhv
PJgP7+06Mb5EiVd/FW3U7EKBmytDEDO1w4cIzyV8SgutpUvkd4Pbj/OfOakQVvxv
TdH9weX4pmQ93e3931gHSVDi+I2041ixSh9kcU3Jw+6wierzUo3PoNIAzrC2ZCmZ
uDT4bWeAIjeROi1pOiJw8BtydL6iJ+YvHyaObHwAOovEdYfxr47xe9OmbJnwSMWP
xbz0gp57DuA532/LR130RQHrr/TukSu3hhrlc3wFCRnPUGpJtRLoWWHZvoQLaSGY
bPBulb4cMW9UMxIP2k++KwEDBzKe+Ve9ACJwPKPomxx3s2OOot9aLyrEhbBoBUAH
vhx4CRlaltJkJhA5OKxFiLioEH3RxqtOzGUKvFnhVu6dBic/wL45dwiAAHUVBO3h
kvKx5XqsfIEleo+G4OdxJW9g2Cz5w3W3mWd0PC19K/ymSAnO6nyUsBzsXUXujX3U
hw2lRgVLlGy7N3fxdPb6Vlj1d4RBD2BBayEBr9juxDSknruORDgH54MqplLUFWDO
EvHAatTYTtRRFUvSLUBjj10u/xnNgyfuhsKJNhlMW7sdoMQwj5R9Nl5q7/hDHevv
Ig/RaT1J21vY/NhD3CAUIQBNSO3HgI2vAS9c9E2GeGbwnApnRM58PjHmHjs6Fx1+
0BDfMh+oKY15PvYXDyj3vx1BBwsvG+bevCLplMujnRULmz0AsliTzCPkTugmzsZg
jIO/fNMVQzYGctphiqfJdk8YLM7ZhmqdS8yf0rYlTOfkN8opXiNiS8TGFKdR5ytb
HDk318DPCCALW4LrwXvOaLI18InaiyqOrlKRBAN/wrMAwuPUdiVNfj08CEnRKi8u
vjcedBJSgt5Ne+nwK3gz25qvpTnMlmfHuuhoN4c2WuoZeULkeM5d5V6Qnkdt1m+z
l/vz+p2b/KZVu893/EghHyVIXE0zzUqhgx6GyfkIw2euKgOmh+FSX5Eb+lQ1uAUE
uLJVRpELpBlXDRv3jwUth2WIsbIu9f0OHCX9A9cU7tgpbckpYwRmKFx8uMfdnXoe
YEbyBfWjquJWAEmqnTsYEa2/baVObWe8RTOwQXAx6ijU5RXSWQTFyfJCF/uWdMeb
lalUoilJfKz6T3S9wUaCZgDzP6IALcWR0NrRGx6kXiF3PE1qBrrMHqt8DAbOatHL
IDLd4/aUQwtUhwJ2oXzYXbF1cWJCTWNyR6TwxqnxzYpeAzuyR5e0ufk1E9SLHQp9
rvOnQOLxHWsCevAJMK8TCzKVKB6ZoGB5PTksavaVA2ng2+w6uqTsz5lUZleb1mHb
65euRe/SdHjlQbZVzH5CWsboCJ6d8R/rL4J0ooEMnGG3xqDerHYGbQO611jpfCZx
kKHPoEcBatD4IyHPmu+aEvHKDwiOXrbzTpS14qR1R3DXJcf2aUUthJ6vynZV8Fmq
pYJqLWRhWK1aDonaIaVC99QHgjRjJ/D/YszLyr3YIQpkxenj0KcbyOmiQm1mPtFA
PiZgYgNW1QthvyLNdsBxZBWq/QK6SvJe2MGWHmLidk26ORLyRBDUrUDk6jsmcCJi
Q1ssayFe/NVts89VK8NyOe/6FBQ5JVXfjB2B0EVPHWg9KDAWUoL2ZlQeG3QPwIUT
kEVeLP3roN1RD3swi6JEmBb0FJvQxVBeD+VxCElp/3s75C2YuHiGw5cEl4HC8maO
90qWMJiOxFnxiVP4YwsJj6KN2lPxcDnBMlkP2SjJu395n0g3Mk9/8HhDvs0sUMnS
zfp7MWB2Dw/KBkxFpwk1YF9UPWl7m90i+ocO9SfqDNNS6QCVMEq2IKDlf3l8HIOk
MrOWYy5dA021fRSzWBylzVrw4/kPstuys8tRn74saFktjzUnB82RAseentaVa04V
ds2HbXXWRN2PMlrtAoXPs7qhK2M02s/P8MJ1GnCrUlH2lUhwF6gMZrl1CYrfdhnH
zbV30jKDBbk8GLuWYcvBbKc6fi7mVLO+d8pyVoCeLEd+aZE19Zjy/aa8Sl4TPY67
nvn1gyS+otdX4n4Gh/SShpIHZCLEEskzA2sCdnyw5T3WQZWsOH+GbhOd9LU7Xbli
H2kNT+e/2aPxn0+iVfMg55FwqThtGnByKkTe5g2xnQPmU4kzvuX6qK7dJbHZfazJ
N60E2y5z7vl3tElZpHWtFP8np5XPQDreYaiuR3WbdlI3yMGtjSPNAfxoIiVFX/Gx
zqg689OwQ/8gf1upIyZepJi6WHEyv36zXGTyEbEe+ah0qJR6vHjjrhdlloiJn95R
x937PXRiWKOSuQri29kXSRfFuQMHKE0cmqLAKm9Jo4ihYkDvW3PhmXhkA86UFy8+
TJpZdUDpdqVv5YzCzZ9a8GCu+2TBOn8WGVsskvxG6qAcRl/Lv1GbrWOO4FKdg5DQ
747ptwPt9+T94D1ZMuHJhT0VgshmuBGQJFdWdJIOwHCih2X4Q4HkRxxvGb9D9ZRj
/sHaBiIztc50yFKoAccnqoVafeGXcXXowAcIJc8IMpyAS8ZBluMoUQnVR2Xkj/t0
xl0p9yXfTEStvk5I2YijR1R+h7Y7D4izdeGrZQYXP5uoaZ1IzoYwY4Q51xMR4Jax
+X5XE+CZU7nO0raI1AAZjM+OErGAu/ny5e3I017BScS4ejvMKyujioGPMpZLRayH
Dq3gDUyM8IWXKkpJ3oLLdio4jkP9Oc5tDtlVJGk3Axocuc/NPWYJnS4g+FgQ8drS
RbcCGOfbcvppdwCuMjXr8aAkN1+E8w9mHlmZj7xLPBLIGFcI+vrqbwS2M03hmcax
cq+Tn8SfgPj0q8ryMfFt7a2D5go9PyeGdHA2q/yPzHhe0PoB/lfskXvpZDi3uJsd
qHDTAF1BgtX9389+eZ0MCJig8Y+Pi25rzFr+05pHmgtdvOn/uqoaTISJW0VtlKCC
LH7IDrG6DXwpiBXQMD+e1kH+2XxY1DCUZsIGfj3i8ezM3L2a7vxf8X1S5k82Tuam
e/JV/lrqJog9USWuWtKk180xnTTbrGKmMuvbOUx1SQXfDsNBUIADqKA76sf0H45X
HnEIHpJp3DVsGPWJNCRPYWCzZ1bu4sbSAqAFnYpRckkGwGpZB6ofpnrWslafPJav
Qt9MAZKDjAS1n2F7lF5ErZSqYRmMZroiZYSTPv+CeDKUzeKIhFn78g5+UfpXF4kR
62AwZvBkP6IlYQbTG1itPpuGoZ+Oy6Smsd9U9lNexffix5ijKE/TuiZe4zCffFqh
iht3KUtz136u2Rc21jIvgc7pXMsRnRn5wmHxqxflXg7+rYvF/EDjhEDnVW07kmyM
uucdbclAFbLs4g3leWE8y2xJx+3QYGcrUDi6e8MFVYsym5v5he3/BbYS0QM2Wd63
7DQgPk7qD+w0cWjuGjFuw1kj2lSehyIovlgXdXg/0ZKmLq59LS7OxoRXj4z09yuO
I1LEteKNw6G+pRQyUfcaE9ACseVEOvtP52gIwYQRP7p1Js2XNGwYAp0fJn6vrTnb
Ms4TbJpCPkeH3+FjxLzxCs29pzDfKI+fGTkwLwTWfkzxIwCjxJZSH10P3vEsewn3
Hx4tn2AKNpE+PV5B2BDqTU4uDhHrKGiE0w3RD55w5QJJOmQcxRem5CqgEzyeZduO
KHYm0GDUB474Vo59O5m3SMLzl/v7gn+t7vjAWPYbkCOrA3hLfEQ4fdh4ntmcxRR+
uXjXDNpoBZv81o5ysO28uYPXN7DRpchXFnmgWqHlaeqyquXPGvehU3uH65nYXXAV
YkgOMUl1wJKLR42BY3fHuLW1FoKZaZROWIvI6MdfHeTI4j4ZWgMgWmA3I7zkFapg
IkrAEmh5+Qr6T84X5D3EJt0np4Ql9telG5lr45tlW4nsXnoGe0KCQX1uBRydaSsN
nYu4Pa1i7mQ+0moVZTYBgMfUZ4eu9CpZpewXCVlS4po/btIYR1hoRDNy1W9XQl+6
PlYQho7GIeEZCvvsl0oXeNJLc0L5MF9WWoZe3c3+xte+WGLmfwkrF0vAj3s9RPcw
4ra5QCmL/BItQ9g8g2j0Tomb7JLu5tPG+rb4SCpg5EVGEeUTCkeXR+l5n6IDyE9u
PG08chwh/H36NgzYLzaCp1BcjCv41zedOzuXcIPytaKSpiP3I5T33O7i0U9xv2y3
YXUh2dBc03VGCkD6kk+NDcdPw8VcH9o/e2SzAeczw2/H42fSALuQiXY3Zpkp/x+3
Mgi5dzNSfFAho527Ii1zIleCo2pIrufwLM2e29j85D0zAo+vY2TiwyXhZcu/MOD6
ImUYEp+hyv52HHeq2NvC9S0zkyiZqUoD4Jt3ejCmx5lwwUK3iwoF8i3cyww0dCHg
zCIsJ2t8cmAcSQJBRbtOf5dpahT/FIntT8V74L47QjVK5iPEuVITYcHLyhwgAaFJ
rfg6XzVyqZ0W2yokSXSUR49WJLhtq62kc76dAGK6Ooip071Pic0Cs8z/jIM84hwF
e4MU1DnPqX+IqZ3m+g/76HQDtBCxGFAqm77ZCRsQf6GazUEJJ7dw4Nc+MVnCzhJa
enE8dGofqE/cjfm3jOxyv9B5kBtubVBpKf3DscNF/2LFxPcxVp2uLplogGZ/QSdI
aNC4wCUe0JC9PFtoeXLAeyemIW9Qttp4u+ShBXXdCc4a8zJCaFogYFBuKaSznUK/
goXyl7Cx+5qtpjJchWuvVqTc2S0kmSeydSSDoWfDFruHsbv3ImkQ3oXsTAOMrCKP
17sIgMctBWhdgHeQurrOxKzUyG0hF9pOgzRWfNRvN+i4BFl5O1jWzAx+HnG2lHhH
0NMXfdJts/J8lxQfIo/RlxhoC+QFGbp98N6Y1U9G9IxoKQOWxP8YNfV4TEJGnDut
6mmu7mMnTghergEOA6lsBWZ9bo0FXj7BSXktMyeuXeOiCbOu90FiFvScvJJXwK6T
hoX80maYCixW5bfV3GSYhBbK74QxE5ZMOB23iyhyZbtewj54SSZ9DqULugkwZ+3M
u6HDgx+HRDq7Pq6U1gyxwnK7ER1GhtQlsk7HNU89kzr9exUOEKHbav4Dm7WLEKA9
iyHyk7P6kHcxyqA64V60pUFZCYPyH2xYctqslbAvt0WyVZeeY9QdLfQgaL7kFw4S
tFmVQ/1BocQz/M4JdiP+w8A1dX75ZG4OAP5r9eptSKsZavFc+02Z+oM6S91diGcb
ngMWzoxI4FuRaDRafg/UqPDAK+rZN6+Rqhao4nOp+zwtvJEUVsM6mzOXBJiNNDJL
xfjXb0Dj84GHgi+V3zd2GeEE9t2PEUWKk/dLqoCMfpiAuQQ2oPAVkQHgrHPcEG2N
9O7SB792e0sUkY80hNOYa5Elk1gimWJ+tkP8I4s6QVDXd/MYoIyE8iK0fgtzUcQ2
qIEZYLS+gfMTR8kWkSewBMACwD8TMhyYfJVYTQg8RMZI9lQW5TdWqxWygfBc6bAr
7MOkskZc19WP671fPsGlWo0XtSnFlz3NXenPcKAXTPupnOg+yzUsoPdGn7779taS
ltdJleaAzx66NtIV9NGh07ZnEws+6nBPMESdoeB6+flZwETJkC/sImrQFnev4Vub
J+AB/g6WxTtJcHRLNLVsaeDHvoGggkzsREetiW4p0FtKxS3HCRcsBqyvleW8u2Di
dp4iUaykyVUtEpNqQ/bNAD08GTG05ScDMhgT1KczMlbn2mxkztP4ZrmiC2oTUSiK
Af4CbJDkTQfKIl/E9FGX9UDRwc4zWmReryHLN3wotGYWqNXmZ62YBD76Km7yqpuD
DU6j28m+zb3TK3ngK3DdUbO1reI+xwEjr0xtHMkPxU4B+ryZ5kG5QspjH2jGNZPV
sFLmaDK9D0AKEyW5vtRXu1kV/4YHkFtpy5WDNgerXwy4kqkH/0SyRtfoun1VIoCR
YyjUn9pornv9T2wTfoWtoNkJ6mkja3GvR9MBtLswiNvFkKH2Cho5Wh72lJM8yCHA
DN3NOn6rr78aJc13L/5NaZxfzwjT/fKMoXQGN3VXdMVyowENr9kSVtOanvb608I3
DrUGyNmtJgQx538T4U/g8eSiWVBDIMKVJu74Y/VdWZStsn4iNrO9ZtNEi07BKOQW
oZta0y8u9aQaa1+0DpIqWEFphOw/bRh2zaSu3pqQ3qtDPza06gUR0SIwx+a5MpIZ
wCs7lhYz00KR9T6V8nxQyTM6XQwfY7D7w56p4gFH4NOr8990OgZ8JkdMXvtcOTQz
RFa/t42U8dFCRn8DJGhbsPVwnAoZVs8AK8GX1NPTnJPQUJ96hKqkS4u5bRUyTMF2
3ObWCBPfZYryf1JKZCB7Pb5hq0jTfHtsFOGTsFLDz4ebgaWzErYYTQK2br2sBR90
EHjyAIe9irrusgF/wuhnJdN4rDURwgM18I00ASrMyd4aW2t8EtSVn9pvdrrdUDkx
J/X/abSgZRm3ReTVOFs/reuG+I+iZ/Is1ZADscvfm71Ov9V+nQUrVHjCzK7xU/qR
tBKWYYj5BqleZkl3LPNoRLtZmoPvGzGU4dZtBR6HeeB58IclAYB+f2Ur2ozT/c8I
DkBn/Vc24nYzCz62cRiobfUO0XC/QGuVR5j/8ME3cLM/1psriLNtINel2DRVON9t
fy+oDm3Mew5m65wzmIuZe4JijSh64TQBLw7hCFIsBWC+hpVZB2i4XviVqXMw3ppz
txBkvP7kN8Fhb7hnV46us2TamgltbjzOta0/6OIBM6dcv6duD+iIIG14gIgW5Fwk
fDXBRnxMx23mdbRG5Ut6JWNcGkxwkt/JEy0i/Ql/w/XLkxxEiAyk/wyDAwASi1Ju
MJCLnSvgDoZ+pgigTCZ407XB0H6Lbvy5aYpSil2tBnjBo9T8vaQrux5NASZQ9FQk
68GAfGD64ElVPebL65i5HTPlA48pAEj0lJo+pBcIOiDM2PMByrMnDXCm6fKWxmd7
ZOu8CcPMlUVr/Fj/gOFAzE8eda5w8IrpXObcRrhUW5pBz377AODsgG/VPMOg/50n
qym8HSMff02xQ1CYzdALxXFXPDDw0YbUFub56EXJzv9JJ7yQ53z7uYtR/KzbnXLE
UOXFvE3q2PCl1xH4fwwVYXlbxp80AxrlF3O/rIlC2pFQFLveKAn8EdzYtFOailSI
d5P1HXP6DguikGT85SKqqiRw04HBm4o9uGlytOrM+88wLVEqrMdamW2kR2S2N2nT
6JFIOCelEkEk0D/6WmFqhT62p02uKaLQ4ittC9Dwe8ozHgqk5xUkQ2ieezDJ5B7t
/SGiNGP12oHDu75UdyuRiAdX7BWWRiwSCs7YcLdyN9PjeJLfF8zWc3yXdW25BAi5
8pfSWqGHfhwaTDMOF9HV7oBxgWVNvQmqfBLmPa1N4OQNdpAbKwg6Uc8ZC/zVi71Y
A3ulcMpjshoAhlJ/HubZ7yCVaCoABGnmL9G41hgoyFz6x2lMdhBOHJN+6LK/kXTM
a9cxTTwcrkIeZv4W+6LXK/85/nFyhMlrmep9oF1CISHkfkhiVW8WHBtd+DlMp/Qz
RoCaYMwDnSjXDobepnhkAHe9mibV6otj5e2UsiiJKWeylhggu9j6XuOd5EdCssj8
m5gcY9Ki+061Z9CpaLHTUvRRJuvVtqwkyOlXQF/hkwJnGvPbRSZbQbHG5ieS2Txg
jipgoXr2gCCONIVGQ/XexXcDZjq7thspKU9SVXZ3DTlFH2QzpIQWnh8wPMsI40XO
VTJaf5bRW1avp1YeBVfgVfZ+WKXymaZIvzwY8Q9kK9VI8oiFOG6064sqX5v3anOQ
W5VCiCegxE3NjiOZhNyzcZl+z5on5XzzXR2qBsRQq4qlFsku7N+m9UTZl1k1psRQ
4JwDLGiiXSR4+mRKmTYFjYErtpdzLDFvcSIwiU+42eD+ZzBMeKSjzV8FCxnr/wuQ
oN2fGydrEN6SIQbPv1HNmZtp8J8WyVaZEWfrQNP42Q01DK8ksexinXLTCo8repb2
ahtUqBYcH0mugTPZHp9uIDuhCBwgz5TwP3AYJpyp+Sw8YBbGll633DkK6gVBGdEq
BoJv6o6LcwJbaayHpWrMXi9OvlRFOf8E9C9EpMxg6fJpv9eRPz3R3VihRt1TSzvi
W3z5rIppAeaaTqhkRV8uQt5vatYMIfKsg7MIhn/Rpf+dxNFw8s9qcaxQXJCdyByP
bY4enzCd2YAn5DDUnFZiQk24GSxhhgjdGrcAkyWgAAhvIt8LxjpB0vJnpKLdwgvL
pvXGt2Hw7HCiU91TwiiPliF8QVXe9IGVD2gf6t3V7UOnzSIsDY3GeEg6BYeTLJdE
fTK1D/KjDMS4w++uEh1vOV20JYhNfiQXYDUefc6obWS/z6xvwArhFRhv04vknWUz
aQXulTKP30j3dWpwmFTTdovlS1DsffAJN9WLT1G0aVW4QXSWcI1Ew2kDPhgDPI1f
mBakCjYnBoEdhy4E3QeiqzqyqXFf+emrADgLFnipdzSUYEzB7tlbmQB3Z/sjoCv3
8HI9KzllDW/eGXhGwJRbrfERD8qE18fd0QmLO3aTdHbsQq3JSvnudrQ93sHgNdm2
MEmaSUFOAnpM8uNLkbcsVKP1ar8Fv46ANlkAnrkB5c/OKBCtrsfbneMSvD3x4CLz
n5KQ7cffVM/k+kmBzc85somBgiiwnY1EInIb8JaSBjCSP7BTYepBIb48awDhIufU
LvxDiDhLygbAxaQIy3xGome/d00ITGKRIEIrkYWfcRU8u/0rWx63Ya8fjfK3N78b
seASO2x3xnTYQa3oiWAa8i2kLL02J/mlDgLhSWWdpCaxBJYYUS/Wb6fN2f316Vzp
vtqSiWrg9WGkvU3H2bVlQVwij+b5HTOX1pWtsTATFvXZHx0lWuwIsadq+/jVIyBe
Mr+UwoD54mMi7hg+AqGoD2fzsNPF5z9Ufs0T08vDva3OjQTN/bH35cIxCvTJ5OWk
yEuP+4NWWrNZQt3OmVRv25AJMzwHloX5u2Qx1NdShsl191gjBSZcjXbapMVuTVjZ
898LGHvjm/Hai6FUEeN/j/JFc6h4DvVm1swrtrS723ixqzeb5MmpIuFLPRA4ES4X
rgsVFPEcWjx/d/T5kZdEksEnsz0hs+5BJTCRVxIC0QQjBBZzZWq7KJhdv/TEpjjz
Mxz7EAxcSL3g6fGQbLFYxCAHM/lkMHZqfige2Pw1yBDVHEQOwYGBMKmsOPhsoDoC
JdUC3meVLaqLMN+Gyy51ra9NpuqqZ2rzW9DheytWZOglITB+adg25xOWM2PgQq1B
8/7YBk7GG0BHXL45uaC+kF7pVRg7c5ujwIwwlg/2PZbNiKTqc/aiU9lHBCXoylIJ
6NtFKQO0GDkDOUEUWO6Fqu+yTcKcR+OCs750VpgOQIM5nn/eBiWPp7DrPvqiHxQR
JzyEWraiDgUMWsSoGvjUIfNA1cZpaH0ZtuF5BBeT5gIuMC8+15l5XxguRNu/ZT93
QnINb0Tl2e30EZkSrukPXEVXlDm4TkynM3jyonDqFh1uPnxIEBk5vMpH6EFcOi1r
ej9GoctJkOrTO7RsINpQXWLP2t7Fg3ScZBATeSHpgJgwWeqqtGr+Bzm14PzUEdru
wUoITAwV7nSkr3h/Kt/gohKz+aB8KJ5/bcRZAXlGYqcge/8K37aPXm+JQDMwHrR9
Gu+LXLNrTfkoZCYXyFqBlh+ANc6AnBxPyfuafi96B1eIfNsi+OOnC5NARTCNGUIB
p6v1bHCa/emhOBHDFy9zq8VYA9rJqL/OjoRNrhn/nTBjDoqCbDL72NfLzDJmwjfZ
HTDoh5p3eqUKt0dXWPoO3dyDMnu3M+P7T5U80DPp3HuTqwVpX94B/d8Cw7rHZxY0
39pWR1re9XVsQ5Tf4wCVMIPqPXLRFPDV6SzWyT4Sqo/GB73A+8uCuGfmPx6BSS5/
2CMS6yW1Q1tdrdLaDQWI891ScqgpbjyQkkg059sGMBl50ReZLr+7VzvjEXP1ua52
aeZofjFp/6pQM23xvSuOlyrguylNlR9XflBMMM6Ziyg73aldnp39yifGDcxUBajw
x/ef40R9kqZeY552f30c3KPH1gneOOm6AjrhIcp9aJyroLcVkXgy1JKIb8DgX28l
wa07u6DTSRF3pm0NzOmtR03TIKXbEvQQrV9MIkliUWZIf7flDQXmQvRIIal22Xa+
kFUicT3rsxhBs6pZD067IjmSUZUD1ArBp0KdlFDOY6VomlydZJO3RVw2um2o4M10
zUYNctMxoIDNz39cZq9s8sJLTig459NhyhdZRZkcU6G3yFKdyAzrz3+D4ZmOF7hH
e55MTVBvmVTj7DIUOEtVfUAdfZRpMDgo/aa39SMaMfr+TJhi3dRrSp3vz8qpna8f
+6dmMxZN+fah+JLMil4Kbd2GvZn5ZfYPymquuR8UCZoZn1kGd5KlpWw5joDGtLkg
o3Z/OOQA84fwaofUcK/emR7rixr9nsoXLnlv9jiJRfksf3uIYEDgfuCwNaGU07fM
FKt3ysNjoGohzfFvyGdWrK72hRh3pRc41o2n1pFKNZQgvszIR4WZCQz4TDp6PtjI
iQVEPlDDBkE2XFhcDWDrS/FFl7CGwtrUm9qfT0mwBgTL9WD0zai9boJwv7aBtenm
5/XzrxVuyxR1fTjtypqH+RLPHGe9x5JkhiVCEDIIU4NR1GQGX7qKOBFXrbNddcT3
azDb/LOtflff0y9HjQBJynrm9ZVs5k+z9UNa6y+Hwt5xV3LQRy2bpDcl3JQLMdNx
FCIM14GRAQHdSOZ8lxeBTTcNOndKs3r3jM6DZ0VnTdHHoaJtRkD26Gdg+c7Qcjps
TzKRouMNsPewtS2T04zIGFZWFW2/oedpq/+O78VUR3oF0blEHRwSKX2MX2FOszgX
P9l4ZwDozbQUqXppERQM9GXVMczUBWuHzphiQMnKt6LK/fIAh8sIV1ai92ZJcqdO
Q4N+/Rv7QY7qVgKp53aImou8ANueeY227c4VZuzJ9xM7lPrhl5yPRcR3u5axNBNA
mTmuxS73l6McCClZtfAMS4Q/3hFZ0JRLAHneHSki0inRqCcYDakKL0b/u8KNGgBB
8L7cFVVdKVeYOjq5bsIx1AxVM5Tf97CAVQ0hI9bLKufa73fThauqapNUHmE21WP8
zcC0sBXWEr9QG3wGcDqLxqsVDtvgDuY4i17uvna51wc/QpMnESktYiyZSDIr2z1n
wZ7anDemdBO7Q1aMSfl9hfY04iMpC2ViI0X1q3AyId2EpFYXllB8c5De3jo87rAJ
R4QDbAXVLG8NPcuqKgrscc0ufRZ7COOPQ0y4Ac2U5DaMqAFdG2q+Ip6aGsew77yN
RoyZ5S9eVuBB7lyhAFFiTDjllwFP+gl+uKasuV0d+JKa6z2PKOex2RT9qXm8yqT+
DoPBFtAm6zlOguUYntrsFwas6/v79ED+El+chXKoRAEiLfsA8vUStZOgwBWFxVRi
BAufsEFLv3aMUFNartCqx8TGyfrQNfADRWRbf/UWh8ul7S+PDLqwVSrZN/xpSaPQ
eh4lT3Is+TTvfqQklmeTrbm0k83P80SpqpBftxaKkm+azHpK2W3npaSvz/IAzXGg
+0IOnvt6BSCuMiFbK5MpZsVRcZquWW1ah2HbeozPzhDSTpsIxFE3RX5oD8HQjtqn
yedWoXDYaB0Y5+IUJUiPLt0zrRzTd9JKVyG1wbGo0pqbMNpNRqywFLR3yI9jnMeN
qGOZdEaYCydVZXl79f9gHPhtwAphghFaO6SXNguFrhdf1Q6mcipMG1/P7O+Heklj
JF0dA/XmRsUd1x2Ed6dPlMYnTdo3o7KKNkdsW7iACMT2eb3NhTiQ1WKFFwCu7+Nn
OJVV88k+loLpkHrTIElv6NR/j3nmQUsnHMuQ5NTFW/mOUlM7+YgBvtXa14Gm2aYM
mDOqBFE5S4tcso0fm7nRHTkavme43gzhluNxCLOFoRTWoaTy/PnYxccnkxg3AMcc
OErstX/WhzcyqRROfR7zh9Rkv+3HWMWmJqklqiBGLN2aAT95xAtsDYRgF5WtDwxZ
5o9h2pX0ETsv3EXOIBIgHafjCTRxeoafJQAloLyOcEgko84Rf/lOdAE/7YbwFm0O
+zS9xXVyN6fHRaJVTBdkP/3A5xq+DMPV4KQqDcJWCB5qvIrzOKNknMSx356bKplj
tX6cxSkyjjUK8bgAAoQ6bdamzpl9NjjMNdojsrFF2uuroGZXRHCkd3dfgGuOv5ot
OMuYCeHjbOAuoHcw1KUwqwen+TWKGr8VB4kBDgCPRNXXHKByL1aGglKVTHrMQk1H
xWW7W2fK+P/n5IRhcxYdPrOlm8TZe2s+BbAAhgUy0eMvn6GqZ+HkqNOUJDNT9eSL
CsAWg6NzAf+3QI+l7pkrReEdcZRHH5kaVLtBUj+B4gc4uGPVVmgo5RByt+FYS7B9
zHHmB6F7D+A934H0ptOo3Ws5Tl4qnROyI7OexO/71Ia7xOSMQjJqVmtn/7H1rzU7
D/H9g6qZRyWSzA55RFiRUZqE1wkttIrk1Xx0D1YPCXG556k9EmrtY2t5D/Xiv4UO
TkdtXT9FNWrWF1zn2G7FZyW5dtcyTYNmqr39oNWXbiieB7Ogsw7ljqxJXBgvMkNZ
ixTghT9DfTeMIiY1x5YRA/jnQ/Qhxh3G736dZCD0z7xh+Gpj/G3H1x4WPaIUngA8
MFYnZD9CliIJIx+NsBDmafttJP6dcMudNDs8SvXns/98qfsal0Hgmvl6brDHWD4o
zbw1oPQ9wRdh4K6P0/zK/OHqLd5Z4VGu/0RZZngXX0ypLbNc8pyseNqlKl1BVFzh
0fyPQiZei0k4yvMCw3mkx0FhSCe6VaNtnjE505iA2bugNuMIG/Xuc3lkTfLmyQfE
0j3NuPbe2ZMTieVJ/egrqz6EcEM/kp0lDKG+nS/aWyziCNZ/IMfmnPkfx/m2frx3
sqczqq87WAAvL2STmcZnoZ1lf8cJd7KZK0LP7YL/w1xf719MhWcxKRiS9l6Dt/Du
Zcr9VPIERCavmimI/ptm2Li+VBECzjCd8BVKxooKTZBC43MWLsaDRs1ZPPPaNSwp
rN6aig8kp7fA5wk5O36FL6EPxmlNQh0lwqO7vgRmL3BXN5TLmoX/LeTckIud/+IY
svF0g5953bx5f8Ob24yhG/Pi9jklme6JDw1duxzrCFdK8FbksB/QDPQS73BasWTU
u7GYXBNRAcxcVpAThoPWMapNLyM2/KXH77mFNs8val54APtUP/aD9g+ftfWE1Xtx
qCuOIsAY9oCJXmZP2aaYCn3yViNKjbcerIECTTFcZ2SqMAOHFaVshK/I8C68RGsf
cEmc+UJVJWUVMFT40qtbKdF+MdMdHjRvkyerAOmgOzQD13y0ATk4jPM/3MIglXKb
Sixfdsj7srLTt1Btskp5uhogFPRGW9+jwwwypoEuAdcGAypMer204C1tcm7q+u62
eRSQMexogZZry69JJqwxCA6PS3dkPBpptRlsQho7Sth/y6s/DDxsg2NZbc8h5Vhi
59BnnXUAUzoFvLVnWANyUrMzSj1a7cOPVfEbu956HiGkec0McKuU8WXpQXDroDR3
uekNMgNeinN9Sc3BJNyWqUNTQjMVIhOiYRWXs0WwUA9NC0ygMWZK5K2+6GXAt129
hQwsSNSvjoVGDIdUA6jAQ2xt/+Pj4AQcNx8/8F9s3ijaE7JkGXBTeVSJYBVgPYGM
3xLuN0Xkf1ABq/xt3HS89kEsVnNEMULsr0KA1W6K8ga8IuQByfhe/WeP2ijvyaao
2XI7kwmWAAMOSPF5Hl9FPc2RH1LeykQ4rLInS2ykQof1lc6cRGs4nxsayvCSd+6g
wWwfKguwJRCick3o7n4UNjNWTITR3aMpbIdbVi08BVxb4BIVPp/DcF/I84lqvC4z
QuVaQse/TOGOugpXxdozlWtpCvqQY04X6kgcjo4f7lQoz9e/n/vTRA4aHjRF6FN9
LFESCXRTbaoKUcRzDmgRlXGLhkR4H2DTHqgzaY7UQIJJsgSp6CtyLSKOTZUoZ0gr
JnDC8ug4+rz3maqVwgP4eON0qSRmYDlW464LNCafc41huptSvAMszPmxMcD7yGt+
015KrP+V0Yw+bdChVBfEZ23HLQU/7OZ+VpOFHJd4l9KD4ux9nfzpo6c9H0FhC3Zv
82zEY6IKLd44947WemksFHKRW4CyXa/gWMrmYHz8mZTL9xSoyx2vEjU4ixU/HbHJ
+N+CWMM0eqE51BAXK8RmeobfVlSn5K3BgJWidJgq6HGrFn65rkcIaAnPby2CpmwW
VVh85pA65zkpejsGCBu3NVO/IFqZJC415fYBDr+fLKo3/yliJR54TPgD7GWb4bpv
wZBiIozxmqFb7yyN4bmltxh0nB7y5r4e63NNxtvmTGn/H29VuvRBfuB9qm/ChCfl
hF5dF6IThHkOSFZlnpxBK/AxSAnsWCWP8o1m+ytS0xM8o+MPC60nuYJjjJNSO3ID
QsM8u/U2J8T7GlBEpS/7vtqtlwYEFR8Urw0JntKPVqPzGWeGdXTFhH/+0dpOX8Az
a8yqxnGiS8SJvOyo6l8d8FBUhLqra82RMwl8rQI65g6T9WPmkqBiEASE79y+s6a3
Lv3t7GoJmyEL69OeYPsEEXmizlzasPRr0Nc+K+TWldcXXNQf4WEOuIcSRNZ/ery8
dLA4BzJ/2Sj402BnOOhgG64qIn4Y4rmO0vGoe+E7Z9Dlvs62z7MtjhTWgVhCZpgp
Te/EdKuqUyP+hkUsLoyp9CuVTg93EhjT0ybzG1n2Xr+F7XacmQQpX62oIoDyaM+U
Z/iWiTuBq1gG/TqNdz0HcE+V7kXBqBX8Q7zujbbUZMLTP78LSRTzqYCb6fj0Kugn
PcxFUDTCthjNjAcbou+MX1VS5rpNSt7Kpo7c/03G7CSoze8bxQ7ZAl+M0UnCAqv7
1EePTTmVep/MDpGks7/taIGT9AVwyxuXXNjBytkdEoMYdyrESWZS5B9RdeD3kRSR
nmJYo0JVBepEno7fksefcugZ/BY1Zm7ahznl8MwvA2KP/gCEsiqBfYVKZ6xcQAe1
d9peGa1o3q55wWsuaInplJo2xiInpWMV680sDHhiR3oBI/ff5OaErgNwEOSndwIQ
ZFDj2BrQXDLLLnjjkE/0hmtUQ5kEx0x+IO5UZDIItOXZSabBiQJE9aquLkm5GQXl
tOupKqsz5bDZR6s/oDNbLs0LKHLwsZ1+eFy+j1nt14lu7w+OsvnOAbH/LyyqRrmo
LHogszvb3QQIhHJPA+osQ7rWFkxDlHDIgbuXiBme+dXLTzQtFLCoob+3sbRa8Uo+
4vv/KHc7B3zX5DWHmiQL3Wotjq2P/FZ8bs0Q6Z4utUYlEzrlSicjU2WNUYHKlgAc
/u979SSwRKsyfut2JMsBH7ZMor253hBa+8OhridXqhjVpt7kMRUJQyiSC7EWTAEo
ErKMVGZy06KpkHoxEsM9w6X2+zNyDw7r0rtEQpK5N4/Z/ICHqKdX3TrZw4BMQ58L
di6T0cOGCEUdaOWre1/axyv7Bv8U8JDbadZeRc6vkM3Z3BrN74q6p/zNEFBXUF3o
mAKEMUMoSXGaFJAi6sVdEmvfUUB8rJLhI0LHJSmtK+/CK2sGX6QzMEx4WDrz6n/j
+MxlI2U4KCyRhZ8MLwOtPV8XNkfNaWIqYRzZReBrHQJxk73k95W1+CyUjvVXx9iE
x2ODiKkc8L8563J/xeH9kn37BgHtpFUxWlXsDH7B3OSfPLrhUvFcddiN+GcB2EuW
i0ebm2h8WAKrl0FiLrMXg0Oo+OR5GIF0fIncZ7qe3QToOam4tOqTwz0s+h6AC7VV
XQvO3F/NlaTQN2e2csU/T3EmflOCjR61CqZ9LYP8L88CUKQubHhWjvFsbKR46SVk
kMgHHcVFOWIpm00eCRSY/VDef1PVslxC4kN0po+sOyX0EcANhpKaCj90iPs/9h4T
UF+WAOk/mqGhwjEAJpql+y+xZkOpfD5PWDZAcsQ1U7pw0bb/lKltxdWUT9C9b18a
MmlLaThFOXNVySCmfM9WFDcIneRZ6DzNbHdOrlK2vjOAIGGL89msy0Pcf8ZAdTEm
RixZ2zq4f3wimf2+50LuLMVpk6j0/kiYl7eH8A7DJYy1gGrBB7v3Y7iAOqxoaPcT
m4DlCw3+qNe7gn3iiHcSjmCjDKDZ4i8t27YNhL0hzwqVivD7XrMwG2WQ5vI73QBU
Ss6cSsSRmo6jLnATQrTzuRGCqL+T1B/jrxdXibdxa7u39FLrymlaehJwgIq3yJGH
R6dGqNI1ew4dVyJn+NOsyptRIpcW+IbJiAhCZK9qhet9Wba7Dqgx+ZgvSR+zmTy2
AdfPrActtr9+vnR9OJALmZLkhMpM/idDK0vyIIpNh9G0T9svaQBUR+I1E2muAmhK
9R3tv+o6pJx6TKYBUvCbPqMGaRwAQIql35SITGeGPNBBWb1pD7E5D8TPMBicXmXU
cFZSOt145PvFzdx5kQWh3ssAdlIAm/pQk4jLDqqfLKHLN8WdI67CCR3vADWClhuu
RtQ+VQl4SWllplIZAsXIbLJ+G1Mu9g/MX/9OSirJ/+imggbFt6s1DloW/b7dBW5A
Pht4tFau9fwfPKAaQqxXxzmxc6mU2gez/3H5BSY8w4Scu5u6FyiW1oWYljJ0psnw
xZmD/O/XJ8QM4GPJfUpOTFplleT+qNjTKDvLcYBF5em4W4JjVFRJgaWgJsJpJp+s
HDsn2kbNTOkG80aADcifiwWPzrzSdFtd5nHAMMDm9NauXL4fQcXwhOZ7imuEIknq
bnHZEicLiAlHQTNN7Gr+TDKSc7mfoLWF0rBY2d+3A5lKgWsEGGsKE3IJYQ+fV+sv
rrmwiZRkWNo9I4IynXjo5n9SEpCCeBbxoIvLkTW8KlfECjpQZOgjOQahD6eHMA4+
WErfzxT86iE+v2pJ6viS/lB8TgFCs1DSX6FIQpLBY95BODhZtAksXJGyv/YsqKHv
a9tTG3v9aAmGQDO11IIB2hyGXgrfc5fx5XN3Cg5dZhN0knHC4lsgfINs8KAjEB0J
oFiNBulHjRTtzyvq2MXzNbKnDd1s2iSOWQeEVIQ4NACIQ9Ird4Iy8IBk7R5RmOcR
voDKmMQ56KBYC2vl56omZdJ0TPWwOJdIT6MF/MxaOAVejA2Sp6HrF2Aaz1jh3waH
BkHLHCRRVxlBV2vVKYneZV09H7SGZCxJy7/bCW230q+t9cRw5HWRd9E1sZMYUT7B
p8Bxg3IlEyhbT/Z/BCXA9PAxm89EnNXMW0EwaXtPa7thQ9ONozzstN3MLQQQJxtH
jCMQ2+qT2rXC9KUAtIAV7to7By2/tnq8i3MAwmo39l2kdyXZQYhQzbstgKDpAH5+
pf8et7S0cbK7hyHHfdF431QUjVsRZYmyYz2P2TUY1+VajHJCD0NeJOzrDAv4TfCQ
gQ6RfeDdRHL0duYPkC1dvJvYTuHz/TTFtvCYbF8WHO1Y2pX6oc8pr1z9xgrSmh4i
rAWPRM1CJgYiQWdXD9QYBuTuJOO7g9lxWqmKcGzlFpsLlfvMA/mUcnF0Vc+JETwc
Lbggajt3n4f9RrIpFdihU7JSvDpS5Coe/4F+wFDIwS9rGJPTVZeh2MOio/LTC+VZ
LjKU58puoFNz/nLDSqr5+XzM2celQwlBiOPjkziN8bzlhPSs57FvjdUJaQEl0T3Q
R/82rKdcTzxshgN9eo17RQ0LqF9cgWdrnGX7yrmkHloQMyMHuFzhcrNpAqW5jTJn
/3V+OMToq/ZujAOT8jiJZGaS/L2vGnhwg4JYlT64XRvu1ofXPvAwwW5x4FfQ51y5
yBp0Syx86z8DU6Mv86B+ARudxsl/vOHWgVK5hlnqav2UvM6l9is84R1wHqVw3xKL
cXwGgodf2b5smoUCGiMAl3lCEy91BFw8FxJuXc0HHtFEMLSWlFfl+de0SFexHXlR
WgCHJRYkvW0geFARhlaSefbMesqP2UU7ZvLRLdlFhU4nZsTBEpkTRyGKL7ubRDI6
0W+Ul0Q0gZ9/WZo4BFJD6hdpXdhkCKnRfRmJLbwmb7pEyvlC39kBgRjDnREp3jKT
I/0X+45TeQ/x8WvklybLH1A6v8ar9BDuk1F5R2dA61BEhAooyYDMoo5TmI5gtBdg
OyUj4AEhqVp6o9VxWGIPP8U4X9qn5aAzmUjjKDq09f06z3bWJQB1fulg0GODV3/P
sYhsrStQMca3Uw2MS0B1MABAJMxFiW7LQTjnrPpYA/4CR8sjMyNPdHEvftkW5vYZ
Kv8R1OV/MxG1S4GCJEEorKQ/K0xapU2ikXroLZrlNcjaBvjVK6Op+jNvV3TEltq3
xPiylWdMZtNjrFRAyjpcVl9ui2Ql3vWTH9z2HQCuc4YIjqUQq3tEgMvayJmDsoiD
a2zFJzCHWU6XLxEUnMNTZc5UZ3iphhKyYyTarw8W9UMnahkRRwwH0HYpDz7xTFwq
dg207jMyXVVXfOlIjort/mgcwYao6oD2xLjftMFTm6sZjF72q9aA4FImgcBpH2ap
Xl1EhraMtHQfu+V8chTvfqJlTkxsFFqhdVBpnHP//n4ldYFTB9VwkqduzF+l8Ofq
T1PtFkXmNP+QmaIkgpExQVBjcQZfbFpZnrggNb2vb1SKcZWMKZ8n2jFho7ZOE9LT
aksnhMYx2afZsNPgD9Vwesyn22GSUkvAeTylvIs6PuF2f3CAlMF8HP22iTWvxRwg
aIUDxTTafIS2APusjDiuFZh8ILsFIpn93vEnEDoCPfP8MkSLeHYavkoHL+Ro2rRO
gOykDo8ax1LrsDf8XLfaF3wMs7ByrTobKxlsuRx3xIiIM9MsnxEP+pZ0KYO0QbJX
T3K3TLC9xZcXnkVdbA8vRz64879VbA7GSMa/QOKWpr5xD9L8OCfLBZQEjGq/jbt8
KuXEyMYeEfY1PNvGLBRLMxdJRNecYr91km/EpgeVa6JT43LhvPlB9RXqFS7cb4ZF
EmIKeB2LlN3c3N07Tnc5ZYOCT+nbLMSio/ui2GxSyyG/dxVUgRCBa9qdzlbapZmc
J+1WcdeFweyRrqjpAexL2aCvf5PReiGEQvUbqqbmq8OATMaBYgPzn7q0r3eH1nVk
X/zw8VCgXGexTd04lC/9yxbZVtxOXHBPn1eD4PxwquIX2OypKu4O1+Nk4DlsydR+
TlTWvMlAp4UlropANPcgB7l1kfQA5uImxW2V7Kv1z7dappfhia1/5uRAQlYSHBni
5aCGF2sdmxC/EFX+/RZDCLw89p758rTHpsZ3qdmlpwDh0ZKC5ZxY1Lv8slX4h7zq
H0ijdIjE4ys36UjDhttOgrdjRO4MAhr+pWoiuYQZ4qY0rBnT9vTz64Wdwymyiwue
g52M+w6SNTm6RnrQ9REHnSMigj47iAQcoL0e8SbK3A03WGUivsUhZLOgwUrw/ajZ
mYWeKmtS7Sg0BNxh1VfQzMuyzPn6P5K1oY6UadbVrW0BeDfNawAgdAcISrO3dtei
xPX7qrAljLOyHpPtBOxHYDefwD8rHYEGx1n5OHXpt4aHJLgUY6KDc1qwoKuT2q+4
EPcL1SaXN50RIIBeWwnaejDSo9YtCQ8TobtPKfiImu5yvqpOPvJM5MvOwxqinHRs
VgbKGOO9T7lkxCy/MctsUdb0dLvE5VEobiuvNMq3kZyPDV4EP3jt4NW1PX9Cb62N
EvLv/SEu89hBHyX6yLcn4YBdpAwyhdLqrDr2GjH8AP3z4Q6LKpRAi5+ckKCvGe10
4TYqPyZTTZ3IAss3EoQWYdb1wjDadUt6lSsFtnw6ccDG2lUijb+YDl8Yz6B3SDsI
SsdOBKazX0jF9dceUSsHEmAAMlj1CDmNZ2ILDmkqOZzekkqMZyFIlP/gzZXlUeZy
pVVldE+l0pHfCxnfw+ETfI0nWiCSug21CWV2+oM+js/bUs7VOH2STUMEgiafKeEn
yzZitDrxIw+ZXJ1taH6iF4pPgFQz60E7qFJdxjhb+etJpB3uFXKxZ8zSxyEQeABx
S1HuGNCcXjifp1SvUXq+8id1Y1s1maf75n8sY6cHQD22Rr4B7QqL6NqG0/1ckku4
CittkFCqOPmRZkh09saJCinWhklX+a+vbnkOiKDhf1Qjq0vxo8Xwr5VgbWJU3GSb
EzcINLGzAxAfUMuvmlYOnHu9669eB4OpskDnRGZDKyTIx9iFt3Jm1dtG0IkSz/uN
XLtI5lQ4ov9ygDp52iV/JCblt4SqUD96mOGo1F2PSpDaYcgZEDKvoghcVJuw+LCQ
qrSZO+YVYUNFY2zO5suSmwfkJb1c5wyH4fPZ0Ui4UireRzPYOa9ZkAoomZgC/s4F
jx/FUyBdP1lEXCfvwXMTMUKQPXIFcUQD3i1lQ0sc9Bi7XGjbdOmvgQdqmlpMEt/x
cOWIbayhgp3ohev1IHwlxiNqdK+zS1aQhPya9jW2Q2J/Vh8SEpTxdsRTcQUYG9xA
TwQhkk4Ek9wUWlz3HJkGMXlti8N9nsfPmQn+5hZey6uVJgy4MEXMg/etD7w0KH/z
Ovz0AdXFgzg6HTlBFRiL87mbbuCZkxTVesETZBaMl2JuMuIjAAHd5j1JSHikTF+F
30a+k7RfyixXJ/amkctDvVMPnEM2LLvAyNrCMRvHfQCOl/qYXha4468NFqQzIIDl
3MEnyatgXLh9Is429RLNZcD74Ma5sNjnRffe5vBQOv+WvAQChfmeImK/1KZ9iaoP
B5Usr59PJDYFWaUdzLG0mWyErh2/9dp8tPOlo0FkBLtfkbujFtGkzJDxEfua87aM
sel++m6uMGZcD7QZeCdYYW5vXHs/MfF8MmclQ8461QEFTbo6cI5iDQ9VjDaY2AYG
tjER44cdhTAF9dbQElhOkGeW9PSdpqQeCoNlOApIc7TbckhxN+tWWhlS3+u6+vqi
lOs7I9Mj9lha6i6hAV3GREJzax8fdKhRokVhbPBgJ+/0V1nlKee9q+qB2AUo9mPe
Bvl/aEyOq36IwNvgEoo8RdpcPEmZr6fX0mla/Tso/sL/AjAUJJgGaatqV6UIEj/A
2m+kKUnykKKU3LoWILKSgFTqMiwIlYiNXQy1lvOKoyBqM6ybLgeulv5oJlfGA9Yn
7UUUlhEWxjNDaM/ekVgJbTM1/6koI9IMQfjn6vgKxTM4ylgVsJxUVLTbJFykoELO
cCSW0mlEwp3gt1IDwcLcXUoDr2Yx1M/RnoLoCduEw6azk4ymiYrjhuDxhYqmHHKV
B6r4i7NN1kd4ZQSEPqrZ5peo460bZUT1GyC1PKkFMEam3LC1KAZSEotwks9aQ6jp
AQMW1n7SXNhe+8p8LkVtG2GkarI5biqTw3nUzkg6qhld9z31r5DYwcGVODU+f2Gy
GWA1llHYfmdA+dWjv6RgPHGct6mNW6URYohy6TdwGeDkFHJmNM9eRg2kUH3NE99G
dZvKv5aTBSWO7KPROY3laOE6llJyPGHmC7gROG+sMJhVM4qDZ/d/qyZMwsqhavuh
v9B1Td00/iG4ey9u1wEkoknJhRGo3ScAPRvIenKfNI+r8zrkHCo3U8o5ZCNZEJL1
gk9eTMB0L9XZsiDfW2pkZSsHe54DgSA2B81D2Bw74Xnjr+Kzw+wRm+8qbgX6Tvdw
t7SWS1+suryyrJn5MJqmE8uceZAC9rSRM/0Y6+PNwDTR3x89hG1+xPA7vAvIEgqS
xGxqOTEvp8631ak5WMV0486w6eSPeJsDgmDV15ww/S1F67Ss4wg4/iytVuxHa3d9
FI41ef5asEWpUteV2/s5usBFWJcI3d3CO9aD4HunjiL6f8olCScKDLa8Pz6xoA66
ZvpaGfblTy7/cwAU/E4Bw0UEo/0sTcyUfwLDtDg7bfgB4tDHxvXhzkQr6afJoMUB
DHVRPMOC4+pBxLvP8OesYqnAXAPhf7matIxDn/rfz+DzCU+eoxfeLSEXy/s3+Xfw
X71wuoJ5PF2cI2FgPkP/6ZxFfhfhSZuhE8i9MO6OApwJQJ5S9cYtlhycycc8fmFw
Ii/Q5R/RCyTwTtP2gjYCL9M8JMBHXdvab0kNqiULgB37Ec8YDmzsiVppJ59eePIS
w3ZFCNSxftqXRAaSkUY3AosablnfOQXOOqAwSnICb63Lh5WLjMBZGh91WMiqKikJ
8m+GTQSZWt1hZjSTfmg1MpMOAmR0bikRFoOGM5PCSftBJplMvjVhAdnZoOuNBCok
u8fx2sQeR9J6D/wCXfVjqUQIPxVhSO/A1G3sZGD0cNGMG7Dv6UDY6g+tCN46eeit
jW8KbuofJsPseKlQPNJWdyFHgMEqzlLw7FcjQE0MRFArMEknlT7o5zK4SB6CSU+l
6bt9H9vARtjdh0iLt5J6ygwfpa6dqhs9FOG7RTVxBXhJb7WvYe/alny38wNwIrt/
IPfGXwdpVwmQvKhLgiDs732NEb6RfTJlwYy0huXGKdqRMkSmh0D+iZEzvl4C3FHd
+DZBZmw9chrSWJrnXJ6flQVCiaGN0Q41hHmQOtcUOocbiPaifaRFhEYuRcN8YkPQ
AJcmhO6Lli70dKDSDxXcLK0blV3czwG3c/jJem99jMEaxdqkWb8GUVEMSKb9xQ02
ebr6PL8GE1eRya2HUz1r1NM6iiBvSGFVa+k5VtSV/kQ1q02EF9k6vA2EBe+pT/eu
UQn/5haTK9Iq0YQAu3YwCm7hCiEq8ac6RDQkIDl1Dc8Hhk3U3lBjYkAjAt9c4EkU
Ie0EwnJQWyW7kIv/dFnb/qMRwtGmsCJNyaseoPunXinirvmn9Dx1WCJEp1CYbOiu
76Jjnrr1QIj6r7aY3GjE5LyMQJOx1iHMkzzoC8QVqI5U2Z5Sw72irfhaejSkCohj
xn2k5CUnBumcNZGMbeZoUWuZp+IOwjWsuF0b9JQEfsaXmDHRWd+9nyvCdfSVsZPL
89adTSZSPHG++eFgDSjaCXmBDjNUrmaotf8v/ZIkvhg1YCBGafdMjIuVK4AEZl51
zIm8+I6cWjf7v6eoYzcOoKUzaN3O3N9Id9oOeI8rqLj68MLPy1eoNh4cKG7OyLSk
uF4JOhx0fFY8D85jFGx9DQ3d6m8mbj9oVPkRRb/rkT3MALZcMriftdOyPo23NMYP
0iPjGaqeqKgttG5UdTGXwDpDheNU/oSqT5eRcSId4DiJjagud8zodd86LSQJLGFq
Hsdwjdjj4w9tO0llwuaw0vkTiMApqNyxKUHrXcpwdrPefj6Sbbek6OpLT6FGnH0a
onxkRbTiZzVUjShG1fOO4XSUw80qwtiBK7XbhuGcUB67ZoKBnHKZK+XaSoD5241u
CfBrilkvFTRVaf3JpeVByA5DOie9BE1eDrUJ6NaI/spy5lE6e0w3ueKjkDiki4of
Xc4rvgGYZHJDQRNVzbpraMCHRoV0D6LWMT9t32OWZJjx6UVee1D7CTPsc7BFOOYy
boXnIxRmXdrORYoq19XONpR8SDJN1YO4cX3b/MIwqcnkVAwyaJ0gY9bH/FBUFQGT
K45wrIzG5pF3fS+Xu/9XZ5gx94IlI5beeNobfNbDW/GLHdY9q4pG+E0ySewvKtv3
y644m7FphmyUlw+EG7D+YBOV6/EYunLRvQ1XueqEQ2mnL5JSTWat/NEec+SOQJZV
vZWaSThSNRkQ+MujMLcb8Fd7t6U3FwH5aPB/XLnXfrPjCMOWPYsfxbXvlgxBO/0D
oYY5X+stbT4RLQu0ytL0K6cvUbmsLZjalRofX/mOyaMo2PcvbE0Bz4pLpU6yOmVc
f54fT1zxRtiBrY6CP6egl5i5yxD1oKPU2d3OKMgMcgKeazRXOnuj1/rmohfy0mFP
bMxJ63SanQXUNqvT5EUqr7jWPN109w0dVEXMnq1YhEr55D2TRbCPRooDh+Ql+9pI
dQUDDcU1mbFncKo6qHxnYSXSeXJRwAqlsnkde8FJw1wiqXHyKSl6oruc5AwmsUzS
QaMMjwctH3clhmzGZIOR1INgEwkwM8WGFV6w95DhbqmkYtVtjNEJeE0rT3S17mYf
X/FyWEzzS+2WLD0gjVKP7cCh5/fc5AMEEjT1vbp29e01C2ocQJDkSY5binusfcjG
fKHG6EtHWz0gz/HoCI4cYYq3/ywSchZeA+TG2VgpX6ySADc+C4Bx30UX6dOlu6io
lILg3YJvKvyMslCjeolFvQji51L94NWOJyU6lYYW8JzaiiE8xrnihPPl5cEQYNDq
Q0ID+kbB8gN2iE5Sn2L9cOSafbL2VRBsd3WDfA822GIJWQt+ebw17YUSP0hWCHw5
16JTPz8FpJBx1YhsQXb8UEG1Ik2lCbVQ6vQrBKB8CB0PRLctGf5mfjdjsxY8SWly
AxlodHa/AZuvC8+aO2qmOzWUjs76R+0lnVx3DxcYKq/Rph4npJ4u5RUDQi5ylk6W
MtWLbfbClfil1tMSQe/Pm+PsSXQprcD+ZIceD6XSbd2Rqbz7VjTmed3zX8OuSx4z
8I93gL0CVCDJOATqP/n65NWVz5pD0v9KYoBAwbqjpKfUSWLNhTEBPGQ0h9kN7kU+
DCEiBrhgS/E/WE5EwaKWLib+x7T1vQ14qSJbhaTq82DCibprnzuRX54AbExJN9sF
FVtgJxN+/kpyRFEDMcfLBaymAA1/yxaGwV+bv8bBwlfzOhDpbksMftgS1m7L3FrW
on6a7yofVmeWZfLnD3CxkrRxdkPJkEsWAm0SwkZ6d76GvKUHpj7jXg79tRVRB0VX
saIbzHeIi1a51stBfCMc7JCJDqnQtW0CRSHPSS5/8oWJnWfyiMsVplED3rIlqbXd
Is5KHgbOgoFy2W5g68vV8VKsv7lk+yBHVdHRHBx6zgvi6qHv5aAvF/I2Ci42ktNH
k6GY7m8lUNkeHC86EYHtqr6QUlEwwwCeUedB9FDaQE9Ai4Iyowm83fudXF1QbN8o
GGjw0l0njKMb25/ivSFStxzqXNof3ay0P9I1QoD3fuO8wUMQQqztd5PKfmBCuLKT
JLsBdSZgoyadfeBN0zkhEd9Dgl97+VwbuoWV5U8lUf5TUsyup2EweF1WPhapbuJM
m0gEtdJ9zDX16tTIBXOdTSXPAB+LTLGt38218LKQwf12EKSZF0hcTkrDto8EhTeV
wiPz5QfL3ZymyTJjte5gcBgcz7MdRsTFVbdSpkJrUEcrgqrc9LwMxy0hd2/hrqVZ
AfbDspYVQRBFJSZkvsToBwTQQ4DwZMdOezdidROLLWg7a2ofwvDBf9vL/frXOJvz
FXIMxi23h5H+n8Wm20CACfQ8RwP7ncAXSl4oeBt+3rGtgZvT3thBfvJXVeopwcA1
fex7qvaiFB+zqmNPRv45xR159SjcHlInUxMxYlDSlHANIsKgaKFXmHZ/YXqPeckR
00eViW00VgIkcXiXuprOSDqKFknfUlO9R4J+xk0dEEIYyasyReuLdKmhsEmVDtit
6e/fOVxAEKBEW/Rht8XPA2GFNyLpA6qsjNuq7BGoiIMPjBducCgq/wkLAgp5B9fR
z9MSjhkoAht9saXIEI1pu4huZ+cTCV320v7Z+uORhwPAxh9WqIefuaIBqn/dEi0Q
7iLhGmxRkQLNUjghf+KtVgtBlVs/Z5f4bin9mQo8WoAkf9VRJm0aEzD+KUzHoepd
xE63NPWbu26ma0qeDqd/6tgh2TgxEzhQHqrE9NaQw8ZSj78H2+1D17/nq4n4+mY2
YEzgjgyR+oh7b9mffrb2PLZZevndGPSUlookIdPTnIxcItkPmiGdUidu+V6/NtU0
ynvmMr4XkseBPjXGV32ETXzFk+cxDg3HFcxbZBeASdhV07g5gfe2noPhAOxKwk2u
sa64/zZz0hGsXFgiQuYwkXCBJ04Zbj3dAyAqsidDSH3n3OeZEZR/YpiOXgzkdoVE
oimXQs2JUH1is/IyiAEP2pP4sKbRu68t+UfPvi2jaLeUEmIX10rCJTIApleIj7vW
PsFXK/mjO6fvVgBD36DLKMt5iaDvqSiAYgIvtsSNENKOfAVX6AVdpvZp7vDMfpW1
FvFbCxkYGGOHjgaXB3ixswlNqGUZi1SxkzUZ0O27S/3/oCWzLl8Ex3hGJz+0BMkc
q/0Ve6ar8CusWO0BDLyEs5rV5tS47siGM8h06l+ATO+UIjl2Ddwwap65XbXB2QJo
EVgO/fEtg3V6VM4zNxY6vZ2AIAgQ24lz5BFcaaX0AZr8heax9zA+RdO3Q0qdVyEP
4P4OcH0NLdrS559HGuxKabl7gmuC5jNrN5DkY1+/mDxIMSGKF6Al3DP1Gl0xBKjz
Umo8YZOMDByHKETESgPvSDoAgQ4IuZpJJIk9uWnKuUGPwWpj5co5GU6DAXaFguRX
frA9nb9kozZNDNPSJjbgeOJ2Bz8DKxivT5BXAuY+ZD9s2tDUtn1pWEFUCT2B7X+T
Wtwa0WBdBp55ebemGQS8ml9xbeXLgbaUHkmW/ylF5fK7wBITDq6A/aVu9p2Y8cbB
hK67JQcoJjq8rELnZfS9z3Y08nQ93/3FfSm0IPkaQzQelHNE2OZohs8jQ2GT7At+
8gYICx1SdYzo/cBWGjPGEnZE5niYEbgnRn0y34i13QxllvG4nMtVQs4DMoDKH2wK
Jf6YptUAv8SInFrf9dgXKFD6DuY+PacXO6Tw1Lex9AcWLGJwvMkmP5iu5ZDhLV7q
OscDlpoFgrTHFKQ1NX3d/6aloRXMHjIb1AzKXENlzd5al9yPpZ7UhrTwEnPedt+g
MEW7doj4rtQWwQEmrKn4mfUi/4qdIjGxuDuR33FCJ8sipo0zBQxn3fNqod9SqDjs
+coPzQsCyJqWT6Ui5fyDg5Ylk57+edCDS7WzVu4xYnNMHXHS6I7S4hjLBnaRSMHd
W0aj3zNvGKu49Hd9YXam7fpF6kt38gVOPi/XBz5xf1nQayTkemrGfZm/3cp3Pdzs
F/bs80dFxg4XXNdabA0VkVCYPXzBJLRbwLpQbKw47cJy/wVuuEMai/SPTZ6M3c98
qyBnWVnfWONbQwcGoRW4Aqjegpuz3AbODTvyjZY7Rvlkdn+1zKRTRGK3TM3RIcBl
pTv/wDmX5dlantN3JBLiz0FmlK3cuZpf6VOy4BFVy7OYkf4Wimo2hEufZPNoE3AE
6clNrMdfqNj44zkLK8ZTf29VNhQzBnNB/7t6Q9Or84SUfHV/Qxgunub3pgYwZs6C
tXBnNpmce6+tntw/WzDqXd+2tK1H/O9LxvMDSsUG27FWQdNwdllvTmiJMguH6uS5
KGi1hCa0TV7F+7ss+yE3AzPfsr8FH5+vPE84tnBOQAzAuj4qGL2rkaWBOFug/IfN
RnedfR/orVAAVN4PoQD8ZRE7yGJFM6tHOq+tx7rYMp+GUjyJbDz8vSMVc99NXrN6
AlMq8hqT7O1U8jprRnoosOV3vrwMVlxCF9QnqSxMzDCQ2buhtOhF5OJFtC1qJBwG
Vet6tn4+vEk+T2syoXK1i6vYHu6xabftPqNIy0UkvFxHruZ50SLaB8o7JWauU91W
kzr4OrPNGfKzxUWmzfwbjXKxo74qmTbsUXrc0ASgafMDF1ey0dDtRZMCfuedpArU
OYJA69YzYwt2ErfiIQGwtHdgOAWYm+N9K34Bdg/2Wqeo89FBk7SMx3m4GTbivVVF
Vqd8XFo6LCfE49Lg3Ik81GbHYigLdz4sUwNURLHRvHIJKFkZMB4ki33GtJ2RdD6N
//SXVti+vXFjITYahNQYyV3FeMjOdRrH7d2clow4pnqd4KC+jnGx24H9up5IoJLY
Hjlzf/73wkIYJrr/eaXcxKBfpWB9B/7SexBExLjTmZj+lP7QnBNNwOc12r2y0qRj
WC9DdOegY4dzlvAD6hWJbjcatc2dxUMVui+ATdhMmRcKixPbIaDV3vixsfgdaFpv
gWoEGENN2UGaxD9kjTunm3A/dE8AGg8avmeKYR0vnJP0/Gb+elS4bhcALXJsTI6b
5/rEpguQEcgHkBEBXVSjWIwUVyqy4IWAvrIW/z1I2T3zuWl5VdfN9ywSVTriVf4d
HbMG43YiTFZ3LaUuftErL9WxmFPS0nQ9b9IpURyYrpP+nxp6e2y+IqyeVIjvnXk6
mRjN6WQH9DZg0ub+AwhH42Z2A0tyrZRTG/Jl679Mym5G0tch04iBQOWXGA0oL9js
QAMkiJ90Iab4ldqRFd9yn8IfFdzZbUghaFm991UUbvVwze8CRQA5Ohv7cOLLrtCZ
pCZm9iMB7gb+bDZcPBVjwgwqZS4KV3xe7vPskf2zo7a2rui60OA1jaQL/vJPwPKV
pdgDm0wvbYHYzVxsOuNKVrKpbSyLdYvMXHoRX+l2AMlAR8ml0qKeM25c+b346d+R
zxUXCRzs6z8e2nTgTpzO+vaBBtsMI2lnCBhNNC2oDLalk98AWSb6ivp+jW0Jyv/O
YGBjNr2+ACU1s+SgXn037H+nYx8AR5MiCiaXl2NUEUHiuL7Tkz12rBz+ukaw6QIa
kAvB2Y5RjR3JC1VlSWNCuP6UY+vZNkkZbHbKMv4djTg0hZOp1Dd/GT0FSwqjWpHy
lncG9d830FGMQwX849rEfLoSmFGmtaL8FBDwbNxJW53iSXDUSjMzJ05S66aV9R+M
HPUtWKjeuaO2oqctf9IWKZouzzOHP1YkshrfFd5em5vxEwPTpt42bVWoXF0ikkdt
sIfIGglcpsMoibKib8JbIA/nv8mS3JCu64vabN5cVmFTZHimqMeiafWKI2Q4WuA0
DgsXrlACgr7117gEmTanden+QyyYs2QkKj+ZvULJJT/t4Gyx8dDgLXv1GL6/eiev
yrg7nXDiFGnxGViU8p+23ZnjBBjIsXrmYQu4L01Qfw08w2sRqFUArbpgZfy0nfut
Sp8OMVkwghhcOUfuVJVHp1+UJBneG0NWdgRm43RnEsYsZfkjIROGvDPU0yojkjyl
ZVHAHYDnfBiVw/CAc35OU4/iFBXupO+qd5m5iFmMobONPYDvBCN5rCuJ1JltRVFT
gnOyonE2Y5mHuL3oQOq48OzPvtdNuWhPjoW5RubIvr+Ja0FBvL8xwjgyOQnVK+xI
+oIhjvSdF3VKGhxFZEMf7A+oBcl6Z88DgC/IlFLp1eTw0ZiivpMqG9fHqTFymsvH
8Y/nSgMrQnIXXi5BmM8agE9Q5DDwEhulsLETmaaTD5BByKh+w7qppnmw4XCq39zK
zUGDRjaz2PaCTaCBAanHFe8xTdxur1AFyAKKW49pFTsCQaVp1J4qMX4soo4K4Tj7
Hbj0skLTWxvZHQOtfIhIU6KsK8Mqgb4asyemvL/TDY2aSGQX0DJu+iN03P6XtnRX
vgf1idMuVsFisJQEDzIRNwSWSDi4dGq4RdxorHk5ikVGqNNtzqzQZ95Zpn734ekn
oqe4sMM7eReGh3Ah0NILzJtDMPpozV9ClsALcd2rwBSNYvbQuyw/XWfIO/tYw0ui
lFTvaxN8iiPuo2PjefeG/DuIfroW8uA92wDJDHwcV3Z1wnnw0H3yT67TZiB4XyqC
RxXmrId6ydrkk61yFkI+EMAlwNKkZrNVUwktLIAv5SCKof3eSM6ZUllK9Gqgi3pd
kOxGXRNnmG6HFkKkRvO7PNfOLOrOkc5sBJ0+gHVE4TSnHxuwt4aFpERSFm25p+T0
db7ehwX/WDctDBZ8wSjPiUThXovC1rxhKCi7cMf0ni1hYzKo3cMH9XTBLw5V3bpB
D1cLg8eyN19verFI8yV/xbnKhui+mhKydY8GsyaJlL8jCEvNbYLy2JIBRHbwflTX
yI5FVSGEMWQqzGQ+uY+rxtJs3K7VBHAIiZU1ZHOmRd05VaJlevSfGpuMyU+hCkzQ
7b6zHE5vDjmzZc5zM22au5/WUghZAIQk0iAuePaddAtQtlIV62Fzror+5dePhUbZ
zhfKDqoL38j5cB+NuV9c6zJ9a89T0f6nZco9bCkeuxZS0to4pdt60PUBGGadH8qN
9KBbVofzjlLpZ+8hreDfFiPoGArjORO4KLLajekBNNXy2QAAJZfPw5e4dhY6/5Ho
y/gITBRA9Gdo7x7u8LaUbz+v/nxrZQrXCF1K9M1xBTUESSPKO8oHyN8/ZAo8kByB
C6ICcRThNNa4Wjq2hCRy8OJqPpr4H+OzE/ZoFEGuNps3RJ6nn4D/szrUXktgvMxb
wMkmCp6T0OyAAmxMBP5ygJ0m1L3m2ZsXuVnWqFmgIhyX/GdB5IIQ0U5ErdDVFrKP
zCiQTdUAm+E16YdPor59AB7U4lZqMp9L1//tKXbXBqKn5R9/Hk0ySy5aone+OvOI
SyofFbqqE/zMfIwsio8dsSziAPet7mfB9sKL6HEUFUsiQui9qNA0W9fqcjQFbIs3
ntJLAlqNOY6R53/B2+7T9bJTgFkLgIhZsztwPB1gr131t3y13IJnzVLlj4VBUX6b
bkEee+2C4MUaRE2rgtUk6NZViWFqZ8KRaSC6F6EUjFhbBfao+sVcIf1vInQAS1ZF
vpMtbBdZAD0A0FAbrUb98N59hyOFIW4xJ96fdcH7wZjpgtGehiDfrJHolLp/SPPN
lda0XjfetMHMEkd9TjzM5lj3fEtyEVzOTLnPw5YT4rzkVaQ3StdmII8Ur3NJd6j1
Xwey8xInJfNzdzOwoPLlOjQudzQMyz4PqQUdF5H5PsQe4yRFI7IhqTiY5NfEJhr7
QG1IL3L8e+C+t7iBTQ9V/cSI5zB8FAVtHnSDWvPJTZ3Zt6MHCpX8Sxjc+uRViEbl
5CTRVQCMmA8WPWoncXVr5VS/XHdyQE8irfw3lGQj0s9KGjEaqZKECzaxCjB4btfg
vZmj6jgV+vsgi5hWcIedu54dd9nThDDVwaotm5IUKSwZ7b0H9b4D+vwnZ+BrfQtn
sXpyjv/j+hAGj6FztxtLVkYmacHyPQ818MWi6jSdYJhSVUOoSFQnz5DoxQPUe9rD
oGz2EDn0qVnRKgt9burUrl3coF5VMHyFHQmJZmFfmy55W5W2FOqYq0AQlE/Mjl+A
09lh09y5q7tZyO1/TuYdpp440J6fRKDGJI5o9EzDxdw1gVc7aIW9DjHunWgMg3qK
KIleYGdTAuhQL9sPmQajqkBVswKYCAw+wb1k7TxAWt28BB+qirqh2im3iCLzs/CX
BO9fjiQ+oM0t29wz8hSofjU7le9tkhXQ+Dy9rvG1RFzLTuOOllRU/leGoVrAGLO8
HUPXBqjqEb4XTqefXC8tU7JUw7DFtYurDpEDkQ0sXnE0dBHS2AIiJL0UjVSIQbMM
pXVIlYMoV566uZXll35rurrHiGsIos/M+i60QniJRqNzrMtCyFqrbNCUVhrOLSHg
a5488rOzyN9MnolhExgd6g5SgXNgY/FVbz5n3g0HU/uuplOzVyIkarRo7Hu54FjR
lN87iGZkiJ9jC5NfKaZ8KIMSiF+dQ0dnX2RqadZRVDmv193X2kloGtFMZuB9jo2X
fEAkt2XJlqdPHYi+X7xEi1Y4htnvwYvLWcNIuaqGRpMa4W8gC0bZPfach9gcRCI9
U8Wh6099scKaZOc9qFlTbreAgC7EkH71ZvUiOvXA2yDj8yScHC5sQc+iePFz1l51
p5KLUQBWOiR3wVzt5uJwL92g6QXBqcbYNqS9P8diJ8UlfZxHQEBO3UXlcprQ5GPE
83Yo8sHYG3XlL0YnT+PP4lp2ZM8l9mhHqxL8GMBlgzTi4p/J8hJ42IUYzTmTw1nm
8jIabFyw9Cj/ldNXfhT9hXlcZODGjLZr5T53AmXdDh2xTtLAr23hDcjITAk8AKHD
Lrou//zv1L33YBz/wRQ4ACKDeiqDmb/0FjLqCalzDEEdPksaKeA5mscNW6p0znrD
XIACvvNelAwcKWHDZJE+8xTFs22u6C5nfFtqtn3P6XawTN7psHZKwn6a1NOqQin9
XfGNcSU24HygVMG23hFJo3tqgKseAK+ojcB8NIYdhbsIeOMwxwoMVXBDGlcL7zIm
2LNpYvN4etm7c9m6i9XzmlQt8tYiZy2De3TgH+EFVC22GnVTXejPOZSRpV+J7C7P
Q9cUsZx7K/f0TkGaJZj2eRKOZwCp9l9419emG9beLbr+XKhKtucMjr9aeSopp4BD
qSPIpof6EDiYFXjkGypCoENr3o12CdcZvdlBhXId1VvEhIHZ1UfsIHOoOxwgTYTf
SygVQFjA0dkd8Udu3joQ7IHKLaKBNHvcpZjvhn5+kaiFzf/OPiP8zlQeoHS4i/aR
3CIYoqIgLTxqiv92egnVlHOFCMoKzsDgnoWyCVWNMNzw8V28S3NF1E9e/LT9Unj9
I00zig57ou81CeKGmmu89Mh+5wvpQK7RAEVbq6lbILDAJCUnUQAlGh3liZqG3QBr
tCug0VeKKqLLzbx3DnpPuIDeZ5QSrg5z1N5xzJQyrupwHiHLLyVPJ8FgL7uR8fx8
IFH0fIYMJYjVEyY7CgV6dPBFR3oaNFLm75ImSKqAb5ScYFNkt9MsTEQOIXMju5u0
Pqd1cAIt13L6qWdgJ4nOVr8w2H8XfMfxPmOApyBL833h1HVrZjL3RnvZIlET+8BG
D7jXUYB7Q9jz8+JWJaEqMa850x87J+KgbTe1SEVwWQTEzJ1yDkDH5fkU4C1ZgUSz
Ak0IH5ovkkvl+acYBVrDn542vdZ7Cz2oaOjl+mOl1k/B+1KZNTH+XZE67XqI7i12
yK+anUKnqgP5I2ypmYTcjOXenQ5Uol7yccJmU/DCsSgxzf7YVSNRitxHjBUsGnok
KsK34R/3bLcblWFYcTigsPXD11UQPOqg/LhH1Wc18kmiRqab5Wt7zoJ6N1ujX2DC
P7pcRy4hpno/xRq1zAV1CPUlAg2SDLlKMtDCERwKijlwbSCEjSo0XkHFN5YibYCX
PD18SyAg1QogO8dSZvrKBSTXk+CR9o0bzT5Edyda+8c=
`pragma protect end_protected
