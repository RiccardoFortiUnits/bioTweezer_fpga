// cordic.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module cordic (
		input  wire        areset, // areset.reset
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  en,     //     en.en
		output wire [26:0] q,      //      q.q
		output wire [26:0] r,      //      r.r
		input  wire [31:0] x,      //      x.x
		input  wire [31:0] y       //      y.y
	);

	cordic_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.en     (en),     //     en.en
		.x      (x),      //      x.x
		.y      (y),      //      y.y
		.q      (q),      //      q.q
		.r      (r)       //      r.r
	);

endmodule
