-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PFDYwYaqGXUHB+rrNjZWCDVd3/RdcDe2Vj4hMMi9/cRVTucpduODjXx2fj04DUD2wWhMh5iZqwN4
LLYajV+VxTiecw8E4rFMn4NZJ+/WF6qnOADfw/6j/s4jNcKufHIpoEDu4OG1xiTgrcmE+h9q6JN/
zvjeMuGzweanF4S1+CJXtITYBhP3qm/4OIl32G0XBGI3fmMxbBYkLZobzYJOQ6A1HNmh2Wiennd2
74sZnimonLbO02jOTyFzdfIi4M351CyUMzVTpt9IHJemNM5DHRm0eBUpFfIVGhkHu1trUZo1wkID
6LYY+thSgPFjYvlXLBptB02+Fs0J/v7+uuKh/A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24768)
`protect data_block
RNipJ+vyK/TQYy8bxws7dq3EDLDgX2MTbyRw02CCxQfq0K4lZfG/iiwUCmfmksX+lBNK9FMaZ42I
j63QMnLX9ds0HOL2rMNFgBcwQJorsc7m7pTuuCWwR2EeePZfNZBisyaza56KT2fAioNOsObUTgKG
Lys0TjpruigVMl8xQKVskDiBu2ZZe8VfIO6Q7XgC2KFcDnPkkUtiiSfeeYGDVqU3x1VVuJ5pAOH8
2n/OWsa40e1gm2Ci9ZCdSHNoPBe4HUkB51ilmSS33FeVnXhU2iPOu9+WaJ70WQ3NBNU+t4IWplEg
cUrjVGcrIt9CnKxaHz3GrFscQ7bFK3gV7EJCxWbQugZqQx+hfYUceR0TW93ixP3DK/LswLR5vN+0
IUSWpDhqwS/f3CQczKEPnYspXlXkx6K732D8cfILRZ06Mh0IZCq3MNSYW1fYB726DyJBGyCBNPsy
yq8Uyd6B4GT2rS0wpGIkpDfHnRQ1ff6DlqaAJTHHwidOYtsx/u52OnQrLkoRbfYARorFXuCpeGwo
AFqy5vUCBmHBvd+hrYf9mOkeJl3rnYHWYgV0sfWgD8hYCbh0LtD2+Z6OfhU3cY8PlhNMJn8VnUGx
ZvAZO55wEaf/rM86Yt/w9gTaoZZKzLg5PfnAFk8qCrhCvpmz/+GH98rf6tf8UrELFqmHLucJPU9U
H4OJTJth9GSnbbf95JJg8v/dwQTh3rG2Td3Gd338SKj0/3NxWl43z+acwgAtRM7lAVkmM4wQA1er
DW+WyNtd0T2alre34Re56L7Bwt3wmidYAwx//f03fqnMX4fo9KKuck4n2gGlnEkywlhFEjBOE4MJ
VZLP7oabl64m/5ZKcvHc66zfnO2CqYTzN9AHr+c9tsSsvB6BGvW/j48lU6MFCkn4rCt3Nr9v/fUO
Rn8Ae+HYkvd69Txxwd4zLi/QAxbWJlD9xy589ryL66GAWecZtOh5ddpbpt1RC3Tx5AxkRH9RyHXu
Aw8ILtQYmNELzGh33aFG/QycF4QX6Zfn/OqY13bIY+y5MVWlB7dRv7TAlWKN2JyOB8lCaCI9W4oi
z57/fmRGPZ4dIU/yEx/SP8Q7GCUm/GgHMz0LZzAgYRbkbdal1zVfCx/6lRIsZ/2XgBH0M+RDxmYm
YXmz0MIE3KSN2agdhu1IokpUb8wEonKDpCWJGqUru30behQDmmZGiBWDkFz6o08QnL4Xu5ox5OC1
2Ury/0Zgx1QkfCPKeFUbX8LI83FKDquj5NFtSw7J4BePMZcstKJo+0pYWL4BV61whkpxHG0rHpzH
mkdNJ/P5rip0Id4JKnKlaKt77iGmuC/1RHA56qELNeGtPnFeLQdiLaPIdNLjDIUjYXNeyTBaZ1F4
eFkzLKRbI9N9wMlMdMmjG+PNRZ9CMp1Tp6DCX/W69zoDnxELXN91TJ3y5PZymUj6CeND1Onhu2fv
W8XH64mC6Gsaa70b0Hxqrl2AvTdz7zt6kEg1XRtIT0x6ZbtlQlFHF7p+mdj9PG6uBXZwDukAm4qX
tm/iEyUiMAryZxujurRr9QtrXi4dSFLwzXEGptG0HUz78BU8iLOOA2k1kYcc4bRfmrG4XAehNbuP
oNsnlqAOkmbYHWyTP7no7HFlMLu7OVR9y7qyJkxCJC5rGfktII/UaR+jtpErdz+FoactG22x70Gz
FZL1cVeViPWgLJjRoapuv/pTJBvdzCyw2PIdWbcBOgc8LxEiBBdo5KEmg82YDIjWL1bXkHrYvo1t
9Jz5Y62TckH4ZRzX7mkebizK6a4oEQO65k8jmAN9pWaEH8ppy+PDHoXSuFzwO/ALlV8CuSxwM0Z2
3KqU4u63DGcTZwQInSmMsxXfETNmK5lgkxlUQ7fFZMThlN1gE6Vl5RyOi/j8nuZnPAsI77Q0vikI
22JHsJXmBdCcBChrH/KZmZiRtW0me7kc7AFftaP8r1CK3jVP2V6WvHcNfygCevrI9Evv8D9PhfID
U6WEpErUaijNAexOkhAzURitviANoi/+i36ux1bJzltv9v/X28Oq0Uc/kabipI3whWliJ+iooOzO
owwoOIwaSPEQQeg8wtZOLlV1Y7+ZnFzrtdq50GGHEimCkNix9TNTinVM5sYrQFHDWZsqORWAEtkQ
+cA/pWyNIXR/FwDnrLatgqXyP3/LV/g6XiFtP0WbBj/pPY1ivRVzSV/5wbpGT0B4xxuJU7i3wnEU
M9/o6v0oAFcKhiWb3NmB1SRgMAWs7RFAS0bpxlIqfSSSvlDCBSWVqBQF2BhNvRbD+uqO2j0+FfGV
SRw14APyifm0PTOgBtd1Ge7XvsRzKEagD5yEztx7Jod24iZ+q3hf8tkJy1f7SVqAK3iTtOzyJPTR
oIAnFJW9NoQPhLOoRZtHASihrXyuNd9/tfg7T7Hn+aCZyAR0H53jYKGGB1uvnm3EwwLkTgnT3qVs
9Fb9So4bZCCuMh/lc+OnLEN/LR3EDTSWnoINktMDpXA0zOoSyNSTFlzlh6hsszP0nvTIlho/WNhc
N0k5vg5gb0tIqdqJDFa+qDNabOcEWbcpevzyZPwS945c1IH8atW++pGY0mqefyw6dOOs1dfKNSJM
nWh3p4/9Wt3FtG/5zM4W3jqymWRiAh/+uX64x5b+iTUv+6k7jtzkVUADIgdt1M07fMuV39XuMaIX
EH+ZfPgzqLZennhdpIghDtufkApRvF6kh7PUVfdXS3we4vYsDKqZ1Xb3si5eImYjUCdfQ/MDVIQ1
ri5dOhoXS1w92giy+veC+N+YA5bG3ggL92f8mPz+AUKPQsISki1F+2bcxlcBueWo+n52+SbuZSZc
C31JJSohJMAR8KbX80AIEs16RqYNOGFh5fTiA8CF01pbeIoUjJocjLClsu4CeCmBo6fNrUQo/2iH
Juxtp/lQtS2wzxxCYP3VUlPMHhzlGS9pL2qOKCHsO2QV6Lwx2DOHMqhhMZcgJxuStNkSw5D6vEi/
hxhgDVIqqNzcI7+zx4SrBqB2j7Fe4ijMejugFfk38FUaIvNUp0wvufO3VnBe50nj52rXjZLOozkE
+wPk9QrjG2ZKc+OLQILuI6EFw37Xkhg1hyunQmjksbQ4mj5SDcUM5E+MqyKJGYN97kWJNRUgN7q/
2MYYGjRKpmosYTfPhZ2U0uxDjcgta3rACbsRDfIXIWix5xZGIJnfjL7xemzsFV26OkB6DSwCYuNV
gKpU1FwhWH70PgjD7GugogNur9UQ3KENhE9lqrRofKNndrdPzSnagSSOWJTZZFTsIGciYY15AOG6
KzVOO2Ia0XTCH+WvVXk4ENih+2kmGEzK5x4lDzrrNIAZAvVCTWPO8B/PDqtBP/CkI//UBEUl6l1I
i+fcC8BEOElyikdBg/eRtxpzxpw4QrXIQh9+Lr0LcG8lSQzmqYMw34lbn7djdXCS8/ZYtILZOYvD
l0spXpf1dVFxEYjcMhngckCP8OX5QX66lvk/ikjB8ftioWZFHG/MZE3mezFPMe8VNKBDEHiIK+T9
dkq/eHEEzyWj6ntqkFoSnT9MamcgIdqqKg3KaPp+PNypsX0MduQkmuty43ZD56LHxYgA7+4XbQwv
Q5vCu+WWN1PhVTHdRrUZsOBNmNPbgE5UIESbFS9c64usjcSdfH77Wvx5wOrZwZ20ZZnBEUWC3XJs
QSdnb+l90onvM6vx7ywAGsEuR9sqblDwrD7N5u1C2KkMa7iN7DpB2dxs1CnikXm3xR6FmdMyRoZA
8VKqiXhP5zbZyoGbcZOryn3QDBb+xn5n1WfOKNbd8NCY08oHn9dkm9gkd82zXO93mus8aWwX096y
NBpemZhmuEvF8euWVRyrKyo5gVg80XrkFq9NO1fgx3jRM68vK6M+NyYHd+Vd4wWNXZp9R2BoFK5D
b4cXI+d9rbGe1BF3XwZf4zGJiXNFLvpwMuRFAbo0YFOL5g7K5csccRT5buKJOZF5OXpH/bSwNZA7
mYnNu7PBCKZLTwgEIDnpRNRK0p9EL6BQD647Lhq/N/Ck15KExwFX7NtPCvjS0rrcSoNYKif62HYU
Te98nmw3szMVqDrLlLc3ogtPAR58FjTXauUALr+3FggNcsF2P6E4XjSh1imw5Pt1ilZDkwx7HOOO
q4GkkmFLaJb9QRilGAnF4eVLGOiV/vlSJuIuLYOdgspRftQNfGh7QFgyrUDEc9CN/LxhT5XeR83u
+ly8pq+KIvwipy+NJn42q5uV19D2l6kzGNtJ479YJMI3CHu2Z5rSPi+Y51KMkq5pJjAIIbTLljcf
BEECpkIv+a9G04XM3XdSShVAAimprU/mrup0lY5Ie0QuLPYALzLWy0wN+LiNKVcBR3ogwH2rvBbT
Zc2Ue4mFSkDqsokXoya5te1g/lZx/6qfX80tPb2jgY0Xep+uPwfa5cVKiMQE4nwI2Z0cdnSoMAkf
D2Gpa0paxwsZ3ePKRM5VPz+vYUa5NY7PKZQJUN1edpDHohESl6MOVFy/i7ldd1Gdr+vrX3Q+XGSS
AsPZoJUmz7bu+S0POUMMuFG/KRjIlNXtr3v21jWWmvtuVmExcAcgccJNT8RRGobax93h2XFE9CSV
PMauIWeC7C7x/IVvDj6ouenCWB+fmmO3WhU2TqQpTecZJr+QqX95ONPZVfMw2VDxqWKMEZQN2qE6
gPIaM0nQyDO88Qo0858nhtrABNOGacEryNNGvne/PY29r+R4wBH8MaIU+tkU0tCxCt7ihKeLKIGK
1r+XPEmgcb/0ChfpN/jXbdnLE3mWWaQkMTHXv9nsivpjRCx5sfuZQ3K0mdV7Sx5F8BnDSm1H8WyS
7xNvV6Z1FbD3yk8nZGeoYAMIchT9A7bqe79u87el+9gWgQ/bCxoIY82NgcVt83UTqd8gNenu+FRC
uW9weeKY2FQd5uVGWPdgXS+QW50q0byEbGvyZyvSjarqDkCMVB6yoj0DKljuiE55anTs+M3FglCo
TQy7+XR7p5f8cgj4I5Exj2ixoDlODcfrL1E8CN7tNPV6GiPdfTxsS0xsATp0J2B+CLpBAUssqmId
iynlfcN+QA8ZXW74P8FBF8D6gjCbCGMCEYfdl4nFxT+Plkr9AFLo8w4AO9/N0r4parDXbRdU4qXy
y15JjFcy4Xcwz/vnDB6aFl9tieYviNl3s/CHXAyEYJi14gl4JHTfCXWVM4oL70qiHTweaS/ZiYPk
RnCzs4SZrJWbXLp32oNMD5AkIB1RxjJCfzQZU/gasGQ14GbFcyGsqj1C03scwFALnIq+3YigzHAH
RbcGg4PzmRHIel0LcA0i0xZSeWSergr6oPLq1WXyRRnj+phvkGBkhXel343oPm0qyaWyC/iLq6Fg
/iL1cYRMYuCmCxnOrbKveJTHMNXWVERS+dKfmRXhEuHwdxEDa6zRqjLBtZjLBnnJNfoU7JEsnqSj
vm+KojSUdOH1hNH/gppEh3Rl9Sf8RYH6DcMe5l17lIjbt50UKw26N3tbVpo33JJ+oVHBKpuWLVsL
yD7GWQY0+WyLN16mnFhnGjRqBJFasFLe5cysdoRhljZ/hwRTEWlpMgQgELaBVmIjBymc/mmK94Jt
iURLGh3TvGwgu7LhACemanFTxa7MtKuPUJHNy88yZoaSvoidTSt+1NO70y9M5kEdk/K0+2gHOH9f
tU7yMoxbDIMpcsFC+sqZcrHLbOp4USw+vMKJQPjAgbe12J3acJUi2SBoXgTqsNgqm+aGG0EbbbKx
zYcL60xWk8N83/WrQOSdkmEKq85WaLc4+HIetcJajTu177bye6vocPSep3AiZK0NdhfUVeeB9P/d
qCyHuQT29rhT0f+cM/O7tUs5zGIyK4q+OA1zgtitYWR5jnvbFpVtqicJkIlhBK6jfIiVH7jB9t3Q
8MpmOO3IivVRFSVyFp51AO+nDM3BYzIk/XPBjb/46QryfL6vF+0yY1qwVkmxe+FYN+nUZKtTALFN
xoqw9r+9+ONyqdUzH5AiaaUJXsCDk5Dx5EWXCv8pIE89kTX/E3i00b9ZTa3vBOut4QFb+15bcOgc
rUwMJm8D74jkfQ+Ir6O8zHwcxLAG/L1oDyRcVHRTHKpESh7zDayrAwwDdwOt0eHpwGUgFHpuAi3/
5WDzdEHjVDGKKMLXwh4fX4dLCYY4MJKOU7/iT3hxP9F3bghe4HTw7PjGqYS60b1BiNOn+Rat76yS
nDLUaJ71SjJjUibOaJ8mJJ1BV9VjlZUd/ubLU5yH8F9kUCQRBrVHlDzoMRQ+qKFQvp4Jq+3J8N97
SD5USI7ia7q1tTR8VEDLIEI9dwTaEy4q+4N1eczQQaPBCeQxojFf2TY/CSYF0jOSry8rR46iSjvE
JUFzf9YjCdYHvxGLPONIwEVaTyX3ayq4AqN0b/ve7b2hIhpzg/GsRrJl8z+3ETQnkxUCni7QwHvF
6q6cq3BtRccD1pMmPmUXkaK/cHp+TLU/y6ChvtxCmC7rL40lgjITkBOJRrrhAF3OyoQFz21mINcn
H51eoZKycgNA4AYhz9Esc1JxLzKhE03me4CueQiLkKe/PCz2e3xet0+0s7Zan5xMqrIph+e0bjMA
ONh/Sf2bRXYnWA2vQN/Xpr6YtAJUqsP3Ig+DjojLyv/P82EQEl7vidOP/2jDIzvaZY0Rh4xe75ht
xEY146sDPOPv3U3lmD/MU31IH0urfu+V+cLoAj7cnee3uXc0zSSobtwdxavpvscS5HUgEBMk1d0u
H0BBQv1J6aURwRdaUXUKmhy+fsx1HoVe88ye3IxfwJgiPjTiCvQFmLxNtwn4oh5lssu5D50dczxt
KhqcYxEY199gYAg8Pyd0bBXwNPVgqAes0vqWL0LpJAN/oSg8HK2pgi8Fg14pCA1DXSrtx+ud7nru
G3j4Bd9JOdoen16Ct1va3ydDI/4IvGpuVWqKCxCkvvzoxg3flryPzp0KO2xb/caLF9yPXwcUNO1L
OrdLtVet2HskE62cI3eH9e9Hc6ki0VWZ1BszPARE0FAIIjPCBYRkdWvH3vU5+NjU40oddDAR+Osd
ZXQ/kXdUS54cIs3hmdUyYkLgXxfk4gubP8AK/H1o3eAe605mCaUJDI/OzpqxerUC/uUpY1RXYzLC
PYIXyy8RQHFAw7+5B1yAZRE+S0TodM+ou29ufecYjW91Ydli0qEp66wJGN1ltrhYouoyRClXLtwi
TA9D8rx2MVnIjamqiV42Csm7rU+aY01ZT+qWlc5UOJS0RTzY6D3zF7l265ZpEjX8ugTw3dMZpE5f
noc6fCzqpApAppsy3BpH91muvqJqICB5GvUncvAiaJtCRX6hx26STu2OTKpzHUg6/wauL+ioVdJK
CBl4bqQuIgm04M1hWQ5+8WWBIE41WVUeVVp1wefHmMHoImav5U5ethf6MVzZLq3XW+CgzIyqzObM
hOWkaXflS0Ej4EAb3uuRvATkoORWSNEvbQZlUBCJFQQsndtGCWKOGyfGQXWo10aJfPTn4XL1o9eQ
TrxPrZYoiZG1AEAP0GDfwwAv0ZWWOnlNApsXzsRgOTrqBJNA+kKstW3rrFF7Hc6chCKcV4GBnWxW
Nm3loR4Zak9dPJsjny+LMxahzK8rCbkAND9gwtcAZaoFVqNynnBPKmTmTFjODGi4Stio7iYOIAtt
RIj7055Cvybm3nHA4fqX1PZMKevKy+I/CLQGlGlbkCrviWiKNqr3Jz6QbWIMwjfrg9ComYxBSYNM
OoowzGFFlJM3x8qSvuU8KAzpwQy2fGNrc028Yp7ud+1K9ArnSFmBOiZBM0mF4R7YMPP7qmEiYbfE
6hSS8DTZUGz6Og5DZ+rrH/x3pxcbaXlotorG+Vi+kDKtZQtnIQjgPwlw4CkJucxihGdx1OcghN5e
HdsKZ2XHy4OlZhlKwZUCLNaIYFODIrX8L4JYGE+wb+NbfTtUyeuA4UAQLq8qZ7NEbm3mpk+KgLLU
xxLoa9wblOC90yU1gPHczylYKw5+Nwubidr0FtW2p9SABzDMUtUuO+Y3FvGhfpptbK0+VQHZU21d
lVNPPNYyIkl6OsdX9LTbSyjtysy75XKUK1SxUZl4YqxUNmlpynteEEqpAnl7LpswWMtwA2BRdlzm
H4AhaBA2OmlS7xbswjYR8tweQLV8jQ8ugwkfWkzBQYmpmlHa4k721xpQlkLZc2mGXLrr+K3vfj+O
pzb8Le19KOdGaPE0dYAD3W//bUXrJ7Pd9DTfTzTDxNknW6ijo7Ki88xnV77LIh1Xhn4/mVYXzqor
V9+Csn0EtgJvS7Stnp+BYPpxx5poWdg69DXB55W8Ezw6DlZZ2oB9H2L4LiUINRZdTqFGa1Lf/Smg
OuRa1ArMiwA15s0LI1doZQb6N0ZD9B2GtlvD/AjUzmsYxE4yekTL/0uZdxriSRp4Tl/8I9IwKSS7
Jd94tGJZneRHkrQryEaAVmJz2vTnS+sMrl3/DiYgexlaNudXwPTTHEu72ZvSP7yuQMLUZT88fF+W
IoycVQmlu3Izv2ByyMznof/CWqblULN0oPosCp9BZahCqUXFyn0O5yq24zOgKCoNQUxrWoSGJFM+
tYvl3OW/SW03CCHfZOBMp20GU+wl7fILYP//Nt5wP8t45tU/W6CsM8UehgMwlHrdb60+l1xJCe2v
9qAVRiWS1040n6ej9tk1ELIaGAvZ48d9OaZ5C9tNNqwDOqzrc0QA1RjYJUfzHhCdfj+1LW/M/36W
JCjnejAqc49EJFuLb2GaNXxPYIim4XjH0jicbg7KC0YoIEYqJwgUTQu1NJU+19nWP9l8Q783zwbl
C/EA+pH+e07H2N/vgUUyWIXp0sGDvVXxF/jjSgcuizpPOZDfystTZ5c3BprsHzsYih93Ads5A1SH
+DRwnFaZk4dIASdF95eXAoHSbJ8vqgrlCjfNeDr3Q+B23l44R4mVfKV2gPmCiREup8Tw2HE06odF
yeqILF3l1LfwJx0KDOR2VWTWo0KrBDnkxat1iaMp0txqwtMch41BxiC5InQNF2J0CJrmrs5Uw//6
ptMzCtZzcnTMot7geZnrYWVXA4w1Iyv6dP9Jcjsv+j5JvSDnne/Ry4YYnaMbQChOCBAfqXMyET07
HGQ09kTGIodnAayWU+H+Di7UF0PlE2S48D7qvAFbnh2tdi+gFgpvDqCTr5RQkulD2vO2BnF/kWlN
gVgGhMpyWX+g5jbTXwy6HSGN76G4yT/zFulODSRVBeA/3ioAufw3gxHmLXnHolQr1xG0r/oUra+K
ZZ165++Gr0SM31QlI3r41Qva53ZyC7kUNEMvkDcHgbkIMQNPblWe4LlfaC/E65Jj0UN41lCRyyIC
7P+zNNlVw53WXlsCAR9fqgqiGjYDhp/A15xPvcTOA1EAiiV2SRbwkZ0OiKK6I/GTG3V3PctzojpY
UrcVU4zR3WzvJewD4g/GfCdkVTZqfk2+z2HydezzDlJMiWSItClHyMok22Rl0c62nWhk9p45h6oW
GEnXCSGzqBr2l30jA8ZA2oAFQM3qM8DxxH9rfbtRZOf5egQYZGDTpU57fByWMaCdLlFtmGamrtNt
5ldCIlpiKtgGoE1TuPNqy7bH7rdlQ4qIKJzmklR3AS5OESupOSVuiJ/uiOjVEy4J7sgEkz8u6vxr
D+2Edq/ZWqtpYVNBOSkcRR5MJ3Ks97a86a8DNbJh7zZKNbvuAoK9h3bXi+73+YAsn4PEnLfU+u47
IyNrv0nE60cwlHEUjswKm7eojrV0ycNLAVTYxDhqCNQ8pCwTD7PiZuhsfuCIqFzNo9T/tPXLebqz
W+UVfD7R4f53PxZ6wRyIfmDhXFvGLcsJby/3h7XrBK/CgVoKG/atgtv1/4XFZCZ7cB2EMzU8z081
Li1Hl8NrbBeHvkDSbwQxSsor4ZdcEjb9AQEasIwDqC4UYaMlabL51RMqMIr+sgDZns4D9PqD0e35
UU7UKQU+s2lg+EVSiTAKY13Fmutj9CvH3G0JTnxZWmGjTleKNIAUfXYagUxAcrOJly6SeCM5Rv5K
SJa4AeiSDOIYCq4ZGTXMrZlhwX73aKZgyUUeo/lODVHGTn5X+aPo4MtiL0JcDSfkjOZSQqjpXyaz
sz40hmWAOO3mpAoych41+pYBgmeslQFkaVNHOZeS+zldu+5LYb+nEWsMnUdZu4bUebY6MDbDPyml
jaQPkAdDQ/ujMVvgQjun72Vx29dsb44aSF1snxYFnw882NxhKGqRX0VTu3QcLYfYmFcmTH6id2Gb
pMXy3H3qPQKOY0z9fZQGmXycpj1C0JI8NX1t7DeYcvOYLDyrIfT187ZsGkezV6T2Q3jtTjTYtlVS
Tt2UPf7STsIc8OzLb4szLKNr8oteqPoddMLaBlO6+K+7fa5sDFy1wCfhFs78KgHdCkcb5VkumyhD
Uk1yyaYrUCc0zQq8xMqZl46+LCWdcwk9yQRITFTBxI0LKgx9QKReE6v3Y/TJsRPuKzk9rYy3Mmno
AF2s1O8egL7CBuUEjgrikUrz6tQPC/x2Wj4qmsvCALQGCA82Ql0q4ViLEA3m3t6RBf92VsT2pzWm
FA8l1Juo5oAy7OZZV7eQYxos3VtU8Iau8oXQ1T+IcQoQVpfyancouDD4dQLUxotjdrZJv0GPETJZ
RpKGSRKiX/unz1O/Gxtc9W9P/jIgi5zI8P5+5WWgt5mTi1obIYAyHA0D+G3yzLHYqN0LhszQmQnT
rNIFIzPg+xUjTPqHMLbCRpbW1hdwVpyGcUexA55aKcq56dM4nZtOeDWNSNMH/2d+FNkc0duOJEG9
nyQ88RWgwYtS/+4qDvHB73ewb3pWgv5Hzgmu/zS1LYz/UR8NyWvOCeiluAL7N6eLYS80ToJR4u1K
JiPNsHgPXlqLTRDcaGbg/Xq5p5DXAXsvf2cG8SVeX7MT4p8Rhe3rdXbGh5Ko2v2OCEHXEWLxOkj6
mfsb13yk11UZ9AtMaS4y5tbgSTaRGqBDdeTPqqS6C9qNxsfYV2EvQn5WctMWW70xJS3XaMovDT0D
iJcrcWnlJu4Eraaley4niaFViCLTi5WgOvM/BWsqSRbjGdB5L8QBEdNdTqCQrrBUZqiSUFsg0m8Z
uisr5pZvm9Zumgo2u/Tdq2ehwFGTrPcEzuiTsBkwwnpdjPsDbgZ9w/zDb6iemYFpy8s/HphdYKaJ
v+XatE19ttyEzoYEyrsjTk8A4QJYx7lqOYnJJBiJ+T+3t5jo+VaBE7aJ/sG0ucTvHDINviHD0H2y
5CklyVALNtDEyHdpfoZ/CnY7Ps8MW1xyvPBO4yWX9vc/GvQPTqq+WGEBcg04nNHYTix+bJ5uw5VE
Z0YiPzwGpDQpagmXRZLfmYu3WLgaQ7rgHTlsTwZowOWAXKac5FY94n9Zv5mcboNyThEAl0ivZm4+
er8zZAE2NjIk1HG0PnTn6Grx3yHvoI9lTm5C17NGBdTLFCZwFAf21hgGDwzfNS/G+kPqhg9SCIh9
EuK1CCSyn6fbgUKcP9ewf1UBO2Cy/3T8/E9XR+6iCcE4xVr+aDan0RKXAm/MP+ZxJfhFsvTV02EM
xpzg+5acXTh11bZpYS8YjXic0BYX3ljK3na/iRiyKSufKSR+NKu4ADKqCjknVt7WR9qGa6iDiqBa
04gdY4t3cve8CU+lwqdAa0c8GztWu9dVZXSax9CwZy2uiIFaTcct/TyxvMsTS51niGsgQpCO5csS
sDazTGXQTVZgq9PX07GaiH8d0whfpdQJoF0cHYHo8mLXJpaVsJ3NHMoK3nVAsF1Dp6w/a8wZy86L
ra3q/VvGFtVZbCFWhD2esXCGBLLoOJU4Kdlkodb8+GCTH/P4lk/Cv+eEwVlw4e9iIsciqG7O81Wl
lmp5jonHD3MGz4W72LTasbYO/oPmMIXFJiiVGtAzU4gp7glKl+LwCzPFbO+UAegM2Tv8bAUTBy0M
zuvbcJZtCsNrc+dQYIzHk3qy+rVL3+fcpWrlsak/frib9vfHZxEvtX6Iy5zJSrZ66y3b8gh3ZA+E
Tt9+6yJdjqNmQLJzLtn7dxZ5mX1Ds+a+RvAJRR8C89tErWb+6j/cfX0p8A96PbW4SD1iu7bA4U8J
vjrwZ//DVJqJc1BVwenqW5a/lc+eRjXro9P4RDkv1SlsZJegmiHvdUlh2ztE3ZeG8FhmIzoIUTMs
mxA+pYNQjOGF5cCxXOId1oPW0sj1qEgUKkJD5qo0eKbhry29fAMF9ROmakPMUH9VUMSwcIFjeG9Y
EmavtKlWmZJzgysgTHTm+TW1I79x0VGN6RCV5gA3AR18Q+5UMbV5oryDhQ8zPwEYQxk6gWJnGGbW
5LQHoxPZPspIxuRyyOrzpNWgyjuOS5j5SLbX4sMzkBoUVjXm2DlzbM3qyLj0chuAX5EdWNPemfKs
NH3Q1x3L8Om27NfDj7l2I5Jo4gcqt0I1jdAqtymLJ2q/1lrStgSDTmKXqbpcqsv18d7uliaBUcGG
C1K7Hd11xCsfekDVSWGP2+U+FvUodg38JKmMdXf0/JJaWD8fiVUSo4k1oSvFQp31bDfzEZ6mWMru
Ge/x59t9RoLOOzqX1nXQPRwZwQ7qRds01FOssNV1fdGDTZJyAe9mVPjCX4tWIqmy7g1eE7fTPC2X
nNeG4qGvSCBb+GoG2VFnBmxI/dCFv/G65AgYyE6rs0WorCSrL/XbYpWaHDjqbSR0MotA/rty9nuk
7bN5g1oMSG4lLqQUYARb8O/XuwLis2Uj7bUxxEbGsPy8ts/Nz9GoTJGE/t1IQiFbcZGIoVvuijnb
CK/4ZG+lM1Tmt/But55neoJaBOUl2ew/dhjjN0b0cXG4nfu4r/aDdl52jLYsmQrWp0a79htzen5e
7V5qGeHAfwbmrkOJ2yYgt1UNPfd7NVaLLMT5HzRuQPVc+2PlIVcNh6F4MG3w18cIVDGjcZLM0XkU
eG+9ZuVmgLAIsR1ElFpfYAYQrdY3KalUTHl/25Mw1OXKhG8ch27S59A/CA0+QNtrQnj8swBOmO0W
joC4xdmvN7j4PYmQ6mer4RAYkS26M5mnJsRS/ucOVk/EP7NXjcOzBdYJqzShrmOoX8aMM1z5bhCf
0X7S5CnpiQaTLk3lYJq3rxrhAmwyu89fikJqkF0WQwA71YSc7yWYzYTcnbB1MhAKeaEmBIWCiKAX
QTAgaTLz1nxYQC8nYyJZhy5mIqrF93dzV5fJtxOSF5/33CIDUPlLnRkC45Rc4wsLq/m18fPU+piS
Y9u7YeDKuLNvp3A3nSnT+orThA2y71h+PqueVZUO29sOeJXdUZKDcBImqjZsor5ymML9+B63J/pU
qZ8Ll9K4BMsmIGqhgjWkp2EP0js0+2Ox1O0z9W4qqa5XVfDzsHUCnusk9ZLi0/ZItNCFBBl1umW4
k+gZYPqCWUgbnO2ypD7gxMfs/Ba/MRp/kmgKQWMGO2PLXG8PG7Q2q6bUWHdT5bz63OWvUVvscUEj
IpdNAxjYg2LVgAuqXWzZTu25Hb6tCbl6pyNk2+n3bob6UGctCnfE53Z9JGGhlGRI5xFTFOoV+7QW
rD/gW1itEJicRxgg2jUPPrBrQih1yFXUEumIjaor08HTrH5OtGtlQroTQ1dzko/5imob5y+nx7Ha
0JstdNbOFDZbIQndLnU7ymBEQXvUJUG7cQaRgMAsTvXERslqifrbjWztEoLctILH5EC9RLpsMG/S
HzyajRr54QKs9nxsn1OO0EsDQOON+QE2hJDcC9pk3NcbYMhRlTCyBtnSGRdbT6jOaUbfKmc+0BB/
1NoMVm0B62MEbiMruu990oyHUPcnp2zZqg2f/to1uSijtM05myMtIDJPMSiew1slBFg4hKEqWfIB
B733xaXFCJq2pyUvQooRCOG0C86GBQqirAgPgOqw7YAu7XPltKlu053D9tSZsCHL0S5HUR5dkOF3
HSICa47O4HiXeR8C6l28XDM2oKnCJ8eZ7BDl/bPCV3xpJRaqOT5iuxEI0unBtyECiBwEFJCcKJ0p
gt+7BGVTUdHOdIIc8iUdk7re1B7inqVKu6121r1WMc25bh84CrDlIcOfBvNcIecJx87dZI43WYYw
PT2FrGO5b8vC3hPRWoZ+O5yG/kCkBrMwnt9KnwOOSNuH5/+eJn5DkfqXJrs1PIaCf9Kl8ZHcmzfz
i/IphUlOAEgaPzn9km/nYkWgOPRQveIDzq2Zq+WCDIMnG4JnhN3m7iU1nzvdVdVnyfjTPmAf+vYj
Yl5yFQQ3U05wvRRvPGfLHUVCzHYwFFVu4rJEA6+iOpuQzVjFdh+JKjFZtERJQ1jPq69LuqhjARdP
YIk0GQAl9m1FRNi0TuWjNf8EX2O/hfatHm+G96Zkw2QlkACjTI6DVlpfcfipXmRPOeOJyYro2DNk
WyQiCPNP89B4U+nFc9rloaqsKE9TeashOvqfnmzlztV5M0MNQdSZdHF3J/Ozm2uE7MrSWu2GGYiD
KxXvpJdYVSy++7i7Q6Y85JocvqMlOGMcCRyGDhAFBlCIgTuma/0l2rne0anMCRzN9gE2ViX4XVjN
VzWEsR18RkQPXpRP8GY6NvTRblSb9vh8ngkC1S261HFofwbatlTvBLRs1laK4myLyhiW4UQE9Q+8
6idQscoSR8dA8nkHWK2VKykjtmNXZSBdAYa1bj+buc3t/ucTQCmMigfvzdAY5csl7Re2WPGEj7ys
e53rzVJt0pRfo3uL0fIC0h3jkrWIcKH31TXjagx9HHjHv+o1AurfySoRrb/c55BX49kqiUcGfkAq
JfajgHr+USfXYMVTM3dEcjk0M1e5CEJID7olq09SaewDrGxh/M9TTdkvGJBXkOQuBAeTo3NAZBBf
Q4WKLb2eNPt6aOhj2ZwM9kUIct/oeMj1FGFRvgUOmwdB8mmQRK+dfgi9A2OM8GGxUtX+m7rVVu1L
HgXWXczEDfTC697gRmVoEOI8X8lcUILhIra15uSkqW/reNR2aQMZdEMeAHDkC3Cmfj05of5tzPmU
ETxfpluiYZUyftO+QvsqAVcnREzumj2WxmXKLqmLsL1DeH47WJGyusCVk2YLZVzl2BKahC4eE8mp
rUvwrh12LtEyYWLOqbEqKIQRVhLXc6Mv3PFCXqBIqlkB1uN91GWIddnoc7Xg/tj/f2gsTrPJ9gcL
ysQYBOlaC4x5IJQ736YfQH/VaHkSUicQWbTCyvq2e5qrvN/JjGATg20q040WKtlbH/cp3M7IsKLt
yQY6n/6+S7wgKKivssO7Q33D/eGyhMkEUPnIMzSq4nqVUygAVMQK2oYnHFCFIhAnlIFRaELeIHka
QoqMdB6ajjDe6JVLpLkv1NyccusDzZkr5PaQe2NKjs2QA03DR76jQESz6eFicXnUDk2ALU0rt9al
b3b6M8Og05oDU2Qiv7jPxydvYgo8Fj1qi0Gvj2oCSBkUJm0Gu3hVJAcI9OqshH4eM6AqGBxbCppC
ynML0aLoPCf8PzCRFnMgdRmJ8LNcD+gsodFFiiBaSJtapkJr3030FBPK82Qnr+63J4RE7MP+HRuN
W8/6Fi3disxI9XTmfv2sy4YH8qjMI2UpsycvzNcrE6n4s4bRJ7tiNqgINhYYqnfoje2Sjp8Yyecu
VmC9Tl8+URVZU+50eSne7R3nSnRkLuRQ9ceQcHtbjq42nXAYn3WVjIWfhKs90+OQAXXlWYPo3V2O
ARBeRoH6l1sRxPetn+oDkFI41+tYh1rUIhDtwj54+bpzP7oR/M8r39d4OWFAYPhW9JUjjrFvzYSX
wyqbxQNlN4Z6hhiQVrzivCfsHubhhRKHW4hWxVreEaXZuHqnWMbA6gX56t1abYMEAznVcQsOELV+
NUsu8uvJv4v8kD8JK5HJFg/smqhk7oAIfbya2DyxmH5JZ328eIJlTj1HhApP5/okISWAYbCQo+sd
mGUN5BJvOSF5ipQWjebClIP/0h06BB+B5lrQF5NBh4/8fzxDvGPo97pEVaQSqLbc6FdHuI5M8+a1
7BpDwpWMcb9UP4BEodcqy3tJHo0q7U2YMpjEb8QBbytz08x3T0wOE4EIdeyHBScqYm8bkavQeJYE
dRw/jb+3hxT9rrTjfBzT5x6kbLYX8Nvvrf7HSoKqG13Vfw6Cadwl3EYZCIcmz23Plig5F7yQMk58
vTr1YrurQugu4+1psqgmdtHRY0zbDBB68mT3GqJ8x3kNB3hvVDXqA9nUjscKhKly7wVkm6hGuVCF
XghHXkJFvTpFxII/jnvN+53Xu0Pllqbse6iRQEc6Go6oqqEjMQfe8GyNK6xS2sAS/NzpwfssYWIO
usboRwupPHYKul4ugpVBjy6paWqf/F8wpeEhhcmOFWi4Svzj1EklqLIy34mFjz2eUk38NxJ7RTzg
NJgC2F5RzDDJoQJxa7bPPI76ucQW+kEDzVy+ZAy5YBr57gGjuKn16+b73jVS3dHwtICOEwvhJnuJ
GuMziVyAzrQd4yUoexwmxY3waD/834E204ZFZqF1VIT7MnDT+9CDxd081RWXLTwqRFiXv0MlSLkQ
RUc/GfkCCsw4Kb9+rgWknT+ug1mi+8NzsO/wXNY12nUi6r7tTT2qK38T4r72OVM6Qvn4KoEAQluE
iPg6LAdaAABmehiwzhrfun6aTgEd6P/dncP9MvIgBnh5MBzJagG5NQafseAycR+FTzVPYtH3zzU2
UvqkkzXZAiZeX8JbTxwRU89hHJfgxHGRTRuIT4a+rNkWw8i86B/UwrqNbOyrH3WIsc7vLmDfq1CH
+42v11K1P9exZBQ5jbt7V4pnwFYyC2F2IA0KN2CnaBIQJgILDpT7AiNP4BB8tTwjVCA+B0wQA9t3
oWy0IecfMupbrhzxkqZITZ/eFN65bZm06cNeMLt/miwN/BBvak1VwJG+HdX2/aZIOXRj+GcIW73z
xC4H2t3dELlLxqkxu8mxNmqEUsY+dQpL8PaQHajiPyH8fBoBca2bw84JQpLr1kd/cs3XmCmdnav+
KXwIZXGNLQj5Mu8vgtCL+UxN9Mw0haL8hrzS1iIhv96B+jJpHvyBNuoTQ4jNjDh0XPt5/RDlbiG7
Fq1rRZ3RT/F2QvI0urr2yYf/I0/7EBp8i63wsMdN5E9rfRoOBIDbpT3zSTwmVjxlwDK++8aBZnG9
iW/2/ChwYdKs+dFQb8kmf0ayZdQ3DrTE4RtYZKCA333S/2I9dcBup/F8zXvdu50WsDr2NmbgIm+b
pHJMyuhb8K683rCgOEAWTPeSd05cSLOp7it807x+aMAJsbfiIVMWJw6vbMTIi/2BMBZRvLTxtTLD
o43mxOr/3RPYlk2Aeat8rdU1rFhYFWg0wCS4dzPGPJ6Ee2ev2EX5JGi43Xz9Q4PboclnmJHhqXe8
er+GSidyNQBaWAYv9s7//MTrjCCfNZ/P7RqWnAcJJwWIZS627bNruvqXV4dPIa0yTL/loJVh3Nbi
PlbRCvZeAiW4lfrmSPZRPBImcHFyNY+Mt2bFWkOI6LOOLsz1fJtwYorff8Ap1n15Rt+pTwzM5F5G
raeoQJL6GbjItGjhDCZ/sGFhsU7qsS9xO/6+wXvl++K55KBVtQyZ391fuv+NBgyDL5cKRKBCZ5Uk
F5I99psYSqL00jIiDI8q48onBBuOj5Fsdr3E9Ad4yMvmMSCZWUyxvCTYLObPJaYilxaGG50GuyZQ
eGzDTxypuIifxMe1EWC7RPE/G/gEezU4aYRp4X+PoWwaDsfRAVtMreMbfO9x9NZ9XTv12ZwIw0/J
MVktCIDC9u28FRoI4hZQpbQLmGPtdjc7wwuzcicbtmDDePcZ+I9cZT39ANMlQeDcK0krOzkPgb70
IcCjawNYuclD1j5UDtuoNCzBH5SN4ydBuLxwwL2qAkXDX8YfTZCg54SgWTHyTkh2k5vkpHJx/xWd
F6Nso3YX5A7uqo0Rnc3aEdtb6M+UxR1kvAtOcQoA4XUfylqSfgzZNVbpbraB1jKeVkYQ7dcIU4Xd
tSZAm8hIeKHLJRJpNrdv0skC8J11q2WEpJ1Ow2Vh3Lcqlsy/aat918C1rB/tkxB10J37Xcxh4F6c
NtIWE9FHtsH1EKw/qjMt+KiUdTFl1DrzXQ7tgiGSUl2ozkCLUB3Dvnm316jkp8YPHeb/TyR5qUo4
BfWwrS5PZDlpfhyke2KolGPWmqX/yL+qhy05XWpM4BLZcrbFs9adqPXbwa0BiM31WIYgYHJD/MqC
QZBxKzPOdsB3ycCzAeceMLjhnEfFefumxPskfbnXHo4hDsprjcmIigSCKPF4etmT5V3d7ZssQRkC
QVklx/Mw+BGsaERZUQHCeJxabR9CPZcsIAoM+iWoPk6plmyWa4zsl5e6MEa8tQ3Kx4REVT8rpoU2
vOHbkZcB3IQcY09LeJRcdGlxmO1bICUrASBxsiOczj0skBQh6jPbAch1ChEmA9KqiQ6ZWoiPVMA6
hxruQ9jmzOlvWOh/aRa56TrxH11QgOncOxTi6vJ4hxZOJa+QeeqI0bsfuvScK+hLu2VxFBCFjFyH
W15cGl+qV2U19vNVcLnBZlHTb6kTi++l0Pzvk2vLJhVFbxShJWfF5RY5OukW3SOZF5SOfpuJ9YXc
CbovV07uIeBp42ZnRiSugnjyAdHX9uw2ECAS0kxOGaUofCwnM5IiEb0w29wtvbZrF0tj/Sq0VBGL
TGMzoC6196wFWD4LKtdPhzYoYhoW5iUbVWQVtUCf76LffYcCNjbeMjyDRz8IhsXw+Gl4D7GW0gxS
nnGONUInxfTIyN9dOSmS26DiAVVUPsU0D5LfB+yihh7si4/BxIGx+gg5DlDU9v+ZJlRZ9b9DnCZz
gRTbaH0Oyrk6VYhAlDhlD4qh58ZWXYtAeLsNLeNqFOpum1bxy2g5Nr4yCFN5OD4L1luwd/03sW4A
iK5sM1uZ/lV8OOUIqmSWl3iIwYwtJXL1563voRtHUsChU0IM6BIeQQ+MMTDNHSidAtvXKk9T9fKl
H5VZfKB+qBExm1iDBrknGnc6f3S1qeTXrcEUtsxoEnhGbLKm6k6UncHmKVSy8EYYZtEqOlmq1tPz
OWl43F8A6mg4twZHZ8whublcnIPf5eVSHgBf0OrsU7/4wUmcmhU9XaT8LOfyRqHteoAoOA1Bs8PL
HYJbFtx/cIzYY0Nlcc5FwOw1vRtKN7raf+sa7HXxnrMvyreJDLS5vFpKSYe9Jn7LVhLjQQubxEEm
+q9O1Dk6MplWUtX3aQTRDEqHBGOR7OM6DG+KGuTdl+j/VD4TEFE3d4QV5yBgyZdKmdanrbOi1YI9
r6Lqw4TgS9WcBZPO6YaTz+515sa/ZZ0mG1CDMMUZeeolOjsQMMOSYl3BdKD4Uc532OsetNocv9GM
26a8JQwHWgWc7CpKL/niZey/c7JkdzZzZXjk12KFEFivhAw0l5zES90C9QzGO0Xyim55uF2UMXK0
+y37aoa43kNJF2rcNyKOoDsQaJuJJzXn8+5qLywG2T2p4Wqd+rKvq9DKx+Qb7Ia6q+GMn5KzKw5s
2kaPULBgWCv5+qsd1mff6uNV8d1bawm/PNrotGA/IcJsZOVk9Y5L8JM8EBnK84LTacOMiXo1Oqqu
jNlCw156B8AtkVA+vaCS1YWRfe1p8OByuip+RurHKNRM+Ro/crNyjfdB1nmrbU0xysrYVV4meO76
8Cu16pUb3KwMwKwhhoRZWjUGjHwE4GzNG0F7MVqPC863mJdgB0RWHhpNCyPvlkfLTrWqTqYLMU3a
TyWv1dt5sgT7oxyf/tX7nKNKZqKj3kt7kyJ6hwiW77OW4lhoj9E+4C4xeCzU0OYNeav6VyHAtJkN
0cM3xiXxfusNaxRrSmSNjKq3LBGJsJB5pMM2ecBOH0aAzcvLJzH/+yg2jpcylEGAU32X8PiotFEw
TbfULdBF8qnwJQ7pSYwaEHOGyTznqysrldkHCx9vOl7XlFPsaBnvzWusMZ64J1goLoZ3qJzrcabe
pBUsuA/VuYbE95gFpTO7KcFWhDRGuHbJTSw9WLlDT2+6QW3s/uhYmQ65YUq/IPouSzWbhaVIGPcz
Mc6liWS48+Fvl6NFs0jPwjEUNjdowHHzso4NEFPd3hxLFd3twH1CxI9V+VigRAxF1sXltrzpWbff
UDWUrO3lEg1FJ0FyJpM8unCNKJSmMzBG6p/1HNWLkEkVrNWQlx7sH1iBQUSvwekumy1FtkuNX8rY
fACryrHEp23ahQMQMW+ChXOea4q5LLE/Ci10GkmdVnqlaleLZDSzpSAoaqH46+ihGgGTnAgGVhgy
9ZH+Mm3DJc5tHPcxtLlorKkNp05JRCvWRGa/yUYGSaQ3uSFV0ae/cOhftwfoRFQea2dtPBVyoN0e
NHZOoPIycooh3JZlfBoqPrLB1JIbZ/SK6tcpovXmnbQ2zSiJrZqyxQWRusx1kRdfCnuTU11t0pyk
8LCmsYeXoI3+eCb1LaxQ2hEjasEi9j/2UuOs/vluQJ2gRmvqjn1I8tyKi6MzWtA9tU2e8DDkYOVS
VOo4Q3LKEM0ccIdqLPBW6YRnObzFbpkuBW4xX1UVgtHgZZoWge+4KZugTj5kyMJN4cxe3v6duOcT
VRvCuR3gPisDS6Tr5MtinwR56AuiOUOJs1YwEpZb4midc4ZZMvt8ryb1pnU9XvVsZyaegsh2r5ta
qpSYfL4Jtdjs8yZiVUFy7v+fXrDOCKpOZVG50qDJJ+3BwG14JCea5BUkXLsWjusD8ElKBI6cR92V
bKAmmZEaceKBjzSAIRHe3k7H/i85EIq2naf5ZjoCHJ7X/7IRCTf2RnFfPNqooAwQ3j2xE/pbsCH8
q5a9Sgexv+PL9EMwI8ozhlIAq6pbYJ04jFg8q7qarp4nVoiJwJ/6pH8U3h9c/30yBREznnwAlZI7
Hip8Ldq+rrvmF8EBqnYIcoopnGYNhamaGYLMhmeMA8NdBfSEYWlSDUY9TGB04XJRF6bjaCZOjmdg
+g3p7k1oaQX0numxid8Nm6a5y4K/bjo6mWQhO2mSPqT3lcSLtL99EnOs/2EqlqFJSZZ/9LptoGfP
0nHdTq/azm7wi2pCxZBXXn+9TrK5SdUNeP38rqjP7O+jIQA32+FRXvknwWAMJyMpf0tG9CzejFl5
IvyzvDbbmpzsrl4vIl+FCqV4HrlKRs5rbpOO/BEOrE23Nr2m+wgu2Zm7bqiBDUFKpnvzUGRJjtd3
EaO5rHgkyMjwrNtgoKLX67WjcoXH55XzTkL6aDgN52tRoM97EIjvugFNeEdvxO7NC6P5e7PsGy3V
bja6YxRhr8/rmep0jXnnOpECsoLzWrot9QavxaRonRjwkx0qz2RS2Wn5S6n9ZMDD5l5GrjZaf0Zn
jCTvKmCkYK8+D99AtSE9GLOM7yS+fDHMI6pZR2eSOnINxRnvb7qvvVTSy6tULpSPYcKX74aeZXnp
1lFz8VhbrnNdF5XLvUXTT320CchfqdZlGq049Hvf/ncTgR+4FhJuxarbMHp78rQ2fuEHSmdBr0P0
vVwhJQa72c4/pBOe/lu+ExPmK5BK957Qow4bE4n3nkMP8buoe7KY7MLeN5M3BSYhamxOGOhF7HZ/
hswSLK+g4k0LJNEY6FiyoV1sGxVJlFeY7lNLPlEg/GkxHGudMZ8Ph01r6mYBhWBkLc8/KxmK2N4L
RLrqj/9Bof3LLCyxaDsTHlF292f/y8iPoUWiUlK6j69k8KIHbnPLiPrYPwDd3+RDYIZsDGmjS3d3
F2KvdQWDdXDJTta3BiT5t/ebFkZ/zUGjNTviblYtnrGxG5SnulhF+Jzsg5fEzThG+NnBvm+iNH5F
fLjMQ4/Gk/CJYwOyitP63lK6MTpEdLzanvIX0QX+jpf9ceeVLlxJnoT75VEYw/MFJQ6+lWbQ2xDV
tccWMhLQlphN0Bd62qGfnLebKHnPjBm4EAl0v9nMK0BZw24rWnGV8ZRtwH1aeihCwvETbuekS21H
35HByKVljJpsR90dXvNi/phWCKbIkKK/XgMsm8NXaDMhAnzam6GZfzhIi8/oiXj/QBlgX6VKP2bw
jm5GJi77JMTUzmzC18GJjSDGDOoDZKnMO/vxj9VyMo6WiTX5to8FjeC/asCYnfEbfj4F7Hbna7BJ
q36mMf35L8ezx8AVaY6i6mkhoAveBv5nhpMryEL660/MYNIk7/tk558ceonl80pGo8ELop17atM8
0vkTHgEP7cBU3bsQvXWpaNULvycjPu87dTQYvzP9702GUyon6WzIZTmGhhc5WnTb643GqJ7zP8fD
WPAvDbLIatpTQ2cxEsNjYmp456+bXKg01cg7FJrMPxsDVkH4h3iSu1hhr323zkNd72HdvpshciwT
37fHmFzVTmK/sac4bb7Tm2ALHMM8WJkZopk+byMRl4lLqsN/bYUjPgpYHrW6lzOhI67972xFxkbw
IlEF6GFC7WFFZMl0+nJQuD6/qqAAqQzsHZSBtC1WeGDx+A0hal/BZrn75KaHW56DYnhOlymFCUIw
eiD7YQi97JyFxQaXeSDG08njp6PBorxEF4/dLlYiU6bOssHj/cSpHzpAJBAJkknhlTRt12xIcOus
JFzdTJjgdkltyUodFPiRr8HUWAPUsaab5n378MNjMSTIN/R0jbLV/xqRG4UomfTGhn4uYQ6q+XQR
D9IzVo9aOvzNPOZGONGrXuoJgQAcxU5TG/u0CRJ/DEc8x9Nxt1QWA7hk7zkxq1VYfIXSMkwC2zaz
E74mItkNBnwYb34QOuvQ5KG0DSyUCYLViu6g/RkbMowLJEmE7E/NUJg3S/4DHgCYOJxnL+dTXDZk
MbQmLaWRdEimkZFYDXrkQbyFg6c1LnyRz53g9D/XPKc8X3Z5MxSbJh8IuohKKkny0axL1lRq8QFs
9/dRpYaGFmU1LRbEiKdiO2XQbduLbA+bDsADcnIIdU+aqwuoIwy9erthQWckSTXQPM+QbsZNKZ/m
KMeInNgzdgAxKD3Pu+K0joR0C+Eb1F1aKO5i3QJyp1BHKrXPIUPUuFySI0p6lk9w4/nKcy4c+MuV
gkv5t3fNVQIzu48NXBybg2QbgohPD2z8xypDzRc230nv1vssFOmV4WkdoJTVPT9tZkkgRrZNw7Sj
WX19SUppw3xOzLU1mABgP7GQ+j+0yZFGB/qCghWCnY3WAul9g3h8OYwJL0HMAPGaAL6c485SZ2KL
+WpYGKySTxY4azHP/kFtNjeb8CmYlf+b0poyl6VscxwTqDU8MGqhF1EaOw5yWpbMf0k9fSJxC6eh
Ffna4oz9zQfXFLcwo8XEgbvO6CP/ppOZgFKcyi1B1E2hHe/4vLQcup3B8Vmdhh5aC1SyVaYdB9XE
gM/1k7N632Hn8iKseqHiK4J3HjFJRQ2AdgHF0OUdgwsy9pZDu4vfRMM1pXezLWmqQlwYPSL50N+u
JAFbCnZetEhmqFFWBGN76XzehuS4kQd5qy2zcbuF8Gzg1c/vzmpLl37OUccHJQ0GhflOR1kLR4RY
wsjqbpzzcHXRIxpXl8vl7WEOz7rIWe74Tofh/4LTmp5WpNIZ5WNXdAZ3fuO9uXd36/WzfFye9ub9
POsuBmsgPKtFXnZuhjURRy2tlX9QzEGwfd0btD4EfFONiURbv1pUGq1rZYX3y7yfDeV8EYYf1ekp
WrfAk15cgqpWKH3wdAlUgWQus4YkSeff7BJhSCJr/izMf8ia9BHiYA+dcOMRCBoG+t8eCj2nutUo
tsR3wQ3aEXcTr8iXIxufl0OrSeZAj9L5pWzF5R8przA/GJBh5Q7CqX087ZGAxdL4kgpjmdLX0Awp
kdMD06CF5rfpPseTwJAWrCsvY5u72X/EH7cDKszTaHEJ5BKPO1Fxm6b9/COMX8nv7pUwl6oWjS1H
p4Ad2W+zpGgngduhjEjkICOYr7gpJZDSx1/blRlM0LZBDiW4ZXf+Aws8mST1rbkvay79fceyIN57
arnzqGBdgt6EWzyjCvwh2igxN47LxErhvsAUg+wZBseK4TKyo/sxKD1zXwg6hAllV6wOJhg+qpBg
jjM8O62Vkjd52uCi/SNvqL8khwpj+rhz3OoiI4soUFnudlPeR8nkw5l6thMKanePpyCFZFUetxmD
6m1USIiYxF+Fp9cmesuTO/U8YJz+s9wVaZeYeE3D/jo7Q9myeeAh5SzfI8jQFN8QnVfcC5HLTYOV
I8QxgQTQ69hiuSO5vXsQ5QdTAQrSL4XrYNQlPly1+d1SQqIW8X7IAHHuFm1oWKUYcxvzhm7QZrii
bkTV7S3mGqtZjpaG6K6C6xOyJa8uUwwks/p7iPKKutpOiC1rRYSM3qdpNtdCUB5pBIzCo+PD91zj
43s1bUyoEZ2p0YauJxxSJtvovaXszHQK62Swm+uum92NOLAecOvCwBqXhjG/Y2j8dbXtQLZuXlw2
54JoTTtggX7HVIRtThgDm3JCWU9LwqIFpYLcU+HK8SzlT5iDFbidaXJzw0Dli33JUmy0K0yBxeEq
uKWoHVBsgsO3LcRxJ849Kvu4lJZlHOdWcFZ7FRHlF/oZW8X65muxosVPjHwR2mJPh+5dWvhROXNk
cluEmUHf/RN2Q2Qpm972HNEVb5yZ58FfT19cv8/Xqw03KJyVQ3Kw96jg/wfN59+0fWyBm1oP1czD
3a13/KWAHFTUUy62v7DvDoZorpm64x8PD9Nyd+zGyYHPVGmCgsxMCedlqxl35AcHlHSLapj68dWo
IPcqpE3XMepunVWwlUY7+KC+XFwl5S6hqVVAlW2JfF6aycaIjXzDQY6c/aQAD0bavn2gLHAf/P2l
1vntdl8BKPtEVhP9xlgpUkFwid4Pk9nNgpJzWWQRmktKDeE4MBFeiTxks9o8FxW2FyVx+z7iOYEl
DyQDUPwoAfaTGeu75sLxhL8Q02p6NKd1GZLuExyXHPpmy7CRanEQnf1SGCUPyo6VvbriIuvVVkKD
AuG5YhGttoyLXtT1r7KTCbz1WrV6CUtjxIMvKMbTcG6vPtVjn+f2HkI2pd067NtINIrAvZzx1cwI
iIB3z9c69AUxQmFGDehhWW0ZSfpK6mJQ8EK1cyk7tCgOGgCNgg5Dfo0F0l/odvBwkoERcaW9UVDQ
NBpKeI8U9Vdv7cCep13feCYiLA9UUKdNakgBF0uHescMYpZHmglG54hAG0f/VMG9NIIB9Q9VVq1g
zSa5r+s+U82/ivB2cUl2uChMjjZpzsXU4Gv4+LfvSGRrWRcYsX83wk1uTYEr0cH5C9qIP4wTVuZ7
ixDwGBlQXUS8KAHTyzhtEliOiw2wz63SpPO4IAKXrWtuvwc/irFoEUvpQk5Z9FYQwOnrWQ/hMKbJ
86KWtSnznxB+vm832KKSJXy5gfwW8UwR38oP6/5LKlH6DX7KIiGlLJyZYgeljUnanbTbqO5EJ4Zz
Tm8mDwClFRdhLl4zY0/KYHEayF7shDZ1hBlqfk3FUd5XyHOJS4VSew18swV6ISBonWP6hrw7wo1x
SSTQtB27YP91lip5vwLc7N3SObXO3gmGKtk+C1KAQ5A+7XQQiT1prlguxKgPKGZQfdBzDywhV8R7
nZSDdfqYVeMsiugPVbRx29euxZwgbJP7NCda6Xm5I1mWnRAcCUIvczCJ5Pg8bZOS7SlxWiYhyPyI
idzooGch5ggTZBsVbDOxRdJZ2ADQir1YQ2WTGfrwFArkMtiGgdJTBDIK9zO4N4w746iaRgl4vooq
hFLiLyb3AdLAzF/yf3oLvFkMYSZGS9AsIYrI2jWh58CnMn0Vi+O5wna1uaLCfQAsJE4g4G2oboN1
nxk4OK1XvYVrc+WooRbT2uKWnXomFL7VY1iXbLSrmtdWxGMTVSdOwK0pzrzAk82/EUQB7KBhOnVr
fQFh3eZie+6rwOrk1VobV4gZ4jogwGHtrUZKAzuLRYPb5fF6BUU5xN9PBDe65Ch3UCwphh4iOXnG
dVfkoQobXRud3nOmXbh0NoxjRCO+nHLrgAjHjGf30EK3x7XqTboB6ijo1lxKFsB9qFyXPDGzlsGn
85G2WEqX6U9UjaF2OhHECLmYE4PmNzTODvL0MY98qRxbWAwp9tj60dcfp8MKfLEb94rMOjogwFSh
32WwibMSoB7RQ9CMihmnQLBcXMJYvHoVCQJUgp0ZzFn5hyDcTODomlT+2D1fspe4/rYew72jfQhx
FsASt09gfy3BjSniFGsmRU5AZyGmBEU7usSHAnM6I71951JU/gIOaBmb0QOp+7BX+2hFpM27hCgO
gHH8Kg2v17T2sg5l8v4qnYDMBl77y4n6UvBmx1jA2cdAtvQF/lylhK33upE/gS15yjTb7BKojdjg
2oWaQ+qcTsnKG66QCUnPbKDdx5IwbomMdPOJftPxxZzbR6hz/c1lUaukCur3guAyy3ii0zgohknT
Rt3tNGLH1v8OYjOJbmENuhnybXajQYmJx4P98As0CDQdah2jbntCSxQDeW3CqG18Y+TBIQdlMoqY
CZuTZLzwsZevbKft92VsQB3tiRifF4d1aQNUibZ6kTEw3SLXSf4qf3W+W8r6Rc6NjrPIVTL874QV
I4JLPXEb/8/vJBfGpcPIZ9pVjNOtyYCck6TToyN/2vk0seeD6NaQhwf4OHwEokFRyadm23MINFF4
RIYmxCCQPzrE9vTCJkDWnb/IORnIzWFoEKT1RO4sWRdhVf0MlN3NRYexQbIV+qV+olNSB85q9WcB
ZJ8f95yXmtHK0DWKKZGEYkoxJmBSNCkWb0Q4yPHEFb9yU5Iat+7/QWnVsMSLqT3+qZStB86GBcSa
TqDLxMq4Gw9gSdVJAwqoT1tlHcGrUDssjQUFGSKUYky6ERnXbzaYTHhpVgLNVh5/Qd3F6Ai2WY/Q
NBYNtSVSo7pN7MVlaIadVrONPz+2p5hZ0xOgKS/FeRMDSjuis0n1Y7SjMz15FJAuObpv3DsMVA77
bgfL5hssiH7PwAvjoOcgaMwsX6fGCiJYtli7SjWHv3iLxkZ/5HqI6zd5gxxSol+N7RY24wK4NhZ4
EGEnH5qVIgWGo7vPk4Mxuda1oS2s5gXxxZ8wL65KQ2hErLdHLHazZHr0//AYmKBbLi8bPzCKoAhQ
AzGqlzjxYmeb71J2tUzQmMz4XestoijF+buxvHIWg1VdHgkUnNWrFoH+6HItYmnNj92kQ6gwjvsu
gxMLXiG4B9s8xGMC8aGCqanUQR3apoLaxWB1y7/issAdwkTLrJmexE1yzgiDAMpwdMtjoZIdAziV
GmbeqrIHuLU/88a7gZgST9po15I8+DOvhZjm/pdnP8NdAd6cRjLgA7h24i297sRSplQxV3k6k0Mk
WqE+O50zF910hrsyeXpVS5N97DSI2R/uT34YuPxcMkOd2VUrXTUkri1E+dO5KAPW7gYaVmXgYQB9
dpSs4BQFZXlv5nZmzKHWBiha3UEAH+mEdQXPH9gw7gMOKfhW5th77fEVwSA48x/JWirmICb9+QIg
C+pNk+iLA1lzzhsGAdSerXhdQ92Xa1r2KqJP62Re2ZY0jMYDOhWjcfBPbGzK4lXpp8JOzsmYZvts
Zgz5Q2nN6LqJN28Nw66s22mvKqj1s4AxMPIq65Wv99LDC4DjFz56OklEIGMqGBsJzi2njqWMVajP
Z9h+F4lhOFKb5C3oAa0pulB9hWPSHXDj9JPeLktcQTdsZIS2fk1XXKjamXyC8FDzPhJUW+u9pLwg
jIpCMCngK+HGA9h+fNgal87or6Dfk+AvDpK/vkVyuvTGaaOzWzq+qFNahFwPsPewE3XGVEusZyiy
D5ZHUv2uQbHSKK5ZcveNwRra9EpkYZlkMq1XTgEEr362ESJ5hGRbW718uree/wKfxQc+VIDTJJMw
yTiIjL8NpZEKyKdCHZ+IE4ntbCe9Q8BdVE5geWYcCU7sVSH678QsmHzv9RawkFr+ieMetrIqVynz
V79OuhPaL3fmAq9Did4+7/jZY5yMzEMvecyrtdEp6KnG26MFyKCbaoNeWqKQ/T0+txDcMp0L8e/D
1bl+9niMyO3Xg1tmfmfxBKILylCdVzJG7MXdHE95j/sdJU0FQKzzknLMqakTCPk8BaOaav0Viqxm
b03jv5O8MDcKDHUwqRmjjb5UfmxGLNx9rldeuXUOapRJnCez94uC+XPDDp07wirCo/j8IvvO/xuU
UUOcPDqub7Wu3wRsQMV8Z/Wrn3+emgLABNsFfwtJll+VkTB81QfEbH6Ni7KL6xmnvRXmqPRIgnT/
Vg2FS2bChaT0szmh7djQ2ovz9zpJHJ9krtnHaQUrWtw9Zqj192TyPapKXyVllPVBE15UbMaC0fFr
npW1Q66ubCRBXRobTcEozDIQTUdzMKPL1GkHh8AslIcowVor2I1w/IiuoX/YYrylZVWAXoLATuTW
R1NNtsA5BuaRNuWES5qS5crznAXkuwR7wKS3mk9gcpHZTcbSRbtLJBYXQ988OFufe8XAskmVli5C
ZvSgJ2LBqv2vb1k+pCd3/0axjQZJq+Qax+9BO1NcLow0BOBKpiPjoIudUcIoWJ5PDJP+VNkWEBXM
nPEJ8eMMPvLMqRgTW7obb+urH/KVxAXZmyJbgaYdJ/XH7aWe8Dqtpx9I8MKG1iS4Y7tX+2gswf9k
ZJfXEnEChl7YdbKY1PqUQC3Q3MXc3yoNWHh38I1Tn1mINfTRqGk2fBRHuta0xt5zKJEPlk9HZ/2w
YysMxAfeuJhntmzbiMBtwShRJxmATvWi8ZfL2gTH5KU1Cper/cFfSFnQOxf9Q8MtLKcbXMMlXTg8
SUv3dB75S4yqCQI8k8DejrJb+EAxpUJKwGmqAswc1rsOk1ViX2Jwn2/7w9WDy7lPsPNAxVSimxYN
hIT9RlETfmFPQOru88RjM7IJiOiKPpPsYcC1i96WkwnOqVEcarW3C3LNYw0XKw6pxsb6C7t81yl7
6SSh3g+EZGws7cRG/T2hHRF4S2G6QadiVr90ZJfpJd5pnOQuKvnlnU2XqlRer3tjBepHvLSKZpwD
TWIzMAmpmZIrMMD4vgv18HoRpKmjO2CxV7t1W1pbLvo2EvCLV8tcp+5hscjGBjoL9fMg4bS/kAef
O2DBJGeKrE3Gz8YyX/lIihY879Yzksl4iAP9nfGwQL+Wn2O+ccsZHkwIZZ7CsMZxqtsOegUy3Y8j
PmMPAkFaUtiDZNqr1ZTCbyo0juuqLTd7bSUHkbuYsfRYq0eX5tD50ARuXV7nw3aPDgBTYCxcARsT
xRC8CORvc3B/mCff2ubYa0F5T8V724XlTSEjbi1TX3Wsdda2vMj6KxtpI2ahDI7uXOMhCxCDuXxN
V4LrcLECweAC6g05yxhM+IR1C5pYC614ajLA2IWhXfZyRXG4FR+E9Vrw+1w9ei1pJb8sLtSkKXRJ
sjNq7CyqmhKOECfNjWhMf0AXrjTl+n+SbSj7/c5zkDumBtwx5HhyXCINQopkMiORE38x0My9cBfd
PB+ppinVZ2ZB80RerZckc38ofYTjKbi5vxP13uXzetGVHL6Ot0THdhI5FPdKgrFq1kEN/ZaI7iLD
iicoA7+1Xnf+RQUdHLfr3cWVEGBuKfQHFICPrqoX1AWfqOTP4+rxiNZveShcoTNt4m/f4AbORm2l
hkrdlOUIFMZlx4Qxo3pxNfpLqUzk/A3WKElohKPgqTGf3MO1IbHGdNjpIHb6YZlp4LbHvr1Ko4pE
s+HcU5ABmAHPlKuTgUl+93j3w+GX9UrV/OOvwfQjQzLI8U4ZW78j8K6wghQjMhbaQcitr6WeMhkr
oy6uJwJg5PJKlwZgiAaff1FYe4UNZnXLF4NwrKjNwDhaDLqQkm0Kto85eFIFgf8CJifTH0ff2OA8
lwduSB0UEIfbe8v377Hh80KbO4Ac1e3cuZfsoXJ0YypHP1mxMxMxo5iPvM2veo/QLl6r2icJu349
Eatp1bsO2ai+Kv7R8hf7woNtenhc9rcb83Xl9c1foMaesyWtkSK9wRzkbqH7VP7RthgkvC2I51s7
fpDLcSL1bGh2Yam946nA9wgaeYTDHYQWzuygTLrPgXD+je43IWBCEsiVOPLShKAL43cseIuRRX+G
2YVuoNfbLgExOgiU0wEDdaZfw9BsTcMte9lxhc4bqyzkY7ZdxyhDm2WqNeJA5Yd2Ebh7updPYemw
XKOu+nsvy18zcTJvPFAZdjYxSnkZlErsocxk78AVeKaoo49btn/cJb4ZwcKvQrlVcCUBWXnRNYMn
2s0IWACy8lTKfpPX3FSLgcKKJwLWz2rJudKyHMhH146yh5v6O3OC1JEbesiPrOKOnoLrJVpkqU7N
CpD5uunjeHMSS+uEkMjv++vAhB20rtDOPyx/qChm6+2XBoZ19LEFTS5kDxAGnSCq4B6o40pK8pGF
+AGUR8hLsR02tmPE5VUQwyddNnqtGu/TAqaIyqd8ipFYDsrJv7j5QkWxzmxlTV1CYl/eZ6gXg7UA
Ndc71mImiRmwxSAs2aRkZExXH+Ks1HaprKA93zId4vYcVY2ZDvjO04nf0s1EbI4VbavXeUgjbb2n
U/lS4EKAWY1eogPOnfLr1+lW8SEslMvmDqpscKMnO+ZiIpXhVfVRBvjDNwdUZytZk5SMWI51u+W5
FavwTBLp5fqbseXlb5rrZ+M+tKiqBj3raqqTMF+ptQC58+V/9Xo1TqfRii+svUWBjpYUQUpwWqNY
9aCiPr4reNFHWDUdYGZa8iEMG8KvMQyNYOwAjyRK0vX23tw1NbgZCckGIavLNYVy8QyggM0J6SDx
InSy8Prv7mFg733gXR2RgwAdX9YFrJ0DmUECYvlq2GhH6XdR/WQ9IAgthwFpvUzTWTzR/1rbuCk3
vPvxo37UlUZyM899CxH3RcJMvDihlTkTH++sJ7XAZ77UBllnNgkkUy58ZzwJnr3Cxq7XqfKrtcXG
fGcCHXPiWVXIqhiaR0reww4qMYV1G4nHInm8bO13QBOE/ilcgAmyprHsxSEVp1fdvp13OQRYLCFc
tlD4GYjwnq3vlVVY47OVwmGI67SrHULkcM1dfz/FiJ/D0K/BZfPMykHnME3THvz+3T97Ev3mXJeZ
w+EYxAyIzF5GCdDdopv59H0aNyPkQl0tEpXJHFSLeZkjcEdhz+RnkD6abintRwqlTqB7sFAp0gEe
yQp/671bG6KhmiEGzL6ptZ0zmwBSp4LClSy1HpdaqbPBwe04aC/o0F8Ambya2uVGryLzMO/+di8w
GqEhM7iuvrPgAYNL73mKhEEUlVg26qw/8+aKMQ7hrhqembJqwh1Gctw/j6g1s1622MxAIEX+4uXw
92d7HTrpKyM+4qBpk+0kAzvkcNxuSbxSH3upYG9nVIXEsK/UwCpclsn2brNZ0eF0ijvfcE0ncfV3
I0DL1K0Sp/aIWqfE6dlh4NewqwkfeCr3OY1n7CedjA1GBy7weEYT/L7redsOzu6MFZRmFfcA+Lth
6Hr/EVvSNH9F/qlgkSvvOdbDlvt2t4xZLanzWC06VELCjhx3Jz+B9ikUrcPWprMs8hizJ/v2dWpU
Yx0/ze8ns6VtQNA75bAObk4ajATFn2b+s4azE3gmTkf8QnMJGjDgDqaBU1rRbUGHYW/Q9gkQyk6S
rgUm+uksydI+6Cawftcr8tU8FzbEz6gpch1Fl4llKST82S7sdYGqlA4kgK+LvI3rRjBAMBG9lStw
HoDtOoIm7e/BvhSNtRDGpVhdpj+rvHt6x7RGjCNLZzohYGW6MbjbUJpyVQ8Z6yAX8SM+K8fVTzhF
VxKOAD/eLUn/RGi3Y915s8tU3yY9UyuPWKOGDIS49G8bCl8Fdwutwzd5kMlzTIV9/PfGPK6xhqUd
f+HWJEIvUi6iAc8KhGodsY4yfvLWlyMDKxSNqOvlqZAWUcAoP49tH5wCVf0JOG/cpgyZmdhG50am
QutiVPwrUhv7a+rwbuc0IRBvpw5i4E9MEhN5xZaZ6Tw9aR/a37O9u/3mRK6lSb8ZTO8IZc/wp/Vf
6Owc3LqRdyFOdmNiEHPbIYF48/Xx99rAfdR974mdS/JlYKgHudYY/dtl3ssCRFOCkqHAHXyJv+Uv
4i7yet1B8ib0xIJVT2xvII48tJbNDUOlP2qVEYErH69u/GpJltAQyZIBvpZTTpNztzicZj0K0VKb
RXVZD0VtJLQJIF1ZI6FOkZ0iLWtrUP0PDaW7Roh3PnNUelOrNXB1yYDgnlknbdmjxS9pzNX/HU/f
nm+8smS9BS5M/b/6GqmdDoKAkXoaNlqR10+lUz7Vqfs8X/73kUgbK6usQ4/4CjCO21Tm7M+I00FW
qbhiZk2LYC1bU3uBf70kgqPsaAUt8V4XLSga00t+WqHVFLyWOXhYLSygEs+fDC3Nf2Fytxgd2ap7
oVxy4RQk+W3y5lnPfGYNOl2ayLE8aZroBe4uHGaNT5L5yWbhzAEpZ3k/xqG497eLVW54MshFbtd1
83DVc+8szuon0c7CrYwz+Qm73NcRhvA2JmtTTMjESMhtK/t7QmMMDH/b8fkOc6TF8OniPoFa7DfF
fM44yBCfgmdoao3d2F2v7U2WK5tWW2DVww+V2Dp5TCMbnXqzDIJx6aaMIOYt4dr97ld4ElUvw13h
61WwTW2LraaFsrmazwNKx8Pfq1s+ZAZSyn7V6yufKZIZ45f+POHgYo5glaVxhTwdxidRcJ95a5W8
Gx/64U2mysHsAWRRROEjVh3b4AfEZ9VG3Smaaizdly6wzvUrqxybqBrphbkZiicJLRxybrnCZc3r
4Ms3mS81YTw6PvWbutYDgjjv6OKY/H4cQ9FZdfHQS9iSfLkkp1z+01+K5v4pe/sJfumK+hJx7Kxc
hkQW2NRkWOEWu8qLXLD/x1WbMd40K9RRqURiL6lmKU3c4LSoshhBZKHpp7hIspeh2u6oa/imDGbD
HnWBmF7umwZWfpPhqfhX0HYeVEfg+Na7O1cvHXZYj8bygi0LupLPIlszvNncJvlrNM1xmmhdPoY0
gpqmwJuEaIpiRAlrBRCw3b0ZIywRsqwC+/jE9KROzF9UAl/S+jj7K2rfinRxoBRn5JhCKRNhrVkD
Cuty5qrA3CTqeWoCz5b0mDOPC60+N7WLaCTtpoWv0DYRA5WFQkbXryHvZecnGetxo0xExADhX1r3
isWIMjlrE86KshkG7/Y819UPoV+Z0lNIxODQuon+tOvkL5JopdCE+MTcx5i7DLvuypKVqNGklLUO
Q4mE07v7rq4GhqVppBmRfZHeJavxDd+r3ilwzh5F
`protect end_protected
