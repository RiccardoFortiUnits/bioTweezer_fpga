`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LukpFOYmAFLq0bbk9FiPDW6kgnvtEgWDLAOys6Lxts3ODjbecRHAaGLy1LXbQvWD
awCbFizDtxMIzfZZ+j8Jai8ycfOgqdNPoqbnusYdYkVJ1pQLN60kWXjDzAgJPr7i
bE8l51BadZiRHX6/tQJ8UsRwRSoc2/fp8dDK30soJt4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35376)
cBafPvXtt9CZh7+PINyDb1aKoRDjFXrvRHSHX4pRpHgEHkBTpKm7fJtGVQiFBc7X
u5E91BGusbcAuMaVpYk7vLdPKFKfOlIffjfXOxmcrMLFSyWIBE6nB2nDTJL+AEvU
TAvgFbnJE7WhKFqMHZMBcFul4A4oLGqJurdRTiulwF3Nx5xpRC7ZN+SUqOnq+o9k
XOyWswOR/fsm+fZN6maalmZlVDh+KiuvwUMpK5/3M6am6bFOQ/ae14yLRZUo75R9
N0MgmXLTG9DIQMxvU4HX1JiOxihs4gAaYTvl0DzkK7KSE4OuCx6yNGHkg6vn+RAN
q1nTswf5h37sjxRbEIHJ6txRo7yuedGW7OY+ksIFRDINK1uagMKRa4hTnC0FzLoF
n+1bgusPWYIV039giTv+0ozMRQEXRYruTb3xBw7es8eXDYQ9Vt1xgzhEw1NPvQhq
D/2900S+LXqTUCVV78SLHv9r8rUPQ+liGrM2QCKMs/mZXILhsmRVqaNYDlFjLJwY
eaTcPBmK8ATsG5KLxAVKxs9+4+m22vZ93zKozuFzmynx8zsaFpp07/oVoDcRlKnd
X6v3bIYY3EWOE0w77OsRBlLuaJcpfsyKgOZ5uv+l1kDcYBOjEelWSUnyz/lc99wt
kf/ouWek453MrLoeXTcB04ARWsO/1mM9u594TFB7HGdEjBmlaNFYUp0D4kFPGUg1
kCFOlTAhuEAIstfS98c44jXmRusFhwcJtZutvTxhonAbGVJ8usqOhTVwLbHtnhvN
Yp7ZMK0UTnrne7+3ShtAUcRlD0YnCvcuQgWs/jxZso5GGxwfc7WirPl6EpFCbgDE
+yLrpshncCP3Ro6ItBs1lJBeS5DyIO034IxOnXRXTMFKSDaCo/XxzR0ZFreqyExl
Ditt8tX3a4z2kzFaztfPqIxuOJ1e+u8tZfiFYgD1N7YKS9yD6D141tuBYX02aqji
74AEGaPzNr2e38VasnIi+EcIkStJVP90FNjnddoXzKNpkA8loiKmjKUJyB4E6S+z
ULz8GVjWiddRgcZXYTme5R7FEhRdCTGh7zfH4k4GQf9COltoxU2hujhJwB6Q62vF
CFcrF3JAzfANBZVelm0s8DtOQoivesjqJPEXyxDx0DBF7saGY47ve7OfSjreK1cU
m2tQ96y/ZfnVQMoityiqrOyOORXFYDBqNC2L3QWyywVFzsWeHZv74CRx1qPrdwLD
z4dFE6h1yol0hjP8ZO+83gWuTsI9JysFdO5xRoZ9/EI9ny4p0+8yEv8hZoqx8R4R
dPWF/1uc0C+VM7zZ0Uy32TiKbJtslz7qhaCgBiu6Y3xg2nJI8Bi0u2VUX6c44tAR
7/D7bMwpK0NLxnNlaoYKGR80tpYoyaF1Ui8J0h48x7fz/RdwJaYY1GVV3HktkUnF
INqQO0kabo517mkQf9wrxrs2wDYqO4fnsa0wJDA6dEwDtaBbR3AVZUMGNe9yWmVB
QIQ+V/QjUREu7W0ohq/wjEQBAH19staXQ72fYMvFNwknE/Wi9OI3nED0Dxcn/WQk
CHm3M98PxqEKRwinRI1ue3Au4Ddh764vayniAu1iv6N0cbEsfsSmQnWUX/0733Ir
GFfWi6mbjB0Xn/iFH5CNVFoQfUxiMR6EU315yhxpSg2RXDskRTF5B+z1Ox7P3SzP
4BMe9Valb1ZW5qyluJ47Vfmz/EBbGKm4ROeKvy8ZdeiI6UuLy4oUAJ1baZUFoyHd
403kxMZ8uoIZ+NyA1pqRwUaSlPhZXC7ulgnL6Am9BEVTB7C3mGcTUH5TCAUOSywU
BWu2siautm+miCvt2Wdztrbj0aCA90mv0TwS8RSjF1UTvxX8OsOmKFsLKlf0Ag+Q
o/qnrZO7XBlRl8o+UHP0N+j9Ef2WICkgWJdcAXzH9slh2RgGnKf381BtHBFCN5hu
hasQF945yS/MXIUL6ErAgo9jAv+8A1eKgKwdQW57Vrb5118RqBPZXTzoRIEL0OKs
aw+DZJENKXigefVoSRpsKa+7fKYSK2lCYgPDjCS4pKMat6wJ7SuZypHUQVcC+kHu
SdGyJCi66MIPPdqgydiW/FAwlbiTiXJ6ifeKbrz84yfVdKUEi1c/SyXiLrBUhU6a
Cr7fJp0/0EsgdhbxarIP7DgWpPDHj0470TdVY9kQPzo+grg4YhobpYjuds666EyF
NCgZAmMMW4JS859vl7DUfvzqbMUZnkxNaNpL7aXttfvWnl1cgfFPiZYkMsBPlVfy
//vZj2VqoL9YBQ6lsDr3rbI8rHcqC2ll4QqixvxYHtPPJTdVy8TjLquMSgAnaycz
UEiFTcfuhX3E3cc8Uw4h8LeYe623fHKGH24uBhqOAk5k2b5XUyB8HOX9Qr8zz5Xh
Ef4gnv7yQTxcUKgGgPJp/4St0+qob/nGxTzDosvpxuMI3qv4B2Y9rLGCEyFJmvR2
vW62jX8xJAMdJysl1Xyi4X5bvl2TZI9mzoEDTywfwAwQnUc//Feq/CtVvJhphuEF
ktYYYj4XrcfaWXqSgVhBBs8QvZXuH6YnSZrobU7V/H/daj3kUk7Uf5ufjt1MC/uv
pq/cZ7G0lnyLmhoeG4vYnFslJLbU2rtYfxLzAC1nyAvDBlk08ZyFAm8nLNY7IIHv
uFte05TX3Iu0I9IhO6EW4SnnQfjzkIDAi1MIi6QnOkefA7dO59SVfC1r9pAwkIf0
VholKR4ynIu2sIzqqlUo5bxgxf2kJI9JYAJd0jluIeX39pNdX0Qcv5TTfz5xKlvU
jwUmkxP0OIUdLOx17fEhPVGtIKJWnKUYna8ezWsrGda/odJ65TNE4tefGbeZ/zWz
bnIjhxPNeRbKjgs3Ez9YoM3g2EvS+O1NKfjLh+ME5Ragh2wL9dqBMfIcEguOGirI
UZnmYIrLjeQ7mkE78+3pzoK3UNKsDKInY0obLlOvLNctcyTcYEijBkEZg16KTM+Z
DscVNJ1T5PGIHgYXfuqqP4p5iYPA8i/iKH9xmeJ/CXRNj/rb2PxT1geM0hhczUJs
ePHbJUrPng27Q2Noq37ZfbEGN9rbKZEst5Q5/6Uts1/bbGrSOZRlUDIObgIdCYMB
D0x8fw65V/q3m2r3Leaq3Lh1Ru2fxQ49o2zEg22FeksG4Js4SgMv2tDCBGyaI4v7
a47D2WM8QYLPbkqgZOF18Sg90qyY5N+hLDGnAWBDTAq3z5P2gJ8y1qCEgs093sVS
lZ/MlAvGDPb5Dcuo/mCQVeg8fSVdo+FH6lmUUChnphwHbr2pqNtg5PyzaiLFbRx7
53hxL6F7q7asUE7c7CmFnS17fZvAsPrxiOWjbz3URzDrWcHUOm+Y7ruAEMxcoBLt
fe4uWe405SAb21ilX0LQ5YZ2MJ2NdX2/oZm8Kmtv3/4xLdZaKTBFNoUhRqxgbQyF
l7m3MnxKKKF2415h22GTX1lNwO2oI2Xut+Oi6t4F+Ng1g4i/a+SMD6syXcfTUnZk
hqncDPSGYbjrP6NCDa58Ddqqqsmfmo3hPd7fNWtguDXEZwfwWf9YPVeHPkMUmlWy
cmNtLdA9+hNINwF011GgwXVEDvHcbiwQKfJMFr6wsOQ63fRxqA9EGd8BAT4iv7zc
XgA7R9g3qT0IHJtWKlR5z+CiPf4gli4gY3UrqGtazDY/z9QVZUMTF841mFNbX4pj
MKVoBEdf0E++dmY8o6pd23J5anT+I21w28m1iSEXDq8KujgWkGyorrx27jea11aY
H5ioWnHN/IohEOEm+Qb4FTxI756/3NEb57swSn1MPlN8WTEhYlTKLnwTwQkehqeG
QtqY53pWbEmfqFxA7AMu1QAz0YcVBCYRtQcLLVQufXGbuG1Dze+KXTLuFD5Fijue
qoOuQEwrinxEGPx67gufeg39LPc1T7+Iy5keXlt0s97KMcSPR366FaEmK3jLMziZ
vdqClfUkuiAROinPRLXm8ooJBxT5x+x1oiD6RTspIApQJNAfT8YaRR+KRxrvDF+s
svAuCdJFft+0M5ftgLXPNAVyC9YAq/HEjifKkvvuHGBpSgl4FERzZwHofyLfkPX9
rTAexnR3OMpq+2TnPbllBd6NXlKdKs1crXI+f+gt8IU5R3s8Q+Pvd8W5DXILv8Yv
daq/6sBREkHOfXUS/aqwq8QEndy76u8UEbRpRGNV1SNy/tyqveaTkmWEy9R23yl2
afoHuxeBICDRc3x4LEeULCj92qeAkS7hpc9DW/Xy5y9ONEP3kbsA1ecWr1+Ezk03
IvLdNsqIJFFg3v1Pw9znDBqG3ucUQy36Fy7ONdNME+Q0bZpfXxDmYrhyR6oYbGE+
SUyd7DrkJJcvqw26v20EdQLuTxnkea1ecI1bhP5rEaw9h82RtKfR9DQveSfYVD/s
wT+hSfXGK8Ww99gMtwEvuTd/sMfwZ96NCadWjH9diNBjbyHz7x6LeBN/dgLBa40A
VFFT8E0uNLdZOhOFWUZXXPRTgJHIgeBFnGGBaGXtRj9n27EoPnyK06ZZY7T4xlwz
02UuoDVGq9wAdHPv6NhTKTAFImWEhMk5fPCjnhbrWZ74UKM7/Q4DIeq9n0+ccoEb
Gb8GKMIsHvtrcZAo8vYi8538D1SExQfLsq53WcXYK6dfU4F3NN87jTnNkgRNStp+
+cUjATD2tj1f57qwZZA9bigjOaSLKZcMle+aOTbKTj1wl+SOmKv8s9VyoxYYYDq+
yXdng8cBdoekk1RQ9gc9GzWb47mAGym3RKR5YwmVLDzoiPD+NWRDbafVRL5VFtWo
47HwxRS4X2fCLoq8O9jmB/7vMLKOFlDYC9ZDcHhwr5yYapfwqsaeqNmsCKOy4/Ob
C3Ir1CTSExyD3QVxysaFZzqKXi1YJU6HB5wu29oYlfOwgpsCzCyFYnBz0hKIhYij
VkRvq3PYJgAmTARToWiaS1dxYAC7AGvIiUCQXdN9KEaEY5j1WZiWTLL9i09aPlQh
7EcJW1sZshKGM+PG9IXMaY/zHFk3bU4OE/qfIQVmnWvrK7HpvY+GIl5RrXWjIEBj
vuwTrJ0taspglKuXXb0oSsNARqIkjNq8yoAlIfLZSsOj5HZaO2hYEaEx3eAchOuH
m1/UzcuVcBX5Z7PnsRda8ESgYAxiiJET8r9vtpYRO32IgrhTgLCe3ztv0cudeXIi
fGy3GfeMJplUp41TeJMSyPGh7dNA+tPjJPzJd7uNrqG8V61bx93yDQu2hT2VWF+K
zWFPpgfl7pFSC17e2QA/aZQmarzCdPM6q7qvZum3F9qM5V8Qxn5hJIbV1RKeZuif
4dl8ftlkIEsHcSQAWzbk4oSZXCBVrZCCQTL9psmfQ5Cj8Q84ig9Z27XCpBUcaSFB
R52HwRcyO/6+HM83bqZdYf24ZEsHO8Za9wD6CDH4aZpxejIf58Hzuw0XPEsMFsFs
XUWRT/2vL3kGvdT7FJZXjjb1wh15AKhZrEWnTz4U+09Ore6Ol+zkSxnzVdDbf1JX
aPV4ZIjD4AC9IyHbYIHuG56mbCIMo0SCYDemCzesi+NaXlVnqsiullFAyTbHuvJ8
w2H5tIMPvZCwKrpvl0YGXW8s4Dx7nXZP9cVn58avrJBuhCPro53b4RmcBK4hUT4d
3mSdv25tV0CHGtdfAZ3AcBgOhp69xAn8a2p0JkKY1vnve+8kVF9tipwXREWeiWbI
Ywqkp1iX1u9yuVwvzKLKod59vCGmk9HNzuHd4sHpf9nebHYLY1TFvm8ClYOuiDvA
/+AurG/9zP81FT2WSZ/V2k8mJc+LE07W2bGi3XWC1IKz9PLnz4b1NiuWkk00vCKY
2fGRN+Ay6CbJL7MuOdp3+ziAovUqyQPSKvb97kgZAAOPiD4uK2aTpPSHC8fAZMB/
qtknspW+v7SzBaiUQFHiQrGuE1iMi3/C9I3AWygSOHp5Fq/PETADqkcfstsPLzZw
cjraGLEJcI5Q44cSmGEGJm67LxXqTTq85U+ZVsF3jGLIy65MjE7hh0OSbgW5nGnL
gHs1m/TjbOr9Dg9Jdu3qAWD2ihJZNEkwGJyDX1a19+N5U9kaJz5E/ofSEBoah7Fu
nT2kQ0R/Q+/rZyawTtZkYdJzQztdrwHdblQDk6zTyjmr9CUALbmNRUZ26hB7xMlM
Bin9AI7hdN0Dd2mIoRTu12hexqY0lgkm8diBwKTga6sIxk7msVT4vXl5q5UK1p03
I1iy3gmSnlW2l+55csxP6Yk85bJALXmVHdmgZTTScoIYJM8DrKdXjcOB/YzwT93j
CUlRcpz6FWHCS2OZ0QoXDRg0MRFDZG4+LheycgVO+6C19xMsF/46AmzkBQbS9Wvv
WBR7bnbqGeY5dpnI3aHTRVvmYhvpAHTAastkJ7ROiC0IOhK47miirwXcV6ji23u3
YmXCOrCGtbRPy0YadNVcE7UpTTglmH4NUv8Ii8QtTqnYUeolaZ/lWt+8gUWYdO/i
aYVTosdUDvqw7mIYDXumL9RqhwIymV3NO2kWZm3YR0uRglXfiTzSwGMkz3nw+ZFn
1vTqjMBikLhREHNYZLBujfx/0I1E0OMbqsFknKx/DfJKm9+dhdjlJ4T/I4oDt+J2
5dq2yjQOtIbDTMPweiMWmGwcyL48Yi9UEDOqHVC9GIg50gOp+WL3fzlOJoPqmUy9
2S4itKZsbNd+YsF5WWGRKXU+7E6otMyqtTDsamJJ+wdzKAt0CDTryuQY/MQGBE3Y
8UqxzJdZDTJ3UrNTimRFcyahSrQedRFLdE20kUKNTfinwSRg+tkaRU/e/0mWhiDj
dw26LmszKgh6ZEROZG4jsPJsH0Cbfnc+enlJwXiOHsbHfz3H+q0sAfX5rm93IyrY
pQc79UnMuzXB8SIyUyZZiEg1ZR7zulQ/lbqmDsZxh1s4v6uHYJj8tbNLsRxxiICt
YKF4U7M8ofw8CjRRjGGWzVth4Ols9ls0/Bd0Eowi8ES62IPYzeedH5GZowNRsBvz
9cMtlNv/31CLqTAgHMHa5OTX/LWYRy1BQPloOjBh7ATUmGGLuybWuvw84Uy2SRYa
s7guzgjy8u6/7sz2c+LMZu4Ngh8GSI0Zmrf8ifL7ajGic547AxGDp4B8ltXr82CE
lp4nJsKFC4CaFbgkFwLj/X+/KdKVURvuLVtNDXLI7vQ1+Vx3nOjZujA66gspPQDX
pJRlGOqfv2deD/Ps/Y9PC6fWH0u+fgkyWC93Qy+Hc9PQDbaETtsYcNB/IM1G6lj/
zgwTrP6seiNMZmF+mQwX8j3VYQQ0MfuzsZCDslqsq4gT8XVhNhIrumN+BL6ZKXrP
SKII+1V/EP1Vxnmv3c1mMPV8BCQITCdLMjZ4901eiHiYmWk3v4V/UGDlRvZbuf07
FaEIbTCh1dgRPjokd4cDh6yoRfoWiz6pskJYZpm/0XyJAUkMVsweYSncA6k9F5o2
vz/NOt0crnstsTaINIzos2I5tEzhIUmw61JvvCSMgciEjz+pwwLsk6iGOSSOQCoV
7fpQppmxMT7YAs2avIvck+ik5CdpKI3yeQX9dSMuXL6xh9IWhjR8BUhRJZNcoOYz
itAZSi66NCt6rII7zRPm6zWYJBrU4MV8/l033jC24DwGX1OqyNR7rBv0tKA2OpLf
5LqAYfE6J+ayB+NR8Ysudn+kUsd3mVK8E23BkeuHnGrLDV+xH61Kk1uZnWOiaHgL
UEQMzhpnQLXHdwNhSc7cgoV8egi0sWVnkuvs20amG0z7SEsmzJC1vdLS0HzwLf0o
yG12lJlgEC+fGM8FVr/aFZtntxniHVZ8ROHccUGcgFQZ/4fJGxW0unmT9X2f+pDp
evGAMWVVXAsk+YxOgnbRQ1YMxICFLC9nw5f9DnGJ1OAzxGTi2r+egPwRVq94SCw1
Clny3QoFOHrUdtyqwRwFpwHhkEeRZd2A14mJ2s8CuMjg2Yw03HZyg6EM62Rq+4ES
dBWgVNfTuyRcrpA+vnzvfm62FfOR/BcAWWp00gcaZRVBwRWNuRyChNDcuDBI6D7N
5+n+vUrsxpKM7NBn81Qv9SyNKaBU0xbmxBBrnUMOYEbN8Ov/NPt4uY9QCVpmQLvg
+d5+NddNSkf231YCxJvwIIXeV2Esar0jDJsxH17vRlUqVlbE6mGgK0cHnqG9bdnb
97/m2tY6BqBZWa5TQ7ld2G8ewmQI+iRAvprJPdFrO3dWgqFVulvDpTqjeOTgRoyA
784PZRoX2bW+R7SczcVKTVbhSQvuPLs9Ktm2ntlxOm73eB2m8DbGqBeI9lyIzuVV
O6UG9lu8lRqzRUBqisyjIRHBHpd5CcjHT2U2b3nQHEUE6KpCnnmBPnBDiqIw8svu
KTZKL4hUq9ZMvTb81FYGNnSiAtXFdpoRsGDjEvzZ3WBpoBjdOUVwS/XbJ2AN3OpY
nM8ebp/Uz0Ygq0eK7wBroHxJsRrx1WnrT+INQtwwrnBvtmY7TxlY7UkWlBws9+3n
20yzt/3rZT572elN2LWp7EfNz7khgXhFEOfkhT7IXTsXP0gNYYv2tjrnl7Re5aE/
+eOs5u4dn3RdbvB8H7o2TpNsPFVSUn/ehkbQ1KDxImt7gq1LVwe1LoOzkf3nIv6P
oaH/mgdgKdB9HJZ5Bnues+uJBeeDz9Wcah+SMgH+wBwJ7WbjyLbVkTz89pNSnd7n
ORGzx79INhZf48JfJ68UCI18wN8vmniuqXlv4J3EWjCnbX07xSYPW+bdp8CfzMkf
lr891fxnSbwQKvf4Jd58sT7wS8ZvoRcEwAL4vtuybsUJsDb+EoNEEtdHhzqC113M
mOPtuq54R82CGKb4om5tUWO1ChQGPxfc0lrYmEBSI5w3GHIUqA182MXvXnqlW3QI
2/07uC785EdCaXc0tLUCocAHlwr878PCF3986Pfk0Fx12cFx4mgaGV1rIf0gHJ7I
4Ba+D+LaSC2v/Tx0ZJev4m1a323CxQBhcVh+IaP5R3q4AjfXBK0ayReg41FMIYdl
fVZt0keB/3stY2wEMN/ATJa0iNxhw4Bkd2vGGh8j8MNSMf9OlTjt8mXXnreOSAJo
aomlYKJQz8Rk8FLm60Bq2OgJgVkdvsrMZsyZExhFrUv/2EY9t2hiGcnX+EWU0dMd
KjPgUSNiSAalx7OVyqgHcZnnHlPMl9KCimjTWFnVstEOF38Q3iVM+LUQCZ56Mn8d
pLNPmLGn8G41GeM/8YO+iLT4QaLZl6SycxzcQoMX1lLar/mMgmiYC1uPgAixg8Jd
A+tnDf7A4p3eG39O16IW3OTyz9y3+La67Vv3IPxtj2rzhZirht3NmPGZjDO4xV7n
kxLKYJAq9ys12j+gVasBQE3qO03BhzwakbccwTWxDHtvopa7/Gi+lML1uodICsxJ
W+WsYrUurJ3W9oE7RM5ZARGuzoYcZ86jUZL6kZSpg6g/08OLRfGhgORnchAIepfV
0n+tIMaiuFWeKVirtHo3yqJxwiAondONsZaaXoo/Tdhtk5wBpHBNi2XtEcdsNg3L
xNk/YSnlctXqfZQENF20yvAYLO7O8ki5R86TIIY+sfjK+JtgkRlv+gvzdY24k4Jc
+Dcf6xoLvnFhvjWxmKaXo2rwZEeAxzDPQYVlfEARoIm5IDUFlpF9o7w9/Wk0ReaK
syS9Quap2ARdlTcLmQ/Ic3zkWb91ykhyQDEkkhhNdKj/3O+537PDWbbGb9Xt0DiS
enIypSSR699whvNPFOMb5T902xO/m94+oG1sneZecsQAnGirXNBX6+AjDDGxP/h3
y+nmpot7ZFo3ArHWlY0B9y/fZA6TS9AO044WvVsSgyj1wMxOPEf5eTC5yw+5irvN
fQ8gduP1vofT/gsNgPOhKHGIns2VcURWBihJ24d/OZe6M2JcGGmKBVtAAJufaaeP
LsjyGl8wRFK8WTEHkjVMQDXE3VIa/VrK8z2h5G7bg23qU/H7mt6wZTPgCbNlvuuN
O80BMLtA0YQGMVTllCGrFa8jesuzkInJ/pK6QSza44+lHGr3VFHOb5eTP6zbFGLr
kjzjhLc2fM7NpI4mggbO3S4jxubA+gXE+sxYgVsV95G7dX9ubJrVgilj3rUl7uXo
h69aqB44pTJxtvc9EZejjAID+d3h2FbI6OlVaDWlQxCgKS6TUZPkXnUfjk80a4Z7
d6gIC3iVzHu8gliNdQNFsFbhN4x0YwJw9UHKM+4X7Dmh6JCILOZJXkeAiBa3xqA8
PXFfbW1DsiN+7v7JxZTExfLr/wTckNMK9LKoJ4jic5RwL8QOdpxqGUuK7f28Xubi
qbqELj1PhvbTetiWM/6pyhJD92RSPAKFv+zodxHHFtlpLpdHnugxvZUqbQFIxtvF
Sv66WBdDwE7fprq6Uoovlw8cj1g2GqvEYhg02oRIRO9ikPyOLSBIPj+yEKctskch
zHBsXy5bI2TznUCi5Bnjw0eeTh0kHWmN7QcptPpQxMS3YNDubBAzZ50F8xVEhgol
rjF9H/OWrW5bRUybB4shDVSvj6eH0WjGYxnHdJ4XRjLgmDVYV1/RpfDVbcmGhfe1
ypvx7oI2NQEja5E3wZ0xB6xoLNIFKq8CqQNRRFPlhYFiYLDrHvc2VDFjYI+dYw+a
L1rIdL4/oQAor89q7OJkifG1WE1gUFiWvX8GDZ0IwcsbsAi5uPlJAiwtBdXnAb6l
fvUPr2FTnQd3QFjdyNP3ooeUulKwSM/a6PbWWz8Cb1Am75GqAYsHpNLAAxB67NpC
H99TFs6tqyGWH425V3cIC+Q8eMULqEgydEqgus3KijPVF1dy+xFElCkqswGdLZi5
JzvzaGYduLgaG992o0tKegKe+E/Q4yil8zlqRxI9QPljFUfqm1YiA7jmTumTTDLf
x/eU5JX9lQeitSMG/R5QwQ2zg0bWohl7w6sTR1xbhrOrbG05do2wtyTKZKYBvQoL
c4PjSzh/Eb873cACB44GqJU/mDI9ZVJR7czdNgZZnoVuN9PGp3v9VawU8RTsKP39
GaRtKQVitRIRZ9M8qsFDjThXSvLaqDD/9nC3ZR2/9xCx/Sc5xIj8ALf4jAF5mY3y
0ZvfcEjjFhR4kXKLFm98qU7upYCBQ+NeVydg8YIAMXRKnbIGlnW0Qnx3DtQUj0Nn
kpJjgSPaAVWXR73ivBMfguhI0o7P+L/IiD80OIUhdpDBL7dqOiOu0ZKJx8LUQd8d
fyEu2uBDQg58+hwJEZHWE+0SNS0pqyLJTe2D/UZOqZ1JEKFJRbYvf93YwI1kuF/V
gxJrCkzRlwRmeznWnOwrOj8pko9++wwfkrQOFoqTPLaGoQw5yDSiGaPD74iWAtAi
3LSyfkoP97ST1t+kjpbDgbAdclWMv9JlEiQvVc6lVPj4h9nfokA5jTUkLWlrE/Uf
D1HTscDIYq7YuUvNU76Zi1P8F4PmN+V4xyxFJHFz35EgK8DgE8Gc6B8+1dKGKqkr
d5GkI2sKCQfZKriHEMJs9+9yS3lOiF65F2W8dcdMPUtfipgkLaeJGjzHmXloxRuy
sct5DmlRWSgzwlpLlgzEtr/1lH24u3dQUK5ThqwYv78YX6FRmrkAqEQIMYSkRE+6
bCYUDEpYCgwOTJA5d7GtbxTmok9svgjZRGnjsrczZ82pw/Y3rLX4wZp3WDF4r4im
aVksnvGac6Q4f6EIeYffdP7aSGI3Vkh34qfXuXomFNxFevXajy1p8zmewBxjWSA7
qD5bZbJXh5XIje+apsWwajS54xUylQ8HKW6cBhR0iZo9cZ1jcOycyzLw5JYIARjf
5TkY12wb40PjZLhi193oKOydhlgHVWlLoADT8BOTPrxknz88HOAQVagLKCDXD4sK
ugfaZLqGYfOGV2b7L9qB0xvLzIS/8lBjcm4UNfgLFcv37cDz1ZIgrSQeCgy5KpDn
xMr6swd5BpBbrt1IKmL90M0SfEWcxN7972t12yGn5bPlzdKNybBJeHtBIPjGiRv3
taSdMMeehExvCAjncbjqsoIROxYHl1Z+pz0CEf8Ne6t/i6KCX9/ghHu3TjeOi7Zo
JbmU09HmQmx0E5OJYpssHbnrugs8u/x9xtNaROLqZNI12olWudPnaFZWhqADHgO/
Qfzus9Z5M/m19/cYxb6aOHD121HDEkbNfzpL25NiNlf4DeqyToNcdBm0UsUZBDEs
q2WYq7RPeo3n9eXIMzZEzU9TfcGgOLItmv7J1e+Ky7cHnesSjbPjJFfWUbzHmlgF
+rrDmP/NjfZEtE0FI4PBr4bLbyReBKKeKCBLuI1t/LmiCYFpxM7iw7WR04ZaFsOJ
Ju8P06PZgC9FZPpL5e98motI4AI2hoiHGEYMwQyNMHsQ/m0CXFZsRMhMBqEb3E0h
0oqGca6WYw8ioErEb5UP/2Os8ll+CUzW7RRyc8/fJy8kZWTfgAh1V+CxRIOJbHzG
JEDG2zfOzPZOg+NQ+STO67guKGMFw1ePTg15v4WYQ0ICi7ojB+Q7UxZ7iny0QL/j
KgF0R1r/d8O0mF+5vEu9f/8ZJecIBFHcO2IW+LIOYIJdM3aofzpul2FZ6PO8Dcn3
AK6Fx/3x1I22znRmXeu4sWD0C9AV7O6igBTv3nhKykhU1UdkN84UtM+yb1h199jt
6QOcL4siUChMCefc+rimg+NXHbPKKy2b/xiEDOMxb81/POJH6LuOwlPgM103C4ak
Sc4+24+HnBzMHkAcyAZ37B4lXZ6dvR//Sa6hyh366wjaA0aQ1VoPGhW4SpYpzfov
7IpfWQyy+KK9tH1Y8G2g/Jlzwgvk0TCsI7OOThExq4EH5g5FzMMWZDgfxQhohb0T
iLpnAhQTW59yNZhi4vWFAPGOnyEzDAWXy/SFvUrUbO7PczlBI8nugBsS43iWBLj2
0PcKr68XckNxQGSIxxB6eyzg/etADPag6MFRwjX4/p1UVMVBff/1VSpxsDpgwzno
iUQbxnf4XRyiAdWcj8aZd5kCHRhOn8JmWDRQaaWqj6PrERDC/Eddm+K8w2OQGO8K
tP2Cy/ocngwMKxLpxLfeVCSrCECwGM6dq6f4dNr6FlZw4N/QDGvIjUTY5uaOrGa0
XmR9lXXpBNrpG39mPpyzgrm1rYLoGWpt6YtH1voYcoaqJY7QOBz1DBC2TQ8JxYR4
mJOjRORmev+NvAjCdD0RFpRNDVfolhu64kRjFivhR+Iu7zNcXkLDOM8wJVrbR0cr
TW2jPAst+VfddOY62PN/oyOJ2ccQngb1mnVwZ9kCyFeRwer/Ieg9aSrJJvf4nVUA
ENpf6sXgq5TYtHNobVZG4sKuOfANbFGQdp61NUZekVDmCLVglXvgMK/jrGSXtOKS
n0r+lTQArZYD9RQ/xak/xcpllTglE7uO1Vv7DXd5tPzRW5QeTn9/hNA7tDMdxKbf
XTYtWntzRcW/Czfx6eUWSZ/rgVe7K2JMMWgR2mtKtM2ZpPIDF27xaz4VHGzK+qjd
NlZ75tp54BXzYljrOVXBHyxCWBox2SxYvB+uEteuY8qnS/Q80A7Urmt8/kbFfx1y
swH3a7E+h0yUp3hBciVaBjWxtQdEL/1FhA3/CMMrVVndWHyI4brpZU2ZeyBJyiUW
vdipKyuHGn3VL+6xwkRIxrI0A4Aa4DodN/ZhSWfGcSlyZ72m5+MkzgqXJ58faudx
KkrS251Vz0sBxVpW3LyD0K0mMtqhDxFl/15VC5EXeCDN0PLyhmdXWPvxMVPqxlXO
a8wefHRQ6IPTAlT4oFHEnUhSeRISfOc3nbmL7Xd9c5U+Lfr98l/VE/P1uCDEx+sX
cy9jTp09McX3ma7giAAsokug7xFWWKryVJSh2rgOKR1iagUp1dYkcfjJM0yiWX0h
SRi8jUCMDG8hK8AYtBYIPytqQRSsc95zUcjFEGN9qM1NBTRGtumrzXHVJfSh63jL
zeHf1fFfguTKaayZ3JcnJKXfq5eZXO4WPS32043nmezxhgR9zaWePirXHZmHtLmc
7+pVp/omFX/PXipWr6QoPx3FL33dz+CguYOV3S/5XI5gGzEikmvHmnjSJA+jbRpM
JqiRsH8Z6I+HVUnKJXpr+CJRhZ5vmLkBxoQhPTuWhft3nYmxpHuobHExtokXiFsX
vXx43yMV+jpWxBArE/XX+l+clri2D+DyVasI5poIW54Gu0SWpqb6A5kxdYIBVkbF
fV3rus8zaqd4ZtV+6nWRRsu5c5NLK21zA3COlD9jWd2OmE3Iwv8Y29kJlPdcMrsJ
f6hTBFWQT3WUzgp8AZ1fBa76vTd3ylo3Tq2HQl4rbsqSgDMxiWm7UoSFByVg/3xu
maROKZG73fzg5AKRCJiEN3qcl/ReyXjmriBJgdpfj+HMPRRB/FzdUmMIpUJTRjNi
mgvsqcrC+tzgIEM2oLqKlHqRvYc1vZ0aAQOZ7Z7LZYy+x0Q0DQ88yj7KKByAjTq/
9QnFJKlkhfvsUEgbrBTo0yB8+ErqHIu8A3O+n/Ip/PfJ2Oq3QuUNaPDXbj+yFv/4
vXMGmnoHrcJvyxMYvhzI1WbqKdUvQy/10GkjfQ9SpDk6VS2dwSziyUQG3YB/6n9R
Cl67zGk1Wol+rLtdbGodmjnIPaITGVoezIW1czZJP8z7SByxvJKuphBuPXwS/4Kv
2myyjCaWq1QB6kNE3yBqlVBKH5knUbkaqNegHU9q8Fa2VHehRQuKDPTzNkSjkH+P
CkVLp5ky/YI9PYIIqQX+PHxbbsODie3v+EhiCbZYX5RqEFEgevj+ceWrmGivwo62
tKWcSRq308maBBUQQgEzdKf7ieFpGkJrQ5KGoy5xCcMdqSEqYSlgIMvIbJXrhVDo
toqo2GDnzwxMO/mzaN4DyuQaOmbYxrQqog1qHAMlNx5jah9WsrLgbxWxGvTfsu/C
qtGI2/iTk7VUAMD+NZ566mPWs++e9coffa2w9eRAds1XxREd4JqdnvmmDYBLxLwM
0AQYmb2M1kneSRkbXwynTuEFtWyAEFi2cdArOL5fgNFm+YUYNg4m3M24yf9Z7qi4
6cM5bId78+lzN766MmbPmN/S/JBf/9QbHVNPFvKQZY7vg37Kis9K0aA/WOsgVjJ5
X4ibKUGh58Wxjto3aKpooWZF7/QzmxMVJwaz4GRtOh90NsAfclx5oGDICa2Oc3mm
OFDri1OedrnVX6Amb+2riuyLn7Qr7+GXsMloBEi/jErsBN6Kmp/vAjodX8+2Xd0v
kGzraxn83etZUSdBSEgKmCwWvCUr8PnK9KyngxizWGBVoLKRxok2EQeXsZxIEBVs
+cnsFZltCmxPgeOlYMiss4SEKug4w/M+dsGnC18DjvHNa113+977vH91l+BLeL8+
rpHshpsooOCqCdqEZz8bCWalFBVbmhA1ANrwZrwPvg8ExJgwKaFWFiwBvnRFsQXU
yhoAGHxDrVqerMmY5q6JN72rFs5lwef7sfHX21tbwpYrqojIOvcbVQtURL6iLMXE
IO9tn17RyAw8zRcOAQZM0ppl9NoSo2N2+iDK29pgOsnswqXnZXWBPW9fI/SC9eMv
AYQIZZBPrQGWS5t+BCpYMOt5UAj0V0PZPrMVde4BIk1pDzDP+QoqGtcZuzlZjBhH
su9S4fUEJva0F97mBaYIh5U8Z5vx2OopdTsFEDILVs+9dBQlafz8RbAv9Ebbucrf
httXVWiOk8hEBJzHzXhsbhXiMhcd/SpSO/ZPh5bn62CqHuMOeE4ah7/dPVJQq5Us
QmQ/23Iwy5aOVTiUDaCdZmiWvglTZ68tIqzGpe6qoPEjV81PzifB/Zqmv7hSGIx5
cILXkloKF1lDuqB4kx8NgirlE4AEmkVBUX8FimcmMjt6W95oRXnIgJwugRDtuBMh
km/2DEfgZW/9u6PNajNrK3HH+2qINw0WeufgfRxoYYnpH6mvig515N5IjabMdePJ
AtAaPixnmOMyfrrdBVGrGmky9t7FxD++IwYLCPmCiNgrwdsx/DydyvfrX65BqpWq
3FJT+tyMHFH7LxBHSGV0Opm5Q2vQs8GZzIbMCr3BPpIm3UOYkjotmDxNmRA7IKeK
P51bIs5kPNJGCNEkXhcWMqEILXQYb+Htnl5C7/ELN8uA2VcdwNREjnk/CMFh5y1q
s174gS/fj3af2RRr3eDtcixlt9cAy4NbB3YsRtOLtR+iGp8H5Hqbs/S5kpeghI6g
6Y6MkJgg0dP0881XGQv0X+QUgAk3O9nvBXFdCKUzS0rOpgHrlJc7To+sbkmtqT6+
E+4JFFTh0z57u2C+xAm5LFqNrKZw6i1FZtSpHnVTdqJ2s93sqh1tth7aqFXzPbw6
h5ILytqfNasIf4SC8CU7nIF+HPaXVdbcGnTQNF6VqwzXJFe3QcW5qm/sIp8hpYcn
Zv/zNxBricQnNnYmVCFcM+3wprNFaeRNtWpgJHwXRVZEwZltkchtEKx3O16t6Xtd
RRL6HlaGar9e+mBlpNEAx2Qgwyr/IgvPRVJKpwvTly2OgdnI1toNIhIeQosVZOR8
f3giz/kXyce3woMj8SpPetq0OQu7Ndrgmmizrd63PNHS6Yo+xg7s0ezhBa6oIsHt
Fyn2vo9DtZzynU7jpU1VeHW/2E8m1oFRh4RYLU12Zw1vdcJ+cMv2qfn0a5cM0swx
Ad3W4reSawswlO9cV+BT9tpTes6g+eJfs0t+QXniqQoKf5T0vPoTIpKyI6/sOJnn
tYZLJgNX32ZqKQg/UGmTaGKLF1rlcrpv3L6IRNaFHl0Ds3FZgg9+bROZS2qeyxhh
BcB052dC+6mVowK4reKL6v/H9TWqur60Uer6xjzsxuwcCxU9eK4GBnAeIUYYSYsx
Xm20cJ/insdHuK1+swtQ7mD/g1xexHU4duh8CZxhWpxHg7i041nvNJpouIDCrVcG
GWUdn/YEqfT1aVP8S+RlAUvsTrOOLXZAWT8elvGggWnLA5jQG5+qdQrttdhhEFiR
dGoMMwbDqKD/4vQ4pU2XyhOrzMJDDmdKrXhhzMJyXJmnT5AKwbl7lGBbU9EgfGMR
IFU1fdB4ZgThwJERFpyEOh6jnqJMa91P6+tfy9T2iD0Uhif+vMGAyj+U/AZOt0Za
6qCmVWewZcWfv08ZX83IbeKArbQQz70606j6yM5ODp2wI+MYKVVcwH11mHfDq80I
2EtpeUpQeUA3bmcmXa6SXALHvIjOQZdPIvwZQViJRxG74npCqKcdQhUBlAoDM5fZ
vnHk85HZadLRd+OVdWOL7OQyU64JFlypHYPH/qTlIf76vpiMPJJYJilLD3pNMtxi
XE1SRHmx8OqmuYUGX59U6iOh49Et3oDZ94jaL8n+h6qTks9RPMjI+mpdTk95YuYT
7r9I4OkKWf6OURQnN0hu5G/hcBRtdzH0kgDFIM1MmDzzhbN9hWh84a6v4AeVSr4J
PXdpU4WTOxFfHQKPeJfmc7hn/HIyquA14HOI2tdgxlKKmBlupnLmDWcP+K++mIMC
MT3L9k1CKKpEkbl666hs2gHPWTlV+XJrOnBe/C83ejll8sMzIeWUC8afahdMjn3v
c0LJc2HmIM4TxoMsgHi7idob4PUEh5fsYRfwiEF04BVhhuQmDeq+n/Jbo/OFijyY
pFMuOHV/PkFPDOhu2EwJNzD0i1B913eH2IDYEiT/mIabuAA5TcnkOE9N3ZOnjUzS
2P9plb/lL+MYkszXvk7o9ZJ7ag7D78rf7Z8XPzI6s3EgUkvRFrxElJD9cfktBmhK
hGdGtJmwFNHhP5z/LscUNu5TW7zDXXw3N16hvbspo6FRd2Lyz9BjS9rMCHlQqy0q
bTJJPzy1ZVfKzzRMk5yyqCMCzE3LkmUlDcLwc0c1M/c1INwUGkarRVReNIG24rLd
7dC6gRLmJQ0a9W30kYNh4ijAzkfwpGfS6OngYRlxXzXP3nSd025fShS08cqyPESc
QEC41Y0pcejBLrB2Cmky3Q+eSEGOLPse4/JkGG8M2BV7VZMcBRN0YOuFnvMndMKo
GMgHUMr+DeDuaApUvFFXlHuBvl0Qudz6djje7r0LIT/J6EiqsOzYqwSrOCxml0W3
afc0zsSLGA+SifQY0P97/YqWOZbeA2wlISD/YbcbDUuvng+0fswhSwdlCuovw4cN
+FWGDUkNjQOcAb+U8zQjgNzLd3XivbWRWg4j3rme5LQ0hPgbazO9f9ppXiyXLmdt
gKDcrxdf5yFpqwTpzX9JmT/drC7VQjRJH/bmFKbCWyM5MG+HcVZmu59FL0LMKzp5
Gt7ybCZRyH/xwE/uK4YYysaGeh+7/tGfjplV1+8SpAPWfCfjvNEJZgXAr+urgtMA
OEQ46xEW5c2SMCAF5Go9NNWCQ6duvfFvnv7CnK8iKasMDFN/vP8yHsy10Ja0OyUf
T7UpexCwk521ytfDmtBTlPqsUBAVRztbx3qXpnrHOWkQZwiQsk4fWxJUqhRNnI97
NjnYUL5nX02CPYb6ybOF2XB1R9MwCol6iZo8Z0KNrqgGjp3LHRRnYMVaGCFUAZBq
ZcD/i+RmCnMpz5Bf1KkB/CNbo++if2omkWJoi1pi0qbHOX8cy9GNsA80utJppNho
YA+YtesSbwZSndMC8mK4syWjlcrqqqeYmPgoWmGfW+KPDNv49nIAC8c7p/BO2YWH
afkeYwxDJMa7msPuZ519D8Tag/zqwUvZsgEQhNIbu5nKLSKyhq9OMzRpbXv0UWHG
z7RjjmJWzRqvEEb01z3MDFdgp/ZIDjYtv0xRbTmja485mS8D6A9FygwJcqmNILan
UDEZCyLIgeZLazgkp/xshu8x4+PsjMKRgq1or2nJp3hWDyoaTrSn4AqDnoKtt26M
J+8aDK6vn3O9TUONKbibHGF6EeIpDdMvXvH/JKc4w5aeO3hnlMNX7qGKkzmntqgy
rBY36W629m/xmba88mScwBuiB2qRUeeYFrFpny5kn2QRoVqCqE3PdXSQEqZ9+AHY
Unmocsx0D0kXFZx3oshuauYWnFoA9Qny3TxKRy/ZX1SesQjUBilPU6rbt46HecV1
+2PAFfq9Hqt6PrrVIWbxMobmWGN1KyNX0/OGdc+junOMB5r+TISJbVPLLRToGsgO
AXHFyE78/2/VMVTPpyR/o794TQawHvFsFYXJrr6hS4QbcPQTgEInsfTSpDI3eqhf
bIANtv5SVv2QHw1Cli5cjDc912TjWuCEoIqIzPIGPE6fSH8OegNTNP/HYvd6wS2R
HYz44saS9d66Jg/xil/GdgwPKzR6Kd+YUibj9sf4YshQsPFLpMJsiDWXOTBeYXqJ
oKwbyYRixrpSKzAMMUhK+h5tV7BhuJsdUn9HR3EL2p718psOHUhHXRHBDuGag5l2
dK+ryk/vErsoK9gfCA2N4IYpRnDbibY0gxF46lEBaxYThdbrr/Ak4xH+4xrjCAur
XSdnvnwBNGK05t5lPbImwC6C9Xpw1gkcl5Tohne/4z/PGSN5HLhTmTIZmhmdsLZj
88/5MkJtm7J0sunQb78K7A7N10hJJTFqioykrTUpX7fWWlhvy6YOX/4GmPgwa9QA
574JhU7dosx8LHh4atgkBRVHrpKDfh1i2PsEo9d5wb+q+6rQWK5aNDFwk3aPN1B7
vIbycQ/RuuIF8mefAr+1sVOG3725hwCSJ9XbGl8khozYyBZkziSG/q1qDN0JmoZz
9SUFypEWWMdxtgLXvivEPV3Pant0A4kqbMJcfj/Pe7z0JlKEIM7M8+NgqvyGdtYn
tVCkw4+9pm7QLO7XhNZHiAsd91z3BezSKmrbjg0XG9H3cSOtD9wdjHTPAW/B/7hm
kYsyiWffhRReVL1pqTifT/SYbRaPnSaRMGuTu/P40S7Tx4gJT4xyg7cg/+x/ewMo
uq2gF6LJqLBNvASw4Z9+beITrhZ/3RJIm2Q8DfQsj9ByisCcvEOI+BBONME+T4Te
q3ciC8Cv221N/k7wGfsU2Kszf9bTQjxbsuZeAokBUzDnEd2H/4mGRwPTHHqcXf9m
vIxL1KVrOVrp6kxlM0077tJWDRTuio7zEv+jqwANjJHKd72dXG1nlO/tm+tMP6Gd
Pg3NHZ9tcRiZalF2mqOIl9TIekRbnf99rvbu+LNcogaIgyOCHjAxUjzrLRKhjcII
+o6xBU7tggJoUAbxKzUibln3my2VIL+gaAE8Q3BYe10XoDz/UOUiyRnmV5Ttx4dB
wOv4sR+DaHX8YolXvVW5gl67qMVgeyaJHbYKdIl0Oe14SEwwliusiLjrKpjiuy/p
r6aCjTQKaWyy2/boN2zHgtr/dJuCctSriSSHS3MARo9ZmtFNQBEzNeiHVIlb8gX+
S8OyXBc+ys6SFd9ia20fY70U1nyNrVyfEcQCquIqcSjQMw6ujbL9G52KRJuaeNTj
76i9nnqvTCvrlZSPNlWUqLwjRatOppyXx4Ryff4Qrb1mJMzkZ7VGTMxb2LeFNC83
x0PXqZ7dOFwtp+kCT/w6k8rlEoTUN31wgNkUZtlBjjbIRp12Td2KDiEviZarATYm
hXqq+r+JqLnCEl0rLYu1j3ogyVIyDONzxT701Wyg4yBH9UMQDDgEWhVSUUjsxGar
ZGaIlyqG7bBfiJxqyljpbLYQkJ7nQ5wPHLsacZu9EL07o7y7pZpqsE41Ajw6Ieyc
oaWhhDhwKoxQjeirbiLYgj/EegzWroED32VnRL5Vir/TPc24LPFbpMp3E7jhlQNC
+iQcwEVDTly0dA4Hxh6VzcDY3SXwaxnveQB5IKe0aDiTJMmr1qNKdiFc4kAcvc2t
5EYV1/cZB/WTlAIOMXMhjcOtX4vSRDQmJAaYWKnEikBg8Dkj72fcrkEE8uzPUTvb
jxraYHBJeKYFnrGMnNXL4lv+WbWKvOnsUS0JGw2s75ICCQVWupGff27rMJF2jVBC
0bud8IRgIBUdBlxDfyNmMMPrphbbTtKL/ijAHnK5b5XZeC5nIHI3+1z7WVGKL7U/
ZR1Yfb30ggCvh6jRFmjjf8SqmWXrTJ+HvWwrtSnoO3X7Sbee/kFkFI6+7Hxer2/T
vDPznPBWyDWEN6NeH8zEWyrrq9To9e6krfgI7pD7JesBxVU0C36Tck6yJLdUKWyo
025g8hven0p9YcfXe6ODTtFaJEWICyt1mfDq9/WnWN7CnjbdVFTdf/fIj6gHIjPg
zcmqlny/rA2iv3ovPhbwGWw2Mq4HsyzZ7RHxfnfpceSN5HLisX3Y/NelIEg1Gm8e
+/369xahmrhzwn7JkjStJGKDYNQlq1doSywVpFlUUmSEBWQ/4dcUVo18DJHAO1SM
3gOhxy1PeJ8DVEl+jplvlkrv17pH+HvaprPEcSLbKe/R2D33LLJ78ywL2UI8a+DZ
10OS5+pGzMsxrS39YicjTcZpyfJYSbXY9msjQjzzNnvU6lMq7OuEOR3Gd5YRruRa
k9CdPdwjZ8oRhsOfeFCeZpoJUodVG85J6X1HOEpbJEAPBEF8rrnw2Yth9jZVQAAl
gGgRg02pigcFu3/FELTyfD3zDI3JRsMvvP3/cf10giLMpHnITDX7LK5u4Fh8NIqh
2MVbRFdGzh1IvgStp7FT7UyTVZQWUgIxMRWXayF3B8gALor9g2wkIfj/hskEH33u
aw/rQMzOovJMPDr+qIw9A8i+beSDPVF6jyJq0RNaR46inzr3SJ3lntMVD0o752lk
en2cSfBVOUQ4Rl+0kZ1LqaARVnUla48oipacNAhy8L2U0Onl77aFdLz5dFNIfZFD
YR25fK57slp8Tks7XDGih1f0Vi8D56ZEn2uej2znzy/Orh9ecaNdmMOG8MLdGnXw
HDmv49K6nfk37zsCSeRqGdroD82HY4+LmWzBzzSBtFNdT65XUVTCrJmtD00wphgQ
75voVp4CZhW2poHhlqYP/R6riza0mzenup96+YcxcMsZMEqW6rmLfLbTs+UIltTJ
O0bZLlZt8Cq5we1UwILHdhjxfx2Bs7t+Dv/5egW9Nz5VOxBflmiHbMyipq57ac6Z
t/GBt+Hmdp9lp7xZy4lrSSiqicYyUDUd6BBPE1oeACjbT/k7djyu1yF7IZH3U04u
RjklML8j0lK/UaCD9FDNDXwEvyUtSJIWH4U3WKG17pzQI5xbQLZEMe+2ccS+NUPB
VjykInIEiA3n+VmJP76I8z3WjvXPvqZH2YBvYj7xBbRGsL97wBsj1wD/T0slio/S
YI39V2zRTTtR9Jpc6zKNr9IFAHaG/1TJhTXUaFDtFZNkCxmGGvJfmByX14qZZIDN
Jfvw0SShRu729kARfzEnh6FfvTPFO4/sXalFc0Bkx6ybSNTgGJiNWCay4jZkyCt4
hAKqrP46yhmFR7DhnyWeMn3uhoK+w2McsCwnVWIgVLJe+4Tli//SvhPQsW3M5LxG
b2xZGS1mEeN5NV/BliwiKTt+y2FqH/kqYVjgQjzeNrcDtnOVkoiTxsL2X5DW5tq7
H4D2LJ+n1l4IHLPwjNlcZvE4K3ny8GBtZGn5Wv8fnRjAOHAzQS2doW23wQbrpDY+
+ENohCmczovQFGaw1Z3H7TdLkcSYTDGYuhzbG/pIeFMQydBs8lDyWEsOBt2WKO+H
8p1FYSFmE1/NIGeDgGoQaPGC/vmhItS5dEXGL0mxKObM65LQq9ibB3/jGX3InIhs
Vq741QYPiNQy3nQH0PpqGsSfOAdfArPVohvohHwP7xd+/5mx/HGg8/6FXhmKjkc1
jT7thJwrO82biGF64Ms445sKw50ysIhqebXyjvQ7qtUbZVvarEmKzJD/sNWnGgaN
9f/N2ZU40WcJAH6lPaN69SEbJeYErHI54/etlF+T/iBS+E/QpguKL9Dd2Zj25N0x
mAkHmdNvYLke4jwqziqPiF0EtX+hhcu14azagrP+2v1PImM1ANC0JLbpduRAQtg+
aqtmFrcxKVJo56eaJ3JDxm+vu4/Drblqr8ZmaA4vnNlxJ8Qk1d58JZtFZRIoQ1gh
uXx67jpxxT0owa+ioI4/Hd890DPcxVS3zBlRfpJvacx5M31qcBbaicmE7URhBUFS
m4/AV5slkZneowkVeXfExKeOdP+0pvMpfIf1fobscTCvrM/bU4ZEyTIOwtGYikAk
uNmeWCwO4+n0V/9SyTsPGQyeDBsZfaVQ6WecrpV4KMi58cirzbxcWYq3tJ0cRIQb
kDCkeY26Hq8cyb11h2UJRVMEMhychQTX6QAMUJdT2KC7iQ7ZS7Z4+801ni0Pe8NZ
/l5CHguXnLsqgJSWlUCs08K9B/6+GsC7MXZpzLE8baF+eujohmn8qIrixc9sxUun
iEjcEOdlzIU+3RyPk+EbnknuzmccRmfmlTZYAj9A4+tXLkGB3zH0QcrO+jii/j9u
6iGc2Nr6CKm6b64/YoQR/ZkdoIFR46vSO0BGpiqO9gjs8MUsE/kmx+fe8iGHW177
tnlB0bswldCZdfMQZMrPPsslVHPO4RuA1ZHJZ7wZKztEt6S8NQxMCzUte7Kjk7+e
O84s2JvreHjl4Grm+gKhA1TF7rrN/R7nGZE4QCwraYuZl0lRqRGffZ4Qm3Edxjsv
P3lH1RGrQlabFv2MaZ5LXd5Shi+qDHXYll45++oaI9oQldGPWY9e1BerkV5kfRnq
CDH5b3gI8vVG/w0S9isZIiudkqwqKneJ6ms0neq9RC3UXdAgUyw3fCShQNMROYM0
G4IbP/s7dzG8Ot8P029RscCvuR8d+WVaw1GT/3o4KbKc+b3ymJ+dBko5zAMVDeC8
fMJvA1TMqH+BxS6wlwXE4kjDtc6L1GtHTulykEy9IuRytq9Jj60RhK4Y/96KkfN9
HEk4/EXi3a4RDbfAN1SwBHz3HVU/cGlgkEvg1HtbPJgvGKGxO0tACNVbY2vQ+b3y
IQqQyLO6DI9bfS2k5Xa9Ts7OM2xzz/Of/YUBv4qkE+wa5w9WALW+nKknKEtwEIAk
i+iOCnUza8DVI137+OYOvg6Kt0uJgiZ64roy2cz3WF/f0rsbSRKRqcIOEqRbQNYs
PEUxzUhy+N17uFhnWij+kIJoHDpuQB4Vfo05WeZQlFtiR0iwghFAsRD2aXoriRSx
D95Z/wMuromy3OXcK1By3umHboR4eu2UaW/pHjOmJWTxzuSV/7zW5FiKIKIOpuX3
8comQivfC6WQNkL5kpsjFeDjdR6A1GBLw/dPBamTj5ocP/Uhx8sUrYkTgqPLifBt
RUdOr0B4cJ65FVzNFpyz6FFR/UHw3fXqn/ZQNTEz65sIamMD9jGMqn2DdR6zl8Gv
n2Vt42D4LVdfwwu9tikhKU9fhL7AWNJQnXxGFP5RlhbYA8uWz/0hE3uoRKYIarEG
ZDoBWqMWpUwFMbMKsBiTJPmZHDNsFEpNT07hGyeZ3EZT/09qqf6eZiSswdW6ZBaM
FQeVrTqfrfveUeFlFV7XKiyWIzP8SSYPpVWtUkj9FtEdq1YxSAgzSRFTfgB5CljP
Tgm/JEmiezKTPXVz/YZi6AbVw0wv7ORk+GnjYgwC31m9+k4RwnOkp8Uvgc99jguZ
8UyVEsrMgMCNJmxkgOiIvjxDusxtXtEG02e2aSg61scVEqvp6jF8qI6OuIzEbjWU
wl9DO1e77r5mEhbl7Guh8Kz8s4i0sSN6xPZRJo9AGqUqoKK+2WXFFQTHtfWUtXuZ
N5q3W9c5jRfhUrjXa79I3+XYXChvD0oyL9HYpc53H2nrsHwzqIn9eozyMrBcmV4b
4mWvIUF0YyLJfpNaXgqZtuTmJXnKeZe5MRu2uILPExLiqhVf4nhqwe5WhLZn2aA2
/M/33IdVWFsEIRi6IcBHwgpI9EixXMSJhm934rvfNwKBvXaM0Z6aghVjKM3jWxS+
zxxHW3d0kTMPZq8VLZy0apeyxLpiDk3hMft+/GveJqtYlLAW7DEjmo4+HSdyNk3e
k2iMk4ecUr2IDz1T62Cic93vLWtKWliG4fJRDTfBlEF7ij6s+IGaeCzEnQY6EXrV
NXRTJ5aao/8hy0+h66USIM9TVEkYQUZ/GWoO+CCXdLtvUGP5jp5s42DEb5yLlGJ+
NONAtOJQwtAblyxnPtj2aSPokUpLYsQvSl2mSGNDNTpk0U6CXX3DY1MGCSJlzXu0
N8lwEdGvJtaKKaVSKRHfX37IFZJH3gaUSVt1pSPaZDTzR2VJ6noP+Rev72+6zS6O
3s96ImDGRVXfu+oS/y5lzWzv8G/4MP5LrvS79+IkkYZTfwcMcCvJZ5CD18zJ2Ekh
LZ5MPJj7yMLHU5DNG3es7OptboyCEJXsQJnYtNU/1bWgnmrJDFaXuKua/8qQWT8U
LVl/w+nstzFIFBwBNP1UMi54YWFB4tUlISaHNJ0K8jwmHrIg1Zokdh/GtkwX23su
EcqFv6pLXblZewvAGuKaYKpBCJXNO2+1gi6vs+cLrxsPdRrdjjT/e0Xf2iRpDXFi
LGbbUwRyUToPB7R+VqYO7IuANuAPGjWgV/IQ2zzm0AIzcYOfOqRGjuLTNi+FPTAL
YKcn/H1yIWeV5klC8R3eUkprAT/GWb9PLWd2Azw1O9DDoTyXLSzYRCVykdPKcwZ8
QNx0+bUiojfNmP1v8O3JBa4hvC22MHzC9A8xunQLOS4K+MCMsqLzAJtLSC7AvQn/
b/JgIuQ6+b8DseHDNr1SHptSdOlPRG5lqtRHBouJ/9VM0/s3ecpMPq5o+OCv9x8F
VqdVxmYK+Z/k2HVpB8Zh2icBjaCZI27pVTlWm2EbeFzkTyFp01t0F/cmqnCo58wF
YqYCpo9EnvLNHqp8z6ynAVkvM8UuIAXk41opMW5iBNEDyK8nTy5VaYcW21d/KPfX
tYi1dJ6g1gpSENm3qrZkXYPfIH675yGyj+235hdURumP4PpUGVhmQiK4ugozEZjz
C4j5Esab5LiqJv+c/i3NN+nH/PtqRXHeQ63th6WJ2TxM1ddXOvaIEhjpmqGmCWzl
+ZOrJVKtjNRzbKrJ2jsxLg4tjMX3CB2v5fZQyYcYNA37FFGDhjxTjUltvhTCpoEY
Adj+Lgo9iJ5jrT8fm8o94flzDzCaW24Csa8pssjPz8aPmw7m7RM4EC4ErzxDtBoZ
rJvqTglvMbfqVC/HPMgmHdbiaMeE+MGd0dLBTPK+hWZ4M7Kk1K54yfTZjg8e7HwO
l+ptVD+dkCCyicpliKxuD8EnnKie000Fr+NWYvPnikFMTDVOhagtBJ2GWHPUo8Bq
EQ2vdvF4lO8AqQHx2OxkoY7pfLNYA5jv12jjUZkOgHEB/6JXoenmaWuXPI4bim8+
MMjtZPA5L01uEtLfX8ASkz2JHn58L9HQ7qiBnFPEWzu9DtcwWfBUEcQW4DD0edA5
NsW+dj4XZktH2U66SU7NiRYhTLrpw3osfdgXeJwu2wdH3pdMs/hCvqzpu+ypnqgp
7KjiLHT9YYtOEc635p75uyQ3HADVGdbd8ajfip0WcgTFk2eQYSNEszlINq/3iE9V
Z7Gh4CyHqKQ7P44I0NP+IHI8mQ2xyljYMnLUcyE4TffRnGC1YuVVffGA7HueBBrY
g2lk11LTIAE9Ya6Vfso66wGVWt3caF9W+44OJVdOYTxMX3k1mQV4h99wNshs82BS
NYUXm0DWvkSlma8QDvHG3mxxVltjnMw6SKEIi2qxSgRAfz+yCrqvCGZX8hi6ICn7
djUzQ5sC6pKg7gld8FWPuP960pB6mhTZrJblx2Dji+2CIVf1V743k/gaJxyP2hYr
ky9f54JmNgPXnICC8k2Yu57jxD1+ns0G1n34c06y06IEcqtSlYdfQLEKTzqJ0tsk
CGsLIc8s4yje9RS6bN2A7X9QGqVKPxifrfkTucyVI5tDoimbKFUaAxeT3Zpn7MA3
PoJ3e96GJaZrl+MWA49hvhZ9JpjYl54TyUU2k679ah0YKmdgyXMhq5KhZv/C3/K+
UhGOI/zNWNmGobIOYskdCAdH8hAobvWORGlm3797l+LYM/P0ffxiC38Sh3/ztdbT
xW8pqYlwIi1FH1ElAfJ2wGwjzQlp8GWmKs2IfroX3IQwLDw6VrmoId6e0A5/hLAS
Ciy5tiCOnR1sIe3F9OwnwSDpZuOoapliB7R+iAMuUzbnFdM4C79Y8voC6gmRCyEl
/wN3fuZT/p4AfwJtkvdSkrtOBxxyETuT29wwJZgCxLAmyhr4yvBjPsTKOpUup8R8
3GXSyT/kjpgKFcYgFa76bORd9prrGe7LOVeGq6Ju/uZ4+HgbIroeFC0vjnJAwNUp
1qtSPxPUJjxTHf3WEhoLxW1IoNqYZbCfQRLR5ihboqkq2UbwcpjMRATCIbUUvFtq
Z2SUKa30DtrHOxCEPAzYXUe7i+ZcffbccRg3E4l3uLn16mwVF2po8vGdciUBJtiS
NIGEfXfjmpXZWRwTdIqfJD3+vmnDqJ96a0PsGE01RvVkLEo/WZ5pWATpbQwwIwa8
XcMKNIxtiAPICeG3zyvcQSwNAvvciCA2L89e2KXXOef5ygH2zNenQ0mtSswBZtj1
00u06EhbMka/03yKmf0W0pvYiA9ahjT4Wy/HKSeJEcCb9NE7KISmZFI7P9+mwX+g
J3quRJQmRR10p0snQF1eWcPPkqSocVuQksmusGD9K33WRtxaU8mdMy6NH1QRm5rI
oYIoXixQL4VD151ONLfAzJUIcKovX43HB235Z73GzrWjYtsrxhfN9xMW2uPovuqH
rGHZApAtHAdG/M7CCqziWwtNKopmFaChvB2/KzEwClsaWpbkp6vAmsprk4Y2VlBb
PokUMcuEs1Wy59RoMrjyZ/9ZVH4xTw81WDwE83olYzY/aoHyvq4dwevq4cSYkfVP
2wbin/HPxJ7f4hFLnI603Y4dp704+P1AgAQ+0F997E5a6OIrFwIfMNONoa8E3tBe
RmbXOXmfeD+bcP/48O2Ur1CaNllKbfiolXhu0QKpPR9HcdEgtp8Ug3no/IdoEz2z
cWVPa/jDIf2XdqvJ0IN9lVGth/+uzkviFtSjvhif3O6g8klsQ4xBEBjZwocp54cR
sZ+AmqcqnKM2thQZ1rxrwbWrxc5xv58W8Ja1Y26lBagsy4Ufa7SumA4kc+aLB59y
m5G5k4CJHJlwdXZEVijXU1CtM1ga2a5WcXCeXFbXgkQ/JokEEW3StDbFYpcUDPBt
ksyY0Fni2HsZ65VqvlrwfjK0IZNCqCnuimmJlhA4eErYn0exuMUoHGT8YpTLcsLT
BGoYmZ3CBWwl82204CCXDJAC0mPaGF5+G+7o/iljubWESTtAx8fVxuHLZ901YR4B
P5MnFO2yFPFOSreGV9vG3CEa64mHlUE2PiWg3rzT+jBh/pS3alrozfWNuaMW/YQN
90DQKFaAMelwLh0NkkknvDFtlvfIUQCNYlMvEQETpeiQj76tdGWhntcunILIQPUG
uD2plvagGTN52IJHxpKxvZzIsFZd0AdvvSU6R74geAfIkejwlJsQbc0OGTKdk6ln
XPgTlqG9GByrz37F7zjrdTXmSPkJ25L0LjIdAr0hOx1HIxcGdn3vRMGfsSOJu3Am
xYken2W2+9AR/haWNWTkPT6JOKuJ0JxsKz1rfra6IQhp+awRbyhwmaV2mQqMhc5H
duTS6hfWQJGtmuGkOQJxCGOK4Ir53wqs5Fk7M9WX3KgtZWULXZ5PeMpaIJfJ6ilK
SFlmm6I41Ty8xHz9BLOqMTmLqiX0xlrQM6X7pJ9XDw2inR4goctp15/h9oQ9lsHO
Q62eEdn/ST2XukuxDuwA6vs00OTXCO4bRtPVxLOqnpV1m6mn+ciztAJxonoya7bH
3aixxH8439kfbDlw9Qp60JTYBVzYmhV4GMmQ1u6kn0sEIhGkQFtfJR2pT34DXuHH
i4Oc3RnKiJ0l4UEYqBRp6SHmn2GNHogNzAVd5//a4oNJ/PISe8K9mio0q04WO1L+
+wxtHsOC6q2IG9B9s6n4mGiPWJv2wLzmAze4uObDOilzVU73t9cfcc2pH8w+3O8Z
v0TxRdNPFuwFXfoMVxf5pPDt8NHTy9aPmW8m+zH4zqCs6j6oWd08uhziIKaqwThO
Kc9BRvF7FFVLT8UmqFW4r2RSxR1ERZXYCQDWemnZo5s4sxMTakJkqGrX9ac4ca/R
UkFO3IB+IrtwQ4Xx9O8iqvKN6iXHPwKssXv77cTAP4lpHtBb1uBKm9pVa6odiw9W
yRwpa66ZbJ2SK6i6Y8VuHr4qc2vUMLOugsYxqPYU7Hvv2TLYiFS+D6y+QIflY8ox
FJ0KNYQi/utAQGQuQKqGAobVaDUSw4kUDjQggvKsxhxEn9sxE0c0jKZplM6Co7iC
B1jN9ToWgHVDTHsJBM09xh4Vus8FRdMoyrXjA7o2p3akoi+DkD5mnsXYuCbrWKYY
NygVakTNI7Am6xVPLI1eJb626j+SJwS7KnC5knFD5vTaez7ItiLGOOt3o1K5GKVZ
y2mvm13Su8hY4dihaP8PNZsjasR8oL8BBUcrpy89PiB9zAKIr0BEnrEAkxdSYEsY
XkZi2kxqcP+Cpjhb4iVV0nj+A4VPauqOE9irJun1Jozjxeg/1PlhhUTxSPKG6hEC
fvDC+A0+gk0ikdd/sXVw96YXmeZTnJqyDoxkEuNiNUZvSEnflYrOEz4YGGY0zdCA
EgesQvqTD/8eOMu/L4P68FOuK32vnMIEmYVgvIeB2x8ECi/p8VlN6LahykqAlXSv
z6mP/J8G4eBr/V1UzT0bM3XJ0eJT3sOBLLqQpQnPFjaeMX2+j9JjjATCoGbBbliL
pLIh+ZaSNCZ/r7RRu+JlXdtS+FzS570b8mZgo63jVqucQhx9RSNMvyGPAh5yFR1q
rQsDCYrgWKA6GNTZfPGLZ5v8FHzK9gXPt7IV/AqISGowBXet71Iz/lsLU6jM+Xwm
9V3ezlLSHHUfJIQXyp+MKUFJv2ReWxJKTywfhdMP6t1FfTvisLojkdK6GNQzLY8k
Ai19YodbZSVUsslBvA1nDSrjf5khYjvcl8FG9zKMmu7gcTxSWbd1PmITZryzy/w1
Gp9LoS55Pap2to5enmw6DuccgtsAsMZRiKJEvOGnwBg1mrFVtcbphNa1L8Yu9ZEV
wLLUefSO/eed/YR7R+wwnGh0fDQ1OBAyQbSZ31lOq6ErroNYXCxsCABRt55yRKcc
8ivbKNKh9XUBPLajHa1oHcFxtXJHIeyIJg9jNgNlUrrZTf5vK8v5tzEaSQe8zRTV
lqp/Yhow5edISTRhjQaa/iT1SY5TPz9dNJ5EE/tJJV95IRE+UXGJk+HIJE4tR1KO
fS6r6JqgKkdtfazcqkFLSOHL9AevCYAhB+G3Lo1MJRowONrjWjsAlnYwLKlukROe
Z35KMmDTr5e4FTI5yhDNVge5dYA4BmVR1RRneOsKGhK/QwgOVcxnQaqGWYtAZAaW
4xDcXWyqrhRglI9F4kREq18elgQ53cTtn64n1nVWx3JV/NAs7j0UsKJvPc3pCrdQ
4CpjyKDDlWxyW1inFHwmuBEVAHvot14yvvqVpdHtIAUvwwdnauV/oDwJTUr7zwEi
r6Nikrb1IFtCQnetjWMOD+0NUPdfsq06Q5gK1TfX4syfApLYGf4vhJRVziVB5Th7
Xzw9TCuU039FU29m7I6uprVGksHFKFIBcOMbJm3eJbmKQRPhDbFGPJV27usInX2Y
FeY13wq87soEdL/xIAwmCsGipP8RoBqLLEs55XEsHHAdIiDoHxn5ABxNKvDavHQZ
JyeVo/QJcA9S7elM54YXe/t16WiwconT51COxPmch23fecFHKKOrWb3VUvwsj+ej
jaAZ+IAG8CPG8kH01YOxfCL0MqdoymKIjEBNfP/rR61OvXf2FgJz49V92YDmltHy
ZIT4aqjrbXjFoG1qWmy5StMuOhqoVeXAKzWJvv92B0D4oITQjK7SFmOfmGfoZr6H
tHoowELN7TILzocJAp2Snpq1djMrdhsfbnjmIVkdFbI0soR9FQEjhwZMcI9o1ctT
rMYzRuFrMtWnQOobJ2HmC7YZKbjkUYcC92excheXh4u9/apFen9sj0V5bIlHSyZl
JxLwEPKgoRlCpALYIa0u9jYQSYbQtc3tb+RQuPLFNRwGsRLiSaNB3TwASABzIs3y
KvfnRaPii2oow0RpZpBZrI4GImY6KOMrKSanrE08UFwmXKS3d7PSDJ3jLbVZLrHC
h8ToN5kBhO+71NVDEmAJgpeIgfR/n7AeaQx2mlwzmquEd1JEQKNmDFrmDAVnyS93
iYAtsNfgBLWBiKTWgvH8hLeZX6ZiZctiR4s2zCaw5kycTMFg4VGKv657LBYEWc7Z
qUn7IapbjprsUSyB3ScM1g2Lgtrim1Kty3u4mOt/boGviKJxxDWoY+GU7D/e00Bg
iq1dWt4BVxAf1M/ng0QyFGa+P6PUIQa4N22psCkt8zPNV4a0Mx2QT1/bSwbPkcZS
hBYOjL4DkbOazAXPq8XwsaLAtRcwAiKno3sUjliaBGlUn+Sc7Rm5UAMdc4hOuSpp
Nx8WWgWZMb14uLHM1kp3OrdvuLsQSLs7cg1LHp8bnMvMOWdsSnCSLy0AmXaxV+dR
ewsY8SLAeK1LYUf2v/Q8IM42koMNu9XQbEReSpdkmikpOqyvUvosYvLzGRgvrtWb
2MNH7zAM208kCmFtJ99JiqYvhL1Q/B2ZPRR/U86iqgie1JPEYCJ8WWNFFBZMBlfp
uLE8wUBmkERaIU9Vvy0no41EbLs+Jtgxxv3u/3XB+JeKAz1VQ/bE0tDGH20EWVvl
vpq7Ffd0W3RvPUva7mCHbDa3HLDlwbE19wHXa0Q6XDRBf2LEemp0exEWRw9EQYMI
zbGLNZujEnlToThKmDD+OQeICHVPtyx0k+d5fLcL3UwkGbQeh3AY2FlWtYUpVs3K
f52bhUnP+65r7UbaBVUh/yrvh4Hfuu2hCJJ73j/i97im10y1u0QHKWSiKd5LD5eE
8AGunaR9hvFwpMFfKLjaK7SayZMy633hQBZR+K7cIP/IlVvLpSxkezkmfkneMRL4
57+F2YAXZFQC56u612yS2+fvDM7+xI3+aSLVe0iM46/8HjAY2DG1wrchLMg47y2C
vOPgD4uRj8FZJFFTOIJzINBX/lf+3ynJkF/8VlJGIntk/7iPpPsmD9h7ZuRTpbOu
g+IGv41ODOd/LPkmb+1Vc2qJZooTfOELhFhQZjyTZ640LPn9RtO4Cm2pFA57hNsd
IImy6ZC4jIJRsN4/HDQf6KT+YTpq2etrayIaUeCHSS5x4MLJx8+Yv2XwLLn3knIs
KZEBWi0zg9O7asJBoD5IfofHzfFKT5CJ5f1Qbt5YfasrDet277IKuXKdPkhgWtC5
YjTH1kSKFBOc+QbmSU2F9//yXGwG3nzuhzbl1v/uHGZBVD8zuuuOhHVoDvIQd/S/
mT06lrn/QnUIXbtrPdxxyXeNmegIkGqFinr/KgYKykY6yShsKG7JiIUefBLtEwkN
XT3jAPHXsultrb2TGW4t8xIv4vWz9O2zMC/pa8KIpm8+tSdnwf9SBB8t+l1KY2YZ
V+1kDfesJKtrvckmR+PpGXIAbEiYtJKpRfpJUrug2InFIRG+PypeJCiX0slB58fR
lmGFQDkAoNcKGgoPp6T0OekeuHaMp+pYNG6UTS7n4mdZO5A6P/uxD/PMOZgvAi3k
xCP2dEyU0hh+nyIhkn3mZnXJFDGWFYb93eejEmHGouoFa0BE3UR7fjAA5p/Pt5mJ
cKsIUBnDbhlthbwgyErXiMmUGHUzRnuSsJjC0V4VCkxjIIpZJF1ifgCd2NEsz4Zu
iFa3MVagC2tQQuiybkG3wL2jDEGxoDXMjKiG5CStiV/GWwrMyMN6VtDwJ7t2yNmG
xPo+tBLvOOwrwYFREVyzZqLfD3K3+OzowJNa4kCtqI11xRVrZL/Ate+FytW6Fq+E
9sKy96qdxJbZ3o0x2reKLw1vSnXZckd2EeY4k5YI0R6OsGSJNPBuVAI6TlmcDrjY
Li1qH7kFbwOpZhf+t8/KRZkhSzpz50sFSQ5y19eKkZQVO3hSFL1GlrX7RInA3xaf
CNVqNMkMFPt7nHbcg4fGCWT+3mOzjlHU+nLHBY1MmbCbfsLO5TUsxOD8XtCgSUXn
vAHKqqHpXKLDcm+suio8lbIH/XuxY7Yk7qBQH+zqkpecQNzZO3mp50FzavlW3w6s
6yTgUzX3Yjc/ycflPH3qJK5xceo4BADEjvkxos4Aob49D2dkbfs6UAtXdns+ZMPI
u08nigoeIMZEwmZQWnqxQYy8ZAsgceogh0Yt4AjaYWHNruEXlZYQVJHyYWQUi1nb
XUn2GwITiCYFTeUOK/4Xpc/dNRqDQ7FcrcCacimQWF/YHMtlpNo4x7go0a2rBKNE
9P7YLYcc39E2v9H2NigxeF2bqdgcU1Yi+Uye9EG6to2D+CHuwJRhZ6WEcO596uL7
0PTHXkWoTi5m9GtR7vcfXsR1UKIkwmA+VlR14GTsBw6wqyFbf00rBpUA8Vd3pSG5
Ufaj+zYChbUMvaVcWUQlhrPwoWUKXabObnn+EIkru+/0rp/VCHIeHwYn0xw1HKao
fK/d/UpO9kfizoJwCXDfhJuAfKSGv+6To+uQ+NFUs4OSdXMpHhgZy6lgBAdB+YCy
F1D2Kxzr1g99FrKh3ZdKURKOg4AiABLmVVpgb95KZ1fbdxT/IKzOl/sNWmCWVZk5
11XkUDbkMD7k6rw/YNFohSbaoogPCqWale1hoDCdn8i4dGOoU+/9Hw7Gi1klcQT5
iSVTy57lwbpJuOaEosVWBI6UHLPih1py+NOzF94E0tAGPmbwckJDLzhm7MhZPRF1
Yn7bZyEtliruBRoBfIUXPOkFJPVBd0GQrVKmn9K634/JEjPl5aaBgorfPWYk+ODt
+C2AY6Oht+8cYyPfjzFW+vNX6u8lLZsOA0BXE0Zzm4mGnCUKXonBb2tE5/9OQGgP
XKemmRMGQKQ+HwCYZyhQGi6vQJR6B56vIX9ycJipBRaovTozgsNoBVWUj+1XSRA7
7I4RcvDCpXSB4CZaxAUs+N4BHxrIPG/Gb8gXuYfq1Yw+f2Cg4vA+Gl53tKO983Na
4akxbiAdS1Ll/2DOWy82rleCczrZhYJ9wXYDd6xqSVPCxePjxPQ4beMkIjNDX+wZ
mJyH6rxLpDq3jm8ltUrWcawIZuCnPRklrEJqPtmkYuaMwaicGV3yO8IiPN6mKBVS
QMuHShAoPNVS4lD2UMs0/PWPKql86lLrUyfaF+M6jkasQB65DQwOsFvdBKiqnNkZ
ETUYle86tXm2sq4OhqVmtM7HvvaJhFI2oi1F7JsSIHAG7RYCTpONkD30xjott3nT
vtaWjRgvMAFtCG62qHPdEvRK2cR4CgbU2dYkFfvUtrnKr3JsovKWMV9cBdhaEkO7
78qCldR6rgTFwAxOe9AnVz/Ikwg7cqeUKYRs23EByaR64tv8gW+khibdApnxyKtz
EYBq5/tV3sOGKaJtE/dg+9pagAO75jzuhB5r9I01PEOb31WpwIXyKHmGivpHR76q
TELqwg8CarOYhuzQSjJ7gvOmq0mOTIUFR7swX+Htam/7ydDGXrIEtrygZUtffT9O
KuMmqMGZM9l0TFDiXUpMLADDwGuMZmxg181VCGpHqY2KBZ/1nhahDTGWtdCdCy68
i0ipJeScb2BBtSnWCx4xr3FMYEzzzZFYVIKJZygzUz+5zgInP6BqrRqnFdsd/83j
aaUQ2JCMS2QYTFht23qTILwlRXNuJodDAK4RQEex5OZ4bE2AnqPgEBzvhmD4LpoK
y+0B510h2OlzHfd0/PoVqKGHO9Uw94dwBuHFmZV5AqEvT41rU3KcOSfK1VEiqP2G
Jpp4HOi3PYkTplSdWuYcp8gM+QVcpsJv6kb+zj7qmgW/OBDmwurtk+n/I5Twq5ll
t/UvKJ2orxADT33J/f/glOLFzoZdfMNs02mGF5IP1KFohc/zESjCtyoAA8vZ0fjJ
isKNga3imDXGIQ/fmyIaF+oV2sMNTx381Th/cHuqWEAJW88UJOYStZ94UGxF1QQj
FSYnnlBfv2ZygyTgkXReYNVUa77z0MBGYabJOVHY8D9vfgK1QmQtAJaOMunYMbPN
as/8C28OgPx6jnhQ4RUbrSPBywNO9cLDOXlopQXTW2rsih5tIXcHCEnqOLZnZsYU
l6wPVtQ2zJz42cmLrmQI/20tnBDUOfBESIZa92PIkAe0c9V5Jlz7XN+Cw7IWwRPJ
sXJFvNUsjUt/7ZwfXKbroqpMQKLCv+7EQqlOkd27ssvnQJqDiinqWo8hO+WZ2lJO
SpXT7H7U08acSQAq5DYsiMzE/nqGTxh2xvL/r5dtvwBSWh9y/dly5sVpcqnQagLY
jEey1/eDeqg0MwO9fh9PV5ChTnsWXZuYaGw7l1hLPKsruIlGnd1f3xjtg3UrjxTF
Bbh8iQd+7VOBw/FuMqw0+fj79omWtjEn1VpvBUaG4cp49p3dAPw493WrILxvowuS
7jQc8b5PZosPwxitLMeKAp+i3ZGye+YmP1G1WlcXC7zehuD/6nAvGibvZRS0vmXz
fF7NIeMFMjdo7zSm1rGI5NwxiK+/FsIkwlpvc6REOJms2xlQ0EzYf8BuVmv/VlcZ
jwh4qT4lEhJ19vZwxMLzXDe3v2tsZsEojOJ8sjzD8ETOpT41Uq3FEhFFzDc+eLro
ySQdcIB+fYiTu+0sNj31EP9A0TMWzrHbldkZl2f1VKMPIWYniDrIgKq8ntCydSpY
ZwbaP0YS7b2aGyO+SEDT5OSWltEKZbYd26C8Oyx8aklIxTiyklFd6PazWIdH4S2g
IwLUYhNTLEjPwKXRGi5rD9aeCThFaQOsCM1x8UELJJZfz0hHVIGB6WslyLi1D6++
jfb81Nk240+GWdFyeoZW+AAFDwU5s90qDKPtYX9W5E+651Y9KCnlk45kV1xAA8By
s8KgqsLtNllIQi7Hl/Nv3cWHlK/r90n2bQ2FHqgI10bf2baDLBkowdp9wedziVle
1WLgOQbvjiTk/nN0wp4pBvpM76/P3x8ktQB30kg2TksjKGjvmHpny/k2yH4cJJZY
fW1J+kdEPRx1FSDSFi2UhR0c4piOsaFzIdgc+Ut9gomeP1xmOBIVJdQ6dFjV3mNd
OkjAo+/WFvMzpWGz4DIJYkYvNGJxSSMLYl6KDsyqQToscw1DXCWDBo9fqUgtj7IP
NEEYtasPhOHMVB6WwUAJpQMNaCPMmJ9WAJik4YDhP42JLo2jLsJrErJ49B1JjINR
NosTGMI8iMdSYZ+jljF2xo3wDX8egF+blVSG16PDTtIiMmaqW20trc6xpyOWoEVm
Y12uPpJ7gY2J0sS2MxOmIfvKIj41OGUqIPhskvtEbpKkGeqS33xKiKHq+aO9V7oM
TLnkP7KdSyczz9NgCEXTbRqYT3+uIx5nkFFk6uRaTGofZDXMHaHXDmfHeDYCywSg
8t4Zcahry7PRpZt6j/DvIk6oJ2r/rveLt8xHy3a9ubeUU76oGA4Srp8Mm6/fblYm
0Mkl+H/Pd8oaGVexGLQEx9byJPa4F2fOq5X6nWxcFfC4UbNCFDpgz4cSJ9mm/sRF
kPGtI/cTdQd9wgy3NC3K57zC9DlnBfX7LOQT4LDlkSO0C+sd3lX8E2TGrDjOjAL9
4xb9qrGRd6yJNs/Aqj3J5AGMltpLwADsA0h1hIGG4hGFKz9xiuIJZKC7CZLMieUi
/u7DGqJSeMOP60kx3qamSQVFB4X8SDz2o9NPXhzk1SANP70fUyQtBQhI+BvGNtpa
toW4w1ZiDJrWLSQ7y0/QUqXpPPxy2FSWnme/h0a+fnfyIA1TpHzZBfSuM33Bkcuv
T4YyRcyYbBCrnk9WBcMORRj0gUIsDobhutqj+SdNNPuydjSSJeZNxGtzQwETqBgz
tLCSgI5pN5dmegyr52eZCpKgw2o0gG4UL44CwQ1gxxNNCflvDwav3XYkgvmqyAjc
joULQdOQshHlRtJToHdHMsdqTEGPxUMh1lFFWlOtAFQ1EwS5ZU0pzYxgLzmnDVsj
Id7pWwS4JgU4zE6IRqn5jhnV2nBdUrGHjItqRLJwKzr1Q3i9C8PzPgHpXjP48Chu
dJdaIlEhKEAs5Db9j4/ep3sHBAiF0HVKBZ1ECro+5joEo+fGpxeVzr39z8yZ71ga
/G2itweGRRIKHxME0sMFuhW/N1Ae1FNLZ58pVRi/xKfdhWlNH0ED2hhqGCqaRDE2
CxfjgJ4w0MU6YqGQHLdB2s8zRoGxE9vf8v0bi9T5/HrOJmZJcs6xgAGVvvfKg9dL
uwGwfkWqUd6hYRxodlUgmMGoBojY97ix9PJPEcy8cL1wA+G3SZ+1Xuih2K+y0mZj
URuIKjegr+AyfUonk0N9nUe8RfBvu3Wbpg98/18CPcVcODXsSxw9hQ2Auvg5hpqQ
Cjy4X3Waya0n/F8zFp+h22s8dmbGWzC3W+UNmOBfCzjHd5Cet6stkWN6RUEvfytp
tK6VkE2R067JAaHlKjtm2SiPk9F6vXVRy5EkMR1dW6T3jn76srsitCp8F9MR4KBF
Y3z4JysIh6y0m7Wz2OShOlXJ4uzDv9gzS6TSdEOZ93e8pCRpEYVq3p0Y/sBqgfBL
DWIgSbJsmNRCP/OLiI2s+ZIfA+gJXUsLJSO47XhNps6Z/mgO7M1SrkHfkwBfj6SZ
uOgYtwBoYlCPz+TIbo+/RkHftQa7fwKJygjsxhHHx5vcsswvgTPASPdwmRoxpqXi
7fDjlQ+k60+gZkdo1CCGzs5gsgojcKIYVP9z7i5aNricK4Bd+iczal0auLNeuLIb
GAcsh9zcNJ66rQFdKlxdlO/VrU4YvkDszaj1RxKz/z4M7XHm0+ppzq1uUpVFgxcv
LWJNjRVmtlwHKitGS18D1nzp5Pj0+xHOtAv4ibE0267V7DdDqBEC3/4J+XjGEAOQ
NAJ+H2bFJZH/a2GR/5QMPTYUyU9A4izHjqBLDzlMq4nNAlsdLyciL+DhIwXJNqTz
1qPM26XXZqyyLeLAhKQJza/y2KRh8OPlRYvsibMlLyhC+bBmWl1kuRP6UNmerI4e
YYBMzo60aE6PUloi8jJDtKzqx1nUtmEquTaErNWRoW41gHAnunJndgn5pPIrKzuX
IXVkMj6YGzWc25xhM/k/Rx/0tusW4EZ/7Dwri6zPA7STBc/noZl+SZT7vrhML69v
ti+Bi4jv3vpp2kDNIbdmUJQwsUn2yVugnaNU5ATjqoIKy/nGTxAAVLhbyErbTebn
hoqVmVc5k8SbgMvrXyIb4dgMQZHeIE3VwIpRhHaVokBA8aE6DJ+yWcHyUouby+Iu
f+Tant0iTK85G4HifwM/4Bc3aeeQ6xTS5nZWKkzCxr2sRpXyGSfX2upQAiSkS3GE
1JVhsHF9vHsdeNxX0vtTs46IkbR7N6a0CbWdWrtxj2/YldGSpsY7y4LeIjmlJy8k
jUTVOiayOyTbZifB/pA9kWGfp1/Z661hxDwBDiCkKgWq7B+FN3GNyFWn0myN/K66
OXRb/8a4C9nyhDs2oI6EIy6hxHrq7XmRKBfZ4Way8YKsdU/4K9VORl9KFcPl531J
ZfokLDGc/zjzQWHomx2nccCiuJAZdrErwQp46QVRrCbLA3R4/yAyZodJFD8ZmtYv
CvlZlf8DzpuhhabX8EoSL0by3Kq/jFzu8e84ke4ZK3bSpyhhouQ8nFLZ9jP88DmA
3/njgEP5R8j4AMVutoNK6QBzRDjzsqBv3vz/gdEimvf2+NYvokb79ghCFYYX+N5o
YHOZ1p32DZS0j953lBop6WviRVFkgKzV+yTJs/9o4RUSTTpoWWHXEcUxFE1XjYui
xZqwBSrdw3KVlKdpwWFFCuIrYZeYmaXFBWaVZfPVZVzxSREHYGK8h//Avntacdhx
vXMdo0j7UHLuiJYlmd+xHSn8GEKOmYRCmpkZxPsG57oRtN+u+eiFcpWEHllYLlbv
6Q5vf7zDNAqtn0suexgKg0m5NU2T8IYBUnDFiPHFmbzr13feEpyGXJ/Hj8j7a2WP
h0FuGYBvfqJSQ6J7+G5Og1om3J9+mM5Od6iD0jR4t/8t1d3q7Y+Eywas4Tpb5omb
THbnVUnX2LmsVGPvgI8G/8KYH5x/0tYseeCNRPdVj/aX3ScepBU4OYicqIzHA8mP
+KDh1fLNtBZ4jWRtvejkeDlRPOuk5VwmrloQaN+axpFsgICoIQxl+WqEDt9eVVm6
p1Sqyhq5cxcza3+teCd2qEWLvF212vwgb+KkRFHG2xFbFiregfulNxjxv7JzXMBe
oo0YOnZt5KYGUEFgO26co2K2mnWY1PRZrGFjTQl+sbOODCiLplYpNUgkn6szQW61
xUjSBSMc/iVcHkhTSiO3Hu9sDMxTz5ToA5ByHiyiPWzuYRCemyvcayG33CP6eHpZ
WY+gyVC3xyunwNgnq9HWoMsvaMb5X+QR9mXvoTvbMaZAAfy+h8+zaez+L8vNvbdw
v9usrV8AFyqHYcM/5/hpuQ51EEdRiD4ibP4SyJRhPqOOwLrMz492fxR0haiUVJjg
H+NIijIvwz9nUl5YP+jY7Mpcs3A77xBkapz7uGnwS6Zr8vG7tWol+NGZbk69GJgb
f+9T/lqsnh6/JSGSuVK00oY1N15tUvUWsQaRnwil5XSs6xUJnAOzR5qWjLfc+UGU
llhWtSfLVdYZYkX7B67AoymyOum1IKcd1WGhS7ZeC7lbnOh/M9SGhU9K3S0YhbNs
cmRJZu6KJlDSqiOUAKuC4dMtV5seAd4EhsXLKyO+rJIh3FF0CPaxlQmQK9gkKzMe
r1hXvxfx0XkaW4snTMhnwxAqRXqnzljywKCHXNhxWMNDxJfGfDlYEXSQM0Oqt7x4
IUi4f9Cy23Nf6icKb3koEcqbxIefeV33RGdyBroUtLs5VxB5FYwRTMevEOLfSP+W
LWZ/S7704bAFDImDv0mpz636+MygnnRmQlWZVF5pqaICRt82h9QfrRB/7eFZeE9d
5rTuXIcdltOUDfOzKuCARVJM8hodkqsI6qX9OF8NS10G9KV06GoSwaCsF/fF4pKu
PBL78pkoGn1b42Yg9iZvoDXGl95vsI71f6C6kWP+/HaKoLpzqFiuZSIsPGOqfCKP
yl0fEtxZA0T9BtoEXbYNENb8zc46QwbYUDpehZt4+ITgDIv/he8ioJbCXHqQnv+h
rpraOaURaz9tqB7h27542MB0E9ZMsolqJi0rydupTLbXQEKDxZ+cKxk7apd5OTkb
2wwfEC7Hd18dVHTeeQ4fyJkSOLRDhZa9Yif8kQvGJvwC89yu4Dq0tIpWV6dNQKwW
nukRoLPv2XinFvt4HvKs10T5ChOQ2q2/ST1X2i0koSTOS9JZd6hCWhEY5INmTndM
uPd111+eCtDdvYUtAjKyyBvx1bzHjoci4NkCC2bX37XxO+PP+Yl11zxXUvk8JZe3
shjvrQHX8usxi+ViYmgkhk88CGvrJQlhZ6YgqZav/E3AHHiR3NOuuN+rhlBi1xl2
D6WQP5sMRIfcXlfR0V1UXskohxu957QgtRAOCE0tnWLIDWDP5c6At7L4VowAIXup
uLY2bQlJWo6FSb8nFMYPDCt0YgGhgApLDmFIFI22NzuYU1Z05VZNy/kFfAgN53ob
BjV/yKWlNKcQjqbCLKts9TMkurHxQnDZWPJIfrAAbY0BiEXz5xemCLjbMflXE9+b
u481xFVC3txMnfZebO8/ma9yI2q/dLKYVRh2FiUbeG7kXSTJiq2un2F0lcgE7MQU
h90+5j9YRpbp6AwVB53auI46kRNP4XvCIBOOggm7/DrOdi+cHJ4X0NGKbzmCDpKL
Vwa9KmL54OxF7TBGTu5NXVX5XIietaU5eSSBV3KjV6Okw48VPzyMYvMvo10mkfZl
Td9p/imMUVJDiIihNrRnPfU+NCKstSXYl84yohOtmPcf0GhU8IdBR1GIOS84qMmj
yTonTPAdWaZ33JIsBD2LLeo//sU+oyrCQJkg00P72sEOSLqQbMV5mjchjVqT3a4R
mZa3X5KUvE0n8W8ANOQSakk7lqrD3NCMDeaN2KRVEMScNk6o6G3kynHpOUi9usAE
fEnBx7Kd+N+ieVQkvaLs/f3qiunVnWH/qJ3VDtINHdhg7Q2wiSYhLLRURFy0fdvb
1mN/cA4E9t3LI/DCWVcjRy6SihWoFOon4bN/QFF7VN1jzD0/H3l/5q0+GXxxEfdh
oyhH0y9957ClMHToO7JUcmRRAGiLHCVTBJ+XTtH8LKabMXOgUyeMiGydyMmbT0OC
Ohv9EDazAqTVzhjJ6KnY7wDmZpY650SRI1f8+xX1qvv7Eje33TirXw9CokriS9kf
r9R3RgKc0GGIW1CFqMy6PkNAj577Pt+2rIaj2Yi64EGh0lGlrEHiRmcQaF08T2dr
yUUN/18LHH/yfTWhLulquZFCTffDz8J0Z1I8zwkQvoWbLI+ZOmKnT9eN0oJecbLW
R0GorCldgqduNCeEQgqnAqhQeGaik/+RdVJ2oPj+2UWDzrF187wLbJJf55lCsu5r
vpu6m2cv4uynxsQqokNskuS/R1m6hRFOX/Uze/se6MPhQUnIlqiy8to1VDrOn9w1
tl1ceDnaWWB5QD+XWiDbKjZ3tXgcXIhgn8N4gkl87+/XZD4yJf4z1j01isi2ZfZO
z/dRrPkddP23EeYKcUaCwTgtmzM7iDcfLBM+NG1SHKTANNyv3KFNLX6YR5Oco5IY
y4j9xvIzegxu+yLJ78oluZiaPxPgri9tjziLkv6FkObZHDTTQsyshmRxClNRo35D
tT2LcoMnmE3mUYNT3aTy9fSw0BOTJ5iunPFITa8VAnC2QvtSSMkXtoWFSc7NyVxN
r7rXjOtzAf5M2K1JdrdP0McSkwquLZOP9g5ABkaeSR0t8fybb97QL2XTGZmfHlnA
Pibgyt6tcXdRKAawq+jhgNPZkmj+A6OSF92EzCXLA5Z30Bv//7QwrUHLf4+iVesl
hQp7yF9BbldchRfPrKC6gvlohHA5eHgLwL+q+E2/KU4blvct5A1fw6g2ZyecueYv
wIVG6SWIERMGjOSJMM7Lv3Ah/PhbLcGy0jvpPSp0Ht9ZOd7w5Iw6Yjg4z9lsPiyY
U7zo7BCt96wNOAkoyFKLkEomT/vkM5voRMyaImD7t53w+nXHbC6ec7QLPQJygGKD
bkQ60sfblwzrvnK8uESiBM4YJQE09Ph0YO9VRZHVr+9LvfMqR5vYjvmWyJhI3b/F
EB0ArjJWsiB6ik8y1tKoPa9NS3I0i2Zyi1KdSRug41sJRsEbEn/KhUPmu9l8vwLM
VfkqTrwHOFuMs1F3RfOUgL2aB+mETB41Eu6cjlTY8mtwhGG23XsjJdOJ5VQ4OsSz
LduS7uFFxp7L+3j61AFg99mEh9gvHTL8r/OwRhLIfyBEe5Tfizxk28U9jrNp3dHV
rThH2QG4lCjoR3m0vRYqwY06rKsdik/KqmRMYW41O/7I6zyx9K//XuwSYAhw4dLn
ukl50ZHzIGJbptiPUx5f1R908fqHZfitwneOE0IkP/WR//jq5KtlYFePtbMVHofA
dEOWwBmo2wWsbKo/wWx37ARfFuzTWIIYkVduvDJ4yVPLjz+4yITQai1fWjIr75Mu
3D7yHKsm+wFmE1esKilqfqIkMyocKcogVsZpgEntl6W6EePmKHmmAo0KmlZ+TtKF
FrC4pZsjfVQKAE7DWurt7RTKAic7EckyLZN4Hx6neqrZLWRDgvf8yI+1CgQhBDaF
H2b7yztRebF9fYlqbVAealIyXznUXqqffJpYoC4sNaWxx2aN/wAdy8eTIMOgU4xb
v9J67TaE10WD/59Juzo4c8GolYbtxU1uLyO+uM+Be2kL8/8NSkSA85iO5qzBmt4w
IWEqbUZBmA/ucpuHKzvA0m57WEXFCT3SxiodF6ZBB7Eeixxh1k8pZb/nPX7PF0vH
ekw32pJ2U7VxGR0Zr8rmusB+GlnXy9oBVpd0zpGhf321uljtMc5inL2QzdPmLaQ6
OWCJIvlgDebrGXTezKOunthZFrBEl7QUpVRIRSCtyWTsOB88SGAj67KIGjRohbnm
FlY2hoDFVYmWngwGEP/DTRAnyNKGN94h84nj0G3PUPZPJg/dZqkHf9kOk4+tlptY
C0pP84iK3WMyFle9E7l5ycSUxXZ0h/WWv2BzEwv0u0vxAVS7rdjLtnHAR43w25w9
CBm7H0oWztlDUd/61ca7Vx6XCzOoQaCkBZT+xi4cLPiNSM46CG70UREvKlDqXlx5
pSwmxVT9zBUmXnEg4JLb0FjR6Xp3A5kPYHMmTWt52Gs6CqmYKvexGxzAX85D1ezW
oYBmoRQgyT1i6CFOatRgXOB20loa26tIghXLm7vg4Y/u2JDMI/YHZbhni16hZeU7
5qw/VGU6kgYoypewXE/9DeRg2R3MrpeWo0a+0LMktx3FmNWdTIOCFByfpk2NJWHG
VIJpVSXh7MXiS7y3R00IhSUWdXPeYyvP7TtjYRPkl/b2lj8f6rHoC61nPzTxeUxj
sq34BVhcVWOKf18OMRka/ZoWNm65i2ra2Bj145Y4O7R/bw4i25h579kKgdOv7GMM
MwMH2CVDInIjO/wenViUxgm4lJX/UqdlBTyZ5AsDwXJ7XyTw/6R2qLrfO97HdtOg
/SQPkgFObRUPodOXHXFfr8XhZMshs8DR5mCxHmJc8g7/KrwuV7tekIH9UukuKAZh
V7oyVNaCa/9tG02rZLBcNNR87JvKd02CULRAStQal4cWHsFBMEYEr/26qDqdumeP
FM6JcHC1OUYbSuNWGioOZN7uVdAvXN8NqiT/hLFbSC6A4iqcD2xj/qxOsbyydN9t
YN+BDJRgq9xT/0WJDy/MkD983MEB+kq19Y2NAk5+A395N0FPU6lE3RBLtVml+52j
JgklIM5qcsKZVgWBPL4UkUycPaknBI/jcnkD5djQm9L2Yz1YHBxynN2Q2MXvEome
Ss1xqItADKFtIl+5FauDbF3T7jQaUZGEV19lySGvYvpNa6sPVPB4QBbAzxbh5o/l
xib40hUw6ISczxpgP74YAGDYo36XEviiXmjgFuMKyheRaV8PYAQcEC6H8wR2Uv5k
sl70y+euZxJwQsi5hcTvcPNjbFeJelXYEtHUmJJBJjqZugVnVAsl39MFxf6RvSzZ
61kELNzBOxWXXClalnsbRpmoB/b3l69ZiYmWA8GiCYxgEC9jgt0H+eFmqidNm7Rr
2fZpqrRkm4IVbbg0qGExDVYsBJc+3y9Yi6TcuJvD+mxSzvXu6bzdwpNt6UAXTVAR
5kut0QssbdDnU20QnIo3Y1tRlQ80f8W1weAqSQv1UaxTr08/sNIgKDygvIKVDJUi
lcXAf87JZsbg+nMXxe1zG6f27HsvQV4wGeVWgDC3fU6glWv9pR9sSnLcE/yvairN
Wt6C+rdb+7gB4692yEi3x8kr7TUXGcYiAjYM+LjF+QA9/tn59YdDZ6359C1BVN65
8P9H+WuNt5RxRjr22yJfnLLrEOjBXNiSu8lwKAjVXqIhHmXL0NqBrv+PwLki0+bB
RdUFeTXurq2TVw3uVWrDT+fqAGk5kk3RVAjAP2gsHyxyn6vvjIilSicDBV3awwwD
AtfdN542gC18L96DT0SLLjUI0ypzeT2z0gP2hi/wZ5qzjiu/FzzAiUo0UlbC185P
UoAc2DV6zeIrxLYdu6Mu1oG60vDXDWYKYb8IMNNtv8Ohcw23iLhU/BwW38XVNn0M
3wm/CSddbKfLb9WBF9Xdng1RbtM/cSM5K2LzTVdUSYb7MEqbQ0M1CMcxfU8wnCtq
6rzg5LPaUFyYr26ZXxOYF04jnDfb/giVBsfpr/H3LdHBnupB3arAwOE+XwFiW8xG
HDq5xsZZAfWPHhWDYMXqeJ50MzpbMewNKjM7bmV3CVvPsMdzlngtsFfePcUGZWUH
lBJYnGz2XJhDnNbagz1HrpRUH5xn3FiH4K6765KRsERLW0yaBntysc+LvSmQoPBn
Zcg07YSdA+jHTMv88fTnAkbbv70D2wZL65k5eN1O+TCoYwTmsg4XPXPl8XnneS+7
S8UfSKaM23bwn3Kj4KWNPldPyV0yCE0EfcfHQsR1Pe+WcZRj4Yf5ms8lcNTPubAD
2lo0LiIK/psGrzOOy5pvUAfui9ZqOdE+dSKzb4UokPNQCNe+sqX1cBLwMKPVf8de
hCln29gtEJh2Z86n02EosLDPl5w+1/fSeuopJGcbZacqiVnHBE9GoaUB2sJabH4y
ImHOPOPcPLBK7DFypR8HLcvxtlc1d2LZVR4p5p8ENtg8Np7nbh+24Y2WcntnnH3r
Dwku45KP6vGw+cTStzfxMvbarMDpkUmMILGteW0lTBZbz2jJyiZMvYbzvSslxxW+
24IrSbAOskxgWjI/QHNUr4klWay+QALe3KcCsRlvsYlgKt3AogqUUi3tCtFfTCvD
uHWNgwxkIUZZ6JtSWt8+og+y7atKEyE0btYdP4nryLX1KT75v3141Ba7rTcK5rhB
mCKTo+xVDe183pEr96eeHwI0eevZoGOHyzjlbkdECEGOZDDYcig+UAzNIq1mySv9
OviG0uAVJjyZncqchVafaHZVIkYopmInC0H7PfUOWdvRSlwJxWfy6bWwoJfwYUbX
Nls6eb1Qx1QCOJ35zXo/6fSBQ+McWQLvMKqd9sqRDz7/UFTZyrHbwk+N4UqNLRny
bdud7aAOC/6Wt0+PLUNXknvterOM7bcLQ+c3YpsuNmbbp9ypBPh7CZ+ROqD0FNeQ
NjScgB/AQPyVmn85phijGAxzzTYQLlfhTZWU0v7NIBnm0P/wQtcYgbsKdMYqh6g2
TfLRiz0juN4OuktOIyN22r1ERLBk8VPUZixmAAgGKg0HIUARH+3BvlH8Rg+tF+ZZ
YjK1XcQ+V315O14fxU8Hyo2zIJmM5kdSZ8ER768iRjusYp+vB8TwzyPAXzsyI1pu
PDF/JNrqb18AM/OKku/lX5NnZyzQCT0TmEhkfuwLINrgrrpDRS8VnXa4K5eBxBqA
1jS6xGfTfsyE/2U2Ae43umKE6TuGd7/rmN6oI9SwnTjYW6M46jsFW3QLevLapLzb
69mcxDe9V0lZVHXZmsj496Q9cf0CkWN7g2O4DLEQBgQrVHFK0rSpIY0/TajmOowa
yIQ0MW/3TshyXf/odBFC5g9eGTWoxiyClj/Dib2qwUdOqWhoCSi5mokmUpp8DdIl
fcXaqF6RLYeRUa7WrHt6vXX7K2AAWwIwIYME32b7MDBz1eYJmtgNJBzZgsWoPtUO
i/BSI97G+ar2QRMS6h46K9UwIEZoD3q3+AFGjlkmPxcvmeH4CMU/Kwz3txuWXrRP
Qf6ofP25CfEM1evT2h4ZUIFD/vOzUoy+iKKI+P4tp2UFxrHVp4ipQD+qUVWmRRoJ
7yBkV2NjUd93ZOx+kgU75vEQZ59R1x/baedPgQS0eG/N9CzXQ1vID93UYSx9wjdr
2AgReCrIKlGOVziBKCtbu7Jpfy/BTFu9mRtaIFqo4Xmtgza+1G5rIHe72t/Ke/+4
O5lx9NUsyG7hLo6Tex+mrJPG+s7U8Sc92RGTCkevfvE7kX+afEjByEYbdsmOYk/8
U6pcYTSGdOElldp7NUDYVVDeW/hpmfz/JB5N7IHxyA/amJACGGv+0RxwHgl5rALs
Pufer7wrZwlfE4u0XgPrJfQLMR6zZnvZw1AJbYeSuh9tS3UISYWTMC8hCCpyOQXX
jkM2C0oM7n4vfKAPcjT85zYJKr+eEmZ7qT0FaKefqUG3fE9z7GEX50I5HsFyJQ8A
mHWMhCqapUNtRMB+JDOdQEQcjD8q5QNURMR4gw+FI1mgOzDtGLsSQRzeolr3jBOt
0pIdTjmlXpiwpLEro49qU2ZrzWJYliqF7bgi8hA0cijBbgGwLAJufGrVf4OrOJDW
vL7iCw1cQSGkLiCQava7VoQf9C0tM+RQlbb7Q1Nw7M1NLEMSb9ChhcLZl4dGT4f1
beJLhPeL5doygz3MKgIXBgvvtbfVICO74JLzU92+sErQRW8UbEmygom7JyIajFN1
8lEaIGb0GyYGSZf3pgXBKz9PAsXa/OEYMw7YZ1yYF4xr3MiBaNSLIkGjqgAJgQuA
ogepPcV6L/UrbMAnumnzBCNge/B8psDWKVaZ3/pFsE4kVeDvAJJT8KWeDjGDtqCO
QKIxMe3JySUS8sm//3mqeDSglF85BekCkc+hND7N8bmWkPYwBlWJEAADSQFGm+C2
EVE4wk7NCv4ssd2BcJLT+ah5Rs999SuwybXx7g9/LJnhiPQzysrF1vID0dzlcqsi
zljsytDvCwaRwC2R5S2g3fAHgBerF5/QR3jUlen3hUi2ceuwjG0uoFkGQZoKSTow
Uwo7rFJ/q6Te0aQeZ10w4gu5U1iC1ItMna7NgVgDXxdv4QC8RkHv+ND6Ukt5H//T
f2iPsose7tPYSFdAQYdYzvvhHrLNfX0AZyl8cT90YKTbwA/qmFrCR3lSr045/2ey
g7DN2Of1I3PW18l/fkE009r9CLrwpgkGVz+RYCnyLl3mRf1KcgS8SBXXhIXutfdY
`pragma protect end_protected
