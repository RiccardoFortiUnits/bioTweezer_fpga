`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JBqoTEEaJ9Xwh5akotVEeNNZwprrbFl7TbrUeYDZs6IFqSOqmQ0yAjgmNCKWbJj0
vlZdNL2bLu1BDyeos9QnwT+NRAbBw1VKn27Yfn0LPVz7y1rBbf0Nm7A7RcHHozRJ
yD90YfpH5/7q7mvv3NBkN8p2lIUDowlQYQ1POEZ/nIk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18368)
GLNr5rZWQ4/XTKAXN/43kZgWEbAKa7qnvQWkbrljqqMC2Ycw06SunKs+M+U3AUjH
KTpNqXypKZEXUa0PUMC3etFSPBqupX3p7+T9cSEbzRu5k6laUl118/Pij313D6+o
i43XppCbvPQHfhWrIYqTtmDfXvpRdj+iIHNDR4C7V23hxqBCNiiHrFWrj+ynBQrg
plVKtTrgV0byf+qj6QZl47wGLsNqktiYCoAyRnr1EqHM04OBgQPBdk1sTIsPm7oP
AzG4LaY9EwyfllCnW3uQERZFy5N49jcKKR/1wSB9+QwiW9bhm1T/XDdczK2QPv3t
2j6XGDHE/ejmpk+I21uwnitENYgJzhnAg0rXAbMMNPXESvnCQe0UFZuyVDqrzPfV
j+svWpcJhX2iqXrIeTaCDG7FZndZkuvKud6ZwMizE3LgaTWKpiSS+se8KS9yoGfk
/g03VqGPZ2WkxjgsZOvSILRxLUfeDDuozrLYknFh+tZE0pCNtvEvuJvnqGV2IXDX
9PhPfwMd9n71aIZZYq0HEnthyyqbbzWEvdS4ARY9O5rwNH0NiyeJ06F693n4bpYT
fAa2xTrxeXQWe9Pq9HypkKqFZNhQtc0nsuPRw/oyOhkMsmXuniX1qvHsefzbjMY7
HfO/pUNRlW4Vl0ycJg98JWVNkBlgFx5migGOrAHvpeacdM6Gbr1eKhxK2mvyohDJ
LS9god1t+eh0LrcYyYxQ/RGIRZykdMWtU99SOhfVpC4CQFwSs6v7ht5b8j/VrOK+
yw6DFXaYfLN99BNIR6MvLLRShvL8f4ElAFXSGsycbm8dd9YZ7pJEHnSl6QgthzWv
Kf9GGugOIdhA+pEjSsWbg5EynEKJY6ehBYbf49ZdQY82HgQlsQFCvpT/nrzLkoJq
/RaGK1rxIcp3ldmACEKvViPlST4FTkPmTM8fvW+gAsF9da1vvOk9KiwAdlQkcyTZ
/jccfDWXmJY3z/LWjvoL5ota7iF1fraR10DZpma0J1RGerXCoN8b7F5OGF5NN2nT
0RbjjKrxN0iNU7G9AsrkyJh4ZJ/iJrpTag3Ydk0amPHbfov7evtjkQfbEKGdMvTs
Q//j676wfL/Z7vYqOYzuBpJu7vGkPki3tSuvU13zriBTVDs+0qB9e6E0h3lxBKQA
KwOWWfFECs1YhIgbIfT9XD0ZlRTKSIBH3RmmCLrX+hlRLvUavYedHqzV9P/PJa8s
qkjwOSvvtVmVD6EAKlRL6GWpZaovFmei8iQkAGyZ4fpKfMRsQXB3+XgybQuMgVRS
Hpno5zGNaKZ+McFabYbVwN5FyC0hmIewSJqua/8LGfvN/Tlxg8v3H1IujUL3O37i
Yu00H9S6jmbw5Ln89UvdlFhhuE/WqSqR6LoDI4GvZN4Cv3F7JYtSemblfOs42CO0
MLgCx6eFk3L4WtePag80N28lcr7lDQaEcnkvdd/eBpMUQthFpjyd87OGYKYfkVaL
ekvsYSxvkuHOQVuNvywDaFVEu3rlrC/2ho+h7rhQqDd742Z1qk6+ODG1+FUX9Zh6
pdos9NZWoYhGuzHHsGOrMqpsPu+vnr1SZuqxCsZ7YDYhvaYB/RRbF3jtl2ZHJzo+
lSJGOQ8mqxkPpQcr2fvPvJY5QXhPZABjhcdYOOPapltb/jOZaB49JViq1deUrzVi
PvdUx/J7gxYkjYdzGBXwf90vj4y05/tEzL5i4Ju/E4NBRw3DR3UI11KU5zeJypnX
V8zq8h0Eh4p5mOKHxl/AqTaNtE3WdW3czmqOO1ukfn3scrKEf+nmkKN8418msdxJ
j4uDRfIPlVVdc3R/X3SBZi5x0afB/0FdYVljJf7dRRic100ysaouT0LlCIE4mAq3
nFua0fbwBuSioIg6Dnj+PsSkSdsHGYueg7nFmfK4AXOsnCE1ZI1N2jcDc0rrgDbd
Km1+r2hv34V/anLunArvOjq0g4k4oTIvdZ2v9oNH2RqeJW+Lpnrpg1oHVVBY8o6p
erWugTADU5PSR+G9MSpTxGMcs+fswB/quw9RPIOSFlH4hEix88euLnwdUrl7ncP4
DEPgbuXGWhhE1onO7PdewJ/JtzpwXPNMPVWM6Vjwon4JgAJqYDUnBq6uSbYnKwfh
o0FggABu0EoCQwco8YUZhJdosYixwLAMA0Snm6rwQeEiW6iZJZVT/ew7hqDwfRZi
r3080j6hk0TefNNx3oQdBVOjMIQ0bxsZwtbn6KKnjJ+UnZRZy7LWWwp/5zGATnQf
lqnELHjIz7T8f763cnMhyrz44L50rtwv61X1t1k/AFSz0VabTFTe5GkrjU21p1FU
SMnV7S1gPf/koNPcWv8nUclEAml5ie06QPVHiMOANn8DlKmCTM9ZWhGUiiCd6TFh
E8nhunAhd78HVfYuJGHaANEA35QI+EBDI31spGXUyVfglqzQrJAOl3peGRmIutvA
fnxUIXzhT/VuyJm/icfijD8V9sWB2SfTxDiHzd0aCmo50cyZTCnc6RXQ3H9q/B3f
wYN1NThsta2G9UP0GUwM5SM0sg7DNydqdqEq/IzanO4PWdoPwXgF7LLuGnNQjuN0
MQDuNz71tHeo6sEicY90aT4ECs52Hd85OiiPSMtqo5SWbYg6dbqBBRjfb4KZbFEu
x4sEUefAkJrTwySd5t3HPU6qo0+9fD+l/HvSG6WX34bHrPM88W2WzFS6KrHyUCrK
2MKDL8Gprm/5+jOEdAW/XZIhs1aUard/0FQbaC9PlRrFuJa4gGkcpiv2FeD/yBOj
Lwz6gCO9842IMU15qguqTmJrbd1PPKiTAF9jte2q/3X24OYfFUULDJ5bNWklBiA+
sZGncH9mpbcWEcTyapz9gDRFo1PybiPT8DfwkEum3SOh11q6DozL4Cq51ItvTyVc
NYLWrzfSRc21UZw46UP7Fd+peC6pRAeQj5MbiNWAt5XrCGhkXljHkW9t6pWOSstO
addqa7CLLOIhs9sVQq3gy3/kTN6vfnBUCufD3c5Voem5FfRrmaKECoGOHBbMTzj3
zgf668SiNwzq18e5yMpn56g8STT6MLLR0eyReCa3J+2dFk5YeW5BDAWdnh7jF7O6
ZByOOS4ZXdgjNDPTe1e2Ha+u9vKYuyke4MfJg2PUy088OiURY0XI6B4TZMU4/zZ/
hDMIOl34ANezsidV87MMMV34VC+Bhk0XfvRe/M1r2mqI2FB8R4nhL/JbsIUNKcJL
K4VMvXGIPY9qYUc+4e7FURhaRZjZMcyoUbkpgZi+jkSTiZ7fuo5yippI+Cc+Z8BI
HToPQyiSCU1bqLV04FgHpgMsonHXsbCDKMsAIoicqSQ4H7AH1km0zyKRz9RCUqD/
kTH24Qj1DwydWzRNg6qt4XOIDVddgiwn9AWVdCrK8Y9r/4n/9vJ+ZJOQ9Jm9QHg3
gEAY9Sn6xEXnjsS9zPYc1eYMiJxLYNk+U4ch+mqbtI9XBFMeXk34KSm6Esaza5kT
uyA42akdvAUhujd4IbvBDMS8U/Ml+YoluKAyll6WyVvObI5R4I9cnggNtNAWBvUs
vkckLw2zgeRaOCOd5mkICT49Uh+Gw9hGbHb+tabCl4L5I6RBjFSapNJ8IH7Mf8MK
A8drwij97yIECPa9xXdf2doZfNNi8HhhB3e5rLuzES0fsOnhZm+EjmJqeRZ8E6yo
rSUpo20058v69Zsdp9FYKD5eq/g+youFFhj+iLC0vBM5OKH6l+j17Jo7VTa9ru3d
fnf2wDv3zyaeNlpfolPKxT6SCaMLov1YEz4F27SbQ23+kQU/DoByFTR6UzF02OvU
YTYILRwGTN18TRK79uPMA1ZPS6Bbyjs1BeCm1bk03kQJig6b0p/rK8ScIkcZTKkp
s6IHV0F0SeqMs0pbcrndlAbrbUCQl4lgOTLvjmXH3UGYzIwJmIGk+344+vX1GnHw
+OoQ2wV9LjoGzPeEN1YeR3tClXG2oRjC4IIDrT1+cf3luJ7NjAVlI404Gfinz3oV
Xcw66hmgn19PLzhgiAvIHM8kzJJMV43YzyARCHyxynSWQiI1jCESpsXnmao6ib/5
JV+yREVG356PHkpAy52aYSzGYFUptHVCIhlvkBTtxlt0PyUZUZgARZE5ROEBfolX
mL7bb7febKCofPW1dsfjwdEeLYmflSogRYHsP5Vm+KXLC1ssCVOmTW/kYuYtmv8J
RuiaB+rwuFAwMzS29tf60deXX9p6kM6dPQ2EMWcf6sr48BlHD25pc4IwdGjWeUmp
YM0km9MxUXsh0YMKu39s5IQZlOWhceD/taHVi1lG1mPbh+Lv91Okcj2gp0FHbLbp
HLU+ol33fD8HHG9cpoTpIv40Te+SqCnQyPTHxAygiBJBk0sa2Z+HU73rifAgo39U
I9xtFiWjE53MrmiiHlUX2yUKgacU9kHlDzvD8zJIyooHN5K8IUQAON2bSOi7i8ZE
OQfNxu1IljwXVy3+TTlaWyou8tUPkhc9BidyyXV07CaZtIcmUJEdVFQ3lOAaInsV
SyaHg1MfSgaXBJt8j00vdOCgdHAK4zGzFNE2ildYERb1qs2ng94/M6XrU8pS/MIm
QPIUNGZMyol0xHKu3Jk+l62ymgblLxww6I2I6OipnrJL6p2XZIMSLJ+9MqsGpDOo
ydVo5WOLf80zEpWs9QbLT09cJ7NO++12y4BBdUidETaDg3lCNAgvnCZH//kMBGio
YOHZBox0r5aZ4Y8mACDBvBYfarhkkQ8OmGX8Nu3MXbpzNT+jJG5jaFvuQcr8yg3a
vpzni9BdRg2h14c4x+9xJPAM5vDIL4ZQ+BQy+84ZyJny/fvqpD4VqCF/jFfs5w7m
i49ZKA9b6WqsmYfZZ9ew7JP/5NOGUyUV1QzoHLWZ8bJnKoaqMSYy1KKaG4mOHYII
CSLGA6r/wnrQNZ9LR5QTJo7DAmxuElPaPbBJLu4OfJlIOmpGb3rRHFoH4X3BojBU
yNYV4c8WAQZ+tF2FXoWI5NzUaN+igvonz6RYOSHpsGBaSkcTj1+lTVY4dyUxfTqH
pAr5oEX55sdUh+wP4CKJRJ0WHcaw66MCHlwVbzbpfmnRDz6y207pvMYkDL281HgS
aKaA3WxdvdruuvO8Wm4kZqWogFx9KhGhrJQcZvYJqZ7EQypYoLBlTuentvpr18BO
tHvZLHE6PH6YYCglLhoeSXBhNJ+JTAjXwhNGZIwrPdJOnT1DFQOEkP5d90j+Hsy+
KVyDJYrhdFTl0FYWC8oDSgiiKHtU7JJsvH2iCh9On2zxvG6pTYHhkiA1/rF6Xvke
kRg9Qxbj95lu5XNszFEHxplzqLnhKQ+QjCv2lz+JQf5vVmq6M8yHxVW9nEhfncW0
1g95GZEnJ13WsIU53lmB6+71EhucFHFpvIc7Nt8NfDQSef3Yv7c/gvxpHLpGNwHi
5IKB54zw1oJKf7rshnEAPWFxLe+MCj8+PlBDmpUWcwZAqn3y9ePn0/BFOjk3S8Hh
XSvYECBvsb2mDlqHgm7m6bx0EKYOGetELrdthdmVs36FII/bod+39xUCpRUr95iL
jawjt9CdEAqIeKtbhcQT5HP/S+kis0EDHmxczD3XU4mIaaVRRQFS+ekerkef91x5
VEQOUj55kOPuZWzvJDgRQfb5AX7fzaPeF4HSeHcWbByutUd/OjH5GhBQGJ34Y88w
H8IsaYif6wm60gL4CCv7QLuo9EIRbHI3a2okbJ7ts5pBcBba3SNjCfXeLbusFnSR
jp9YwMJjjOB4VWkJ7pyiJ7oXqgc2L8ZivMJctqlBAtx62KxYZDBZ1v45zgV/PjNl
7LfFnPm5kfKv2GvGdjKCbHnrwkPGFujv6iVVXHzg+Pn929TwQsYM0UUEztbyfTQ6
Ny4cG7yIs3xX8m0jaLlGdCZpKXAc46xzMm75uIn7e8dSAGq/s2klR7C5ZQF+wCZ9
krgvk1oFACoACQIVseuiUgwLHYeEChT/9omN5tgR8W4go3hqhmSfuZWSjLAfpKxj
kO9wcxj+l7LQXxttqSVjoIXrHBuLvYQ+jXFYFmDNHRpfVr7ogN0hLpgwfBKIVVb8
4CldF3wi2kACD7Mo3/dFWu2gJL918itX1t4Rud+TpWDwTERYbM/tgrHIPsNHQllt
p9y7eJqv/yUpG3fKG8cdhCeRq64Vh3DdAnc+RBpDUrZZ0ILkJOIy8m285ZM/zJ99
GifMzRumT3Z5/hQxrhoKpEQWJKNBvr0ubTLmUbHY76mXfJkbLLvZR14Ul3vQxmPl
zY2ytBFAQwzYo+Ncg4aQv8ZYCH7oqZOCy8XsL8h0llN4P1wrc8kNUuGaalCFCbls
x1z7s6ecLLix3xXr5El5PI4lFuA3gLHhULjFg2bPdkezt8mV1oEkayBtxftD1ykT
TG2Kw3rbqnqliuczi8rMs4AER2ZLTRbGdA3CdtEqwBQhEqr+fuj+pLlVPxtJSXBR
ETAYOCs3gweLGcORVEb1ncJKHGAonh1hpFIZBrIFNO6Ol0Fjp4If+VBPpJSGg0Ja
VG25E/ZNZUaHl6Tb8Et7PDctpIRsnSDd49fOqd0JyT8i4In9Srx8izCMM0qMjbFd
uH6Khue/VaKI5jmYK6OrX5G0RkwkOr50VzZymB3pqOPgRgOhtbemxX5aQMlt75Nl
+HqC+TavdyN7TRGnyhVjQXECwESPbRxTlEHy2Z1aeH+QAyWawbvPHsD9+T2HwQSb
xvXPqHpH1HcaxyfJs2Ho71vlV3xfO4Gweg9ucnNSFtgKCfp9OnIy4Z9Bz5V8jbXn
ruTqOKyZBh5v31dyTAeshJYiEP/rdYpgPVlQw+4BPKoR8LDUeJH6Hw0qm42AGOT5
PTzuwxljzXucfODNboeIkYnqbQ5uifR/EjQEsCKEaIubiFvL5x21GMrvDIprQFhO
Fe/pUxTcq4qYxnmN4PaAbKl1I1GR8h+3hFpVzQ4v+WDuOnvNKsBwd80OUkw4mGtH
fRPNzwPicUr6oIZGWpV22yWbmyUs8inYcHCRhS3evS9Pyi6oWAJQan2wQnNcvBG1
+WC1duCEw2ACi0M/8D/dE50ya2ZqZ8D+VKLbyFzICvcZweLf9rSWMsdHxRq/rw4s
VDt5e9mM2HnmwyWmIv21HVCLjFU3bYsiaZk/hFowdn0znM3UURQQicq2qbVIxzY5
OM6dwdctNWsvyIyqW/MVr9wtw/nmstYvu7QMpkwLoHPmEBBEH2QmB4bNB3sjRjmW
OUNpCucJmQwOhb2qdqp2sJizyemP6QeYXPvmwX8b2/+zVmy2o8Btci3HZa0kBuKD
gVSFYlIgg/3mC0NzvPopAl6eQcmc0pNg2aj1unuF6AqdJjnbNbMBJgzsInbnL/S0
QJDkXo0o60iOhL2VlNkpNALmCdxHb6rB1XPDnpjL8RxevFmM+OMfHndbYjVu5cNo
AwL5kLXeRCUQq8B3d6noS2luQGUqfTrZ4OXVdt6U3IfsALAVtUszbX3mgKV+0n3y
Kh5XTEGlV65Un8NjC+hKG+JMWplnbxsVMH5ItYyc2HORAondhJXB3DAsYUaq9wOD
fAsebc2a4iWYzlSHLw8AE4dauqLGvVC8YDBZpP6U6SyKHjkvNYw6W8Vw76ju5uoC
ZjdQpXGBcFbVbtMt42nuNlqovhk8OUU7Uiac+5lcsFVb0MjlhG4M6BJfK8XoYqTy
KtiCwBpTgfsQsgSd7Eqj3v/q2rygoYJIiNqLF/pipd3ODQRx0e4KD1Iew8M8DFNg
DAQ8Vpgc/0dStxNMa1h2GbkAZrc0NMbmcrzvGEUgmRlA8524C2O+oAqKj0X04aeC
jEZmwjLeembvw6DOMxa5oKIehXiocWHeItLjvYMxcWjTePI4wnUV/iqmPTaBjm8Y
yegp/HLcYpFAXH8Tps90zUTIlTWpnOqSH7GQTHq2ngR/vhKI3fFQ+ZK8c2e3qQ7V
GnVoexE+jHO3PC/CyR4IFfQwr8XvcPfsDwqE/YXXCF0uZegoVrLM7dsTLgBCVM91
JcLHpOYAj21UkB3h5l0xq5uOP+GZsor40snRJpMZVi32+L9c35it5UYEv7xZUMDV
ogThLUH8MRIYS3eSA5lsrGjr0h2jf1UPENRpuqZZrO+aCxvrLrzSw9mFZtGM5vSu
CmEd4sJ9qR4a3m8gNjkb7OyOsWq6fRCPB0++yjJWDk708WfxqCBsuZ/TnCzoiE2C
rq7D/1z88LTDpp3oFCVaRI0VkmBJTnJa9Nqm9Kp4WnspXwYgVYWZVAcnZ+4+tkH3
zd9iXTh73nJXIvzSXw1x+E41msy1sQUlJ+6e575x1QLWW7cG1E5l+JIhFC0K+uJ6
8mIHMGGCA0VRECeyQVTS+uHU1++cKHPe8vzDMKgtbixdbb6vrf43p/NwqevQMlV0
uUUCMkWxq02BTzFfWFaO7ShBQJ0GCoOEsftsa6WlY2cOlgGsa9ZyCmAbo14Fp7it
Ow2/ukuepFTPRtmefMDLp49O7ZX/J2/RbleM0xPDYX7Ob793KiNINe65XKJX+dYb
pt8ZhE/EWdnvRw0gHcQ4xkdpllJs0Czflv7i5JV43ufdihAhRFd/cNCH3068aZG0
3mmz6HtVTcbc8LLO45rWMXutcaOIJf9QqAcW74CPiMKD+xPCtL+ljdIBaNm3W4jH
jQDcHLqlZ5lRFLNO0HBdmg1gKUAsWLX7FDurnSMouaUGewPtLivfnFTJ7IE7L/Au
pJoFxkX1nnj+SZeKeThIH/7puDHzY836cGs1tFiuY4pr23cds1r/bZqdqlBoLqpB
6EXYv7HYLJWQAxuac3ovwllyrv1uVptP8PIIDQ+/78ncQD/w1O0gux2GPnTK3SrD
RJanOH0s/4Qd3TodKNTEu5K8ICVPYlGIphYoy34FcpZcxBGtXifyhD1vo02U/f10
9SVbk2+wYxO/n+kuWd9V+1nEv24XLzmGQjnFEascoTnjQn14iqxCwxBzAiwoj63Z
1S4KGNzdgRoSNRxFc9Yb2uRjzLALizfELk30SMWoKulq0+yLIPsDffHBCJ4y3Kei
tQSE48Re61jgI8FR7ntmAlQJVqOO9xdLc6MqWJI5wYusypvO2Wki+xWcdetfFWq3
uLWIcDnKI2VFevvnlIZtLfxyM6Bxo6ckPRycpBf4Ol8VxcymrcCgLK2mPfURddQf
qfC9lzxXt+/c/2/t43THI8143U6LwCh2B80jWcKoGsCA3FozE3wYXNe7bmuXBw+O
3TgmaONWK2xcI5FNfSWqgmFXQdvatJk/yPVfnq8i56fRZO3oRLSiGNCq7sx8VqdJ
REvoI4zFtMojMUE041AvozbZd0xbr6PkiahlmB65d/17HB9MhfdZAcxIEU6ts2yt
j3UMjqIljkdOhO2CMThSuJUIsSapv7bMiDQkVcQvW4oJjFf0b/lFMGxPAOjbouqr
3/L9G3Q/3jDW3OSBD+DiiVgYasTzoYYf1BoPpLW2SeWyjY62E9ceW2BaSFODvesk
0FgEMTaWOSXgl3M84Me3Xf8Qt/UnADMqgS+7ilm6tYRDMm9fJ66Fce25pwSIF2LS
wAAhPqb/Ibh55mIvqow+StuqFu2tPk18jpMuTEQkYD2g/FC/hMXk7sdAsQRissib
GuVD/m6gKNsEsOMvHxvyrgoDr/K09SCRU6npKqUALDwFGaQCuRYLadd9zX2iJq1C
muWzJ9TV1f2l3UzbjRMaqM3XmwOJTGSEDw62AQMNDaq8QRq7wVbMGFfUs2NuOurQ
GxK+jkY6wgqpJ45NhLzVPc+ml/g4G+23JpxexOkeNLvBMxdhN7USvZUmqvd21m+W
D0aB+3rKS/TH2a1p8xsIVtpeXYfxosk3Msw0t6rXWhjuBBpvMs5SYQxALGbGFEb9
+SYmY0honGZJy58if2nyNQkY73dwSeHFzxvd+KQXkOJ55a1nTxNW61ckhYb9bPyH
lzNjAw74nkmGllCKx54SJIJGP+5ea1S94k9OcASIw+EomQkB/aI4FqhMIpFhCOwA
YG1bTJ5JOMh53XChGopJ30tMC0wCymn3MFSVoWtgTwjDGugu0SUwz9S8bkGwasRh
PbSY/1XsMIgsS0L3d3egwit8AyYsSepRw6XDjdI6EyMjURtF20n1ImfjxP1x1I67
EKLaUDPsAd1MyXdfGrlsF7er4hxzcRW19On8wGd3pUeYNLiRAmIW69q4buowB64b
XK5B2igG8Hw8afwdufs0dancX7eiZ7o5zQr152yZowy5jrI3+yhPDOcDCF3+VWRe
64lTtSVlB+mX1bt2903b/LHwHZPAR74HRCk154JO6oYAkpzjVGuICMoVX+6IOvqg
iOshYa/dQ4HFZvuX/TKwLy4SL4+owFd0VexpVdWEvSSuxNKF5+2XTmSzwqdQv91f
Q7f9Kyfujblz7gYhL4RlYk3eaRpO1lr5WK+qGOhbElYLD0qXJGiUNOP/Uo8zbLCH
v7E6Rl5LKeHlNQImW0tQDBansgvSkzzv3X9YURKXyHoyYjPwa3CDJzqo/XZ5UmlN
C/d8WPVzEPL+GOIzuPfFgi5Ae3Sp/T74w6l95z1ahQD0ozfTTXFlMqMN3vAurjG0
RdEUoYVbQt0b0ZjffU1Gk3Rz0oEmNIWftHddpYd2ejrGK8o0vF5OBrJvR1K1ivU2
dD5WaGu/y8fPvx6dcFj9G/s0yLRdDf0wP4ISkbFy8vwxtja8IXVvPcV7PatzQtAQ
mvY5Z21nJzkR/Zu9km1GGGEk2Sz/FNqdlDnzefzfB4//RrH/cbau88XJgJDrTmG2
BQcKNh42Glk0OQBHCQc4R4A7QdSA5+EuhyYuUFRJbMyiGxAG/H7WBma2Q6fO2oxJ
Y/vqfLUuUCnVQUS7b7T7GXpWowZJjjav8+U7fF8XpIgsVN8s956KWuxHaI5ZCjdQ
zK64VcEQZV3geHJWt63r0QC1q9fhNHjsniY5eLJ3nIbPVV18b3GpOMPtxFEY9A1u
jRfspZ9M9WuFdoQbsP7C6qO3csNDoVoM/EmKrEoI2obRGny/8QQ0SZO29+ucnM5x
Yzy/N2vYsnQH/gnHllkzM4GaW69wyckF0sgDq4PhdnWO+MGDqo/yEn8Kr+bdFtDE
k2bXb129BIdimrCYrtx9YR3wr/OpkCSzX479VeaaxqNP9pmehY/cy/m2eNNnPYdi
9mTVabA3JTXoS3WAEwIr0Z/zWPmnR93wSKWflb8tVdTni30m4t0wirQXwNhlaHX0
/ORVvydkmveMd5TBZsoO2rl3TCAazvfbF+JbB1eH80jGVP9MNjvN/uvg9ZcHX42K
LBY3ciuFzN7+IhTMiFRb6vumDvAw1tA5Dm1ZDDOuAsW2p63Xn0rk3nIFWlp1NN97
ZayPEKZdVG1p4UrIuUaG4Q6/XPNfBjJrr3rcxVEIYT3nQkcg1FpJyHmRU56acG6f
EttF+xxMCH5iCj/Z+rIjYTbC/8x53kAff6uqd4zdiBgbJt9of351BibR01P3CfTG
C97QRgsi0uHRcPoWXr6gwOlBgOurX29dU9z9XhWiswF3f2R1sTAgMZ4yml2YgUXo
eyDQyT2TiO8mbCgad71K0mh6CMYObmp45T/zpffNZzgk1QOJrR9fgzHv9Eu/XG6j
L0x+nZjn/R9f6znHzNLdg0PJyWoZhsUY54AWn/mWnTW/+lpBHCMwuOjPj3xRPpfe
43VONPnDhgkuy3wyXDn/YznPjZFBl2+60LQ924fjGQ8FvbuWc/b7XIe+Y3IzgSOs
CbiKIr3+osgBaEjoFqcAUOE/s+f3uzmGrNFI9lizCvs9RBJp6jSx10GAAYp1izzT
eAJQyiEixfEeiTWjfvYXe7lgz3H+s+ZWvj5N3GboXUDLuIrE2eHofNobiQ2wvRZV
9F9hBgHnArDMRsv4TuM9U2EAWPv452Jjm3mguffiD57mzHPr4XGBM8BPEjLcvhSW
47uiHapuGVivkdKMcLLfUoLuyJhI4xydjbXsNgkjDSAoMu8F7axNqh+ooX0UUYJR
uKh4KpgtqpMapd3449vETUyv7L1Ykt3xYO9AEZTXjIbTPZrHDSbQkkQa1Ieki49z
w5k2lanx9/iLFlDMsguAMA/oeJWy2oy7VHsocxxdGLF9N2eRIfJTeZb5bZGSS0Ui
j1WHOFaEw37I/eyfqN819zuO74+4b4ZXn+qZVQGJb80h0qUQvitNDQqNjguv9ZDE
9XijD1N3Zqlj4Z01prQBIWD/bI7QVWaC7H57fi+NGm35flr7TLKLaE7tV0HO0pDK
fLMnoGUt7AHHotda7CjhshMGafec1UFr4EWXWqSnWv32UeGNcLBE2JhRZP0FySo2
RTjxMnofKIhxZsStzTy2tFzi0uImeNvlGp5OW0w6F7uE7y09RW+E2kSp+j0dtRBf
zdz2/ThFo3KEnMJRTE+L2r/fgU7Sa4yDlVbLQS3r3DnN/OPIJRwSR2Qn53ruF1Yc
zIbw0QUHNdek9fMkn6K/9HgmqJKyO9ntodm/oFiJ30RUAIfP+x3ijP+ZE7N8glXm
8ttrcKRioasPi03g94/NxD12+fh3sxq98STa5IXJ74x2XPNsTjYWs8dF8Npq4GLQ
BBuVWV3H1nErFt53WfmWd56oO7tWFjfZboX7/GMBhL7alVA+ZSdBo91V1st6d5RV
+m/mCcRLHU6LnCDfWtRziyRIqXX/RGDdo45KC9gds8HwU5xnSVKPXHSVR5wMkGhM
k9nAiXWn73zgCAa5HdOGqK1DUwiroxK6qprvzQgsuqYU4Ad2eaICPmsNrUtKk47R
jNqdA04Xqrl4KXsmRsEDAehyQC7jxMYyzjnTF5H6yp2+Ta38TvfCAgGmyiauf7Cl
a7+LSJ188tBhFOIlcX5n1IeeilPYtK/wPHkji2UOoDsFXRy4sN5dXhcA79R8YpOR
OO8+BtbNmK4PLklRr57UtXlm7yO5VxbDROD8lJqcClQwJ3+v2Xwa0jeDq0e3ChC/
Doh/Oz5s41abMdS8SfgvFEQCMP50GXkPZj7KjtQpCo0cOom+nwupoj/OI4DYN4bp
S2Mm3f8hM6gKn+ItfUz4E4yxm+zt78GxUI+o7z0E5chAOk+YoKcHiaB2kDMjFPqu
l4uyqbQERsi5w7fanZIhXu5DNuYIlsLOBulKm/MjIX7mAywF3VIfhoSxpkfgu1Lq
Nf6DPRtSGq/o//sE6sX7h9VqW3xOV3Fae6AczuYXMYMKiLRVTI/H5XT0ylQT8xu3
U4PzkOMyxPKjF9GS4rk4qejmyQWQ+yDuaLbzWyuQDL7yydHJpS0aS4uNqTvnUnMr
OBDGPCuVsihjPnlvlXNYZE0OkuC9Sb/GZie8RLeHvP214pYO74Ik7YMcvl6Fh9Oy
znZ39fM97OqotNjMw+0ADQbeHh1/u8nlWVynDZKXdwV9bPmUEc3OtRDTlFaGVxen
Utoj8WR4aR8OgC78fjfkKdhqdzzwTP6sjL6UOAUtwa4QYiZvfiaFeyvvEkv63RpW
sT2N3KddFU5ggrLH2ixaCUyL2+C5cNLJu6jzD9qS81FpKDJcjMVkuZF/Kpa3O51t
orSFvt+U7H4P19RHTixcJcVdmOVraO5WN6HeS/lKt2JXH5H80snRCxbT4sjQZTTS
PbwfPxVqT9ornPdTWAfzOWGYjkp5NW8uiKLl6dgOsr472bvsO2lYyhw/MGBGzXNt
wXZKCNiHaCilUtps+XQyTNluCQ2Pvky1UZa5Ru20Mof8CfaJuObcM8lMDcUvWyuO
+vg1VydOqMRmAmUqYaReW9V764O/XyROlKB5EofOa6/UXY0yqxqKSmlQhBiFnoTS
CIwGqiwngZMxjEehYcNpGquXApYGkNStB82yUaQug949VIaPL1E10Vt2jZNzdj1t
nq2vN/W7SfouI7reoqB5Tj0WkWx7tNSmfCllOewCXII0Jw3T/GBd3piotoImZco1
gndDowdzwXLZThA7SpuepTcJTK8kKQgFFO73c3f0QYPVtF/H3edZs2na2+TIjdlP
PhbloNcyozHv7Jvrg3NeUsvkD8nBIfgr0PFpeyKqJDPIqu1jbgSYhOSgWaQos51Y
+8wjeswI2m68tLNoGx0fqvg2Eiz7nV7OX/H9DIUIVuwx59N98ZbRlTmM1M1PzGmr
aJGsI/IO2PkTzr6ZH17JsnoN3LCfu37ksZBFPTYag5YQa7F4+bQJKL1t0ujXHZIn
fnioadFvnTxEJUjzALQJQlwuqICU3wKk3tkgKAOikkCddQuQsoYIKGExsmX6PW3l
82+jJiTSwW28ucCr35RRNsS5kyAbMKGXOrPbSurYqLkp8Buw7tMNi3NBa4X8Hzq5
94RVLsA7QiLquyYpw2WntIWcnC3PmM2OQnpX/jEYXlpLVh0ttyRICm8bTnMe/kmF
6xkIyRfvdTysOFdJoiLqtDxon1AyXi69Mbi/ZRno1yWNaLB3E4O6dpbxYF/NW97F
+oFmNtoVsrXmx952s1gY/m1Q1pFAWPuGo9rmZXK5s68EXO9vQGpmDmWoIbAazdoB
8UrbOmSCGgOWoW3sh4PllpE2BwJVSNTTk4gpNI/D31CmWR/ZhSjCYXPv23CisOme
nPTXT8Vw0pvtNoByOtNc9l0p3vVL9kVrML58AZqC4Avil3spQrDWYrNyJojMugED
62WNprS7bZn970Pv4XPABAVByOiy7wHERO2ktYWqk7LlHtnaz+CCK42c2xT/v6kx
gcbuWvNHda/0avYdwNndPa1cl/yxG7KEwzCUnZomUZp+BHomVUvmyS4Vi4O0O9eF
/mBLGQBPthyWNsbo1bDnFv6xOYIQlZ8BruVA6FjKFe+JHpID8iAsOCBeafeMvCKb
sWuIF9U2DCkgsbvMuMd8GLECXGw5YCchHa7GWLCx80a0kyGGSmITe3rEZOsVmlPM
dX+vHDQbHJqh4Ii+zCOoFhzN+zAl2DfeHIbTBzCB7Mr3voF+PJzRJBG/wSaiOlvT
reM9edwqQ3Ub3EzzJBFfYrCV2mhL/LVkpF4C2mloY9OdJEDPm3vgzFfv0LdcIq2i
5bjK+PQ/VYdDA9YTiWVU2DECZTmlzEcZF0huWxRcem+oUoeKElVtbCAmp8IzhTqz
FdTak13WjGnGq+5WyCNosgbeBVAg6E+Weq9YhBz8dA7tvJH8e7i3u8t0d6vi4ciy
pHMyyzH+BsAreIw31gqEkfx0h71LNBKdGfxlDP0kdmgKismatpE9NZk2YMXgmyQ9
N07c195RDEMJvUqO0QYiDJXfKRQ5qbu5B6sz/1wvCcdUZn/n3PxyThqhw+egWDi2
vPusIuA1RC8UcIsvwg/yGtQs9Uto7uzrsAvzzZ3fLmnmM5JRTFoCm/I/5JWWN8Rd
t7Zj+LRO45tWce3LVTlAIz26DEb5Hh6bHnN0klvSdCu7BfuChocGu8Os2M+3ooMk
ZrvaMFf+PsHLlWEluHZwA67EtwUVq7uhRN4k1EX0miJG6SKCpzlVILjVATg2TdAo
aLSQKH57omc3W2ZPKQCuRK15DRkkBjODsJhKhbywo7s/nK76JcIIEJflWhD/ZA3Z
UM2j2tC9d8v80Zfw8x+LSNPm95I1Qs2RgPbiVyL8+lTTGqfoya2qZhZFHFIR4GNl
VkbOpKkNeYx0HmWHRPhv0No0S3QXdw94Z5nD4EtOlymuZg1IhpclTEZxlyiPIL9g
rPbI5TRhpwvN/E2db5u8yLIj9k08VeNuobqIaow5Ae2sdW63lvff1Fp9EZplZtHa
PTTtjYRBImdjo8pOnuzdLMGB9bOuD8AfbE0LcuGwDGTjOO5VYqJx/dKhb30AgA0z
jvglQutt4O3xFJmigEH9VjXwmJnCh6Ss2bBF6EjNfXbeFe4CB8qcBSH3BJvYZwrF
xWqDrt2UAsIBO4lkfm52C1K/Gney5pe+ESV3OiHP617MyiGaAhnemixJpMo4EYzi
9SQCm9Nua3b+DV9hVAOIpsbmKuUjcHCfCvTIBIiDsidvrDok2Ad6g90AOydgNE38
8vPUAqy/KoGj2XYqq9vvGzCHWBzW6ruADdxNqD8IsjPTKjL2q4cBYDVTaQ9wUJEs
Tst3B4F7mbsoOrHczLr81L4uzxNqj8Yg3p0aCdoB0EhfHOzxo/hjh6ERrfmHurpS
MHAiPWeowcCUjogtVn5WXLaeuhRlTwEujB78B3xFk3Ejr4QUdGeFo9ZWeAbu7JOE
B8N0pMq7mt5vrr5zy9I7bk6D/ILS9M6oYcEVsXtzoJJoqvBiE0TdZEQEeAi8mfHa
qAGc792mI0Vtq8Xj6lOBQvO7GBh5RPFEuxLWzPMHXQ5LSlFrA72RAtMI1CBwzW0M
72g1s5HF1A1BtoJ9rLoaIowAZXAdDfTNqVF1D3Ipzss3e0KULm/+m2pAi0wB+4Nu
+Vp09b3RGVlVPnQ4BLcVeaSxLM2askZqdjKM4v23tcfQB7BXFqLzi0+eWETYB/Tn
dIjEISw37BqLwBwVPUxgWIu4Q9G6i6o2pmTtUdKhktUpl4uBJzeQIdiSqjLNZQ+A
ua+Ja9DZSvd0dIBrv8Z7qHzz68UZdjPgjzty/UyJ26r9e7B6XmIQYgzhT3fR/wGw
AtXs1aLFoGUU6Pb3SsL2xOsSJq2DCxcsW2eKz+6Drcw+caZVwV/Abq+2vLBXlPUS
zjLxPN1rjLGSpRmH8/IppGimX6AomkgrNEbBeuUDLOm6a3gAXQy6/NAILsFwAGP2
CO6lr+vWcEMCRfvfE8GJBCJPmtG+qM81gviXwJFIaqWjmh2XT+dQOMnWUbKDFx8v
RyZOlm4dFil2FR2OJ4FMzXM9Pi2/1K6H8Z0hnJciKbt+R4OH8bZWdqnCUiNZD9k3
UsvhVYN83EeT7FZqJVBHrzF086UudlmP6ia9VzspSzD/lFS0lcmSQ+Y2ArsrhTB+
y7x9I1WgnX3DVrabyLmtZUxi2B/IqCo0uFeLfGPW6plAEYdHJd7PIAKeH3IVI4Z+
qSKcPGAM1e897ptwMRBmVOCT2CJN6VSrPFfn7tj50wVG3s/i/SeV3uz+44iWKDry
JDSwFCU54nZAChoqf0ZJGlh6DY/E87t59Tw/9/Ea/EJvhGlfucaQG+9c4gWPRS/c
I3A0eiyjtwKzD6VNAA17uE644HIUdlfzpKejlbdxYkGl+ngOOi4lPHDUBzmb5g+Y
jOACLgz2HE57MyogwVacOaIgZhQTt48E9qtmmd9qVwnQwReOgFxuYevsam922mN+
nEtBPKKT0pTH7zuzaH6QBcE2XA/+xvNb7hDeOYkXoQj786inNJ20lOGroamguk6Y
kMXlmynXiA043ql3P12LT12r96VXA6fib98qYdE5Gi3TT0csgFuTYGAEumDw6A4K
Xs72eTWAtHTorjuJKkOXdEbITWjqraHMhe20xZDkdSm2XegR3n1sphH/vWJhztkp
PpifDYctKiTj08p3QJpqXvtI1i2CfJ9+8GUp3YQBZQr5hb809rAPgXEFc0b6yKD+
sjMBbMiur+RJSTxcQLUne3QF8A3UC+0FACp3Ap7LgVsLga62alMO+yTl1PIf8h3B
cCR5NHTrLG7kkEYtAx+Rdj1YP0bNOqX6szIxaB0cAQrBfI/LY1eajO3HdoHyoXlD
GPf/8y0bx2RaTffHmOQXgkGOL0UZbaZ0lajejRGg75Xb8Dt2p/a/PJlRc1dfGECQ
jjlXJg1V2bEEJXm1CHgoOPZrwIOLep0ScCbUWzFMfPj6Xk0W3hZCraBzOlzzwwQ7
cvAFctYjfFWMu+ao/Du7ie/5d3umYTZ7Lw+9PWCWKUStq1Stn/TjQxEE1FTsEbK7
xqU6Kc3P8lNSKLbfE+8lO/KKeOYtgGIW28Ifmdx1kSjFMxI4Vh8fRUWjuHvheCap
bRP5MS8HSCtifeS9fe7uaDiHefu4+szfXEIXUS5qTHTfAxFzAxG284i0miCJL5x0
Bp/K0DD1Mn0x+5auChkIwKv+9fAGX74O4KqXRVEsNB8V8ElNmmzvc5XjCkNW8Gbx
gInNexzWJYXpRFTfmCyV/jasq7yEo+Kv1frKpUk94U9FgY9uh3CpmF1PZEHRYlLx
Y60PUlsk3Z6kduS9GRwO1m+krIdi9yla0JI7QU+RiR4pwip8XawJjNoSFbkjDD3V
trO0ANIaeIEGj2Gsqfcr4brK4+lg67upN6EXJ7KkecoTuNfNig+8BhvEJnirtbsP
Jv2jYk4NdK+ij/rf7dktzLFDjye//m5vTas/AByNMHnalbjE67if6Fi1W5n9EqrT
lqB31oDlgS2Q9ymruhfyk+42RNBLtgiY2oGjGxLSJkvxsx5g2uU0epHr/Luq7yuV
8Do+XwGVNt4Tnz54sMlyWGjHRbf0RdGKhfqkys2WqXpAGOjxZMPd7BKBzu7EvPY+
q7u5LX3q35RU+jZdfag0OEO1CkO9m0weQBAUL+OInwy9LGd0+6hooqSbh7XgprN4
PNL/oDJ9yYUhEFjKPIdgFp4Z+AE7M3evR6SImAsbhoJFSfyI+VtTt9CJioONQ0lO
msfhNeWLrs9w03B1hQ0qxXmdOgrt2Jviggb11edzOWBIsf2/L+aHYJXDH+HMiJW7
d3IjtEzjDiDbF9ippJ4zxGaP7j8pF08IQ1RXrLvrABZr36txcdvmGxLYxUv/LuJP
iQlqdzb9de0F6xs1xvFWT/zpN++bP673ByWNUmWijkc/mkkUwpsr5AQ4wvKfjQSp
szcoRHHpCpC/ffHLmySDxnRk7r99bh1ac9cuLmVI4UdSe3rh08P9qzmAry21gzwQ
RIPktAMWnSL3g3QBGyd4zvxExHUffa8Upgn7TQkESsBWodwAmOrEEj/LKyvwqVsE
R97X1zaXzAZKrePVg2cp1/S6psL9sVvsnu3/5h9SP0MTXFJjheqgmGTKWawlbl4U
rTpM79Xr3F/ridVX2eloBfgDekAolfGcDfwULdq1AbawZjiQsttELi0gBLeFLvGR
iEWhyveL/UIGc0DfT1oUSm02rHnoRHN/3nietU9sNOR/shwI1nZKBRTyopGumYn0
Wrvn0QWZREP1x/pl3m9o+oDqd7cD0C5bMpGehMCUktGa1Xp6oNLihZmZQ+G7Gt46
zpshFLejD5PtotmwS7t1Zvhgckart9Se+xrCz/9i+wamRJ5Jw/WOVovVRrLNx9B2
qzdQ0BFnzCbWPn6UkCWho8bnuR047811e3Bte7kwlWDhztt41IsDroSRq3JAjVPK
KVZyPUA0rmYASgpkNgc5p1Tni1sNMiMxY/AHOPx1pWpAUFqjYm3Der3sZdIaiC9P
ND7SnS0dDRbzEJqHmQb6e4VCJSHuc65AWBRiOVSxDJQF4UO/IMfucRAjD/lEmuIY
evVBzT2XaS1yu2h4lCBnyoAq02AY34vp7cTrrzhSfBd5FDD9P5GIfGd+KkxfLlpt
1BlH9bQVsZIPSPyuRGcsvpzl84pO9feETS11XARkeRrbCz8achtawVUzNbXYIQf8
Qqs2xAkZpRf4IVcukSxBfMbnwoZsRxrkIV08hUVdDeVFarqWMiRmUMFEpkf4aSfM
nNpyLRbuIfdaQU0S7Yno5/RGBwdO0K4Kar9I62SSwH5vehLc82mcd/2b8YS5hfhi
S/DXS7R1WUn8299PS5HeyKvwBGRXtRR1TWhs+/F+HpaGm9vJ8gQ4T36BfLFFmTcY
qA7hv8kbbO1CoUhsMNbIc168LzEhR3zMMF++kzj3dmRWzDLJE3pdyfso3tnfOyZ2
J14PFiMwkXvNE1d5PsM/HSAP91mc/OQXtXhv6xOb2MPnIcOWVZGMF/+qbfIZkMME
zK6zYqM2K4SSQ0VZ0sR/YV54skUwhrtj+9u3JVLS4A1GZ1I/CtG2O1Btnu1AAq5+
NtiJ7FdAUDdHMHrUv3kmusknyv2AByfPIpjCAr4K2z7Phs3I7uALI1n9leJ/dXAR
py/iA7YXSJLFAOzAhLoRKlu1GrdZp1tG29RfmTKUPDnXBO50Gk5S53kVXsZlyvba
IpQaBHwvDfwsQihp5uBJEHxdhHBo6ZEP7vipH01KuZAJp40+lhwHvAZZCtUHfH5f
bS/TPhwMO8omoCeIIBtQRm1SalnrDLzqXUXV5zlfJhj07u7+p4BNVC+3idlDCuAz
9ud7CJ4REYvTG3VO4+LyNJ4dS+n9tPhWfSzlorU1TZAk9Bgse6eufsVJ1Os8h9RQ
SSwW1eMcEXxIYyUVKPy8Ltf9QcQgImcwb2+SB+ltP5I/iJ9JkoBTHh+Tfuahn8gB
Gvonk0DKpKiXoBXPT2wmDUIvsrT1L2XUBiGtmRaXz/sqaPQmnNbLfsgT9qETn5cz
IvFfVuwPlI+vl+651bjl5owpJ1BFK/4KjqVMo5lzwAXdLm1GAIvn6qZ3VVpcbj8M
RAWoqJbhKqvtJG9+nR4vFm1TFWyfJwBDOPKAMClyHjD+BfuEyuPAYzv5wh/koTce
a3kMp7vs4XOqafrJI3kcf8oQHcmcO1C76pgvn7Sr0XP7Isc0vcU380BsdciZJvus
JbAGpW1UGmCvPJ3qEFDD5ntIJqIy+OfCPloOdhSiuxuFmxPA4MtKQUkOlrRQdbCM
TBoFeIfuVzGs+M0ydkcpf5VRRfc2j1X9mbm3bCForIPHqYavp7NxnFn0INYX2E7c
ROisG6aEiIQeYZHn6dm/aHBnG4+x7kK9Rc07yigMShlBUF5UWmU9E3I9d1iV33+C
QYINFoEAav6jhODQxrzGvZzQ/QaL8lGBADVkIzDPa3QjKJDGjJrnE/YhAyznfs5g
X3Js3gO5Ri8gl/aWrDyCkVAgd+ziZP3AzLLBP4Lnqy52H5CPOOuuPcQfNPbhOvF4
2I+MJuZnIVO5nayAbc+WU5bO0R1L8WXMwo6b4/ynqosTFXeDTjVCnyoV32LE42fw
6TPGNMIfc2yQlPLQ+KnjVIazwsZSnPBTAmkK6kwttM7w7k9ec+W96WTQ0pG2AT4g
sX2ZbUn1CozoUjDmakLdup+FChfM0bmy06IySicmQfEBnJLKXwmnyVxFRbhugFUz
d1E1BbatsL7QUTdYjIszSTPAiq05Ic9s34fADEHyOF/sz0wzkO2nXoEGvDOHIyXA
FNzbA5Ty5HHGwZv7MJXjZ76GyscAPx51EkwutiVw0UNaTGiFj3lMJUqPF81tPMfU
hw7rXHtZ+U+8ZXTaTNaEd1xHNyNvKsphGrWNEetpOYqXlUhIKlbU/ooLKgRJy8ib
CLsHBTSaisxgFLmkr3OWHNbB4NZyolm123OCE717NDOKEBaVTqO0n2hLxUVJ6l+s
0KZjPTKMzUwxS3XxoJaafGu5JZ9+4j3o86612+BrXTlepM9ZrDgQzZNnNHfW0++9
BaTtD1w/e7a+flANFV7wUcNCGJJRIY5WwpKBGCUAg035zmzS8PEQGhUOXsyTAC7h
osL57Ncreh8fQ/lrnzSmKejBPFaoiVk78k+UNOry4wkieKpdZz1SMhFsiMq4WDEL
wx2OTNgtvGI4P1dVunA5FYXPUZQ1tJBpPSkrcw94rCnD8CDD3XwDD9ItTHm0UOQd
e/H2p4GZp9oS9Mx9hCyOTZrSZtYuaMs8kC7J6zKF9f42yzB0OuQOzMddSgnmdK4c
seRqZ0knxYve/tdPNPZPY0HIGaghx3n2NzoXSHbHiEjSzQa4R8+Hkk+je66I97Of
gtudroBQi9ndUTlRA11uI+8YDOFSOWZwrUhpSp/xtYJYI9Ngyl5f8D4EWriXyvPn
saBZq+sWDTqE15GvJcF2cWtpBoiezmHWBd4KXNfFK64nB+XdnGhPxPX20nftDRiL
RMHxNxNWe1l5zXvNYArUjl8QXjwLxIp6MEF7IvPCHrsubIY6L/GQsaBIGPxFwg2f
dwD8UiQGCoIbhRB3OgJc1IBi2rtIScJieWHVCat6CTq9yxenW9R3oGAks5www4js
C3s4Ja4AqffO8+g7B0pPEBJlE4uHlWImcafQ8nGE16dshsP5cHZkXmG4HuQDfWM/
IgE7GeYOx8TyVAr8ayeycy+5hzPtICXUzlerP2R3xpnGI+p6gIy6mOcdhtPqBZCa
9WKyaAl7fGcIjCDCeTPBNPv7KCVu5XL7+ZdVTwthgcnMsmLO2thpmKP+ItxQ61P4
AdlPH7BUn4eQxfKSzlv9VzfbQsqmYQTmN8C09X3gyjpp9tz0qRRe+nGupcRg8qYs
2hADBVFjICvLqUNqT9LXfWv72ryIICVsHAzYZEP2PTeScIPrV84T3bCSZ74G4yln
wwzDKfHOXCV6+BFKcuNtrtMD/uwsriJhi0Hs9oWnkavad8ntee0SWYBSz/Ie2LnW
+btFqhQJnXrkRDPjl33EpiVas67zYTTY6yaOtS9HE4wfb6ejdeWAkudsC2I/jRLm
82R5vTxDQJYqA42s9PEhe30xnUNFFyeOiAtOtbjeiG/u4O7yXxY8p+rrdFOttTWb
VNxUl/LybbPD3d3f7y2GEMvAK/j4IRwHJqvZ+aw9Oq+9vpY8nJn9E/pZ4ZXpBFxZ
F7WrXLlHmulduWM1yJjlgwaybHNthHtoAHI1Kd4ehtaKlduy4KGNJMCvte1Y6qYf
7tSX7hmKywqUfETnZPuHie8VUcJMRXS5QGNgz2fBLIsagpnkIRd9zJwSfb1Dci7D
mq+LZWHRf9NzWh8F/OSu3T0I/POgbGa0SYLHEMCnIWyteTVsvQZJtn3Rj0/zWRr6
OzbBxuSNIPNhGOdynU+OH5my9A5/Qt882yoF6QJv54Fysh1t82NlJzlUvRlbrEFe
QSGB8+PzeYx9oL7yE7YGEI1dJX55obYmrTdvyjO82Sh/seNKAb7tJNGKU7rg8C9a
tBCWEBWqAggoj0hYu+GSeeKtvGFTihd2zS5Wr3R78o5dfBBplBoH0WKbpIlD+RB9
vbzn5pd7+XjaTBz9ZxQvjW00C9etiinulPmxie/lk+sH3anjrx76ZrITDgQphgID
uniKoSEG221ZZzBnQA78d3mG7I57dUeCKTAjmqWgP14V+964zgoLJf2rXhUan/4k
1YFfPUGiK+N5n9MRQkcNjuPtQmMqinrKUJ0Hqn4rC0Q16+rKSOsusSmjRZDmmCaQ
3FMFynfs58aQsnCaideV9h2QR2/U66ObTbG5eNGcOXJU0Jmxm2vHIYCd/4SshWNJ
w86F1neIzv+40vzDOV3wkldaxW4blCT4N9oVftVmdjTWPOqQeON/nREwMfpTv7fQ
znQLt6y3bqfHQl3WLEGudv4l5LRAw3je0EKojgarkGNqgtW1JHgNhrglTKY+Ajeu
ccenUpKsj2SdUGauIMGxht/KM6XxUaUJO/xHc0xEkVu1SBqBPHSJuDnpbSmbD+ze
g7Y1+i4X1c95TmT/HElQqUQOLBdpp/vWMvfjT1a0Sqs3jOhknkJcfEj5i1JLtAJD
EettE9Gp9vHRmJPEg9Ho8hh7BAw1BV4dIe6tpxOhBuY37aZO7MIZzY+wzXM7z1RT
wMOozsVIdJ1yjrQrOY0uMFKJF33KiBaSy8A85pT3vJfJMZrovs4+iSYvAIwLtfNk
LhPI981lpgtcBi0luLVMfajvY7ugTWs6uviICjmwifLdN7drZ3HgtySuZKAvDWPC
wmnMhymkvhFXcnRdvSIzbjraqG8XbWIn9DRvuK2GFsIDZe9d6enpf8iWpCG1+mKx
na8ygRgw6UKCiPzsy+oQfWlm2L6BysDEpQa1U/hB7eneYEURNSJ3KblvoGVMIX2I
fEqAYfJOCA12bnt/cRrvw9Inr+bVWJiEzRF/8Dzvk4qF+Bfy4x3n5SV4t3MGfwNr
IoXFbI8k3GiY00Ap48j7Q42yJCElyzSSQETqduMvHn7Y3ZrRU1MdKWn5MR8i7Fs8
q8XeAlje5q8mj4XDG1DZltAnsQB+N66+J6zuuGkqsxF0RY4GyIVVo7l1eN7wfESk
8l+u2mFKHS3oEfIe6yC9wsxFV5UFc7HrFMsC17H+/9AjbqDASCsNNYzP74M8JgSc
9KtsQZMALswQTsKshpZlmwZO7LIJEulqDDISpoC3Chca+G/AiKoiAKQ/4WEqMuKk
1sOLhD2Z++asIS7yYTHGyHEpv2VeQeWZCR7ksybShdIX1ggRZQ5rMtvaEUlbevLO
bP1Cjw1vDJGS83h/bksLZlXpWVJhcLJdY0cbmOWo55yckuUfTrED7sVVq1Vv5q2j
35ymhw9KvHITKdqqIt/04BNs9FthnZpif4ggajbeOTRh+N2HXFp+4bX3CyGzagG8
bC6/FJ80+1OczNoHne3lcsbOVsdiFqyYIazZjA7bYAeV2imvLaW4hdwh4aAQ+HSP
YNtpUn72KC6+dZ5za5KkAzbX3bxbx4oBbtH3FJj/9snW2Oe6JwAZrEpdqOYReb00
hfct1lfdDWTR5OtY3B4QXwe7G4VY8mFZdo6HBRE6+ltug4WYM1DLkP2O3wrIuAqS
uneR6w3R2X39Y0DNYVKZiiAM3+DwmlybEIU4QJmjpRiNJjMm/ZGxZ/VBMyNYBtMC
MI0xC64hE5KW31gWzxDYNqZHcqEn8LciFt7Fo0OPJu2JH99s5ofSmJvmu6sgW0bz
t9F/LM0qvnxzPZVvS++9kgvluaD4N4SgUbpvGzwCjxwJis3x83uRRJcuf4/1f3o3
ltXfXZD4MTSk6+LryOjExWThtjW8SS6A8EDvMD6fKyo=
`pragma protect end_protected
