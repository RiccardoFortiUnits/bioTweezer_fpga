`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hx5TGztkyrdQ9xAmvUjPX0X4REClp4p+JAkcP5k+0F0MrNGd9wYGlEWUz6FFnhNy
iOarGiv0qtdIjxiMwtCcFsQMVAUsRkaNKViZJcD8MVrRS/ExpwiRLo0R5iBgx1a1
afAcshLU6+yk5bDpJ1LhNdodJxZWWbyIpJBuiWnhRco=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5280)
Fkjaw0uw14/pI0EXReFfXnBkosLCkeh79S8AxzSxOLstBrTQu7UKkNnCkrwpI36X
mqKniTfLSCtAp7z2Hx298xW/OUEDlqVUvhz5DrQ6U6+b2kIHiq/fuN7a2WMeuTQk
jeNCUlqXzpadd12zpWopsq7oWwtrOvgvKAMGgQa4bHAZzJsXAjA9uLQCG9MvV/CO
BIRkJNeLGDPbxxYfr3QR68OpyX5VNLnuNTWjhQGuxVtuVRWQGPj+US7ss0PS/lrA
A+rKlVi42uYIlbjHE6X2OXmA03TjjTxnwVxwDw+HcYbcSC/tUrNiSKd/kh2qHBwq
kFgz2Av37OB4yXsvpV0xzdPqDyFwdeCHxwZOL8iR1/1oIpith30nqKO+SU4A6rzw
/evmC6N4bBvDLm2xbkzHEHiaLyuO7LZIAC9WsmtTuQYcFmItguwUuxN6EA9J8Vad
+jFblYPI6gQ/FAQyKI3zXlHmVFhoyldDJ5JjdF9DgqW4ZpDnsAnT8pvo6ik0FEWd
EWdobf8mrk1ZQQIhIWkty5LkUuVjc3Ft78aEjHzVZ/FmrnzKQdsByjUw03N9voUn
QbW8JEk+2jY6UFWK64K3To/Jz0nSYWKSvK7y8Nym3kpbFyAPaw8RQltq9Gl2nLoz
cA34OltI5C7heOFqnX/6sfhhXweZS+BngwcJpciINI7ZZpV6n9ww8eNQnqoSoacK
Cb60mlkIDOseUL6BhOrrFBrMWLelpdiQCdM/jkHfvPWOUbJ6XRbU9RdhQGv5MgM8
Jv1FEhqMhjINLpshYBHtUrSZhi1QK2nIvF7UQP6SZ19/jUVLSiXgQbPQGZO6a2uh
q8Ogam1v8727FZlxH2fkJHzk8EdHXvOIJxej2LKV6XuK38fh+E98EAXs8YJ6G8RH
A0ePeaSx/ELj/wa5KvPLQe1lLa6piIOazFcv1iHVPvBtMJ2DcMht9+undPRR03XN
sRBOJXu5BzpvA9kT/FSBi2ifiL9URAHXiKxj5zqQjpNmRYQoYO6tMDsxTHPRsCDE
O+VFyIk6/48ooPMPmik6E320HRPg1kQQ7fugLaFWNrBFWgMsVnik12q/PrY8Jp8t
ROXRudstZbGBs0Xzsbsk9krC7c7LYE1JohOIl9F+GVrhybS6W1N1XxvmsWmYYUT0
+tV5GfsWWOKWvdvVp86qqH2EWvM537obJ9MSfwo1xcHp7RD72jXJvF6YV1k2i6Dj
QIlS/PHyYHmzXjYOlnRlzm06fVSNrpdEAChVF3ygxtR4V5dnQIAPBb1Eye1qvcBq
77/WV7qDbsfFE9aLmR0wVnB04DU6mdKA9hU/zZw2wNj9n6q+KFWcxnxPgny8VCp+
yYZHgBSSK+iXvb+cVD47WxOoE7TWgroRADc4K4pTfMdTT7UNJwQbOA4ozeulXrt0
WW/Pgufg+7ZkFfpGWhxi+W1E7NLc0h0w8qpA/WqzRA3M8Q4WIdqUKrAJG0BYE7At
LfvKyy8IgS1Q9G4sj4qBsU7vZuSYQqFPNiA88v8/FYBafjTw348IfJ0LSw3nKBWv
R3fJjVAE3nPShp3Sc8US/Q98PotEDG+z59n147PIGhjGlLszsK2eQrxtgSh59H4o
j6WVxRqz014aNzoK8h7EsOVCCEW9unONanqoalsVU7aVY1wJ9OMX4yDhjRaeeMFW
3UrCDqZFPhhNG+bUedTpn/Ywyt9mrC2jG/9C0ZrZYUE0/C/OOZ0YO8n3ojG2aijA
X8oepmQHX2bVmUXy2GX+vCR2QIclNHCzocYr7Yrbmct1PL3oRePvgmgF+UKi47ga
UPG/PRZCGkOPj6kQyQ3kxO3tjJL+Y2Qu1Ji5a2MGut7qaSfQ5CHWaqownGtlCEmd
frssjJjo9qMdG/l0g0QvETUAKQLGQ4xOW5CJ2bXTyfpXGeQiwVlCXx4CLuRa9qTd
FhOd8GchmMVm/T0wjhYzF0JU/vP1y8CMZkasvtEml4em36EQdaiYyP+t6/Yv6mfi
N5EwOftZPByku0luiUvKEhVvgYrZ0LgsN96Xl0irHxGtrGFB+kUomXcW9tjtzWUs
oZ07XN3Paaw1gMwVBRAWZh8DQJ+ly8A+n+V9HSQndNZSaJq4gRwncHW0bfGel4J6
6VWqLhxS3X+dGdGus0BdhVTdymNJpXm4h9S8xQdxywZmcvyd46rrW+j+MLK/4NAu
g+2YDu02YwwVxsWZEssPH5+mdJVJfdkMFeAz4kDuFe09y5jQfKN4JmsTkZXdTAiy
5pcT7q40NjEGGbGSGSbMFqMv3aec0VHaih/EXpbQ5HufLZwiSWDPB9IeGhmNWxu8
987QaDscJXO4GiEv/xFBkuKzriICwuCv/SF6ylZen1jPVSAuCWiJ2ij/bUXc1M2J
M8RL+q6tPikaUVg//Ip3+C9J4oB2JkeFW3gosY/E5X4oAEMe4N+qRvbiXSkKK0sA
3duOvNsVGpsNtlFOCHIGnmEqen4nivF7mGpJ18EkPjNfh+nAEbmOn9/z3tjaA7tB
ltIl42JydZlWwp+ohVAs8m/tj0FquCdFLAki36ls6v7o34sl0twOOZ/qD+6Rltzs
E/rtvUtPhpzNxJ/c/lo5ky2nJPJWnK5k7ygqUkMFFkYlnilrK8O2ELjDZL7OnUnv
oKpeYfRw+ibExtDuwdcDoWDMKDIi2z6cidmdSDtE1jOPgg3RNkBEVR894cgH4JRt
rPxsbVF/SZ3Uq5HImJnVIi/JR7ZblL76FOMKyvim1Bic5TUc29uqNIJ65fLzlCuP
Rg55ZbMCSc4hyxcWzGhkh/JW27o8MmWvu6RnnPhC+mJJStzKgIv7j6r+76MSunj9
5NcX+fPG9YL4xIWdvTiYhecZtDkymTK6IEqGNiu5W6+cHUMq95QnePpd3tPzCL/o
6mEV4WtvoabQ3LTkZh0Rn9t0BaO75z+/O4Zmf/63cXCW8yWfAzcrqbdtqe8ax6TQ
fM8aKlnF83EGhZpEOXhoD0lVPBugzGkExhphf3u9AbBAPLrjNkizEp5zB6Ko//Ii
O9Jm6vQXS0c4uFD3KZvcHt81TrIHTYQj7/+GKIj2l5XQuDOB4l4Jjthj4F+YHWQE
X3ttkW9V3SyMCI/PBw12M35TKf7awq74inU1AK6wWA2QA8++09UXw2KBv2QJDn5z
x1eFVl0AlkoLO2Ek/CswnZ7yyviVK7ALWknH2gOlGOpBEyhuq/xjlEw9YKTE3AYF
zCR354/tZZNIve5zpB+S6RV/S++IoVQ8C3Wn4NUK9IBwD3aBgRd1dcJi2ZP3SDsn
Coq4qqijSZenSxzvWqgTD4lB7RBZDUjanUwbEo36MOLnx92Y9lkKhUA+oZJ8kXbT
mWnfskNOHPUsUv3SDyihC5JaA82AAyNtc7lbtvkhluC8HM3mIdCCK0dmWMdauinB
f72dTdc69TmK0H1/jwv86cuOcgET6LYgkA39R1pXEyz/jiaYbjAENY3zG3r+aEB6
ZnytUEzag2V8XZgQssFkMiJgdk+eMkA0OANNdylhwqR/PYl3KEcrto8w1n8M2hZd
aQ/09XVEpGqUWO9DTcG2bQW0Ze+jlwgouQ0I8rcRTuDlISh2uZH5YOJAXpk4fARr
JRA7yjZoKzK5mMsl8BSdNgxptSgonXOuHyjgc+UL6pewJGC9quXqNNCaMpdIWgaU
BLaDoMiXh4CWLD1XofPvGBdX7dxziYWGhYfZ65JcD2utZTrZJiDvZzXa4mfuPw4g
nn9+srfj+k+lBNFWtb8EibVaQAo0XRB19pKKB6TelCW1F8YMHCvCcMIujt25F6QC
vXzIUC4BmCnyJ1QoCgvgJ9sYkZN2sAnLGfRhStha16pPsxH9K191Hup/LoKvc3b7
RjSvl0V53EhbS4s8TNBmolKH4sm2S/VXVsojbW7UYNrDFn/HCXNvwd4aX8ILGBvq
R4x0PZH6ZYMXBbvIkAaZQrI7NivaANkUHOUp2hpHt+cP+APE1J50GJS5xBSyTYbZ
EPOd2sTaGFhZpiJlE0B7RCeDlW3FqpEWYGgRMWpA/4rO39dmsXGKeOxizzh29W9G
874LbK7AcVTHgOMsQpKuKmX0eKyVEYy7sjrG/XzQawUucO9SueyJGd19VLUTyHO3
YZRPs/I1np/iSeV2lIE8NjDvtaE/lIngAi5vNvXr0x3+FGcUawcIA084bxWzzpKj
sblfvL/ChTMdxkNgWWquEfMp/IDEpJzjkmVqBNVt1A6L1COtrrLMR8+QRruJHyaV
Xx2OWJkwSqlaogRy1emTon8wLd5H+qxHp2DgPK2HhlhapS+J+B+V7Ak9TJ5WLdiW
LASn//PVP403VbC99vXg6AHfsEZ6AffGBoz7oqSZ8FZ6H9HbqgbOQl/ayH+UF3OT
P5foxf+BNqRd4tykGRuvvndBoMd92EQCeLNiVQxjA7fbiO2I66TVvmPZJQMuPA7/
dCh4vRS6KAzhAuqwPrq4w8etAwd1JrMROv/PxDqqUyPzSQqQc2C0HlZzkoSt3fuS
epdnt7ofyhS0RmqG+W3NnDfvHR0++sp/EMWpczidgrp7ftFXljEATr5s3LF6QhOb
nLQsGiDVfPC4kPYYEpDqu/rfVgQ3d7n5ZnTp6aWCFf/8S0ajEWOG1aRxu0YPoitN
D24c1FjblUFM2yWl3uOLrl6GJHOrDPomyi6bIu+6B95/17aG7oUEfS6CpDqkhon1
XtKRzKFQME8qL9uRY+ohXQBu2B14Rr7s3QZkmWEWqWFByb2O9Juq1LVAY6YbSvRm
Bp0LUp35J/ev2rrrxbAOIyRprwNQ1gMAJMdsgmTrPT6XDp8+TfjRsTuzL2p7qGKX
VIG5FizpSsTI22skGqz+wmxaxv5agtbOrQQpALw6TJEmqSN0Xah0TFUVd0v6MJj0
0mRZBCqI/JqFpx6hB6emv7VisucR/M+sfZCzoyBKUK4cebJ9Iuc133psnxmm9lNr
xboKm8x91ao7kZR5rOIkdGcMF+aQNqsi2KgHU2Js67YeObO+UQRAPd5YyLeZ2WEB
mz+UjWt/1/Y+T6XvVPkwEGTqwmVHkUEYAU3XQnWolJTocPevrF0IUN6TM8yqmqPj
poCDAdKy4heNvmmjKI4IXAcTWAMSS1jIz93/CErKhOUKdt4Px4r1M6PWnDHzbQ4n
ywnFip8div3tSQ3YCiA+waGfslrp0yq/O1QeWDQG0zcPLNvNu3HrKAGHqh3aF1W1
s7C6yvj9oWATvyNUVU6RdCr7+8CkYeyqiBitOObHWiTinX18ZteNW0lPuFC+kKzq
nJ5xSW4hVcvxit0K4SAXYDMASE5OGiWa51nc51NqawLL/ucSGgqqF9fsx6HUqGUO
Ch7ARkJcN4VTobP9L0zvreyzc93GJtZKcWH8wAtKEK8Xp8buNUZq80l8A4mQViCD
9yhdb0w4os4wU2WLtH67k2WfsaYB5K3fsmiEQy59cOAvv5MnBFjMovsTGcvz6er7
NPIYaunzS9mO7RoRHAmBEtH+tV1QMhR0Ji7kcAjL0DzNyLutJNkKVmrYaQ/HpzXn
rjx4Uys9VLF7I9wh7F9xQ5FFJh2rKgNsf3tzMw+VhD7IJUd3oBwDe/oQXs/3mcBL
qnD209iPnFhpWkqOBcxYQCSj4kFPENkAidx1xGPriaNXAdQ47O+ZHpvlV6hqFTpS
pQZJsrNxj5KGrQco93EC8l4wUHZQQc8JPkrKfIM8GDbiGyACDUaScIqsZrPS3llj
xdHQ7WXnFUNq4krXa4NUcbBf/n/xnFCpECjZPEZYHOs8ZbNa49DC0xYQ82rmL4Wx
LXaRnY25wH4FgqBdJDO8eslQvZzD1G4ys6lAy9hg8M9PxAfaOofnQoi6T8nh5a/y
GvsYTOsnB7Wjcb3S+IAnIsQR2gsYCwwlj6woFjIyxqXpn3TfIButswoH1ruQeDO0
Kp1kkgTT7BADbscitAjQ9WTq2vQNiXZ87vGJT9JmY3fl6taDBM6B+X/tTx+GYEK6
WaRrgYwenbFTXhXrqxsy1PtIHRK2qO+r4uUojXR0Fznngi+ubKrXyOrESBDO5nN2
x4zFVMfrw6kgjajLQYP9HoTXIuLnBShe5KQBh/9OznEZ3uTqVpgh7StclfeeAh3U
CE8A03Z6Ep3KzQkwn53kBDst8WCoeeBOKs+53m4Jr/g1TGlfXduKOO/Z52s8Scbe
B9Guh89/15I4cUXNhBNggNWpxoOX87mMfsRXxvkbcvTlxPToyBX3TU/GZQMFvgtG
k9lsq3YDdDlgMQxppogLnDC7YAnd5wQOPy6LeTVyV4Phdb5fNUFHoqI/k5gBI+gp
wDP9leHEOhcW/G24LFdZvsTd4rMFHx5dk9flGeTEHNgN/WN9XOkFb4EN5EZP4fSZ
FF+ATIR1tQBBOQeM9vEoAjRrwMakfZd072qhH3TQDyBMcDrlKFp7KblvAOoCAQx3
pm/fzGTomuyIT5s0uahUwOg2GBqdgEoFiXhpKUswnagvNz1K66IDYbhcazuLbWTi
8xQVzGS/5/6Li8+zM1iDGC2L9l4n9TXaj0pyCx+iSzrCLxtBJE+trIiPOyvE2xA3
hQI1NPDpm6bg3gEmH67ERfKE66PzyzRM0umAZIGcEwQQD+vxjz4x2atcUdhAW97q
PKSyQub///KjXYxANCVSpKtRYMIG4buZeUFp6DRKXJfJRqfvB6Isw9lVbWPFIwAJ
IxHuePFmNKfMg+878Y24YzmrQ2JNoEO4WkFogGous9aJ91oOv4MEbH4MbcSKg4z+
pn473kWzCSQonT+G7ENztJUPSNdJTSzDqQl9+plQeGYdgCKNChabnEdPfmZa9ij5
1NLh/G72jBgvwe4ySt3mXIZfN5IFbfdyxnDJivtS2TilNf0dXlOJ82+fWUv8Sqn8
SBRiVxlkHO5SwBA+PoTTcFlIAkjQIYPZJ6CDObDepgfLeZcyaCOxsCgQgWe0FtjQ
GSbiYUlKDvVc2Sm+lneF5qxa8/v4dFVs5qFdD4246iJt1Q5mJqULJEtOABWdhkcP
2+YeFv+FDZ6nANwJBQFZbtF54ZQ5insmRVRejaLWmBkbXtqueKW3ksQNKJkZiW9f
`pragma protect end_protected
