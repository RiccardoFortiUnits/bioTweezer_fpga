`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Xg1maQMyYWI7p6cCgBlzDGwqGYsVapRF6N/h2s9a2Y/lgOAUqrqaXvVNlP4Q+XFa
pAQaGd1wy0UgC+w2k7mbEJO8zslMDD26QWQZqGOPVekJ0/dFjl1GT8rvgfuDYOzB
98jVJPMPNL9adaMon98PBNIzY/QAUZD5yXng5/FcjuA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11472)
AB2W9+ZCfD70mENNmg4XEMAMx+JYTlJFJAvTrpInq29UVbPbNqN5cSimYb5hb1RL
IjlTtCz2azOpiLT759ey0Gi3TQdTJ2+mkHd92OCPGsIEIMotH5PViGRbxP2fmMgn
labMcuUSwVQuUmYbzBlb4ih54lus4fcJ8VgKURRG1xyzoxdihXiVDc3nz3XyVAkY
oHUTRru6kOPyPDSD9QvYrfVbhPPKSX9sHrdJjrjGApZ0/g32oIyFD/WdjRyqUgHu
XgWC+xIrfZ9vL9qDMHpBFr7Sxg6wKLFt8AQOSC2LfUeRHXwjE74bV91/OL1Qs7gk
HIVMSrhF3V0b9BfV6GPIfyVCtu3BySDTKBaDTQGQ89/Syh7X2D+3tffsFjbRkZCC
KbV03e/ogpvXGqS87Bg2HdhYGNxVUPww7OYBS61SSszlAjftqJK9Afb3jL+76Gr4
Bf+z0zp5tA4/UlXBfxSogegpDiVwdWkS5eWMBom/tWGe69zuASAvvH3YH6w0cP/D
zaJa+i+JT3s6eyXOet2uT59ZqybAVbSNRGb9Ke5SUqm7gSUx1vOkwTGwYcAbO3aK
QnjMdlIs/hYej3YA1brb6U2zvdyP479btLGlZeRdopc/ii+yXhisrh6QtHlqhOcj
A23JAovJgoIMNWJmpMGRIpyQX83F7KBqGhDOt/fKESaw5k8RSrF6Hn1ybY7YVzg7
aqfJtadF7B7rR7ylEcmAFXIw756Kl8h/sAxE/B7kicdiprQyoPAyLwRT4M1X5Eqs
kqcbzxHcP/TBa44njLJeCiqjBv6YK2uE0Ew4U+Ki2Dy8Ju9159YkmYzDYNHigTHS
qod+Jg8r226PNTKfI/RtTjO8ELQzilxsju/X+uNAijsJhnnlcJHcR8P84tQQWO/0
u4xkb2tIHxFWc2A+RD769eEqMeEMwb7zqibG+iBXWC6BTNk75kXnP4GW7+85RRhn
O8+FvCPcmdOhHwROeobSmsuMueU1MQ3Vyt75A4p57mubBkGR6oZJs0BiPkq1P/V7
tP6wk/FGmeuY3HX2GBxQE6MYHl5ETyS78OnjdwPIPaqSPFEFn+KPlRUEAucI8eb/
UQj85+eEpUU5vgYpqFIcSU+rs71U3ozWbuVLfBgyKDZh/u+iGPS2gcVl4CPK2PT3
hp+AHqbV7XlluyWYMnan1ZpeovQPnDLCcAwSOv/XTfVv0JmBm9eBORfFa882P31Z
xuIIU5fUKMR3MSUaRNlzlKLIAhHwsbnrlXM7UN7E/Y4XpYWoNUauIEhlqpHgZWn3
Mk1zHk6eGpMuUajSZFgbfIYgvfabLzblrSA7E7+KR1Kk57cKU625YCuRgD+buJ9a
aq/FK+B3Hrj1nBRbHgj2qYFw3UrZXW7wWRDbqGxdEoYtA2nflktyFNpgtSUn+Z8O
MgWKSs5A4nZahH2qG973BRqfuUHGpXCMXF5KSasgT5Q3XPOWye42xMtefxkUthjG
GV6sRBkudz5zsajjPm1nLWx6zGozylbcXywJd9RMjbBBgMfynRhkkSzXms8Akvjg
1pkHIuf1txUv/1NXQiaGBx417NnGh9V7XZsk3YYsQdhWHSRm7TWpl0zosPBGzokx
wtsX0CtW9fctmbE1F7CVcp5GNQScaGwCIf98axwlt2ZdGmVIHbjBYjNLQyIEt/Zz
A+C5QusKEC0EecXTFv/2DCDfweiveyOEiNw4zhLmZrmJQDVox0SPePs6tHQuLpbC
ndT/lN181At4bUDc7HG0gkrcXEKXRphXO9IPTjvASDfKxojPG5pujB/3LG05moEg
KAGzS3esMnszJztljSnNrMI32OzJpGysBpeLLFX5fHt6L4iuh6USWJuXSEM5dLoR
WUy2gZy4cUZ6ya+2GTMkUbON2O/eo3rRiK2O2SZb7fSAk4Vg2C5Qegm0xnKmOo6w
RxheowsToZrgm/tj+kZb1qcnYDwEU6DAbdNbli8IAY3miGavc1fGLF6Sw6BwKruS
tPyIagTqnPXhc1h7gSRGybeYzVIU8R+Dth60D4WCOZIIMq3EVjIOSaxOfqyaihGT
wJhfY7H0jqJnViZw57+4wGVRjaLnG65991u2AgaW/0H4pCvT6vAqx/2LdAzxb7U/
OhiwA6j7IFu7r2sxUmOntq4cT/V31xPWZnHnv9NFhK/WxZDI9dtABnC0l2VySIW/
8RX+otjsmw3rp8dTeYdG4bQB+JZh9GnaGLp5khV0aatQSmyuAbucKk0uTQIz+yHA
RCAiRkWOnAvvDy3K48Mqf46ywQZyx4ymdO2bMtKTDNW7fX1u/rpx7XjlUO4KUXAz
C7OexAatx7gwE3nXZyUaICdPPotVzjk1GZmrQYmwvW0MUUmFWKmryr8rcex1qZO0
rcFfX5z3AAuaGn5q9QnahrYhVWTWIywZKKx/0kxVjDgiKtH93hJ5y+84q59M0qIC
YNqoL6e/h/xaJqNKmoHz+D7oexWy9DaDTqhTqu5YKco5ICkEP0ihofF2GW4I0EZi
0svWOLXGW4LEhLwrB27Fh7CWXQl/6USxD1XOaACp4TMM61dT3ZcyBYsqGUjP6tZY
q6ajwBvsfTxtPfoLeIrH9cVe7giHarh2sq+/j3fmzIG8fV+G72OO9GFyfhWJUojB
6Arp67z48mZZtai8Rdhjb+LYN9O+WQcOOFDgBa+S6xd1Mm7Z91do2KtF5oI66KRe
ej6J/VHfWzBDJ+qZT/uNiXD2YuCnyywY2hyOQwGuoqZseQafBZJkx7UIEGrAMpzZ
aN0PUc34t9g2tCj3Gic4jFVns9xbV7MB606LwXe1aOvou9RudaNlirfJyWv86ogZ
cLr+2Gn48AO3TEN82KK09ofQaVxgSe8D8FDsTev7QjKnyAoJeCocMLPlJE1RIe7B
xrvRrPdmwfk52GWSHGdUHSa9SiO3uQ4sPTIJuci1IzItXeph6UZlylevh8o22Po/
R2Qba6lpA6RHRzHtOQFPPbZIQIrlVqdjLdiOex/veFQp4bwDS21EQ3Fst9Tt6mKO
Z9f+syavL6pVkPnq115DRkQGGAztTuHrIv/7vUH2Qy4cMecUyRyw9HITT6lKaEVK
ux5GZGhi6+fikmXEuAoBj30u9tECMVlD09SvBJa24vysW1sZbjsdcZAtfWzp4IVi
z7d1ZkGPaDlC0bemrbjikrMsAmunGvR501VgmWWSg0i4ltrILHbupDcxJWZZw+ks
hxwr1ORrSw1oIx94rUsAwGGbGtbSJXEog38vXsnTEKTTVjZWFiZxMOA0ilLjn/Fb
bhJpIPjDBed+Ka6wBC4rvmTy6h108pBOiAuZ10hiQuUn/iMpXjkaNVPFA/yrhTsZ
s9vGjTI/ew3sQlRD59++DY+HKdrV0o9mV20in2ro2KQ8q4BTS+DYXfRtMFkG419w
PBM2Klo/yTws11qgqxUd7FAjC2EVRQJm+pxfQPy7n5IFYck48L1rTBO9B19gjCzO
phuD1iKVmXKTr09KM1FWrApaF1emLDdANNThItkAr+wMYN329zhNIm2sZRznt0nY
O6nEvdNLQSB6p5lKpm3egYpTlbKM8hTwa+EwLIUgJjbZjzAFgikf2aytprk4w7df
9K9wpAqWyOWMqGJgf93cG8/HyE0hdBl/lu1AC5mtJUFmpO+Nd5EAmHE/mpWs6YbD
BczRJ+VwLuBY3jhWTn5GGigYTbskE4R7Gxs9tSoEtvzYaZ3JAgc2rWSC0bIHim+1
Pz22VQdmD5TuYj9ZTQTWg1jBu2EmrAU3RrpSQ2x/K3Hbu6SFcEY7yQnYh3Igq09d
vU5jefsnDnlyBHPTbB2axhq96EHnEfebCAgdwmy6OIbQ7Sox/GavHo3AEuEOPffp
38fhT1nb0fLvf5wfkZaZwJFnIWRT3r3U9BF1Rb/zOLtDifQKlMIaJu4gJ6xVsfQV
3uOmYCcP5UCpbN747wj7J4d18/xTSAo5lCbv3O+ZfZpFYQ26o2L3WvwWVsnW5VHK
m3s6hapFSSwPteTxr/GS7hhH7Vmt6RyxIegBrFfuI6/p5P/Wx6nN/DAsnXS91LEB
845XQz8Wdrihq03TBdb4kEmzWeEgJYkOUa5kBE4RbxZ7k+xphzBvx0AQldtZUH3o
9shFpHhlxxZlo/a5AzBac1N3VqL72ISbkHG9uH2dLwWBpA61OUxIhVgtwyiCeeR1
gMrwIOY4nxCQqWflVSFurdUmC7Xr4DWyzDxI5QRdHFazBoo6mZGVt22+8Nd0cbls
IPctklr8lVisa6q4vvNdxonnAxQzbEWObRe6Waubyfu9YVS8BEllNWxhMQw2kbV5
ZfDsZueIJqU+IvBQr6XBM+Yx3MKoGAp2f82Z/3mImkcev6Stjft/WrU0I9TmOhlm
KVoJBG/beIjoXLglsscHonXEFsGpvfQmzJpVzbAdEaKumctuDpCbDUPhpvAdR2F3
axyy0/ydSmUzCYiVOOCQywbLyRCSkhTXbX2H/1VnwyLYNCco4bwH56OXXbu9npMd
1XleUiDvfnP73SfqVjUFTJEeKh0h9dKBMP96Q64+/LF4aFHO6NJY4c2EE2kU5FZE
9xheGg/usz9KI3LAAxVBQ6D24ue5qeeSfAba8G4rhMfjz3bvhLn/9KjSP8f875uq
uMFFsWTtJQl3DtUVG4SOIWHtjJvz36RkB0zjgFRjVs3C8J7TJeYevpJe4PykNN6h
3QmE2dGfzkylhHBe6awFqGBXDUfdsq3uy74pGYkrDwGMvD+fEmki/6a0lLjnTpbB
zGHP0LlGhZLafvTRqTphruXj+6vq15TSv9riJkrnBWCE1Ljpff0OKis2lrdVZrp8
FWlpjzoO3wokG/Gr/lnrb6StfjpFXyz/oUigPF106MIsarQRw5mtb2HdsisdvVkq
BvawLtjfE/YMpiSX9Tr0YbgjcsRQbowlu4ZvNWVa442OfqUjQ9VsBRFL5CKlBHpT
CFX+rN5RD4nfM4ShxLWPijeJQSBse3KGn45sb8iIucI7WauFND2vor9jYm2id6fJ
uSSiefTZJYjbhabFl5lqubSWwkWiiEbLb2s0Cf6F1XLOLfMbCbIP23CdnYICHYvJ
I0JDGMwYITrIKt3x3FBfQLmR4InB7tC97At4WzH/w6El6FC3cbJHdKBkQ1Q0HLrx
W+ps+msQXMSLKaB2wileGEYFFcOWrDOJilB1z68SDbMRfQyYa/Lgg0COa4ULmJuM
9anW1+3SaiquJZZ0uBd/hnX7quFog2np2t5T+mtA9VBj2dtFxv/lBIBZ0Wj6zxrg
01BLMvsaR4YvU17ij4GWBm784zz3f3jwY8ToZW6gKlsREzUUP0DYrNO0GqiDmpuV
qn/ehE1o7mBWhrhpuocJdc3G72h2eGk/3NDD2dgg5bw14OFWYjANw8FJw5wJGD0h
bU6vmvX5T8cPco9r/yy7B2i0GgTesFTfXeSPuA9NQX4QnjeiCnMNLCecgXCmNIlJ
v3m21iJl9GDgTHsXJg55bfhP7lYB3nkRNDQFqLFhQUHcBr1PL76ss7+nKN8tm459
oKWoYtRbNt0uJIYDVmNWXu5Y/jW3NMQ631IKeUNJWJIomMh8wmzuOoltLDcQW+e+
1tRLEqeV661Ikzb6YDNizmFOHMKILY6RJIQwcFIF/vrw6rdAe+D/wxptobsbu7LB
aoky8CIhOFf85GfXcPHgCbEqkYG3S94cLwDv5yP7JF8iHhzJprGg7Lmi/ydhGlx+
vUGod0kfQuRD9Syd5IUaas8EuiH6rKVbTZAWuosg5B8adIUAI4tZod93xIJmm37T
/xkRKzrPNx0irdY1JZC7+pg40UgHvh/2p87yROTjOLsB07wo1mZxUpH6V72e/zlT
yR8Dr1lNKKBmppE406oZWK79oKhyUDyPs+GNR4yju2detfxgvEoX5DpY39CF9Tod
hRtmCef06KR2YDKJLhGshaLdSrvGJRsmvhIGtz38JSxfYM5Qc4E5ujNDYXNkNqKC
Hj+wDzz/4fsA4Y2f7jcszMLYG3Kul3rn+ZSw94slp1KnfdZVUwhQgKJZne7COHel
uVgqsanxGMtRcX8nniXRpU47igWMdF8v+1H61CEyhVKqNBaCk+qsyUCH+y9lD3b/
w4WIAKnyQuNt1vq5fkRigycsSX4r+qMTAl2vmmkPTIg2/fKeaUabfyhH8mXSQIVb
PB2n/xlo44rNd4JxlTRGe2P7Z0iVGbtqlXwmDOa9McJVieK+tPtKgK7wgMw0uB7b
io+qQcGvWMv60B7FusLjU9dH2RYBqiJqnTCg/Jy2vfRPd3SVOf2c2UjBMwtzvRSi
kH72lTv/Zt8XHEjHZd+9MITlnLvArPKz1rY3QGK3E6X0QFdP1zSjiEQsdWeV6TyL
rUtNokazA9VKYCqO1Pwkw1MvFOL+/VXlqaB6ZjSDDWiyx9Q8B1gKY/Dn6ZRXpukv
Xmsq8nsGZupEFATAnugOSHFE6wFTX0/kI3CF8RQIMOzeB5fv42onhwi5O+PKv21S
628RQFtlumJ7tRgrCkfVWOqktU11DiOXSYeWXPYhzLcs0HGZRpsF96Cx9xzS/9Qs
CCQZ4k3pfI/Gg8mzi4S9tYKJ2OaTr4Q5Igz3cyIL0Mfty+MdoTkLLzBP6+C1MX31
kPYfU22BV7/Lms8w4TmkiULwECi/9Yo5RLzMWRRHOdcXAewwwwNrh281fXSlsgYt
+4gnowiEIpejb2cuDQtne4N//2d+CbfCuTbHOJ9XisW1BfM2bXqCY5NtvJlim8jT
e755WRqHQ+IznQwdYyZt1oSOEVahH827KMhz5QTJsQ/11/AJ1/Ogiqc9A+DKfL2R
LyG00AjVF16KkiDonw9t8ld7NCRzFjf/SZOtS+zdFMR8A2UON1SZCC8SNbxxp3Hx
bgcqlhnO2/tFgnzKxbJbRR0y+S5Xw99I3Pwoe9DDjJ/RVw8YVuUhYOu4j5hniPzR
NxuK09fbdE0Y9oS73DJuwQN2F2ZkP9jb/Md8jpPecDbEOoVjguzIWyePBBeUKD7X
NR3iqcWfJeX1JnCW7tA1Okpebc4Qmr7lgFAVHPQ5fJhCkReRekdWAl24Nj2yHl43
N86Jq1uCG7HH0QC1VDFgnPBPmy2LxIhtJYZwo2gDypWFwt4MZc3iyf1eYaVeT/Xs
AoFMP4gAzxH40WvtT10wzi8yQeTkWpAXngsptuPdENg6HFTLBdZcAZq7UDB1th5r
xSeq1KjtbN0lY2nP+jI2nvRnwLjPhmuSkMxs/HEBV4A7jKLY4p3dE06doeeQ/qjw
RHTspSyu1ndY+CGMHfZVZjq6PciDdW8YMadQJmg4GIF2SfZqxtonLVav05HsUbks
EtlT9vUiNu27WWmYqMXnCEuz6uQgs8zSn+4FJuLck4TdW9sY11zZD/DIa8VAeRj2
AKb8QZTNEnAaNDMAr4Um+OGfIBcYIwgxjVSqV1+Un1IhOBAheFuskxMjWhTk4QgN
LTtzIpKxBuJV0pPTO0cnVlv+ZIpGdht+Yo9mk8XW71DJdrGoaMkY6ibeII93cpM4
a1PpQkm4Hio+rFNYdpjuX+qUEy8MVv3IXtK8fMKBAwjtq/nElFH7PaK6eCHJGNmx
fOyPsjzuQ+Hl1uFKKbe9Ma/Ui2VAxPMOfHJqQcCTUb/9qqMVPaQVsRPSF8bliKaz
NMsLWmMSwIUMdNgPAATi3NjKzq/ukW8Tc8oo/CR6JCsewW0XoiKXyC1mjFGb9unQ
fmk0QTGsPqxx1Pf6w/cdhklf4sT+Pitd1r9j6iIEjiWjkCWzASVkW7x0LegL4NrB
a2MbZZRtEEaiiQk6ZZtFjCYdPKcru0PoPmZ/TI3hrmijVd7j9cWbPzHoEd73R4XE
O241FJnb57eaSKRer/EN5Nz+nfPDTl/O4VdqS97K3C+WmQGU6HYwSrm3WsExKC4G
48oq03v0ET4ebtVU2eKNmTamO0ks/do8IrZ66I+/CDdA+TAuuKp1ZGV79rPLHLSX
VuaxsJVeiXTPyfkpK8xMFMCTZwU71jgXWZOCv2epyfwI3WtpQ+3oW/cgFQtRfjpc
oAf0WPkCfcVeTjDaYvQVgJ8UKeoeXV00FttmV2TeTHL0AjJu/ssD5e2/+UfECh2q
EevGhruZn/aJ5NlaVTXtI9EFFDQXbdMwOubc5NAHueDU4EMPvFFcXaSpLiIsWRmC
p+j6RZg/h6a5e3nuL/AHFKi/lpxJ8i7+BmHAy6/op6vU4EO8hCCBKSieCD7hTSkb
dAZC2Z4fedrIL059ERTyGdoBecuplUS1KkS/ClMEFij6dsgQfy/NH9B/p+jiHUEs
n05HyjsVHtciULbivnS5XGkjNtMNTiZ/ItlwHcfXP4B2BwdCmJSskulKyZdEe30D
B2e/rU93ASpcZB3iPVY/f1I1gNA3HSVb9y1QEztClN6+eWSH6iYP+v9Q8UzvGAou
7CWvA6lJ2CiQQfi/hlf5t53S3jSNcjrLagKwL/hwrfVg5G9qVps5F8D5bzJE69tt
Zeqqay953FLEdwUKYyUQ9BCZDsxYrnXwnlEt4HBcqr/Q9jjYADX//v68uRbGFEWR
IcT8MUVJNwU5vx3zzzdGt8lNX+j17JyO/AxIhz78A6wDzgjwB1AL4YvtUakFKmun
uukg0jO9RZiIwWbgfkiuJ4v3SQvbqEc57ccDdGYUQ7vS07bE1u4ReqTr4F+oM2Tc
YvhBrORdTo+DFdBbhCoyEq5rhSs6YDFHOzVoiAWc9FS4zRA1LU5/FetRo9IJgat6
cEr8Z/Bc0Kx0TN1fL+LzUz4U4EJm/Ai2gtEdtBxYggCCrHQrfd0c4nI4dXNHgOCu
Hhlu0M5yNTRxSQFMKLt3PJfY0Pelzvh2acQmiV+fUmXVT8pukAMlW8X77ypMHRpG
PzuLs0ccUugKHTdl/cvnEqWMBZtHR3uOQ4UcfQ4bKQ8E/ELXm8avRLHubGBGKi9A
Eub1o13rttgRhbSUxYtUfzueZu4/HQ2vJqlduLY2t2JW59UsFN+4XK0SXN5E0rdx
sFGlUmPoC6UXPm2oxl4seh+4BbVP908z734dzkmDZiVVJkK/rcq9HdtQav5PcbC9
ENBCfogcVaUIltrtmpdHX5DjRsim+GdnseeH/E2xP4VLr4D0oQ8eVsbsBQ4q8Ysh
hjD2uaKH84nfrApyPbdnOS4yV5CZXLG7Ivmz7fWJ4K0dpEg8d8rWZH5hXIChSHlu
ZnpKF6IT74ubr9WWb9MlrY6kkJM4MBKAPq73rk9RA33d1Id1QofdpNzAKLSIcvK6
clWEg6sLVYWG81DLhbdCrnE4DfGD6URH3bToCHajnyUMMPUkDQ9FWYjBfJ+sIGyx
Kv7ggpPa2Q0k8JV9p2A0jsTL8H/ot8aOF5XrFdVz8OKYW9YRvfUKWtEuN3th/jFy
2my1x+c0Rf31ToHrqmh5KhwXbH3dJTx4ZwAe6LEs/9le4+ar6EpBZq9ettv/VJ4Y
YXxF5i7tauWNf49890HGndgkqDyWGqAtNMEfcGUE1B3S4OxcNPI2pxKPiYZ/vRKO
AYnyFAGHE4J1k42hov4cgfg4SKtr0xnCuTG0XqpaUNr+Mcx91PslgIvphArM+DKK
LAusehmz3q/02b2Y5LmKlZymXM9yxOzHrlNcTVYI98UiXDLOz7lC2nzpet0J8d+u
/7Jb+fMkDzmvbNOaF7rHj5sOu+N6ntMrNeSAaOqbirwP/s8mjVdJ5VicW0qkxlzs
jutrwI9QWJZwmwo+hzCo3nh06Ednt6nPLB1jvWr0Fls7IhYndE8uY765BrUnZoAU
pxTlj+k6ZSgY8bulqA1lhruSfnBQcCeL3GMoI6saSIfqlZ0MykPuHoRonTIIGjLs
aC7yeu/g8bffaVpkWCsRH0ho8aEVOVtO2vHrQImDH36RM19+oQE+Jht+u5kgPI3l
RCdQc4vh4wnt4pBXJ4D1ad2uhRQmdxn5/Zn7B+jim939T8nSPclL2xoq0ClhJbhY
f/diU6L3rLNfGtF6FQk6FesLMnzNLC8A+esCCOFmCeTsK0xbaSYepofzX0i4osHa
nto8NpcEwevZ0VVCLA/Xrb8JTV2sEsBEbjQY6ugXPIM7gMv/xyb+H93goBxZQ1RB
F9dH/4OO8QDrW2Vm33OqPVEKJCFzbRPG83RO3XB4cGNvx09D3B4rMcWpQxrkVqbX
HQ+gKoMxTxhXnc+j1VQjdovdGBYTsz0zrX0yeidg5YIcfCGU+LmUhj1fdufm35gL
BWMrs949wovpCAk4n3YWdjCadBAOhQJW/nt7yMQQGEfRnz6k+ZXnoFI1cXw8Xofu
XmGCv0EYUtjWLl2Ec/GYO3mqF5svkFCjGdKBSrV9LPFmnvR+DCVeB7dW/TR7/cIM
lHYiOm+GGXxHoUuyq7J3INyZB5zKQJ9dZI+WSr1kSeuN//nOmoA2JsMmvTpNokw4
ywzlJASKXFFnNjnNYXFkS11M+ngEE6CArk59rHbRddSmP4zEHBrKS7Aldl/KTMgZ
ObFDwCW+FsgRMT7R/IRnS4Ij5xc3K4CvNkd8yHjZISqLXu505ROxBmfJ45wPhGJg
D65r+95VqfgQMKfV4S+3c2IwlLT2S8bM3YVcFr3R282HFHNsFLf/lYJqWpoB2uIF
bvURu4A8yo//thDFXzBqR0sn4Wc3Gs+6MhDPkCpB/NHb9c5MVrXcJTFLvn6BJ9Ce
DVGW3x1asT0PiYJjDWHls7Qua22YSh7XtqnP5dXeWiK7hmMSHGgAidGD1Y5ZlXvC
Ny/U8M4Ei1a8nxy5fJZJhzRvcri+ZdakmmMs4OHgpVykkIpTfeqUm5ocQXHfLt4x
/fow0X73zjFTg875vc3gyUrS3qfRqv3vdgsjyXEb/pJf1Ogvkn3yE2G54jPs0tyz
JY7/nSkDMy78soElF5mhhDWzxubWyuf+k47ElmpZjesex+PfM/qbmm3ShtVa4kCR
H13O0pvgGtOuUJJ3cOSZzmTviApK6s1F4NDr3sPvTVxfL+/C0VOmlKxRtELqcs/S
JxtjXfh44G2GfHs7ZCRFRtBk023Ac6J8zFQXSYkNsYc0Hk/HLbqL/8AcVYRCG4s9
Mti/L0pPOcelpRYg9iG9BcEEJyZskI2LJXj/RtFennXFyaRxGa9rV3GvxOzItv65
PFHTw699er8I35/on5ygTebc7v9DAYnjvNVBfrF2QBm3MX07RkXsoVLed9tKGUtr
JgzGnYc++GisqZy2t57EqIXT1qQyNQNXU5cBLiPvVh/4n061hHfvWxcLmPjR8C7x
Jr9W2LhgpdmsT8q/kIk5tIo7P0wF3Xtdlpu+h5zv3+y91eb9+g/PEgp2sSVG1/4f
NAAUOyd0VfAAJsCZQdI1Z2MFfPu/RV5NoVTD04vZx6apgBbH006ULf8HINQclP/n
brSoWfA08NRX018H8Ea23LdHKXv6qE2+Xg5OtJKmtj+MYzKF4eEYSxa7vOmqedZ5
G1HMl8+KuXPbyc8CrIcqUnKEy0oAfRXNH6aAhcnnjBfngB5898vBfCg7HPjp2sj7
aiw858TC76U8rOq+IVTMz8D5G3Kkv1cOB6BaQqxVm4UWlQrcdVbcHovh5O2lMyOG
hSo8jNuSBcLirUw6R0yYftHlYwPaFbfe/S4u2XpnNkx3knNlg8Vl3KV1KY39Dtez
lPZAY4BREnIX1q4ihzqDgE8PkM1+wP51lDunMvloEhGycpIGXmRE/zucsoR93IgM
3sOAbnpY0pvscDvDTyTlS1LA2JII3R3sGjbQ+aB3CsvOJLGHRi2JiL9Dnu5ajyFb
RVT9sQ0NU9QUI6CYzOf8aHIMJLBC4AV0u4qlPXo0t7K1vNzQn/SgkPbOKgEX1q6O
bphlG40EuJ69PannGl6m4COR3LwSKjXAY63YN6ZUs78VajHnf6K+rckgZMovnMyE
ssHvisRzyHs+AG8L65caquA24oXLKxizXzkhNARXw+iXUkZC5ZCjkeEensl+B5nT
VBkUHl8jpoIaXLRcji5Xz8f4CC18M9Sr0W702SRovy2AB8aeiN7hVF8KkEbHzT2C
CdYodEhwkLtq+4o1FlwtGNpm0i/npQIk6yDRIRBffXfzXdTBKjgEJRtfJzxsIxyr
Gp70mlew6WVsa+iqcjIOgFomH5gv+PizwrPGFg4vQY22qLS8K1xcypcxohQyipOR
50dyLNWqAcVGPOV+cbhuZJY0dc611bOG0z4Uk+6g7toj0mCd41MWBsxEHvSupo8v
KM7EHw6whsS/y4WCQEsPUS+u0SUrJq4oo1OQauFqusJiScYZOObV2/Om5+DBjJuI
NnE8wCWzkFAVYbFwk0+zXbsr4HJ3YH2QPYV0IubOmu6v/uvVyiTBcHDu46r0b5MH
UzTMfbhB4UJiSdlZQMaqxYdazFE1LAPIeNPvRIZ+7LBKlpFhi7vVVIzK4lc4ONuq
nMQ0e4H4nyKtqUojXHByks7yDm8VdP1VbqTy2CuaWUzi/NYPqVX1S6M4i1AX4HfE
ql1T+BFI7f2VOEZIIRj7hUwKz/Wap36UIO0x9jyJn18Os3AAMkiFjxp2fImRVSBO
rGU28+4Osl5mo81fF79SPzRqB4UKuE8ycg4hYHItZkn13E9BbDXIlqo0r+DKyn/p
JroMz3pldW7rXotj8RAqNhqRnMXMzg8WtAPMsOdiXj6UDTmzDJah2wrL5QXCch7K
J8cK4f+DZgyJKng56VKaGI/2/oDYGKvgTexN0QjJ+HPNYoOHHHmQ1N3y6WOoDe55
B/RbxncmBIH9tP+WYYrz2jh9o7kVlVcIuG4fGyleIOwphs9XGzJEuJjOobe94DWG
pyl7xIttScD7NlFfKkMb/tHA9HWfrhooe9//l7rlrjvl27SzrHL50zH0C3lWOtcY
v7yD7QYikXxDY+lVuyf8nHtH2B9/nFeyawQh3l11NN1FYqz+RFvUuX1kOve4Ug06
zm1U4CsSFDVGesTTOb3Nanyk9TJbifTdM37Ui7sLtuvPANTfn02woROVljXuUuSQ
14scpIpK0V2OOLtpsazKCXnl/8KFrFc/tnDXD7AQ5c6RqKNV1+UqUxXXbF/wFcaa
MhPSUlyTYzPAM0UI0BNz9Nn5k3U8Td+C8ZAvm/maP2gsMDm0tG4JbC4k3hAssChd
aTtmQITQ07/F5sUEQTQ3XUIK8mR9yBjIMwRHDjB/Hx6vUxBukFRtcGkSEU+ZFgDP
PN1e1v0eBLL5aWvSQBEkfo4jH/Y2q5YgBS1X/cDiCNL+OC6I5Zc10+Lew1fYIzM8
PGiRIUh6vloEZdp4OUiZGU1tqUQO+YjmhTrcq91wKGJ+z7MuR1cGuHAk0zUSNiXQ
IqRYAVXeugpElOxWyEtDeNxsimzZb6W+kHRcHWqjz8kMX1DGddVMTIMc3z8lVIfy
KulySeDfYBHFAVxKbwUkNDLBh/AnZJUTt7b8xxt175I2yB1S8cY7jpCb/jYE06KS
DtsZgip6Xd+7xgIPHL4hBvxCZ3uOJZFprLNqKR1iYLNqpVdQmwpstrv/AgwW+L+C
+UsWbOqY1rjt6HMrkUZuDyk+QfqdeJh0LUeB9fI8TzIFLVXlc6OypUYjjZYAyBQh
CORmmYeu6lPPaFOQI70T6+QugET/HNt2OEW5vUOZJjEElYIN7+26zNr4WH4vSr0W
zf6fLW6fjYjm2z+Q/zoIXeb3p2sOwrKVM5onbLSxpEk6GJ7/7lnRJLHc+7nEtes1
NBkfUSSVap7FuyLALLXNzNJDw04QsIiJCc5tp6vB7GoX/rl+5pcrJAouemO2IVnx
rtH88vbAU+JMZT9mizc/RQkjmhqQeNo9kX48J0tH8VYVrM4KkPk+1w4UMib/1zfB
F7vKZWSkr1MVLOnMkrCCIaFEfqRO4QWvz2ii0IWjjhts9v4TD5vJiiPZ0lz9XzaA
Xbdimm1Yfmi+qd+NPWmA+QyvWqZOiVXSG4NuvYFUHWRWGzyyfovOB0mdkUTroOEa
vpkcj/ddlQEQg0RIrJDyDt9d2V6qtgG7Rr/5AX2fj9Ebw/UzF6UmQfneUIKPHrZ7
CY47K5wHCVEaf+Hu0aDqzJ9/Yz8qMDp3AhCAwKKN7Lx9UcATZ2vz9yOP0RU/CS78
UtMwd95usFgiJfSnvOK0o6hNGFIe0r6VsYJfg57fqFeb4jq+tYGylZmXJYuhaPYT
4Cf6LTni+bvfXUi+oobsDwVaVGxSKwm19B6Yfrkf3oSx9CHxj74cdias8H0uO80C
PpkYH/ZkP/qOpA6FaLou3045orNTU3TDE5zJ/SYrWNlPeEYeEl9YL7WRvH0OnbJf
/GRPemZelRi7HiR1xHqoTmTHUB5Em8zboD2pu6aEfbei6VDz254N3EpPYrgRlA99
Jx75B6qWCHcxO4Y7gLehfBSmL2OylMUSo4spo6qLogBA81Hx0DFjiNMEg8EPqZMg
H3JYdB0AtQLXda+ZEzUnZvR/MDfoB0cnd9edWlRM0PXiarjrvQEf0KJwKFyU/QLv
99iCSBKuOWzSMOhzrClO5OnKMqsr7aEdDDGamXjS0cSLlAQaNKCUmAMB4PYY9Is0
FeHnEsEdG/M11LoDx4Hwr1604bdP70h8VKj3YJAsAzoo6Qw8A3Xg0EKocEHAwvcM
LWIcLPGU14Q71cnG8tK70S9fqkXGzd4X5+kDAb7OYir+wimrxTeYzcvhTHBVj+bX
ZuNcdeH6UAZKKOCqxFX4+mgnkJISubiHRLVpkJiq6wDp6OtH0znclNSc0RIczWFx
Z2y9CTZSuP91s7S+GIUY2LmYF5o4D3Tx9K/w1qTTL8zGDUvXQz4s3F5segvjAoyg
XBPM2viXIIbNraoQa+Y/i/GYkqCzSffJwyRBrdx4LqFVIDGDaL8DFltgB4K6NVxI
xH7M07q8uHykC9pGxpKnFI0UwEeW/VUyZkEaXBdTPKVyAFebN76tHeyPcAMkXRHG
FdA41uznnmhZEIVS6hJwp2QWMJzTMIBktUbBwWx3oymwzrI4fLXZqCLF3ZRxnArg
8SVLDOFNLft4gXg8+XidTOdUAjsY/4EHKccpHLNE2fjucEVLmKFYhD605j9yhL7A
X/7l3w/ffnTdBoebUiK7o9P7z1QDQuT4gax4yiIxBEWTxQbWLYG2YASnMNoz5DhP
zmI5eWrKBDi0MmK4ziYFVOXfiGcfMTZxsIKtaslAmfYs4LDpaLNch2PlOK4MSqqc
LGboQ6emjPeI2UmSUh2yeTrBb4Ou+OenbYimwe/GPqttTzc2aDe838xP3LE4JQlV
vlF++JhO7wvoKYvadiOOkHBOxTxcD5rPuJy6ia/1aXwYCckEH5DeNNKVolyAQkpz
/STFkjGZKnphohuPBlPJZbUOVHFavrT2VC+IgCaEu+T1+mvKZfmWH+UyNrXUqMtL
`pragma protect end_protected
