`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bZEArqT0gwKj0AQLH9tZUGfWH2jGL2TSNMImDXQ4M7gzKlin+seOzAhAiodx06mf
8aHWEEP3vvLNjh6Z1Khwdo2oM4onryutJWsBCgSK+uPrfhPEo3u+2aZv5xABrqLm
y82qVtGVpqtnknRuRInEhysAMo3srXMeAs5QmUxxehc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71088)
jopTV4fzJd+bcpnIfes2hpH+jyf4ajvGri6iyy0twhy+4QGsBXrjJWfOkPU0facl
Z5oElxHj3zTIPAdRXfs0tyMwpUzPnrqoO70kaN56TAHIaY3umaNTEqwh/L6BABIz
AG9H1m9yL4WD+0GucCWyJYO5+x5Ygq3jKUaS5PANBRM0S9xndmK30lK7WE2IyD03
0UpHyRPNwsAWaz2G4Vs5pHay6F6KSl7FBjA4v7N+M8pcf+aklNh1VMqLH1jYYQpo
+ypc1oBCPmk1u3CFU3gui7mrQqFLsVMyxQGUXCFulnanpHe+ECkSib7ni9UCyK5V
qa4/ZOqv64JWdRn23mGx92hCXXkG8hdrcJmbCXXCXTa+K3zWPSXJt9Q3/oq8wP6e
kDpchpcUZME6woOfXRHDWIASJOCdjwMioJqrEOwS++WaaCxai6AGiJdOH/BR/1jC
nxVArUfGPJxMym5jEfTprg/4UmlzX7N2HvxacZMkLUq5PJE2mpRrQ5u6EfBPTJQ4
L571rELmRWUWvOiC0p6Lq63zPY3Htn8CAyVEbh50UH8yhQ9JN/Xj8Spwm+6l99WE
IjPsRkek3z8YgeoTcaK4rNgHYibskSRi70wHoz8Vltr6Ac49IDt/6punhG31MhG5
yvvs5fxOZU6pf/IyFAhPqa75+1BTBTbcRAe1cFw1aZEIFGLp+jxtUAd3UODr0bLB
bu0FPtFwb1MXmmiZTS745SSmP0y5NNdQBDDS6WaC9A/SGDydIhINsRzjMG7+a8FY
zp9qYOsCPkq/xS0cfvKLVBOwt2isRm3A3ZtEw9VI+iLDH2N25TWnVTEqbWF6jSv3
KW72ll+0C2EJt/hc3CO6mx068tUHkMroZ2yJvDaIB13itijC4qIfJzW/JCle2X0b
ADc7PRhLhGN6U4/1A6o6WvSvfDFchUYG0F34ktwrXiRnIEb00n/TrPT4fIeUs3AZ
vORH3t/Df0I354aGqrUHY0Qco7yHC1fRm75bHblU25GTDXcLqBYzvgjfUKIsbI1E
zb63tyvCqAaCVVHZT38G0bt1MZoCNxskHqneAWMcRTDGFJHCAbJjqF9O0SbHgV1k
68cXf0SfVNAyJdW9zhMMJ5Df6sZ6grNrIEmhoOk+T7zEpV13zOeJiwyj8HvnJmSg
2IB2TYZ2Zm7/Oxj226mNl4QtiGCTbWz9Yda98aWCY42eJiaQzBMOuiMfqYvkviwd
KdVCFB6dv1nLdBuTmE74qu+8wP77eULwTVUe7HxfCG6fOhsToCC+5G0uLPDmlZUh
8McAp0RI5g41ReMMT+xIk9uNwTdXsbdkWQqanrx4lwzCOeelMitSvZJztS/IBHzo
kbaKa8snooy+JgWqdzb+1gVH6ZGJXVu+ZTKj4a1B+AYMEdng28fx3HNfwAUqW9tq
Os0jjDTWbjEXot9EsJNL+vN2KYxArHm179hF9ZNZGm3T2c/JelPD8d9njWLtOTLT
JZt1lKNd6ytP7mir28x4EIyEAgoEUXn5P649V8D6oc5oWmVPgf2h/Ddyu9bSO04n
RpbWg38ED03BjgPb+gR1s20aV7+YwYt6zb5fOVVaJ9HjXxOt0uo0lcuVYiIeQJKA
bzNIEolDEcgW2onDn6byEmRrJ6CEPBAvoHstrOrZLcZ2/CE0L3/iuCz91XoeUASO
GJ/xsD0n4xvX5GWlcybx5CStu2+9SKzWVr/Q+uTCPd0VquRM1C3C2A6wtsvkjhTM
Dm1razXEv9Ys4cafgGFvLf0bBEf6aVcRmuQMdmoTcqL+4rlyuzY9HtOK/nRjnJ7s
k6swr+OwOqKxHKqE6DQtc14hyDu9QH1ZXGZdoprKET7M0p8EDI1BADGfU5lYtV/A
buSq3LbKVgjKtpfE1CeLT4AjiXQROiLQtePvghrB+bZim+dYh678knowhqxywpHj
1AaE/7zBhxrvmKu0ogqBQXbI+/H+5pmUfplEhNhAOqcVZlTpWnDiOGwTtPB4yxJ4
kxikmRrWPWU22UCPWPVVxPk5f2FqorY7VADpUrDvRMbLn0YXSBVIIsdgC1c6O2jb
1hz0Gzlk0dnKZqtPfFCkoauZWeKmEijNXXlb/j+YOB9BcsK0cKIeHU+sIbpZQQvg
le2LeGGgeqgs/KK2gwzXpW9GXc5hhXHG+xoW943XKD+dvF/F9otNTw0JN8RMgqQh
jKLqrAHDYdxotk+smVeX1MFgbZOeZmimGkaZ1YK6jU/GqULpfWhdL3JKemN66Xj5
bGfsM5QDeY4iklC0twPYXND290UiJK+WLEZ7vyPPD4OQ0/GuoUnVtny42YaJ3HIF
o1SzYm2higMcjd3UjoaKY7U5kBPA7WRIIVEoCOBiwqjHCsvk6yr3oFnr1IM1r+bn
IbzacZ03ew6HEp6yRk91NLnzYNLeBZTWkUmbbyDK6WI7De4U+JRvezyvxBfYnqXP
zitjHwEViW5wdZI9/5VY81uJ/J163DsbBtkXgn0l79WCf42zeeo/Z6Rur6Kc6aTs
X2C5D9cR9le0enTfCQRnNfjaeoEvz+QMR/E0taf2PJfvtPL73lDZHxIy+Gu7SHJD
xujElkCL9xzmZAO43XzNSi+912xg527k2HaS1i1eCLgnSkanOm2hV9Vfy2gI42tC
20CWNaxUHnCpGbIlBUWXkWLS76BVHN3eh93KNQAUfwk5LB9q19n3ZN/GBGSGO8Ip
88NExyyCC4fwgrgns+F4fYWxW28LHAvJz8oKPHZ5VXt+1de5tV30Xi4spWEvCFNI
Fd5JOeOdFhvoLJyiXL2Ga02hppBF3PFj0vUlUIigmipK+pe3GrZarhWSQK37TEFW
t084clYZnbPbzhVT3CkW/ejmhkTKOA+vUwsLT7zwsLlV5PjWTLwJRG209Pt8bv2y
G8ek/xnJTJ2/Yn7f0x2IPtkeWktCOxNT81UkAMhQARDngrzkWlpn1JBs9V63eoGE
yKlFcj1Vc3+srYxFFDoYAslQjc2RgwuaUiKb2JjnaK6/5sZulhBKy5H4XzgP5HzW
uJHBYd4jaBU9wO5paRM/qpvza9Ia3rM1EY8BaLJ1Ai3c756lQeIHtLqRyVK4rQ79
kFnpYa6X13i+X1gN432rIiPVlW4u0DEp5enCNqtEeepcdAK3UjWpE/x0kHp4yJrQ
bE/pXux5HACWhlVK6rzRaTdJ1gfmm2QHd2nBaJ7VbeGSex903WbcUMOWWNa50hqw
/7e5kJ3d0HqZgxpEIZrtQPRaFJJtwW+NuBM3D855ds/OQYjDRoyzMuXDxI8MA8u1
osAHTEFFX+NEeT6fmVstnqQ+drHi11puwfxzz3bOvSGTPg6toF2CrJJklGJstPyX
T1Ny/5+b6miaK8jYoiVb6yMicm6v4KBYVDeqoSBM+vdZyk4vwnixYXSv+k8LRrbG
g33/gmrCo+YeFtjFT25iXugQSvxqTmKdiQFA1HO7i5PyqkvfZBto9sojK5MqxWjW
9vtAYurnNlxujQV5qFSr0gcBYxZ+vegzMhtMNUDqjYsEvuvTQBTn0YbQHkX8QBpC
PmcPcsdzs34dzERzAMR0fMQkm5NDeKBjC0zcj2xJ49nbmisR4eHZ74ZXtljrSlAw
cN4nXuFOs8v2xNPfBW22r/lmIplZo3GAkxmDMzC9tZkSO/T5FjPZHL+LbasyHMsm
vf3/Ezwksm1TbIsOmurOaipIwA4ZymBQ7JURIMXNOSpim4vP27u9XE0g+kVjEWe/
RHKnYCr229atzWuteKUgUxw0k2psg4cC+eG8BrcLtYssVGsG5cg0diqhqovBVzIy
l7fuhpEW3QRLuvZc75YjLQsf8YmHh7fcOv9Utd2+cqUU0jnPiT1KHJ/WsVXIPXXu
H4+DHV8rN2f5IHfAsTwKxMaEOOFBQSpctkTXdpS+TABDWsXPJVpEqnWYtL1DsYZO
hUPOZLtM6Itv9Mlf6l4161wVtYmNWXOuVStgOmUiuu/zYZlYkuXXfrWdFQS7ibqx
9xvy4pPR1M2lvHnXo1Fcz6Hm8K1zAuNy5/erdntZBXBXpI8TgXKR5lPwFr/azGUa
2Bc3FpoNPlTR8ulV6J+ZM6MMEpo/DEdpxFfTZKptJ8pJdJcim0ZkrMk3MeFWAzss
8dx2KZ7M7qTtL476wD3wwxkd5a58/HhHxT6BoCA9ZZo4RLCueM3U7fZKIowKFm+g
L9tCopYIRkxCbQVQJ3qUVajCqi3fuFKTKWGd2rro65rpePeCQxkVm0jHWsl8584a
1eow3Zel6DptslQQZNLyNvo3rwnzzPU5veid4wvbqP8P1OglwDZG2/dRvM/pZFXS
ds2K4Eb6Lq0B2cOGDBU7i7P818hRuJFRWF1FZZgFjd1pBG635ezyYogCEj75hvQA
tb1W732S9UN0PCIiAzsKPky45XrKOgweOeXDZevDBioRPowwk6cZm+8EVPnrCqRF
LACurcoI55fyClFGjW9tHLNmsl/9yd4GHUVQZlUH2Vice2mlkF8rUZh8zUi5NTSw
xVZbcBS4ZQefLm+9J9zWy8Id/6sWM9FSVGSHJHahfan0B9QN5F54QstLs27nwSDp
pxlAK2gG7JSsScZXhfA7HNRQRjgENWHGexrED5RBow9iBLSUPY+iAEK4wvK/jaxO
c0/2kEppqVAFYY9NOPpDCO6xttOnZCiQzzqq0qhA7GTPBT68SgImsz6U/AdvH4EN
zFqq7uW29qg1TqJGV1pM5YBQnoxLzwA95uPAL/hVvg594mXsD6WT4UfYNB8ZJJMF
oB9hqGaseYgpuRUK80p4XHkl7NFqvZLNTBKpfcaqDSe3MpfvAi4F3Kb4wZJaHrUq
HBUuft1un7lKb/ICnOwztl1uVMvJAE0ufA6jUtgXMNsUXdi6BhktO2TeKM67I4SR
E3s6dJ0Ja0H07HEDzD8C7F3YBukaKqn+fYHdUFr8VkEgUjLxszZlMscB7IPdDtZr
1KKAq8hUIOWseGXGnZJg0maqSSETJqFAWGp7BG5qVNsS3QZLoT9s0W89aqEycRtT
gRT+P9RbCbnJd/1izYYc0xqVd1NVD0vdxWdr5apxHthurDtg42GFgDfJAJT8vzqO
HU3cRZt2xvthNMMO5TyfuPewFpPpqEwFSYijl6GOlAmdZe4jFR9kY8Dbycxc+JaJ
JlRC9BVqGNh/TZLYxoqQORzoF+UbW8PDXmMGxkF8oltpJt0UH8A9f2GKxzQhyDvw
ITN4ytZ3MoAFD15G833GsfuzkdsjJaa3uImP6XcWo7lmJO6O/9yHCCg7IEl7E/4A
ONMqv1ZtYFFxvDwu2j0YlcjPfryGpnbMvmZOOEY3U90/CEiyZ6IVI9cJgjYC+9KQ
7bifTaZizzy4887+wNKYy3FNewhOdlurNiXEZIR9L3eld0DSfoyxHuNKWEVdhWhr
BTJHKLUb05dDUsvSkx6KdYkweBruxse8mNuUKrFBphkGvOD621Fa5SI8GzTJSsDm
mLYB8zUd7fCMMKs9E8+y4dHN1x4lVR+UUMCpBjRLkum6Y9h2LB9CI1XI5btHWOmE
Lz+usT5Vg7DgPJyjRv7Ha9xcnbTl0NEjAgIkWpA8mtqX81JNS01/XjwiPrtY5Pex
begfr2vJh0GeNqBMdbyeCV2jEDGOJ65ak93lM5dQRhB6RCk44s31fneL0ffRcTWN
AuanPrTFs9s/n9L+KMwd7Njub+TUplzur5gWwryWVNTPOr1QMw2fCHKwJ+yXLGt0
UY9f4Y4zX71kj7kM0dn5KotojbipybYGT0wkwAREL/kKDQI9ThDuUOgK/Wd4zVRF
pQnz/fAUuxTSgTISJ3SPiAJJEWNj/g2nXzxOWLazN+dXac11oSA68Wgicw1KhbH2
VCwoa97nBroxeFi8Y8koyDjqGySbIhbBPsa6r62C1MWhbvhwSYYOGt1Wz0od9oX0
41i/8P3k9AMxIL03jZgBrIpanVGJSnQUNMt0t/jYGMjSsuLouY18JG6nNN2U9pGd
aX13DEttuNTKLwY6CBjfbQsFofkI9SsWytGrhACZZPYpaSrFBPoOPOmdEcMcT2HW
R5sADBgnuvoZ/N/ac6zyZZvzjuqwtFckAqBTshH+XrtdXWdwi+uPmIgL3Sq9zhd8
MTX5rYFrxo/vYaStz9t3MjHalbgHCv2ELjHN9sr5Bzpcfu5tYmNNaHw6Zu/uSLG9
h5DZDLl5dK9WIw6tIT97LNeMPvvkuVmy2YjGD3idSeinyIHFZ0PgeRpoqt7KfGai
EG528iAxo8CgRtt1PCXmr5qL9Cg2bNnHliH7t22mvm0Yf2H2sKH530xkTAhU6hgp
md702+JsLkg/GOURJJPBMq16QTySJShE8RNu+4ZeRlrmS49G/EtNgGQwhU1SA97E
AGD7RsCnPrzPZBMD74mcOPjWMngKWVcVyHu3TZmPOBoZldojF4QuWj2SYypaI3Nm
pdILbADoLkGi6q1/Lmj/3M4tiVtJDOaClY9V9n9CC8g72gR5aJL7mct0tc2ed8fr
0JMhRn+Fm2gGRQedSa+VX5ALlF9NLddAnXf5SXW1te1gE2NZk2vpduKmkLTb/VYX
aRC2kEayLh9TdiM7mguFes4+eRsHF8iqVErGWPSyvMSs4lnzHwSLKIOx12n3iYQ/
cGcDBzqly1C4/G4Hg8VlRi/M/qHDUXSBo0GUWjmdAqPJsR/6yxn0nlUY6oNtAgo0
tIPOrQlPNsi2kcsvQHYh0E4Rnl94peYTeS5H1vUYvE/krapaBCdKbY1V5U421Dvb
L6K7jvKinZpQQby1Xf4Vj9LY2GYtKcjkaaQDzUbjTuV3uVFYehDjwg+4r8Xrq0f5
dxWyEDkQXIxhgErivPfo5ACh02ReYliLJiaKl9t/hz5XyzxZEVdQ7Fpu5jeUy5lQ
Z1IUF9MnpBFaYlZ5d7vVUW6Ph10Y6pZw7mYfTs8zH1ihR3Dud42FBpk2qzYH4i5a
7pxGMigm9otjuqKW9HfPgMWa3eqZDX+AI76svWzUXq020mY2MyaQigHJHm5XGXAH
AadAmYo1yzgbNTpuFaAncFAx4adpzg3CfFriumZYIWwLVgezdCgD9I9J1NWQQeLI
voA9MnJWQ3lOR8M7gxpf/8KTQ1Wcz4WdO4BuuPCJH7dBJ7nl3cTT9d6mjJFIZhDi
vTQ6FI5VQeBl7MZJBxbIfYVbBZU0bvf1WwenySvj0ZD15yzBOdH4+1/v5nq8BybN
KGfB7DNHQYVxo2KwJeiBJev3kAc4sL+ouRgfuOXOzr+AvyfzjgygROvu2VXiXeqG
S+z0oDuEYD9JwEndendERzyWQ24qTphh1ApudXLCCBa5+StJpxVOCoXTtpm90VIT
F8zAA5S+8IQXTl5E6nfD1zUbPKOWZ/7c23fU7hgwcZ5yzFou9PZmzhRPgMkZfsfh
rnAwJJOQU9fCtCOfK0hE9T7Fs9dW4Mf9xJf98S4gLK3fhpplTgRwXICAgvaBnPz4
XI2MCBqrywle0XwMJAY3WDdVkC/Ib4UmnXesHd1nmqMtS9oCwa72AuLnrxV8pHgC
QBa4fS5beUfqfcWT9YW9wIvlR3zCfFzSh0i0iYG0Yj3lwEnJiCPERrMstuxUmyKN
xvxzSuhWO2ZPnx6oXpzqyDnINJBBf9xopoH8qNyDw89a9+K1moE3CEIf4KRjme+s
59iNEo+4Tl1rcleTNag0TFQIADTnR/EvSDYZhc5RCtOQju/zpxXEMAzvLX/lC85I
9RVyK4DSfgfg52ln90BWd4YT2jcdjOSppkjcrQaKTZAnY9RYOKSJCDpaJTuq4rmA
QE0CW1LpkwLWR0CZs4EnCUkSbEt1UxDgpgeTSaO2OphK3OwGgkLFclRMmF7sOKbP
5KOddz8MLEyIfINJK+ESHzqJFB9BgwRw828sXCiE10Qi9c3H5SsQQDvVqAx9Tk4r
NIqsG7vwnyqPaJI/o+t+ieCna+8Ag/EOr89iEwKXvrzViOFLAHyJ4/QXszbtUttx
Nz2w8OFBt3j6xtkPahDcaj9+3NErh9N3/5f3nIWAcfcLVVXX64lrlZ2suFvdXixv
/6XTsOAm06gw4Ig3oKgvBVCfbeG4EkFfNMnCEbF1ZBvr7uLVcBfW8ae8OXHveMvE
RWA+sAl8HhM35h8JI+/GjIIyP1P7losOrnWAxKsu1Df5m5MiAxZkjyc03JyXcMEo
1qZr6WGI+6gzQeb0tAP7wnXrn+mnHyaUaO2Svfo6HjjFDJOtX5u91QAThlTAZkyH
vJjL31IhOtONBjBK/MfypLyC8kzcHeSLQbnAYi7GwBN5IbLo50SXwn3kXDjRN4ve
yqwSaKCFtOgx+jdloZQMmitsL8ehml7u3UzH00z0Le64T1NmhH2Pn+CP/SKkwaFD
jFW9I8i3BMYAZ7hoGlzRq9QxPMwvaiAigRKYWcKGInNI+aIMfrZxJsp8vM/PJuo5
VX1ou53rXOlp9Z9GOEmD4rt48X5tNTVxPgKXGpYvT271VyebseXx1PUnsl1F8MRW
j/RYZp3kiXb7wEKsAO6MxxdnaoUG4rmva+paaYKvD+NlhyLpaMSjae2wyxwlb0ER
S5+HA2UiAbMYSaW4untAUBP1UHUFmH6rfgcSx+tug7NRGLXQ7slvEw52kWeprnN1
HO718yQ2WIHpMO0QWP+/QG4d32WYpU5HmTgPiM0xJhkr1NT2DkpxhFddEnbcpQ/h
3QqiurbsdNsECsdu9GDZbnFmMlVLGmJKgDCP6AebMnyn/foqVjDecBr+WR1R/861
6wlAlqkiZkpk0W88+ToDwb2KMU7Z6pg/eCgssjNzrs6+nCIHfizwFT0NBG+vZ31d
wCcDa826tSDNfVV8rvwdeLiWqVB9isljJXI2NWO7otjCE51WEFt4H57BKJcIClGH
/FNx+j0wE6QlTPKgtpviOtdu7UHxDfcgDfhOiT/ytA9aWx0raUzCPH9dU3QV0htO
N78/tNAv3B9yT2nf4UklAN7/tVARaQAvP7x33vpaQGTCbdPSixI1m/2/Nwhw9nhK
SterxXsmgCLQfF6IxQbAWzaNFLpqdl80WPQWQfutNCboSXRyZ2pzQmBdmtEJ7yYg
BkaVVggi5IVjOBdSNKGxNv0Rvj6PrW53cjDimyMm/40EtoNWPsbW7NGp3OXlIhe7
jBMF1R8AyQNi8SL6yfSLqxnl3SwQ9CpjM8oLzfZuXGf+UtF8SuIAfQAs+YtI3cCO
yhh0WuwbS42mSfBsE1W1xFjRHJ6OdNXZq0OLFvdcq1chaCr8iGjHruWyVCqoRc8b
HvNGmszOztPTNKT733Zgh9LwUtHly1RYJlu6xRBq3SAYBq41kOnvpsI7a6s1gy2a
V6HUqaZrkSMwxc3N9aFdEHNL5l+KuvDx4JPp2cl4QjpuDWiwOYzSJDO98a6I8LFz
pyTOjFpBli3xO1fQpJAJMQBYsTr6qcT612bh6+5rOcukgm1di6uUF3v0T8PAuMZH
Lzoq5WsjzZIPyYlJ/PCJJYw/RNv1j2Cm2u749CGZXeWwJI9XhIAZVPdGWRY7dtWy
sdbPeWly5E+OxVKU0Jp0WfDkmt73R0Amf16wyohtc9YJlRq/r2F0Vi8Zi8ZpUH2w
/QDcQevwt4WwH44iDh2rPd3FA+z/hvErzD8LuauNdjXeD1txtT0jvCsPTzXyjrCk
IXpW7UT7By3m0J9to2RzLLw6F/3w4df6W56Zpv4Ye+18VIOx0TBqwjL2UOXOk7xX
omqbklJUOHcLBGbG6y/UfJJPSnttL2pK+qHMe8hi6XwGalOJxUNn/qrRXLquDPnH
jk1czjXV+AtcZk1hx/TsEUHvFLMpt56E8wusbhXTOz7c+NUYEww0UrEj8yYjDGkM
atyzxkrAHD+e8IcLOXUZ34k7d+W+fVqcwIJqWOmkFe3Jx+9yWjrbk304HnV6tB7Z
pmkkQ8H+H2q2xvtq2gsKJciEXNmb1wIO+Igr5YXv/sX58SjHHXiEGtVrQBWdp7Gj
zWTDk2Q/SLv22AYmx6TzshkIA8W0HNOno428QgRSbFWzhH5zZerFPw0DccwiSWAX
sfYVz/eJn5gerV+VckmIME7AaQNq9Cp8TwKH0W2dlbN97H0t6YABfrsJQCQf8Gm8
yzQfJbo3KIe4LIK0sCxa7zz7+jYEYhnReumW7PpB7kY8HAsSXZ1wYA04S0c4zjmW
YY0EM3NtllG1U/DtieUKhiiTpxW3yB56T8nTFhOSLvCBW21vxXzGYce7eO3Nz6BO
dG8XHcGJVDG13GwUtygeW2MqdWiB/BI5AGzWe4dRx7xeNyrYBtgmmChhms/IqnBT
rwbmCkKTqWcQuCUpclw8r11rRcgkizQejnqzBmiRkfmy6F7zChT62r3sOjJ/yN5h
arAaDWceJi2Tzh2pf+mbPl4EBMFi8hUvnWmzAOUgVbs++R1b7uDcXJDGFyu/07HC
SOIEypNh5TU9MN0VQK1B8yYX/Rkg3DYcZUIegTf2cLGN5zqHH6IsVpQ7G+OyRTOg
62mr3jUTwxlX6novxrWm+ZAMTMaveUFNvG4DWcGNAx1YmSjA4VRhJ5543IPjYHPb
EUbHqFvx2A1G07VIxW177MfNPqU95/TS9BGqcKWMIMaFxNPVZT3/TMX41DcnORjQ
PuKe8kVYQZzHdKyFqHZkz04p5fZXLkKwiVlywDqYWp9QlyQ3fFM7gfUBKcWFgdgX
qi9YhWb7qxbU/236OmVX7X+vLjmkAEd/QGuoI0ZDqOzBUAnfbCklw/0fnhjLA++e
EAXtA1bNv7QGgnB/DI/wgj6vW82DbtiOfow2MSPuIB/N5zGPGCTsKtBU47kvkXU8
2zPkjWVfoH/YwNAaOG1iRyl7VTIhR5GifNJJlY2SANNzNACxlFnTFsZvrLPUIGqv
B3M+gL9ZkRXzWSoeIj25NZX4x0V3PN5fwRY9R0fD3w+sLF12dNzjANeNb8KJw4Qy
ejKrMED6+QpzbfOvQMRlJB6INVrUVZgajJHxvEvEvp/8GIcIhS2MMd5NburLRCS6
p/RCXG3z0XJaE5A0snAdMYz+qhbbLrIKU1/MAVgwcsq4mHAt2azRg81utMN6+Gx8
/7QnIQ3eMpONAUHoJbnJBDs3Vj+Z35lzq9DJPZMEc9YhffWoAgZontIWbb5uHyuA
ARDmoARYyMY0H31AX7D4edVoXT/qNf5kJ5q3ToS7sYM5Yx0VG6giFgocWipW8ORu
FRAHv6PdSS3An16tPVAV7SwRNHtuVSl2gekGvPUQLl63cfV0P/MIbrcb4bsPrJmw
JNHLZqH/ywjV96sgdOXDkmcFDhzvzPQn6QbbiIaqqrfYFEU1WKOSNMHwgrYKbu5v
vXPBlpcIPYc3IjFpe3t64DkPjnL+L2VVPzIctTR44qGZ8LD2CiCnCTn9/rua+wcq
lDznebx1T/oUySw3Es7Hty157sbxwKxi5aDcmwlLL04fwLoriMXF1FELaK20Pd3x
9NrkAu/lNRV11e83h6JxCUYH3vn44T7dS4xZYiE1wUvmWLbPAfB/HAm1FMIy+Z58
H0wCFUznoZhswiOUMuazWq4cGmVt6TiXgL7KyMSkFDz6h4A4D7bNLzLsumrOwdM5
AjeD0ZkfJvLofdW33Z2bu4PtgnBfi9SqLYuv5DOM9TJvzMRPdpl1xqfkL/W0EhRb
+lj7N/2yWS9VHa2rvJb0j6qitEWF1QeFy27QPQr8x63KYtX9v691XqDzbz4pkAp/
Mb9g6KlB95wDZPGpC0IvOoanDjn40Co964inF8GuMssu6ufV9jXMv4851/vd1fXi
mdFAajt3JskHskgbmyN4ONce44+XDMMjVuYCO+7DgWy6Y8TWIuGW7SC+sG9Rrx3X
hT+YEHZ2071M2zVep1kk+Zr/ICRSJ/i/Tk6D1T702LmXK6ACL/PUlzKPSdJgojpv
iPQvHdE7hABISXrKloGgSXMdUj6+JhnqGzBct7BGAPwajAfY6V8mBYLYxsK2z+No
jpsrsxi+6dZ+mdiKCZMrcl6+xkghTUTFtLkW80EV4WY6sTMHewlGD9dNpIbtFBxR
YIR3DqN8Lea7a1pqR0jkaUyjZ4tNAK3WhsWMD5ly0BOOQdNwT/E95pPWRNNXWL0D
UqFrS5U3KVA5LSz7KraiVDGWB5fBuqR4vWNLE6W4hIFM6iQR100q2CPCDHql/TMe
r/fyo29oWjUCLx9dxYhjreKvfiMVXuz5BxuMcR0KKNyIHdkYt3pCVtN6+UF7Mhsc
saU22k6yhGHol6Z3TqJWYW4hL3Ez/QtsN5YBcCOHuZpkVGylFvBOYOgJOrtzzSeg
gdJXL8/9gm/U3ft2pY6HxQ8fVa0MZ0fQ8OAkyisKEphOPACaS58OXJAZhIAam1iv
5gt4euNT0bDcDwolAANWEKPL4Tx+yMUyK953xBTyAg+e9hJpqRIQMtiGFOd9Mufa
k95GMGAic3SEU/1cuVCxZQIhfxppT9gWadXNaIf0KtUUUi4sMkycZrnO8QJtnaQw
MXChONljFeOdzY0PHB0O256J+9xI55wKtU13xXEBOHDtg07GY1cUrU3eALR/by3C
ZwjnKTpsvQyrUHo9PehZvNai2oEqXQOVrmnHFcaJ2flqAcccJsKKbcFwWJyS3Pki
wO8bN6O/RsGE66torP2xbzay3/bY7fAr4EvWkIUOJjP/bsHYaZPOhzV7/MRtY4Uz
x9TmFQ6SJzTwT4DUUYGxL8bp5D6oOnn13fxalpAf4NlbFMKYRVtU4y8C0haBBj6K
14imcoD33B0H0t0aq3bgujo25GgENzEizsCqO8ajCdColHx0EsQsM/En0F7qUg2V
JAd4Arqk8qzGF2y+7iwzIOA4pwjBUl4Ic6gsi4E6nDPSCOPSdE0vf6dXqvHy9yYl
t10cR9JLLWEnbx4X0EsiFenZfxhvTRl9S97WbDCl5C/WAVjJSMZxxdCwGm5zU3vi
oV4nxbC0zXGzScKOPGY68ZAznEt3UbgWawbsoLUdTc0mg6xANhiBLCeOYNwKe8RC
mXeIHYXEzonAr9F+GcPLp0a8XMVKy3QfPFVCbstBB35Y3YXH96e2A+4bXjGU2K2y
UImzuK9EHBVL3JIMG7TczFK+uIXR/iexA+/4pqVbvBkJvEv4mtmt25OemFOK4Yzd
FuLZIcGU+eJYJ7ji4/pejeQC9oTS/z4+hOw/ENDlaNxbrhpLhUAxupA1P2JwC/XK
2yId+VmVqS2SeeOS6Qpl4WKwU5JmdEEV+M0wR1e/XisFFgksPm9CZz3i97FDyd0r
ca83etRoZJqXR5tQooikqEJvUBan86lUtdlcLQrfLMP3rzBZKP0op4OiPRAHzK3Y
3lGMw0wGf0blKwoxRVBcH/VyAXQVP6meUpFt8IX5i1Mslc3kd642NnuGY+z4Di8V
LAf90wS2d5lPykoHZ3n+RISGvM0DAEbzlWaF5y9mC0/h50Ylb18U02dZ4e+PzIev
D5lH0i6ie4NRAD1hVvwkEEuwExDUz5DYmJaK2maixWDF0Y2gMAuzQraI4uzENnwE
TXwueLicz0Yng1tJaWd7uXYuTkMCJhoLjrPfI/BwHpvDeDlDbO2IjXqJa0xskFwf
QZz/08YdnTpSFKXtvKB4N1/+sihiHrTMGtDUPeN5IitNOyPNBwLjT3wsvngXdQy7
oZfs39tu2tNvPz4xpiWkgEUzdkPpdtJOORY35hjawSj4BZbEDdhrW3mSb8M7pI2Y
ThfNxuM6H8y56i+l4xkzEkQ/V+SLhnpkIY7loC/+op86TtnWeXZT2XZCqOyK//q8
BAX8mNnItVM1harkPMBRacFwJMMvRR+gnVUOO8TGymgDSrztxVM0jPtdIYKo68Fn
QMwJqC4yiJo68IynIZ/db2ofxTRaDeAW0xdv76qkI2fp8HfrsVHDXmcLr6oln7Kk
YuXzUbJYHQuFZXW3yXEuPHpepu5qJfQxqqoC8SlOXQqvbQVKNNJigOtNq7UKVQAo
t3EpRLiRNp7kDTTtvw/Ro2YXeB9AYzjlYuTE6LCoOQHzfkhYsyH6//bI3jNkfTDj
i4/QGa/L4ZsrsyYK+su0y5tp8pC9iLIi+TJ92oyXKRrpb3frgcygvW1ZcSxbzYNM
RUXDRwsVDXw4/w5luhwDPVizI7I5r6PCx1KGpHBlGI5XcMyuk3FBdI2dxTtPNVKq
uMYGlfFW5XGge7CHRMP2flMZRSFSYvBwat6QQNzUEQUgAPG1TYVvn8o5NIdYR1WA
knFaf+8cqyQ0YP1j15iiWzMI9uilO7UXjMcejBJxIvJi4PZI2WI72BJzRtWwfMGP
uHwyJs7LPHgyckSDvb/vfYXwLqKcXk1vOUotUT0eavZtW8QlIhaNT4P84kP09iX5
35kNbriQomGdVP+nwv3KSBQbiTpq4YJM73kjwffvOyLyakC0+HNm121PRof2nu5s
9C8uqOLEzcPYgc+5E3aCVQ5wK1v6/F0X82IYcWVRuYcZd4QrNZh8VCJkLjDtw0s9
bsH/fw9oKp5neuBreaHz+xacGc+Z4a+n3Zt107bt/tO3NSBSCTvHcuTW1CzyIrCt
Guyuh/Erqfgm/2U4++5w/x5bLUabMtzqy/bTvUk6neAPD55iwQse3Ak8Rf6PVqbU
PrXbOt+MrNbTqSSZb7Wm2M09NhdwcUsAT5gI3VfsEz0F7dj4VBB9s3kZjB4iKAow
QV3LC3H9GNHWFRDv1zRfEwX8jygDZNAkdHkGp0zdxvt+lOjZ5Ec8TYGSLKONNa3E
pRaaHcd3KnAllUs2i50xjcGUjf00/65YnI3XIv9HIqxo5jIJOuXIDdsNhohvsjcL
umLgzhOU5UW0moxwq9H5AHrGT94DVSrBzVSUgbT+JvApVMuO2YKrTcJAVVjV3anh
eeN4PT3FvYV2nDNQyupFZdQY0Ux2oqAL+PLipdAkySochnUg8C8ibcjkh3ZqBT5Z
ks5Q7/F7vU577UzXmYq4DRW16/56CluYWSbVDVKymID+o6+uN49PN6gXAsHyOESU
Gb8pSeXh6+hAhXX223w9hG8XLx40tjtVqC7VizpmFT75gKc25dz9j3cCy0UWC5a0
1Zf3zMVGZCbVJRlIqChQ1Ho0t+jIwBb9WiEuZSXXpYzFLkZtn+e2qMNq96mGiSrR
qGYgJZLXuxO81w0W1eARx6qWE2QZfIt39W5rtm8Nf82qtIZP7D1WE0WK1a5X5vGC
4n5wzHrtHai+4xjq/RnPfbXGFtzX7Wy36C8gBU64Tk5q6reOwo6nxqGTU4hZUJiY
rokhok7oyxVqIjDE3ZpdEGUvR15Pr0CQ4suXQJnoIONEMRB1DxW+jakSLQE6OKcx
anb70MxgpNzDOkIQyr1mUcL7bDtG/6eWetgod5BRcxrpd3H3p8hs1KvTCYYetPLI
2qSafLZtcVqoqbIszJsc63PbHRvP9rvzR9MHl5KC3NlSJoVWu8QBC3LOsmiZ/pdF
tqMbm/DLYJYX+UhRcFTcIjyH8ymRF5VZ6I2DpPE9BYjt+SDucfx/5joOjQkeFduC
q8N1OUbBZWp6hwewbNDBg6OeN7D3bSogV/5uM5LnRm17llsSRsMWBtOCyotj+hrh
CVJtH7HIq/JjZOLmZ1AJcUFkPLgzbmrwaAeicQw4Bgi2cKoQM8RnpHCdrIfMKHqO
WsoDdlWvs3syh+k2jeRvy/eTBzqFXMcNdNTkvsf2eRVlJxJKqYbtOWud+OciV/xO
EpvnoGsZyt9U162P0JrWfo6Nfrn6RCyGOjRJ1LplIiwsr1B1viDk9fVUHbZiweKe
gP1INKhp41zNJKoAMVnam+PWWatogoBOKJrjKr7N7dvDCsarwOH274P5ugEUvJzu
dHJlj1Q6oTs14TNoAG2PnlyJ2GaaX9ehx0+0D8ivwST/tf9TRtHh+7P/BwSSktFD
W4j8Krab2X+dItLcNmb1O6LQD0IohLw7u62Q6ByuUw0GHJUfh0rKRYf9VJfv1i6a
zmoJnjBdxZTx51711+QrLLncExPXr8QK29ygMJJf+PFJrMDZe07LVjlSfrJei25n
8J3KJUgljyn/KFQouU2MKtSkJqIz8LsyIBQtAySfqzZjWyXaIVBHjCnZP041Cah2
OB3I+vnKmlKbyxgPcxuLfKEBzIkT81jyI/KbLetOX0Rz88qykWN27VXrBUfzjWRi
usnWGmp+K7xbR4q1vabPlaz6HYOKqM/ztd6unASynmbzNc/az4FjwXI5byI4qvfl
QlCPVA537KTtlaIUAiqmuSmRBU3cJXKVc2ej8SfnJuYTYwJvGQlvfGq7WcjkhxvB
/xs167SpztK3PIu64qM56MYuQA5uDbEZp4udjmKoMltojkVIsuxTcNuCge0yKEu8
18s0gfY8I44T0p+ohWOeJ+ETD4K7xF0DasXlB5Wb2eiziTvqsXdxOhdidgLt5E4/
FxeBmNoejSFfI3LqDNqMSRiiEc8XY/za92pluRjyKhhJjdun1xW3vRVugG2dKkeL
4HdYZSQKHeI5G/lmeP1DVJYs9TNtjx0IuhcTQrrr059ToDbNykwS5AOweGzTryfD
rGTwR9LheM8cSt5Sz8ku9ERCiyPblIeF7M3TS0DFuHouhA/wiWHoVVNhtseOSiIz
HFWkHAekOM+zgXMwILhg4vAObyxIwtQ/gwVTWmrH7ZgsdKkDdnkIMyNMVzie2H3S
vA35r84cOXGNbpVUU8ol31Glz+qsstKzGREH561PfS87fi+Zr75aoNzWh1HQx2KA
GU0NleMta0qYCUj0gFGB/CvfsJhD9CrZgmR/5pGzqK+M/3W300E8s5WICl5t6ZF+
BOeKPzX9h9wKdI9qnI0y8jS9csuVvAjXDQgDGTbP3AuYlImW9TzSVNiBZj5eGW2E
9BKTsa+EfxyuHGUoGvJ0xg+pWVgDfQ1OX7MDYEaJByaKVcM45CRGmoNJ6wUO4NS0
vqhtP3tr1bUC+rqJAYvZ8xCi+RXJlUKG8WxleryBfJS8lpdx4RRq246dM9HLdRru
ELpC/CiqN13rPZOX5rXlZXhziENOeiQviPMrmpBJ9AMxO+vmVrK4WMyJ88DgFSFw
cyCC07dYQ9Rb7F7qCQZpNGdWKv0odBeIr1SpRkEUx10hfjpvYk37jt653BZBnaL/
yAaxRpSlSVS1Dv5MDbzRNelMckjnIDWp8WrMWnIIRQerp5aScrNk8CBrFtT+d9Jj
Cj7ebMPb8pMzvgw3UmLwA7X4OAiV/HC7H4/fihXP8K0HOE6VZxxB4arCTMufZI+d
+TAfOEV4ODJLys4hrbyZtA18GCnBjme1h88aEWNNibDwsvX2g1a52BYIwnsCsOFR
19mFumbpLZziP0619FtutuHYCnjbOI08HC3skFLX8mcfxFTP6ycm8EWSOYp552cT
39dlAnRklm8vMqB4unCzUqNxOc1pSFE9jFgV9uNL0w9Phm7MD1K5vI5VT416KVgN
0tL1Igp5U3iGFIJjBCBexMfvUrMv3h1QbavCcKtH/gQh4g7c8HS/ihWeUbvK4t0Z
5wSzAjwTsBSHYWJrVIS/rrzgpei+AoQUZAjM3tYEvWvQNIbGGQXATC6+QncdH+eM
65arx3cbPnf4De07Em7GBF0Aw7G475icr6xChQUG6ThqJeX9R8FYRtypR1ULdSMR
qoyq6RlwUAEdAQmwZhPTXYYnEQEXDvUyUlAG4dK9uUz/b4zsOQt4GMzckfkUSm/O
YHbaP8uEN1iU4+OGwVxfT4eFDFTxNK7BkC2nmPJKxz2jsRRPdp48tWCLEckOfqY2
WtOvQKiSfG9Nd3DNlqZfpBctENam+7Ft7SK9xMOYBw/q7emUhpexScGHrAapdlTo
rksx3q4ulusw/7U+NDSjibdMqBOx5e1Yy0QUt46H/5Ty4H6V20oIG3SO6SF068uD
ZGEz5eunFxwuW1+SQRrSDKgumLiE29j/3IVQgliKaUgdVRLSdK8qQtPvjc2pzikM
kYHd31sN4eLRfIDfGI7lo178z8CcGWyS52vWCW2DHrnvJnwvqRLwbWoqvsLIZVQL
Gc6fng1Ahr9+wiVY6lxi+Q+8vezFR4LY24iHQyily30Wzf1acoP7A7l4CvlNVZaQ
7Ye0I5EtPthhaUKcZaslxLMGV9HGPMZeGR+daW7ucDalcaPk22hh7HcUz2uPOWCx
samMwNeqpiMz22AKOoP8V+dTT5LUBIzd72m7z1oeBpZWPHeT88DmxVE2iTXQc7n4
/IDbnAM/Jy/UXIscOPf1/WrnW5ruv/FHngeEVPh7NEecGcoQw4121unsNX+9gqwM
J+D9tBKhjyHjs7Wju/ywqMm7NsuSZ/1NFZi1o6Oxoszfw5qwtQ21BFPTVMGywusd
W/Q9zaYBN+oV3Ekv7ilOhBeJjlY0hANuzhxnN/ZyRppkw4m4xOcF4VGEutVl+WW8
8ype15sagSFU5Is8Zrjj7KgbrA2LMmbKJG3kxLCUQSkUHE8Diej4NlG/sOViZkG7
PxWVG4mLZ41GpRptuCte0XxifmacTwinFpi8BZnXI0/D7OfDhzxXS0YNTbiT8j82
8/nm9tpW6hXqkO7GyWp+5HtlkPTGMHpLRXYQ2l4fZuB0Nuq3vkb4P1gTQvJuzqyD
daxphqu7shmBE0BGC0h80BiJjb8ZNelTrQNQ080TXDSgipn2DRbUGByLLUM+n3Ge
b1KHKnh4Dsr2iQUVn7zWpzXydo6tPmwA0wdCEQVFu2eR/pM4w3DgQTeQT48+R/ZE
w4fhLxFKX8Oinb6nmqEwrYKVEZhbJuCIKZtmemzlG7pAfpuM2rg+kOX1OrONTiBg
C9JWOKHSqEv+hmk+XepSGlmI1CF6IdbnoQtjcU7A3eDlS+E8SUZVBdjOxyS/OtK/
SBFBg+k0sI1M9HD9RSAmgS5FpO1Mnakk8DU9Rk6U6Tuo5bYEsJv4LeXKZrgDo3dz
XuxrA83qgwMYT/DTt/w2SY70xtuQgR91CK50+dvtd0PTzVfc2eMEK6sEcR76CnrU
iw+PH5bJRprW7Sdh+m1rPYlMxF570CV0Rjx64SMOxFKXEzkLymZgP8Nh/gHtzEZ4
I2O3qgSg8PXqmRFFO9XtmTHLAhbZ4nmqmLh+CiuCTtINT2cX7OboSjnmvoUfZxwR
/IXJfnBj6KkHcjMbpWyByPR0qHrXBrgW4Kt5fTTzLTFep0xWOj1vLJUD6s/5bXSC
rbyRy/QtVcL+nld4wa204MYLfRClQlmxH+kzN/UjI7RLrADdOzNUZ6o+RZtWVD/Q
rOQ8+2FvAYfQthdoWiR1YSy16hZ7jzCGEZnp6j5m/3wuHgR2nzr5PC4Fye+Eg70Q
UgyA8/Y3i15yToM5C8VSy2I0VJyh4searAMj0bNmi+iB+NyXJfB+8H1rj/z24nmQ
cP/ZMhmn0JNwoetTUOieTNMuyrue5rPfCRSoiYYxFnfOihY5LqPhLYQnPj3Lotc+
0hrE0AbKWLD13hPyoJaxs1eFso+T8QKPeqtU5WuTWapCKe5XVY8JEg8RhriNUIPA
PiNhyLeIrQL2KzEB7ac1hl8bD/YSlY6oJL1+FLDr9V8X2NiBM8UOjbO2NKxGIo1E
DTJ9F4pPF0VxFnCKkhAKAl5HM1g1No6B69i/4259+h6MmlT5jcxBVnvMBfL8BMKW
Se1vXEMCP/Vq8ToL81BhZUVO4dnsvrwE/CVViqNwE5aZVD+eJQL/FoTROxJPV6C0
iGyWoJH45lLEtHIaA4sZbLCSVTQtqm/vTyfCUKs8wNXcOTawh4I/wT3uJhnw+gJ9
V/FWe9J6fvd+beaWRfd/SS6vDU3iEX9SB3C8FPm9+zWjFcFoAnvLfJ2SQP6Gpj6D
lnF6Vf17mP5Bqo16E1oa3mfYUzJ4rd82HPTBsS38fOR4OQtci0AiypSz38qbyqmY
BPWXeFhsUX1Og2UhueL5tgT0UA+iL0K0q+OLd5rEX1exkxPSv+8OvskONiB5ZX91
tfy4gL/QcZPNAuSaDTkti3PNvWmCVsTGSUZ92Pcmet6N2uPtK8HRmkTnRSPMTaNi
qHzMN8AbrQp2a2o0VAGfGsnF/WHXj0cPlUWbs115o6Paa7tNBA0rHPGScS0Sseji
Rcse3otJ0conZN/0KhN8RtMxBcskIV8M2oiKpLIn3oJhDlXGtMsTje/HCTZZ0BwH
uL1jRZxdDrbJ3FNKX9KZ4TnYjiOt6eoikhXybN5o9WteSFFZaEtf4luQfTpJKtm6
OD6hsiuPhGFYKUqViv9YewuiJIc9tXfYaBn5DElQySjPvhWnkYaG/GR7/BSRU+Q9
JcxFR/51PlHBwwxjo6WKaw1uzs8HMDgl+ot/GCCNAzWnYm7O9hxoAqUeuBPrqp3s
LizGrYaDuoaZ5cAWao5Tl/yPJWW8JI7OpvOHE/piDAq6/NFWOCnJyaGyHE4LWgA1
AIFytMl/hAMWLR/XkdDUlqtzBw9EDtS9KDi3n0ysg7wPhwkIP0FA3d9PUnYk+4yT
ablqgZyj4kO4eKb6ixsJ8Oz7/Agzwgr3X5ycltvnPSrJB8KrzN+X+ux2tLpMh5kY
KxmWJJXUr+nDvCUJkQ6KjgfE098GSOLaRXaIc9gG9PUFgJPabKcVIxmkzi66mSMd
lRrt/GrldujChzyCsdRK3s4vWMt5czVpsZ7StjvtuqgufNYbjHBVmpPmwU51AlZY
DbtKQvhzMhk35QmwV4eCV1Nb0GfYjwLnCqUFRPhxKNnwywUiPOGghXu0wVuXOCTD
uXbggo8zJYJb43tl6VBskS9hIEF8Gi9doiUl/lT9EgDtgbAJG4UeMKOxy5u7IOgd
Xr6Q6qbm4FFe+Gg5Ddi3C4qoxHICeb5ORbIYpLUR3V+MayauqZGgye4bvClf7kmw
1/V1VIlP0vuR0hAWj0OmZ1G9QbfT6cAjW802ELy2ZJkmiykCPnoGbXmOj8lumdbG
DTEHeErEoZEy7hjClvY3ZacSCQPRKpRduONkX2OBS248PkHApgsAF/8jic5t0XFn
H5kV4uqrlmNIAD3vYvagZ627wVQALzSfZ/7Sq1xMT7tmuakCEx8o9YT7GcqM4Hd6
AzLq9wKcm3D2GX45kMNj0tQAV73Leo7KBNqadaJnQXSAj0eIPfwmsfc/IC24QY9l
V/VlqdUUQEThTHZixque0/Y07LxD4w32biGEFwiXRLon/Owv0Oy+TeReVjB017R6
dMoFprhLaBlY7YDdG/7sZZOERJ5FeB7iQPwgvdzkJMTL9+B2WBZYTEOT/wWdPW+V
KfcigcrG202Vvo02L9L2K8ISidySNkzGoYFhUIJNexSNQ7woo3l3wNWl/OXN+UpU
qZMMNYaZbaAmJVhepTMHWxQ+KrI/FYm3WnEfyUFQTD3MOpps8HTowDQ2eIU14xgd
4jp4oKAtRRHHyJVXveqZde8lcRouy5u0vyncnb8hVtfdYf4GCjhRr2z03p1f0x6j
H+EIc6cDBeku5QB14peJ53mkWhyFOpiPx1JkFnteR3lasQBUQfNBCICFsKCo4qN1
EfHk3i3LneCD9SEKGogAGGBQvBC8UNkjg9lYzRGPGg6G4eXnJuaoRE6ulh2lG110
/UUSaVHwSlzMXHYBr6hrFyHZTLqAsyvdurIAaOXHnA44sGFE2FPJ5qSI+VFGQ3Dg
LffSkZIdssurrRULKIcNrOTQZxJoSqxF7kL4H+DrwsWzWZAyj7PLYCg8mGwcit1g
qP4w1smUyxluUdDYUInDKOdQk93y+9b51hnIii1bI8t52eUKRA8wSfvVcXtWFeYs
/ygFoN5d0mRTFkXbminz0S1u1Qj30W3/LhwOpkf9c6yDggi0sWUseU+LYe/ElLy1
6xsQKL3hGvtQJJoJlu4PCsSGmiNJPn6k6KWym+U3+PXSycNzvAyXR5dHBe0pOCcP
i+K0Bdwp1lrFGaeoBmF2QbD2/Nt5m5HWPPv0IERac+1W6FErzkHQJZN95mOe4+ZC
dilw6LF8S1hIbZyz6aZhL18UeAhcHRf7Nlds/rpXm3V7/uhNjHqWQPbZQYPpK0v3
z0Hgwe8dsxUbD4Fy6Gq6hv2Dciww31ER9syPkekPpc8HukALfwltnglNBFTBIptd
hCsWMkXBUiys0NjvBcDx9Le9XXzHkKL55e/jisxyX7tMm160TQ1dYmt8n7dTHTon
bRLxLUYs4z74ZxQs4ahzqEPJQeaHfbnj6UHmDGri44+ue1bEiAj7uFFZJk6aGLES
y9ltAYXLFLxjhn8784E564J+0E7X9e5wD2ev+DYquBql/K9bWDGsoIwAgQrhoLiy
/PzI42LeNAzbhojnwEET2QQ36F+ykPbQlkQ9XJ/bBG0oBUdLYnNhjFe0hf0BQaud
cQu7TjYW8QfxNqA2G092BBPwJBWErVd2vtrzd0vCqA2jHxAV1BtIp/0NgQHwT8MS
EBowL4tameN34NJuCwZLJrf0gxeiolacfBaMBjZYJrTemMIq4GbZccnNX9C84gQN
yANIn4tboHfREpuxD022INRV/xbm2j8qPYkgF3So1VMOeSsfgyEFM8uEVGIvh/C6
cOWBWHOtc6deSS++4OjjyrQNxR7aiFebLewA1jm/dE5uMhknllaxkKUd/IMeb9tE
cIJRV/Y7LoR1ewDMaLm4Yu77b/2GAY+iUdddn3JkFaSlUKEIMJyLKXJZJeX5Vedd
bFPxK+l+AlQyjnKNcpgFBBAUAqWj2RafRBn2+aagJnRpOP+54e2j/NlQMEDrkAis
o5SqI/7V4qLkdqdfxUfnkp3YmWndn280V9wsXl8egpavDXPHVd2A3CzPTfy+Uky+
5AQ1bvN3+f7QAgZh5L7wO1mnHWZqxF5tCQYyr6pxsfO3AXYNh5PNmYaDdzYYUdj2
aFFlTB9XaBebm4KB+oOZRAiLchr3iHlPZGZ0UBLY174Z0TQf/noZy5eVkBLJv5e3
oyOFaP4Vb2++RTwP6tWBeSMEmnOm21BDw4fGKZbyW6y5k6roq+XvHFW5u/mK62yx
HWi92u0UTRKugPi1HT3DWpyKyfT41HulFgOQM0JbQ6EQKe0zfcHLV0zS+Xw9T6BW
S2/CZh9j+HGqpR0hRdc9pAktltX1WJpnAnsFkJCKsukZwgCwcQJkpGAOrWn0EzSQ
nsX/IArE/3IulEwEsCPvPCmkHNMAhJrKiK5ZKXKYaoBtevPmcXkOrDYM2uztDWR+
XoY3/x/S/k43AEvjflhmzyBM/BEVqM5lohcf97s6QtXj6EHDzKNAOxnDCrtguylp
GFTiOWcuzFTnGHReDQm2E16zMbfaTkNtgxjoRto6yALeYus5XwBJ3+krlnW3B0cG
b7P96q8vBtHeNPxB/UXDNjhXFFBJaHV29DQL7t6Rt04rAkTGSLbU6WdLZBiz+Hl8
e8RS+rmz6Tjdp+Y0buaL3ttJw8hs0hgb2XCiO2D3gdoKadMwtXyNJPnuAZ1UEWyz
ZWySSb2kVF728NOc0JibP03BBOy5v4eAUvNaWVswepCkKQE74+AdR0xoI7TfjSGH
Tor/0Zr0KNpCNpafq1fPgBjuWzOgpEA35GDFt0SKjaX10nwaDavOxE9NnCEj0stQ
OnbPmFy+gTMJPwgP63nA+S/ovhDb96NXxORdcfBAOEpyfOFSJBCJZq0VPqgRQT9V
L4qRg1jHkR+Kar37radqNwyVzHXDwFYlwACwluDDBEunOAc+mVqTuG5gC+HdtEj+
HOp0XcADvfeEq4l84dPi4+k1oJwBPJnffvog7eAAhI4zt/j3vDAZ8zanBRBre6f+
wOQemQYQ9RNTzHkR+fe9Gi6dv/vHYuXU/ienr6pFlXUlOojsRdUA49nVBrw+nx/F
HilGa2xilOKadyIGwCf+1/7hIGNnlK0kxnOng+cpCh78qP2pTYEPXycekRLFWZsR
IvclAQxLFAb/xHTSq+2Y5w+LWaQDXRLRn3OeUECeBcBclOPYRdDPDN7NVqN1EgPu
3s1WzjATTPA6DvWZ6vmSxRaVfCCJOs14sP4+QutM2q+QfN7n/zeoa7OikZROKmT9
1HZq5HSf5G/e7B1q50FxYjJxRqyN+c/KP70ICd7c7dlHk4yX4T9IGaaU6vIz7Ejz
U5Hd/EgRQSUVAVDlyPRCMn0gxuq15Iqrt3NSG3EPFIQeAHUypbs+DNmauJyO6Qou
zDN5rHACQgphnw5HJf1aw7N2l3oqUiQuSxT30RRM6EHCnf+uYXOfCf8pNMlT5Gsh
Ji3JWWJOQesQ6WjiGrZvsgV1rViC+Xu2t3tw2uqALq4AxSjUw+p6eMwWamdIGdT6
Q21gZfpjdeOecoAYtNjMQI2JT7UG2BO8nVtZMcVGc1MEZz1++XjL45DeGa4xIYVW
S32cHtISnXvQb5BePSk2RU4ZnKgki2qdXqAIDYEjI+tn6B7NdnPwPI7k3LN55BKE
xN5akstCv1wv3q6Pgb/gXFBV5245HWA5h8dml4Kj88cQf5CaymOZ4EsgaAaSTlO/
qtQrFNbtudQytD4K1TOCiCayceAaCdc+NBzAEfz7nJxoAzoex6tjJgV2jOzYt5iK
Fq41TnoDSpPKu7sfJXo6rL3QlHCTYVuVMphx8QIp/82eizI601D2u709XxRBgL8C
FkiLiItkU3ks4GHlUKYiSorE2nD/n9P7mGKh0LLcb4qjiYdE6aq6Vyu5F+h0F36c
m6R0H4FkChvXLASMMkmFwWFV4n1o2wDKbJb5ljUjusZMO2CNPIq5xgvmkg8Sia2p
VSXxvwkmiwyFnilwcP6Bmx9nZr5tsY9nYFYhCW8aJp0j/L8XO9j5n1yxGDaxLqS8
zsi7N0P0MAh4DnNp9M8DhSXZlXGYHj/fpfXLddc3KAnk6y1x1/Qq9+CuCEsqAyDV
m+uzhvvXbJJyRMXEwAm0ogFI3eM3aIkGY3N5vHKomkMhsgt+zgPYAUniVYxSxH2s
NFjGogYjhKohWPaZk0X83fLNuV//oTmUMyuQanQiDmgu54yTPQLPIQH8CafkpHgV
46hIQA4+yBXlq085ZQF8zQ0VMCGYl4Bi5qXDV+yhONzDd32l/aIoDjYBP9/AXRAA
NUjWxS90rTNFdJpR4kYLsSDQK2J8vbLL4mJ2I2K93LVdDfW6ze83X6M6083iB6sz
Zx5pIGE/UIST+Z1poC1KBtpsaWZMiQkc9g2LvWcGSE4DpslbCaq4jB69RDkFEc9i
pFZoycBq9crpMA84RRh3mIVvTeqTqKiTgI+ifZhOAkOC2F1dM1i6JFRYlS9sdXSM
0aLI7zfBNZz2mnik7nzeM0PyU2XN4ge/bqF5PvQH0ApDSQReOBi3K5hMQrr8nhCR
2dhCcPduSQuhc6u0qyulAYo7sj5tSVb5kojx9dZyRC5TJX6AYLEV77M2Q+MHbQOQ
Blxyu5AXSNwlZBG77KALq/Z+YVYSUwiSPBC4ZHTQXyAu0rucFEdKPkf64m9mb6e3
1p8lFixz+UcWgaHL5F8nAzwAL4xjzmI1GLY/4+9LfeG3gFwO+c2njMcTDlPV31jn
27N4AoPTumwqfeT96a33hpK6iBREFzAT2wWsqWoobttD4hMQNHS3xPfGJ+B/haHH
2Wq7tQpdRXq0mzpQNDvC8pA9h23/q4vvPGDWqd+A07tc8nXYeK+Sdffs75POx45/
U3TLsGdCqF171kpwG4HgsdAB2+kVipLImQf2nLSW3lZ/MhyUdvfXz1DzQ8HNIST9
MqvI/x5/ArF+2wPagaINKyrfvs3mm1yEJMCngRiw19LAtfbtK1zqNLYAlxRvmHDr
H2KtSDJoU3hK+iAT/QzHl1HICOjoCn7s/Bs6zjF7TwksSOS9OZ3JzNYDrT42/olo
BYVdnFt3FEZasupN/CKJKzld2rkg0mc9fDaRLDsvFKbXqFqFKZHeMn+4710lQtTB
1pjbpE/3VDV6zYRHL+xwppNIy5DoDfTsO8axEA3Ex8kRTXuRA4h3gMOu19DXX9dY
EbOR8rUD0S0rZZivooQe2nqzH3uLz9pMQWi0XjJVZzEZasgeK1F3X3DBwaNbtcvn
Tvn4+vP8Fpbnnv+WofpXw8wVLUyYNy8bFKk032p2E7XgVrUMqbBkwsvA1sywD6Lf
kqiK79Tk9EhCtlbi96Gp71jmy5XR5kR2QEfkns8IpAZ2aDX+bQcJGxqiN2FSgJ/G
+s0uxleT+TpzACaDU2s7nVviIFAgjxWpFHpOxSgw5g16W7PNWff3wL7rLARlEvrV
H+PMAPM/rsDEx5IBHNgs5U85TDbw+5g0qTKI8iCV/FJTPMwb7qpR97IKYUDoNJdT
fpvPtyr+btFQY22DDVAbfsJbSOnf3E6PzDB62JzrnTcvp9+YXNpEooguYo0BviZr
jZmJO9TesQRqjrLBGa13Mbz06f6hpK7XydIDxhqdk2eD04Q9SibOvGS680HpNfSp
hkDfTPFDrLFKRJC49Xb68bTtwENQTtSDkFC3hfscegBiKbj1jDNJMvtw9ZH+Fkiy
78pIqZKV+sGb3QHZvEFQrTZcQ4M0zS4cJ2uNiRnuHR/pbgR9fz53+wt09tv3W1jg
bgyN4P5Rrs6eZmcGNBwfjtA+IdZhxBQc3BKRrIq0SVgbQ2Kz/o05wjLJzRxDqDFk
YMOgdc05EwhhxROIqG9So+Cb7stO3B62L8JoRNosJFFugB9CZpK1u4w+pnmjW7I4
4U3z4YeNlmwPIFT6W/+jugYnu6AP5Exsq88IYkJEpYJW+yD73TEyYAzRbLmWm2r1
XzIo257VQDNzVmFcXFo1P4J+8cwPGc6hF9UV3T0i42n9OSfO/39TnEcW5tymwWLS
vKkwquVKpy0EpfJLzF28x1mLWZ9CoQRWT1qVPMlMrsogyrGRETAl4VMHizpws+2P
2tRctnXSZUcrCFOR0V8I0TjTZzlk1ebqmpHcFnEwvPTG2uNhx0iVAgiAgWA0b/Ay
M8MPtmrf1eKNefhb5QMxbH3vwCmoH2lKFLOkYGnHc0WrwfxrnYNMCTCg5l3ZPOIy
0ZAUb2xR2RxtptNUKTg6dzxiXMTYlMu1SMxnSmp84VSHwj5WCCK8ncX9/sQ2IUwc
0qLi5Df0mq4bpT9kJ8qtmOc80quSKoiKznN+xajOzyEp7etdmzl2tGxY286xBqaZ
0ZX/sLUP5XPv+zW2oCTLV6AYfb53pIYub/3rCXWxs7nM7YZb0mrizjf6/SOB+KGv
OTEp+Eb5Uv3l0F8qwfez77XXwhDMKenYuxFEwb7Xe/vQMT1iBVK0eCdvwH0pJfyt
7Cp2pEqVxpEWVhqO87+4f5qzQnKDJkHJBvaxDeJgkHf5Uq58jngHh5BMP0CPggZT
QzI/fslpndLGOhafvR33kQ5gJ5Vvbnd3eNCV0YQFBNqreMdXaDys+mOPnbhUYwFD
nwCu3Q8ofgS/+KWzY3vP9Hwq9EKXFIx8xLnNLLupbIF9jv2REkKbpHA6m2hR3uz7
qXPE1jCQKARfN0KSr3gkMV6AGAiVR6DxBb0U9MY8L7d9o8eSKlUvmFG1Edm6Ie/G
6j3jyvJtSRzP8KSxOPnO8B1ngqm8a1jh31bEhYu/OAaqyuXqIq7Dx0hgvK51/6Ny
yOJTPhMWL488LAZKcrw/gcGsMzwyPoMARRlUqZGSH3QGIinhaIaA6z+mNxwUeCLR
DshTC8DFVRuhWmBYcRkTf8hnfnUqKVqbu3SNULwMVfYpaQGkV2Ex0zUpV5gjyFlQ
Ef1akCQCd3z4mIM3OzakcAaR4OcwQJ2Uz3QCG6sEOEAFL2wuFDbSATYMbzIemy91
ZgPCT2LIRBEIHIv5ui76V4X+0TiqB5IQZD4gcUSc7U8noBejYo1mhlgVa6KT1emc
/HV21YVe99j8jnE5h0hm7/tkv65GqCObNdsMwoDOrBMHIpIlBSr2BWMQJstEAD96
fYJ/8R+4SQRllF4XE4n43Pirz96o32u2KPeRYMvQzp3WqlfvgkP5UKMaWnxyb3St
iqVP+srlFCLUCOtJCYf1lriD7ZO5G22HiVoD1XwK2gNzmCHJxQQqi8IK8ggphF+e
0dW6HNS/BvprN9u1ptfs6ezP98lTEVgyI7iplYnH1oMt9QRW0aFTS+JYxoMWaXmC
PHzG2mPu2a2/s/S3A09HJ6iShMZky5DZNwsuNIMW2+iDdVZQquiExM7TwfMbZApu
2w5FxfcgaFD7XlW1UEAgcFGMhEAQZEQT5iyGWt3KPXIbsjekgUr159i2Baz3/5FZ
KAhEK91cdzEz+iIZ+6/38ha+/D39/SfJsIr9LUlk/Pg/eHrZsmr3nDc4XjrOw51X
4HHAnicaXfeI4PZwQycpk7PONnWx7SGUQX7EwVixhLqqc4CXg+xRbDA5ntDL3FFD
dmlif4JZWasdFFNQ5NzbDeE2vaHTljhYWbldPncEOscVYv/z089zqw46RzoP9dna
l6NZpyxFDyYsF3ZQYK0PRhfmp6hIg33WaMS5y0DhZWOh41aj0EdqYKU4HIdE0RGa
A/Z7yrTRwUIpWvii+mE2G/j9E4hydl7Vs4F/ZSl113Wd5jeZDA5+aSoCyoJ0oJ4/
jDXHycFqpSNn3cAADDW8c+IlbTwScdXURgLZFlijzNMIFnCNoKytO5zjcIbR7TnF
pLmkxz0CVjm09k5LvFF4mwAMnnRcNWDT0hJebh/wDiYgRzh8XeiydJJm/55pBLUN
Leu4HbrKDRizYbLMO8v4as7GwffrPsn5VL/w4Ju9lM+kt9jGErYS72dhL445NOvE
FdIJHwkcgiy/5hkIz90bt27lh6MPZm9J5mN3exsOPveN9rN96nIgMth2lF53BvUU
3oGzholJsQHwKSVJ+5zd0oiB5EQbmmY6dqUMQA9McBwPMsquOC2dWDmEQNRKiUPf
U2WdL2bahkGp3MBBsLPmID1YYwgWK3mmag2TZIfQt5Bj+rwdJNR1WgcvzZ2q8VS6
LcVt0n2CDwRl770k/KwdQpwRksVWV5ZGHFPOmuyrhnddJ3zeIpQ5BIRnWJHPwS98
ZGyxaToq9Z/CQkLDyugddfw3dztCxL8JP7ZmVClQjgNlrWHCL67EaM1Yub6TpeD8
Cl8T+8AGTpqNhrdUgIf2XPA7ULbPDvAu85D+p7eFoK3USuYIIq2yEcJ7IiRwkL92
5ey2TLlmgk7U/vkYqMGAzmzhZouQvcibGobv7DqncqYX7y1KbFFS6GpKnQkRpdlD
I3DMsJ+kLBVOMAyhELgsOAchtCQT+Daf34k7ERrasLONpguUhD7Iuz2P5VvxdzMN
hO0IrzghaiCWLqGH6Muy9a412M53/HmrwUni50uu7r960svVuVw3q1V9bgIMF1Uh
NoK/SyKXejDUQ2WO/02tykC+Su48MJ7MHizy8w50mmM9Nj/k4OTCZJKETUDTQeB6
btasPBFp0GTrkk0sw9hmbe1x7ryC7CqjN88ljoVVpBosrAzLJ/QawuXkq08GuUOw
lpzimgn9poaTYAZQiZ+acNfYz7eaMG4EeVWNVgFwBQEaayjXS0yI3JKg1MEuDva5
P+twv89rjURE7N07U1sehvCuYvlU0U0uhb8/qaLBIcpQFXPt+49ky/QkpDHjZUAR
j4gYbUGFW+P6PZHrETnh5PyXsIjyENEu2b34mztWFqC4NHZrl1e7HbopAreNLHo2
9zbLtXkL9WJ6kvJAEzPQT8bQ/YLCDkSOF4/hsVS45XFmeR4B00VjZXex58Wadbun
ev2LgwCOFHHEbi2mOJQw6GatImPpeTcAgoX1D4qnvpYvgP/nzIC8wLzGG8mNq5/T
B8qrTzE++Lw4WupbxrV0LkI4WIG6NgLSBX7ce+AiwDdo6ABoy7IuQY+BXCZeidGU
xEWTQhQtIWN3apbBe15FtOPgXuSzloIkRWOyXS6aeOj0WcEPKqBC+bRuXK5Cwo85
wRh9robFORWXYkzzRFtRm6MXkY6gCYBypG7ilKMevsMuFUXWmKwm4m+LNPnpPeDH
HLaEyo8pbicbgDL8M6+68Enf+Q0Rx6/i47jmUMPs1ymqpYVfu2ngr6Kc94eJtM7D
VcXmBS2gRnz5YeIFEz3cnaf/jyrxB7eAu90lVHta3AJ/5wHLuUZ2lx0OF2b8TmRA
52P71DkyCq3OfqfbhKUW+8EK3ioX8dFcTSfwScY4Ghy0xjzdQzH+qwNW7y6IYYwp
7oMOeC1tprLp1SxEXwz6rAvykuCUEWLtvUZOQK3GOq0jZ9j+diluz1yWGJb6pHhX
/lqaFxRCc2Tcq+Y6wxMFtnCPjQgVJszIERJ254/Qs0NbR+PTb659Q5eV3GtJ1X/4
s1hYSrqOT+8VdVSnjgeP7T6932FL9a8DYsqh8Au/hVxqjgPNIzN9u1ESb68rrj5N
vgw5uhasXhLQ2Z1M5a+cc5iPpcHFLcnIy0KlrzTmdxD/tV+PpSAZSHgtwj3vqBru
FYbXjuRfLHT0oUOA0CB1h9YvWFxz2g+vX17i5LouD6gY2xQwM9EBDqELm4SQf4fF
ZfDKJ++f4ypfEbaPPOJ3kaVcr0HbcL9NwOUOUNj80wOxe24e+DRbmGTOjAwYzqQ6
JbGWGqt7Wyml/lobAwWWx5iesbAPlXQOBzOnl5Fv3v5l2sVZycvIoHdFVOw9pcsY
WayfTKIX9S1DyPYB3hjNQPGpk8SrINx54T1fQW/jrxvR1pRQejvUWwQ88uhAcknq
Nsy7ICJwKhkfO30cHupNE3pL/xvpWhbtB/FmjrLgfJJ7mUr+8Ngh05bG+9sGfnrn
m/FBR2147YmJuuvxhK9oaSwXaZUJlrzD1oJg+Ge4itsphTKRz5RpT8g5lWJkZH4g
Qn3fkpsxhLbardcIFIheSDr8yPnC8tb/Z0HGeYyLzNfE0qWBR78hf1Dhtw/5jFu8
ThO2NpgzDibITSUmGN3HA0HqC1CtM0gi/sJvMgGATCVPdGN5KoX8qsqMPwsxeNWn
yeb2aM/6vfoqRlzt2k5AOrj+ezKtO2VzIvhdjcwpAFPiMAwcbbwFArGTv7t2kvgn
FIROQgCrDGIYsF69NhLUng46wZyhDSQw8mMupZaXrbqsaZMOnxiroasES3MU15uC
A5uNPoKJNrUJuFCV9uQKOaKxH8k7Wjj29iuF2MJsunzgfqzV9FlOS557aptIwqwP
ZY6bq8C4FjsIxpBi0TrWv8z7JjbXzEl1PqJIDuzkZVZTbCiCQbJYwIXaWZqDRed2
2SkTsQ8/xgusdTPQxk/fjSUxiOCZqW4D8ZzPTO76HaFM4XqK0LAFS85NABG4tpPp
eTdDlWc9rNB2XHkpMvUQH1pXFqLmKVSUp7uHcAgQRcxomsya8Fs5JxS+nvjQHjxC
3hqd6MYcrdOPuunVD/UKsRQRvJcr2+0siqo5giGPX4Zi4jqnN4iPRciBTCY4Anaw
JcaHr1lZP39aZcMDSE1r9vM3Ewfc2EMTigi9vKrD1MbbMhCVPy1n6x6Sh/iPqU28
rhNfLgM+A+8bXO5UrEQ1LUxJcSViI+MFl6y37X42AdAiqs/uvL80XttlbcXPRj+i
nToZnfU0sUYAOTdpxsynwffcbZ1o8Cgdxf3HPOma8YPMc0SnsQPKIDY6c754urKt
YtgUsl2GWNxAMj7RMlX2U1tkBFkaodlyikTMLySQvi1yZ2pM8z42TSHf6qfau/Pt
FiN0jOraKdoUVZ30gFPk1CT4FW0mMrVe0da71IYJrCifYhsqPGafSVtRtOoMCioJ
OTLxm3HffSwjKuYPJArAFePxbCRYkiX4wL4drxb72k86tA3cyKfHMa0iU8NYTjiw
LoHifoiNjIQAxInyV2n9qyztld/MCTjVUFMXAURqWK/2mrsng2LfoJIKag8sV9Gk
j99C5W7rfkxUWCwyHIKqwsvQbRoqyiO7oKWFhPQS7LkyKsCu47Y1gT08hxQMb5rQ
ETHUc2U3DRSRJ75x+s63lJyNq5Q9CjSGJ4FdgL3JlF8YsQ4BfKIHK96tqmJz0VoH
LC9Nd2TzDbLYYF0U/WLbiPRhdHQAw4/c2B2uj6LicKxV/duYmGaQfMDckA31afpg
HAnRaYYjnZrv1EJoPFIJ6o8jlua2qGuBpe4LWpFHgdi4aaR1p5Ya+ZMU0boEaJ2g
P01LBtjpv7hvKW07/0JY22lgd1eeDoG9N0tzWss7rmTDltpppURbCpL3HIRurT6A
nS7NN31mPdFssJwGiQvFq3ELKhJPWPf+wscC4grKAOq1QQXL5/PuJAHjzOCbjCvv
Aq0/q4nIDGjFlkMYbt238IHAMbOd8saIw6eNxTYSxsovPARjVZIIjCaBiNHqBBHx
qQbPZVN54VK38F1OONtY8QTjxZia949nOOeYg+B0PhaC33ZmZVKJAeXUA4S2fiR5
+p/5WiuywZ1SHck0gbzVOf9yja+NMTUwZBThfRPSH2z6XweYS6tk33l4c9VzhddQ
k+UFUhqM7zuOXGJVjwP9pNZlpNKawtPh5Mi90kdbMVPU/y3wPSryZK5rAk+kJuB0
KO0liceiTYGszkAj8sXQCtKmtbxKVpR9+k68DfhUB+l4wL7ZKTtcDHE+sc/4kOX8
1VV0dkuZ+wejV6SC3npxoz0dfg5MVH5s7k+Qun9k0vldmhiRHQygHmzObBz8Ghw8
RHGc525OBeln5Q14vVVwk5qa7jVIGjiowTrwySRCs4rdoSbob7HRhMvm7ZK0N/lD
CZKzT6Xe9twDBNLB3Uwmp3EVVjMyUvNmqJvcOLrS5L3eOV2Gs7srVDX3ip3vId4e
yvALhGwlj6ph/GcqE7zXgRwGZ7k5vFhr3jXvJ555nRAZzHp9iQFieIBTCfqNBcRC
8Ax6orQVGDxXbMER8T0ur5kfu53AdKpeZQ/MqbJgILFeAzNPqwu1eKnELcN1eC/E
oXQoN90Cf/z711H2/7I0vn4K4optV3yxus41tFDDerFfLw6PruRj/4CjTN9JpLcC
eLOIu0beLAV7dCW9LR1yISSCKwd2th14WkhjkhlJISmfn770hKeQYR6myyxq6lDG
YX2Q1hxGUh7R2CqvaSOyoHjqLv2Wst9/wxeTWDc88JUW1cdB3p3FVl0p7RfXgy8r
C2x6Fofb2NMm3hAPJMVsF8d5oMFvwI3JTQ9Mpa/bXhiQnZ40J9/QwZk92bofPlVj
noIMtbK6u9wXsQecUSi62zB+Tm4etdbpwofTxAh/non/HbAiS9cIYoEcLmjnondy
V60W3Mc1749a7b8pHC0qD38FpyR11nzF21ic2e0p5+CN96otWWyh+IeD0Ih81aZg
OdrMmgi51cVrdyK5vco9eGIgwRKRbaW45jd0HgAXQV96TbtZnUvV5xY/oEWNroFS
bL3zLHK9EMLRtScfx+Dzo3d67tnejM0OVRoMNvf+7gcQeL+Uh3KeOx/yX2CJftyR
qtwOIJjawH9pcC4cYuP0DzM+OiPAknsoL+ojCzvG6cwVQVFZ8S7pLCGse8cMeXuk
WX5JR6Ly5xLa2ucp/CBKouvGc0i27/q5Cw9knXpluSkFqJ9UNfGpNnLducvFjwYN
43vFQmYbV8Bo5R3fS60LsGmWBPii/V1iDyXECxQZeJK19f6q3x2FNBkf3dSPw5pa
PQQNRKzJDVoL61AR+MishcxRXAzw5QDmE7RIVjNjuzJ8ca8qvypr2GPfDB1G6QeD
FoAliv++7r81MI7UzgxVg7hdRkDD63hYGl9zL8kW01iTbXRNVxgHnwbt9iE4OOhK
55NJS8g0ML+pBu1evP248DBm8GqzAxltqykkdjocD5V+srL0cU+2Qtr81Mc66ppm
MJS/rYUCoY7ddlIa4LuAFxVthCO6a5aGw2FXVo3mo9rkEP/9kheENPdIy0O9L//r
3xqCG0FAtuuE8X34E5/j7wSR3V5rcUtNJcL/7nV2oZ8lFjc3VV0CD3CAaQsjy7yT
qPSq2WAVH2PMxGho0kXh6NqlChsRp25pkXdvawyaK+cvaSOvQvJA8a9OSMb8nDSf
Y0XTYfJah9Ptwthvyq3amucUzMSKuiDGfxODLCSxombKgo7JPkoCcE4aeYmceTKa
ReNu29OgA/h3R9LDIK1PPvNILdRB+2pcb5K/pfQxAOjbZArG67mOkjmE+jtgXH6b
Dhq1ak0dIVizNJW8lIUXNOWfnZYxuDCAla04ZiNrK7s1F8adv0vF9MVX2U7Kyr8m
JpKLLwf2A6RWQZOOyRMGLmlZUvBXeo7e/YMjQnFpUW1spQ12Kn3J4Y6jjVqicvqV
eD6Mi0VaL7QSl/+sfxAsHWkvzK7z4bk6L7tdncKDgEra/zS6ggM5pEuMJlOrFpJ2
uN1BWS+5iT/hp8Gsoz0ZyLWxq1OKlOuLVfnave9iTlakgB8nUknPW9wdPkRwf6A6
zKCa4OLWjsboBJ0lWrUnjXhHyHIo+DQvNGWX/Z6Mpfu7LARaLBVI2rrPgGJ3cSmR
nXKsdUklM00KFaqdaRo9KT6J7uDDiWEKveHIW9cTr7vF6+hwivZzwrIQnP9zGto0
3YoooQ6PLaqsDW9Ydk6Itmd3Z7tiwVyW4/5Fjx0oFevRVfAxM5nxlAoLSfB24103
pqDteQQwykCyOYRlOyl9eMblRe1IUevN7mudDCO57OP+05D1pLccT8hQYQwDRBsM
2fBw0SjDhE2ylI1hl55OyHLF4pYRLeyCUH8WsqnX6pFSQZNAJXYs5X3swtnFdV7g
o+ZtI+vMXVtu4Ndx+euwr3Ua3S8CZccsY6UDZ0NROnpw5/XCCpR9GLat7iemB2ig
ELNqPm45xo/3aQ+0VXBwqNOu0CvcV4DoiL09U7dSUHUxz1YbaswOvrx2gmfRHBHA
o2P+ujHfn1cbXqJmiNQDJRyVzo1aRh4qjOw8y3c6gTtHZ8MPhHuKFwx22LKr/uf9
65nhp3oAwyoKXObZttpHGOT/iqmFP7hFWuutU5BgvM2AQ4zoW+VmiUie8Dh4nvFV
h9mqVsVOFX/1aBIMV+XKyphQQWzOJ+o0UAdNPDqEtZ1f57M3qin2WAbkCojjj2uV
ZZMB3c/dHpmB3KOY/L6anZxtwSmST+khOepUtyt+NGrGV0W6CovkIc0ecOtCug44
8Wi+0GGDidm1ujqvDVqX9XQZHlQ+FqmWCNSbqrlVZxNgBLb0N2ZhR99BZrN/HKq4
3qaRO6ACLNu/9YVyWVxRXk0CrppyzmdLvGW1woU2sno5Adym5Hc9jpIylEAyGSpS
6/SsjD84HlcDVK2KAWuMRphAi1GAB8E+36HLDv4H70sG+Ra8yI/2Uh4xOx9HmgcZ
gA84A6Hu+37qnnG6KgkPUaIlv1iTlzDLDxRAHfY0yLxyGc7PEOdxfyInsDp8OwxU
rLoZv2W2KTgkFqBFNBUZn5kI4+cWnmc/cerYVAUE9g3udYM8Ks7jKjyzk0PChNur
isFE7vBXmhtXyos7sScr+/V+mz1iV7pPdD1keC5CBk3n+alBBWvO+V5xWSbRX/vb
ws/fUAQceU3cJQSo9G9rGC3clJCZGDjh7wjHa00PMRiwfKJrIEAZyOW4ynyzwRW3
aZ8ERBGOusLEKvIhtcc8DfGbiKaH14QW9+QUvidwRa0DTOABZsRK7oktrLoYVIa9
GIjDrS78zV01gIryHUShwlLitMXPVRLCyCqerEKgRGtV+HruzPuNws/WfOkLaa7O
ySrbE/875moGr1zGhmC0zaoiZveqIoA6zVhguRfXW/y97x8jQwdL2MydLIivKNHs
Zx2IGpHKL/mmRPOnyvWhMIv6fQIbHirwSKmLyAndysmYav7GVkHhh+MlyQKaLltZ
xzph8o+eDhOio+CFqpOqWClD4YGM2+uYW/DV7cP16KJ08ueLWPw9i8jjIdpQl3UD
uNdsl33EJ3R5Yl7/qzM11c/Q0d6sPNsmQLc3mtVCUCSGFpqybNy9vF/vbsS8vbAO
LoCofNnKezzc0f0jx09J0R+emkCmp9DP/ec1kCKPG9pHaoOybw8MrQHL/fxXAedQ
ZgaSmXr7nSkPBkOUeG1mdSZIE4izzcMpHHIBq62jHUAKusYqhmDUvb8cUYSB/cwL
s5CzFkRS1MgNFwYoX/YNuJbRVe8S5siJHFqnzgkmI+hrd5Krg2rCAc6+GLG4TqH/
qxQwFN8U18zSoiwgs0WM4o9tSP6s3PeHen+ymCHkLI/4QmYNtdKj3eGvnUOhpCjh
hY0DunNCOB1GPfH3M7+dtiSEMWU79d7ZEhcceJh1cU+yQtBbzDL9Nra63/KIcy/2
eQW1OhdD56KFzY1cjLdY76htqCcTm8xKqfeTvP4Vhtibk6fo5PiIZVcpiqbVoNxt
duI1IXpR/VdFv4kDjMasfVIeHPda9OKYnHLgdYVqdn3SPhYk+59Dz5iFjC1qdbfK
V7Wlyw+ADgA6rC8XpjaPfIkYymWxiQpmkimdeKLG72fA0wZJQP0WrsynkwUjONcz
WL2Cyctk8OJwOpXpKx4yLnq4zWfboUqltNGBAIyvpt1GjPsEGw3wqFb53FPmQI7E
M2YeNnqcTZaFiWgMxbNEEEPoe1u+7jtEodXxHjHAVElyOZN1eCDPA7uHOW5A+vMA
zqUuhmZQWxXBG7tPdJqvC2s94U88jXxkZPyGOryGSWibgSlC7o51WNFUaD4QwNSN
y1zcxm35tWVQFjUHhY2DKSPUPqe6T22MPXc0rPN1DvJCpOHFmgbQWIneFYvZ6SON
I9/jLxyvhJjPPnmf3+8k0ZY109ps6JuR36+IS78TlSx0pjC38bjP1BhAA/7e+WSB
XxPtFRHXGUaU++Lqy9NLd902IS6IYW1Rd55Wjug5ZVbx6392WjfbaNVSQ9+EZhR7
h2OqCwCoX8TM7m+7kQatbqQVgDUqFPzja7ir8Puaq9xL0w6mjaJPytJGGyADuoyK
KT8P0EZe91jaMkSufrmB92lGMxD6RgaTFwVsen3Ph+fCiO/btG2CGI59i2VZ57t1
kUR6LlYIQgLox7k+hd7k7UsI+Jp3Zzoe7tbN+DAEkw+nZITz1wp1P4g1KoTHAUwP
FC63/VT4n9RS1ufg4FlAvX/5Ol/jLxCqkvZivxr7olD7vO/ZNZ/CO2v0ne28pfM0
ciQglrfzfSQOPqswkBZbsPYvgNrBltTuNZWleaxfPRxSxw5N+pJhWp1zDtCxDvuR
G8FvEEKqJGNDMEQSZt7rWRb117UISFUAxc/j3FE7jt14LulmEhurwCweE6uZJ0wp
5BLRe4Z1QdDERaL3998pZnsspb9Ncqhkqb+W4N/39dsdDYjB7uYjBWys3Kdpow+G
O+NiinOecGDVEcOYI/iDvb/cCwTFbAbvfibkYYY6SKP+KQgViLKB8WBrbSvDgDIE
lHjqwXPJVFO/1laDCryoaA0BYzr56yP/fzSjmplFXVy7EzSMV/RwDMlXwKWuAJVk
UoTf1ajb8zZgQaT5xEtQ8UsX2jRTA9wWmdJEdZysUw/QcQDFKWANt5OrVAAkjpZr
foqOevYLczgcn5ZK1Xz8pgaYJx3RfeZk8eiewk7fXEWB9b/3JPvr6ZpoXivQR7l0
VR1TqGogOg+6uCaqd1MxYJDreI1W3bSWZiKl0iCs2YxXUc5tAT12sABRg+2tGFfV
3wFx1+0ZORps7ierrGNRyYAdyfu1+69SVfGG8UMWxUtTHxyaGH955hnphFY3BHSZ
qN+15ZhxWqcAVQcjqqkzUYmZuCIH+GRvud5sbo1E+bz5mp7iJiNCy0D89ONGFtkk
0DTN3rYjabwmeH6cP/zf1K1lVoIc14G3na+P7yUDROgvI5OARBYG+HAXq3Of20qV
vVxLhIAGO9Pp6yaUNPd3mjZMMpYPMrwpWv/9Xeq/B3PO5a3nGU/TR7SXMgbvr/cE
fBkES5/5OajbvqOAUbb3LDcKZaFcrFQ+jMVt/E7D27/r3stpWmKXQQiXRx5JVnYv
1R752jxt8bkhGj3W8y01uyi1PWvTdIrczo1F2UBB+mJiadLVg7cHaNbOWMIxfweb
DVyDcHmHwR5H6k6MhQM5kKze2SuWl6KWjGif0Hn299p2fA6Ke3whWKEV0I+55eaE
wP0vRQwkLs82nMDWwfIUvuMvlItI1/FTJkEdJMySkAtNUAA1LJxI28AYBTlAkzBb
IZhEuOBRTIs9l5uKx05OsYjgVas+y+1zZQXDTBb9SGaDeSKRpLIiW71r4PxqT6aU
a3KMRf8+lLYMc+w6dpJ9Qngj+2Ii+RXHdZgxEHfNipCriPNcGQOE1rsgMNPUeypX
A3HSvNcuToyspvIGFNcPQpxSP1qx6rMIRsgM1eQkDNdCJeTpT8TZ+6LOnBYVtoXZ
IyRSz9Xtb0Kb5aXwDzZliqCWgJE6K9naiK+z+ZYp1HzWnyb1GpcRNHAICvC7uFGG
KImlFrjYmdcPB3ZRqo75gUFZxSBLp5wS9yjKlbejvoa2CXoe/mjAO5kTL7FWS2kS
Kz+Hq6omz93+S5L+pqEZjJ4WL4umABTptu9z81M+kCrXxheaiDbvufOa3vHJ/OwF
np40wXTYl+eR7QR9QyYKw4p0WNg/Hq69P9BUDx6wYWFqNMYWI9OzXtIakYUKdxWh
LX94zu7glS7QYW/R75j9/cz4Ujx+kTFdefWwOTuccdjXcUJlEFEoQR5k5orUfo+A
lSXQdCiF3BgtsriwgSBTDlOfNtjNsqRO5+hrVmPXRhrwV4pnOjgr0KuIa0lAG85d
ZRzdU015S3W/qBbbX1zphvubmesUK81Pjk2y6db42cRSc6OKbb5Fr0BQwPEez6ub
KeZk6+m/Me9TTxb/f7gHADB4Wx4JR5iySlhS1XybtOdrFNGhKL1p8p9JWolK7Lm1
s4LOxwS0Cvy2wpa6UtLe44PaFzrfVLxB15fEBgueu2+glxNvpaOOJw2juNco+t28
xmltU0ovageFAXt+KdadBpdVqEGl9R2qwM/DM/sQ+9ZmroarCHfczWuxp/8kvXJ3
EWIIBOOTD57M0cg9NDgdF3Yu3Dfr3Loyy6pAV7jLDqRpfPCo4+iGMjVIsV0ziBqL
0LS9LaGMCd9j1tF+0Ar/4Mz/xWBWkGmKOWR4teEpaG3ayqGdNH+w349Ze4C2XIUR
VXECoJFcipwvJuwRx9UFTBuLachlTDpucS+j0tqk3/FDZP8lYUE6xyhas535aA7/
kaz+xngshoVzq3LkIuu+S/ZP2iyj+O/hCnGdHK4tlegkSuERHM7owmgKRVwl/VfP
s3dyLgWD9PVtpbxu5W9qRXfvbAHzq3R4Qn+OdvZFfHIFMIWavysStw27M13detOC
kdOUJxWq1a7pj+Ah/oslJvnobfQtno61t2xClucHufY9jLiO3qTsG2Zg7RpaoI3V
cte+tyGReQWJh0lHERaVMBeL5Q9mo8RzYVqF+Hkvujx5FKcIlP5uFIGPhLvlC0MU
+VaykdyjGgmSqZWkufoIVTlm8Rc5X2miGhvK7qh+767luyEEM2bz0cA/rkfCfMCk
PfFgfTC4OZu+5F5mEwZUAPDixxg2z7Gxx66kCetGLfDgn6BmxP1ef3FiQG99a+sH
6yMNxcdMrfAto50STfa7idJNyaPgAwEaWq0ufm494D9AE2pWWHKvunmxBPKKTiW9
qZwY7sPQh3mAtIMGnqHH/HMOHpG+tGzwmjWaTbKbIIbjAA9TBnjhmOOk0XyZJK3i
e5wvqX9BalnGM1WCFnZa/RvZAE+8IGrUM1FyGKtqJnBERGq5EhH5TlXATzJFmSY+
8RdAyPwHf7FM+sqjDrEQacnyLXCfy4J8f/Jdl8DBoFaKmd+gUtMPx/NkLnWbsYSR
RjXgqvPTS2yGlE0gX7TwJ2MNT9/HbjpiCYBhnQw5d1FguVnnLcKrNHOfOt+uLqfc
xhYjM24cG7mdRgrjxON+kImfBnD5CF7AyueqCW8Vpddy7/5Oreva7WOq2O1mS9bw
3Q5EOTsn2c2vz2/jO3iMERVaWnxxKnJJSb/mELrZ5Dn5Vk2FTzjFXBnWARWuzamn
a4jcrkLDXSIfxMFAIQ4Nb439MJxLQONOYOTe0wJK0QZD2ut2ib2JYAXGoalOhHPs
rkq9sTvZgRNbtdnGfy4OthLYGeDkWScABXJB74ipLISvtJH0aNpejapV/3tC2nVr
+iVbLGc6nYb50lzugBBxgaQwVffuEuBHp5RIRVRFKc0R3OLrfc7mGxm1xnXFq4d2
AP3p7ZNbl0WkM9uDY3DneaEjTT2P27LIprB35Mk7AKBQL7lLfti4r/2mzwIRhFij
uv9zVGyOZMDPvOYCLqm6nCOOYTXUrhDDoQjuDbDrA6HsmDRQmKGH3rErb0eu7zng
M3b+QHyFP/VCnGO9r9/q9zFg/ZeCoXs82sJJeN5ixuAyu1e+4xLEtrOAhBGUvwfp
h1z58fbHjGgOTzga3ZmtikfgWcp81M+Xku192WCLbSwjICkD0Zg2+fpp+DscaeN5
DRSHJUf1yjg4aiiPA7hnevU7Dc3mSGTKFuBKAGaDVj57nnUgWqcARY7NilwXsDrz
6xXxFj1oj7FgfYIcw95H3KwSCfNsSIk6xLtA0kfYYXBY3wPHs35osF0VsL1Zhqg6
y4QaTEUjo0yFkJ/s5etFPKcd8/pxop2ZK2jRgbQ2ihrHtR2ZBvLNkCcITU3AWlpY
WViZB54R2U2DZcQ0oV/2QBTOmLsA2B06jHZ+LISVKEWsYYeFnwgtlJmGNKRXGWqt
C1+TogZYPvZuaNEBWqu/ISz4Ez8su7mxl6IhRIgkcOE5y1F5eTsFSUVDHs3zDZGL
6sbCAit3WqMP8ysjJ9YE5poISehtWduk2x7olCrF1ywWDwpPNt3aTkPFpSP1Zojq
LgZfo2naTs1/hrYS3yWhM5Fu5YsEmyyMyUDzvy73hcO2UXqhGjtU3Dlm9TTb7/2+
xwlEz/cPArrstAA0/fnBfkszImdZLhNsNyLGG6hjSv6nS/6P8jwbZy9LbgZ3SJ14
/DjrbnEXT94ZGRAI3mZBIJebSyoEvfSako6M62oTw6k5i0Wh/eTLPIWZlxcFzra7
qxjln7xIhHfRt/cUOb2z5qsn9IkpCobBRWr9EkW/YWcDnniB4jQ66h0u4uKeWTWE
GEvgsnBeyxssn43l6OoLQrI48Ez+VrZfrIjmBahvzbUKUMDFaMzP9s/VRQoOgqKv
6ByV52XucY4gYjsY0hmpoOqcQ+l1wyqG+dWW4gmvZPNvmutVCgnYgMoRXEiG3txP
FnmGAYsbV9dAFlinu0i8K2zG9knKlOZGrZRmQJ1pN8qghm73nb9LAObOnJtD5SBi
blp9xghhn1uNmOcMLCtfPFFNC03VYhvMIDwpDCIVeAeeTgB+jWaC52vusBfFh8M0
zeyAq3UX7f3evDYahffphI9z5mXaqdfhowj6AIJ94VOkryY6bnfWJaP4k0jHp90+
lypFY7r9nem008f1FZrtsLY/wMiljFq5LZUGkHpbiIP/YsEI92I5CuwNmnyS10iB
x02GvMr5NLePSXfPh/MZoiyyjDUh5DZOagXwnDha9EihZX+REK/c+1S0AY3kqgFl
KxiCja3wxeocG3ihaCs8f8TUdiFWHuOGjiEv7IbMf4eFSpCnIeVUsqaY5pASztzT
pc41RT7sBvM1eYNk44X+A9uHO+HVwjqdvjQ45a7Z1tR6aLdPOpd1Ed+LoiDXfFKM
whQjue5qhAP/QQVHFvU+DOPE8tM/bGh7SKKxyMixM9iFEWFzNx9ROx7eE9PRaEuJ
kOmMMtXQdgjBf+CokR+ZaA16D8MnJBwKFcZvIHw90waidKlqOo50t9nQ6AhHSew8
bEia2p/lnBmnGgWrWEhsik3oz3ETt35Ahm8J+KF5gReASB6X7Yy3Mc20Lu1mzN+z
A0X9lz5uM72uidgSiMzf2ZVTzpkNtd25ZCO7zzdMOAgcHPDbD7L4U6nPaeTlDcdh
Qe8ZVhzN1yO6wAEhZig9z7mF0fVvoDRG+rARb0Xzi2p9s19++zrGFu9BGBUVGA8q
nUHOEd2hxo2aj/8tGdW/lZFG8i/qBn+bSwAY4AhEjssUZLOmxqV3fXgGSk8SDDI0
OX1SeDc/OWRuUhySlAfIA9AKC2hVutLtJ/N9q9P1oFh/87d8bzLFK2NNoyiE0md6
+3bYpDdm3+OZBOfjzaI29APBmnam+A+7imc0dknqWpYOJesR4beJ9e/1FPcItOK3
U8vobITHxlvXWRpfacIZ99rnVpswomh+filoAmaSetLDgiFvGQWrxSjPRjQ91QXc
aKb25d0OhVNZLfdfzBRlkih33TbJ6+wxbGnzygqOxMhGtbLW4oiWyR2AWuw6wfUO
7emlX6fdyLANHGvLkWvESk0YrCNDOVEGTxyG0XZ7349VbDbbJuQpfKLBYZ67C4xB
fbGHQ3mpAKuaUNwjslEP54iDRMA/Mu+Os9kn7jdihm8cVxeSDJuxw43SD1AezuZc
qpTVzcWvAuTFI4fhR+b/cR5rvsRW5quBpHqT7OLKh8CwY9mDHRLMIn0jspv2S7le
Drs3rnG3u7JSz1R5rkg/K/+hAQhdMpFcVI/ft2Ij85fVGbGlKW9ac+hOInuZR+w6
YWlyLdytAOlY8s3fOOlgBLVVGvbqdYHCfh1tcEAvoLkHd407t+xRXstxhJfYCYT2
rZfntSvD4Cp0u/q2i0eTjCeqyh11iESxSMY/PaEtlLGPJvBW1AxYsFykWVJ4dcY1
wPjdWC3g+WWgQcGbXI94qHwaIMOLWIQQubBOe8V3X20hDkJWTZ4CxCFFFQj1JSwa
oCezaf4vWDk5ZTDUSdF83Z1l5SmqL1/YATBeK5QbhDICV8Fpe9flRBNs34PAOVGi
/FUjhvysZd0vskbaVCm4JVpzumEK/D5ct+kdAhhIG7CpLZpwe5v288JNPgMRZHog
C05oPxteHOCM10Rv7kkOvQv5iLWKlGaNukVtALLae1ph+KQIh5/RN6QxAClAgdbk
/c7gJ4uUUvbRFar5xDA34vSm3Bk1KgqTDQL9Kj7vUKSVbBNIsp95r41JYtb4YpGg
nIuhB0VDIP+D0NlRmQlIU8ZjZY0E9ksnfQjpf8nA3GCVCMd5stUaAtS7E7HCCAxL
XKDOx/8pjKC5UVFVyEO7/CeERPK+TAv25h6qf0lx8F+oQtYH86etI//2/VAJht5u
gA1S7brVtyjV96CJZSDSujLppD/uLv54/SmBvB8+TIDNW0VAGruyfTYQrMTSMz0v
qt1TSDhYFXj6l6xGsFavGWJiRKlvK58xaWXsyEf+I+DHayxoiS+meo1ZqFqiNfln
yUT+By1oy9M/rXTOfd6rVyqIayP7ebonn1gMGvsUccSGbReiiazy+2hpiE3Q8Zy4
dQjrmhe8fJTcjj3YBwjCRCgAP4iT08IXjv2lQ/zHqHGriUDmEdkqhamsMDT8tL8e
RR3UF6/wE1pZrYs2/nLPqkfpI9zw/ZusaNE/w/vTH1c6peAqvaDXOSCWNPt2+fAp
JCSn4EFqJDHgsXI/gfGCn3tiXLsb8zUoIRnOndwODs3zNYx+j+0eJxBxEaJsz8Ab
fFi/DgyAbPUxB68WpfBuqg2RRy1KW1pGSObj660uWJSNc80kYzrQAINhqk94RMzJ
wXVPNAvzVrDmIzRn4dEl6LAzOvVqT0ObFY8AhCl2eklLgvwsigqC7qqU0DVf2dDv
y3qo2fzupxZEpO+sZDq+C5RzEpEc4uy+PdvrWg8AjyFX13mm5xjzH3FjhrHptT4T
lyBBCeJGkD6JYwQjnhDD46td3vkublGDtMtZ/EsGsnozMP2fGR8iD2U+apd79Cab
ob4nTMEwBZRGYFJVVPKmDjTC1bwpxG7NB64UX94kJhc+NQ8cH1FPCDByotx659R4
lqURq0pU6hY1aIz2c3XsAQrKqLuF1cnRHI65wm8iji1/b8tooPTc4hoeRAExtFDC
nqLCBIrZguBWDkJ2NajsAORl3rRcTUouLZefr4TbPBApbsAAYcxHndud336GCG64
OwBoTYPqZTciWgbQArunwZtUavokHUfKQGUwcgDHHQaCqFLZq+kZetMLsHEjtasa
Wd14pzUrvJYFlzHG1liuo7CKMC3IQb0hoD1HvQHBmCc+GzY+Mc3Fwfn8xGokAoG9
LxI6IILIQvBDzYFnAeAEOj48OogCwXbF5T7LTjmXhgBY7JQfcZmZC2p2KUHBsms7
WO7AmMjURh6VfyYMMIbSkp+EI6W3N1O+gd+R0K6f0C9lbpxNnUHsUA9CxYHXZL01
lXrIh3e5h7Ub244aExVVGJZQHyEY5llRKLCYjQ4ERNNfUnCyx7WvkN7mxeTX5lRE
Zrn/ifI3FQFOQc7CYSJ1U4zy+BRTceoea8vjBuxAOI06VKBlvJyBSQqBbkuTdyLZ
RHRmo3wE/5f0HuOpKFEx4ULkkq/Hi/c27x7W4GWnU7ko5uwy5yyG255312K/BZFe
s/PjvcyVEvW5OX7CuQ3uhkAekO8pkGnyuP1hPWJWIkJ5pAlvtRt0uKkeMkKIX1CK
C/6yjSXEahGW0ChF4w73hq/jgW9aBg/0/k9nzcWZwa66wLAIvW5mImD98zhYflxz
nEg7nMA12yNMfEqS7ZLDeTj/44tmbHf5ncVM+wC7J3HUxmMn/VRmL2ArPxDUkqcK
n2/3lp4tiKxoxitIo/B+kD9Gr3hrx/jpfkQYXIYcKY3VyJTR+eYUXs3Uol7ISLQE
nMTqaekT8NH6KIm2cLz54bcNp15WNyAoJ2y0aN2JeQO90959hXCsy/Mzx6Od/6Zz
bGDPlYTjkMmumaXwoMGMsxxt5VKC6aF1v+cCK/TjaZyJSweoaYRmiiX1uAWiHnAL
HLz5Eo+MXtzLP6adQNPeAMp8vCfJGHyWJHjdr+nmg07rrvhrmE8T8tpQ0hA2XwPX
gk43EdMVeZUfYE6XgwWBDftYjWHog4YjeDQ8+rEK916XPS9PNTu9MXVUhKArXumA
QKAhUNrt7BLqRGm95IvnJ+smtf0wcoDfVpzxzshbp0hENqpknPNk8Qo5WkkRRN8p
9DmSM2qMyL378EU1V0RQT8ok+ngPZtp1pBIxW9PRIF3eilVKQsOWwNH1T2EiQGgh
KpAcJmb3Epc5kXgxTLpJt8GJabg4BlI+XYrPpmONghKXn6SP4BZYL+iQBaFWhfy8
BG5WvooVgwqn7FEhklYDH+odz36j6oS7LQrXa8SJXsni25SLsR0/0uYnACYFU9Lk
scp8IV4TUeQItbZq0qrLa+oT2OPrrSZYj85pJYTh0Z2b9s+vCSFLnaerYV/4yiZr
QJYjt+N0WLSiCQm+WuiqoND7WgStIWBrCIpyhM5rFOLyBUW46beMwDK1WYYRM2xl
J9d+KqfCObPExrgDYl/BvkFaEoRmKpp7i1QafHfgYVRus0VtUxrjiJCTijyfpgJc
e7D7T7uoj4U4FDaqoiBWAv1NPxr1NQoQANl5TNvOhJ769cwrc4SmIegcBExbuT1O
il6kHZ2EyG7R0VAlu10IoOD2XjgLAvdWlPKk7hWLn/7Xr6zjeR1YdreTnAIDdbuK
DUISqmcpociWv2I+ATEUik5sdr1Mg95vfBEE2qzMNYnun3ZFjA/y3d8RL19FOVi/
LjQPEpPaDsP/fewTPvW3Y1iURB7l2w6GcI+vPBbhNqKwGkR6ChJfMFkMSbi0s1f/
gwFjCZW/WqnQ2ZXGSIpEiGCQH5TqwoXfkxkzAZb6J6gqBFNdc0K7WOIWpSnt+5pI
PaL5vO78voCVjTgRLvRT8Mgmbg+LEVg8zgIG9P8fgNArVay+dmsd5Gn38hrec7my
UOkx5GDBBc1o3DYcnpp8fhGPpuBm9xHAlDsbSseAd/fKPQq8ldNHxuxW0qtFWn32
qQq6XVzcgdF5dvcbYAo8H+/lahYHCe9JfXfj9m2VNAf2oQT6HDpuvpanDXhTPrsL
rci04XFc8hJ0nSe5tQzxycQllL3UvZAR/rF6uj6hocyZGI/jf1FqQvpBUo7maF6O
YwEWkiZqCcvP0liaQkJ1wZQMCid6GSn9TMeJwCOsk61kCXG78ENah9Shoj2vSD7F
j3TRGO6y+9iftgapRVtWQuHPngXcEljUSLcpxHYnZdKADKI4Ol6OLVI7cL2QF0Ki
+I+i9gKJkiAKOEtPTV8ZjFrXeqXf7gqZ+nmS6vvI9FpOdBgy5sYuKKTCr2D5VoMk
avKdsTqCJ0j/CvmqsoGM9MTtbgMZHhNzZzht+lGeHbwYkQJvVKLDuItrOgR7wJsz
A7dslX7JqOn1qR80qVz49qp6AUQk9d5JYbI580q3vCcZIvwo0/Mu7XKWaAtg5cJ4
QbxnpV3CQDKjzXJGYmmE3K2H8YwB63UHY8CfMiTSKEAPPO1czkZGSNRDcBylwLec
r1RKaoxey9AydxM2+xsIE5CKHOlN8QLOVUXFqHJyDGM4+O4BJcqZ6CinKhEHFw7w
6RWYNRPvO9DaUQlaNAG8U9qAEKfvaBsBCGwZpQr47a2c9XpAmrzK24wMZAJe+WOt
+k0fKv6hJw2aFsawUvP67w7De5OoGQfYVt/xy1EmU6Yg3ne65BPAzHvcacGHJHUE
BMSRMmjAb+NKlL+6v9FN3RVQiqzd9rQ/iOAkfY4odOBX6dKg3b59/HJzL1AdTObb
Wd0KMtGIG4VW6lF22cU0qUslWytHEgJ8svzTKQxZOsJgHr9W3kiBsiVfpNH0SED/
lwmuVRH2Mtm/D/Co27gYF+hHXbXkDzPBzmUDkz+CF1ITNixJRXizhFQgxCY4PGcn
bB4Po/4HR2gv4Uy/BHzmObPe0XxQouSwjWZrH2Uq2zGs3c01nYMyOSbKnY4KXklZ
68Q9fQ1o7EAUPAAAC5wf1OWc5Xa2UJfMAjJAEsav+IZLO9LdCo8zkSirgMUgLoNt
WEXeO44QN6urTZw2yIC/dAVAYwqzJVhcm8JLzMRVBXreHJs1Q2bieG+wzeStrl4e
T6u+T4AhaavDsizQxt/9gZpkqXiZuu+fQWSww9FI+1ghovMkKI6evnJuPP7iG0N8
o46nFqkHAC6vXsjziitHbD9S9bRWpfXtz5M1UM09Pg2EqxMTgNpa+IuBAMioSnDx
G+JwHekqM3yA8fv4atYpIxCIc4swKAj+L5xpvidY12xwuW3y6mF82NQzwbRe9ulZ
Nb+fxlSnTy8Ns/aO//lqYRWRsELS3xkP/KxeFGNSEPcGXgLI7Vrg3d1VS6KEydn+
GdA56G34TtYiIAgUdhDFqB6FSyWXdY5kgEg4iNKC6Qr4OXpNpfkHfnpzcALAAMZ0
PHFUzl7P7UgA14kXs96dAnJQDlsFwV0/XY+XIHgaMDAPOeNQEG+U3pybcD+cfevF
92Lap9TM6vOW91tkTet/m+SZ0XYjQKxSS+E85cZsqcGxPwufLwPYRSYXBDaNCFwm
z0vRgtepiS1pXRWZKHnlguXfKd0TnHJfwxCaSqBE7m8XldEIOgTBWLi8AHe0nxgs
27lEHol9oxNqrbF9jm6iscHdod+T+qvkEDZ4pwZl/se+Ht6voSP0Cpet8bN6yq8r
YP3IkskM1cmDIAXzfiYXlsg6wAKzEQLqm5rmYyFuq+MEBBT74eQFXlEYuC6RgLqK
KSwx5v3nZ1PjWl6BTryD3gBDVrepnyFSr05vCwbS+rMblkXEXxR1mOWIgAXiX3n8
r5DNgGdFYagaGQhO2PoecZ60Aaw93IFI0BCMJufSHNxhWqpTNmU8CNLCbnRrt+X7
xq3rY9fEXJQKncl3gejsNw8PRnSidLuKo/zvZoBiJj+UKKaAJyzt9aldIEHYZDA2
4gP/qra1jZTOxI0lXP4oFx/RLDEo+lQ20VN77tM9ZaWc14PIosjt85I7/YRjIxXG
K7jR9NvehQT6jU9fX5iaHLhHCHMDJ2ZVz8vprOwxv5E/afxUr1VeBDJSC612oz6x
SYE1xMpn2jv0Ume+gWeEp/C2s2j33yyOKiwlOL3NvX77JjbYPiEPbLYK2AMkzrBX
XJaz4whoUVMlq9AeA2jJfB9REbheiXKsXLMyXACpvr0yTRhvQeDb4QpwnygNeSF4
U4lRLsfyj1f9uSpXd5JNVGcWy/xNWkg7GCSj+AJm759Fi8HY6ADbswMS0T+nY2k8
W/4BYNr5g3CJH+c4O5XzdNt6bFz91nNqzeR3CiItRbCAC+5xrmMfZUL4MCL6Icsb
vtN2d8fhQmPg/00Yhq2dIVsrthZxxDL9QnJdDLIMP765tt5S4Cjj1L22eeU7/U1L
N5ecQ951V12cZMleHNs3ls4vUkl3tASJNv54ik4nrbpWH6+Osh53S3mWmPRLx+2x
7ZvqhoDqamaZTFGN2W+XLapfdXcdaywC9zQz3fQS59XwZ1hGKU9iZ8YiR91WOPrX
eNwv0vsY7K75umY0BvYYtsoHlYIV1/zQem8z4SLlVeEG6tk2iiyCXKWcPIfaUnIo
G9tH24KVWyw/RYd/jeos0f9CUoHM3pmBO6vzwjgdoQTT0LsLTvOdE8cuBHKHRXC3
IhsUBj2HCIP5S2zwxyWCWPLyhQEmXNDPYPyrJunX82/2aoHvgnDvOVDvEJaNxRm5
ctcobD5K/5FPcdkDjNnEPsrotOYOAhX+rYK7ghSXm4eEU58Rd83tPuM2eySeG0HZ
0cKupf0HUBIUKmCgI9EqAOHK/x10wM2Welh+vd6zi9xHA4jLxI0eU1r8BS7jiK/3
7/idJSDlgL2q6TIt3zLJqsdx0EIZ4rQmaGuANUausptyF9HJ4Nl1pFrDoDLV9dyd
UqTeeiJeujPmhv21Ny+YoG+NPKKLevQf+4jIbCe5DQ3hXPgNzFkWkK/Kd9PSwUh0
FM8NnxsU2+luMOh27zpNVsU1U0U+pZ23egtk1y8BhCCuVVxdFInn7fFj1+aR8EMf
NnjTMKJ4TTxHElseHhDNXaId3RaKXVOpWD0h0UGNGTSzbCbdsp2IINEvP8EFr/MM
iRN/yvZ6MbGV3TyAekEbg5rJIiKosR8Uvy0d73vi6gOcCXhE1gh+Qi/e2cYGnTl6
1wxv0cap/dQVbM36mqL1A0eq4NfyuLBo8oMp70q2wITn9UUtQXfITZoHvCe0/Kgv
Zfci5ijCMDOr1Ffa6FyW0bNv3ZRCMoXt6NlQCrX7326Hy6wEAwRp4qyMuObCgh/G
Wn0nnGkUY6JvoS7kYzFkRDfwBbP8DdEhrkLfzWk/Ky4de2GQmMyB8hXN/xR1H/Jx
7t31JY8G3dITwke7XE95IIcCGxVdaGxuOIL9RZ4xtH4YMhoBPXYRbv66J5/SLRN2
zYltyufxPz7OLWJHf8lc9P4aeyG46geY/9/S04zqAbH05zcVmHgpo3yTsIC/Jpv4
+iOHuwTWqTp/BRMZXaFFelsjDw0hwIqZgSh4hlIeIUtQ0PeQbl58dt1JlMHVeJ3Z
ggp84IJsg4ttu8AM0bsakYnNlnEvK9Kr/4lk/HbSlKaCOUp9kQW3kOvCT08/aoWc
ZuwaYG4YVMdwAneD5rmifMAeZ2imqCc91BUQ9fK/lA7ikaHKLvtLKLkZRu/ccqLe
SwoBzsYJqJXXJYQOqE8VKyHJLySJLeC+3sQSue7/ef8v8hNw0bxRdgQE2BaQR3T+
YqMnVkqnMgIygQuR//5VIKhFAocy6UcctlO6l68rj1iksJ7f6OU+k2EpkFStdW+4
PI9/d1F2jhEJYw3u2lp6VPxYsj5w4tqsNnBly5UMLZ8gfaJPOI4vfsoy+f9HLNL6
TYa6/113iqo2+8fWN60cThaxRF4QBFTqcPN8TmKNoNJEqTuZm9VSqeMrJR9aurlL
5DCwG0m1Vwd4moGqpYSqKke4XEu4y6aD/3Q93HG7WW4bEoPX3xjZAqNpQwV7mOpb
NCNdLfmBOXWDfxWH5QtcD3OMhTcGs69we94M55ljGhF71/w9XbRv9D4mJmpsXWBW
dkjobsSdURxv0BpJXbT08fMOZjVTnD/kdhT4Am2zbHG0mTi5jspQeBJDH1BE6vmS
RKii9tWXGoLyFn6ObSZNZI5Y80d4RTD9oMbE+fqyv6L72AiH2RW7jI5TrLPk3/Da
bztU9yHKwu1tUV3/OZycjyz7TBNFf6VRWTrzaBuviL1m/wuHbKaLHAWkC1mfcKXQ
+E4Vg6CjTcEd70d8RN5geoD75HZjCQIEDPQZ3WxNRqG0jNT8A10GnWGkSf1dFXWM
Huu2i0dDi4OGKur3mfmVNSe5Qv/hmnvX6wDt0fg0RlEfCcskB1zH5E1WzwSHhmsa
StinCsx8aevWlx8KtOf6sm/CQmoT7mhKJ0dYiUnKz/7cGTobZwJvHbNmQF37DU/O
+fZ25WQ6Htuwmmc64COhOQMcHSTOM6n8byKssHiFAvE5QgzT0fwp2Ei8oFPmaiHE
m5XOLn0qzvBFEd169BGSljRFAZQF0SqY4gdmDmBuTQCnjdzDs+zJPkGz+tsIbqQi
nliGt0IxSEow+EC0In6ZcNIERnep0ZFBkEvazeOUsOPX2h0JwGX/Lr4TPTZm4EnY
4HU7Z9EaM/B1bqEV8q3Dz/ZI6ADWUQOlQA8Bim9jyPoCCQwIx8IHc2JFSNvhIR3b
m/4Qn/OZDsz3oaayiydCOx1iy5z2qXKzsMGGQQxQf4In2mZBHk/GDkPQLs9DDImT
kD0fGWvkOVZZmODYiqd1hwXz9cR4wyeElNSBnXwJn0nW1/ikIomRjYRKBVga5HdQ
MSVB8+pdyrkfvBer0Jlc9WLEhXV/qRnYxXB5ijlfplq65m8nP+jeksUmkkjUsQwh
SYkEINYfIDv7SHmcgaipTDtCzsrPLo9llFKVxEOdB2+SQicP2MvogQBRZRhNPNYY
edYEgAfo6viyWhQ91PXuMPmU3do3lDmNiCLHUZmNBYzQFcWxpXaTVzZWq7+4J5Gd
jEnqIXzw594BFvpOiUC1QmNh9Hb38bGuHwRBkRV/q0C8JG3HHcA/3Uvk2U13mqbT
bKKqamn4g4jZ/2i9Dx0Zw4n4TjtEnVGG8FkHecwuVR2KEd2D/M/IZf6ipvwGxS5H
NaI1fLj35x/wlTMWIhwrX0R7UcYXzEuuiFO+gM2zXYyNBYkX8IlP1CuWuNzJRYRc
46+rjWgYloIu6mYaLFAsqq/QmI09GUq2OmZbbRj6s9bxgajLGr6rlHP/hthiRK0y
UAgE0JfLmRj13L4+L3BR9hTsN8zEp+um5i/bvxRmoFx+/8eT1N9fMcvKjOxFw36u
Ed6gTW+8J7M2nzKVWbwXqEB31j9ahnXNFGkC4+4uMjXbAkstEjxDLJ4LyMyrk7Uk
zaIr23mz3wkjcaro+GMYTb2SyS+drqNo8mYQzNtYc6wPtngbi78BKLD+rIEF1i+J
XOSROqS07+ijX7vas3QcNWaw8dfAJ3lU+rrZXlw9L9JDJ81cQRVukP1iKZaDcPLq
TVuUrXyE4gYRaBpNA00Fg5/v4P8RhOMnC5HJyhR2151CYAl5t+Qhz9EXXfkzjELy
yJvaaJjt59gWiwzt8Y7gcaQI6ioiHrfYsGI5JBEDo+JXx6nIO0Ti3GBHxs11J+vG
UFyECSVpx9RmB1MQt1yP8rDoODRGgNpfJC+Zcs8QAt06OXUF+UEmTxJcrDM6iy7C
aR/u2H5YVsH8QOANS3SfrxcrX0L7vtCBsH9CwTJWn/M5mgACNpNh513aYmB39HOx
7aDfiRZtPtz3fm7ovSMbXsTbvuST8uLdK5GAqcnIEPQL3On6tn4ZrfMgnl5NC4Ug
oMrr3RmC2AcvXrw32JC4jOIBQYdehl3HfMQIru4VBvYqldGwMWhUUIbGE7ci+Y7P
6NFQRl306asfPhMkyCdx/O6eWKq/OY8P/C0sCg1sWxsXHaxdshanx2Iep3helYIX
4ElVyXAJYukB1gNtd7V8S7z9beJDehdFG9UM5w343kqEtifWGQ7zIniXZo6FSgF5
uszz5iQgpCex98PoiNOkm1/cbzqVgeR6yVCEs6H+UIuzV/+tHFefPEfiPW4rf3GM
VXlFY8Cw5xggaE/TK17j6FTZcjCGy2gYoiuiMQvY+PAa60zEx4DMMzNDYCEAkWaG
it6y1Br6m5s/4BpgTGSQUK1bY9mH3YH4wG9t6fEWeE8GIUcR9NZy7AvCKp7/y8Ne
J4WoKriIpztXIccPUt10B4HBvr7befRGoYTiX7GiaKtFYwfsZrbPzYJu3BI9XAry
7MceMON4EBvqaKvCmHh4vjDNtelcTjXbyA2ysE7Hgk/laUpLfFZvhmrm6SLzW5Po
DBwTH/02bERASisUBkoMeIFAZzFJ8OBt76qp8GK/VTs8GLfYMmQQI6VcqWn58ix/
rLudoJos5xiixoNYoE60a23d/tC3IQYvpUfX7mmjAHm+i+61HzklQ1BFtNRjGktt
2pWdp820vHcNyFzCbrMtlGnFZ2tGU9vSsrxQcWDaiyJGlOB8X33LwlK32S5XLpfr
m9wiCYjlN+I/H55XY/TJ4OWz0zkLlk9OizdOJR9gi2x6udy/DcfzVbD0v+Wy7nAv
/kJfvchiLR4DPRphOzjfk9hJQqmVIX6mFTPLU0mYf3hjUlG1B6e4GLLOvVgQzTQz
FCPSfF0HcTX1U9LEXW4WrwT2VtFFCjOcwUwWLtp7yaHe0D9+//VZmmXhlqX+g9w4
Wi1bB7uNKO3u56LuhM6hgyEWI46jQdhZroSsoI+D8vS/wYJqOUUyzSRLRmPF+0Pd
wBLqkbwiUFKvWmZrbEzKbqL+oWkNfN0rjHlo5dBbUwGsbLImjKwLCRCxMguYKR//
9MDU7KNmckqkxsJKpBhf16AZSOPx9JIbiKI1/Ru6DzstcN4in1MKlsvlRTn5QzKA
DmbU5tbnuA8fMj0eVfbGRergGBnuSqx2oOZr6UZNJQmBluc4yv/AhDWHVghtlDm3
xIp2TNa+PUpAU/kpedaTE//aWn6Bc/09N3d9JVkiDSUVlaW1LBSgPD6D7eNIozPh
xBNCfSmKiDmvcaH9lIKmP9wsgRmrZcB2F973lG8UBpdSoc+c+EByIGvzUA4+2XJw
ruxJsylE6RYvFvt0p1dhUPnGVaMrXZ38Y/wnkPtEvd2zXltDHO3Vt/KmcfhnDz5K
lEHLkod7YohpKojB+U/7d+Lgxpoo3hbKE38EZYCPh4NJeoaEL9Rk8QnzY+McPvZq
MVdOH6/29XddXN7Z5Urp0UHntkNe5wob48j7Lgc+2A8qvvDqPvLODH8FGAnsm5m1
aa6akAAWsocD56HZMuGmG22TfGQBd2YgTIne+BkHHiVrf7+lvMC7vo7RirMhTlQ2
qhU28oswGET2qCJSBia9Ldke62zEUGvn6zHEISGUi+uas7Kwbjvhe2uodTq4Uz9v
rzt73rByFFghMfgzrpmSQqJ81pu74RDTarYfXT9gPzwYc2knAlBRVzqIxRau8fKA
ibQXwNDryt/3PesKjec6/LKtv4JwBZUM1jfTg31yYHqsV/88gLor+3tILJDzHKrv
GqDmctNiuffWaazqo50tWbtqK7E6Znju7LStW2DsSnYKqNf2UkzfEor4TZ2eO1zX
/oJkgNULlyYQ9oTrhktm/tSeM2Fp6/Mk/uhiIP9OXATn/l7QHaQSQDvSLr1jFwuE
Tgyg0gq5E44SGQtQe6yExBP2cd3F4Hp3amsUgbVJfmJwEH5HI+aPcBI95Dzz6cNY
yhc+BtFiY8dwIAm5WeTgPqOGu06GOJVuMWe+GONElkUxdAO+tuoYgNNTjCMF08lT
J3+uK1lpqoT6t1AprKLgkjJUGDM8fz5gKziaigP4dLcmuYvWsDxhQ0eJURcNGose
yiE6RTNw5k0iaKuIVtUZiKvrPHQsG3noedBZVlZPC1S0vUoLGWTaXsdZca9b/6HH
y5fL3i9SBQer0uU/cfhQWcQS4W5wJTxNl2z/T9xQoZ10Job3EZHN9A6UTeICM25a
w2yNq4UAk+olbtu7t6ajJonPS6VaMgo1p8+/ki88XhzP+7HzSX+k7PdmolFtTaKv
3/O5PHmFQmCC04pF1MEcNHzMvRvPvs/ewgvb8AbkxhfGpxP2+D+uBmuwRBsCTcOW
fH7rDaiBT+tpOZnxFNOmwPLlm48F0dmsA31g7xuIcIIKF+vP9hZDtLoWnhBFU2Sc
4nKmdWWxnwthjH6XTQIYybRyqymRDUMfkWK6fDj//1MTqnTlMrKjMFRIDx0VgSZq
cfP9PX11X5Jg263Knd0ZGNIpsSE/Sda4kTxLGyoQ9WWroIQoYmshpNTufggJJVKr
cNEI5vCiOi5gMe5okJf5kb6W9mRHW8phbAWPp3AI/eAM414jEXY/kPVixGyPX4WY
92UDRM/zlLvC9AU0SnFZpiN0KazJ8AfJ7LKNqNfYHy0CLbGM3MYFnyVOpd0/NicN
/R//WYJElk4N2vZnbpgQwQYP+Oe6wNgMlojEI8+nP24ocvdtvtqweHas15pxRk9i
gnIblSVI01EO9fQv5J+ShB2CWoQoGgr2ie447z4/9UZ7cZXkvxHwOyfggFDfWhz0
jlIYM5Gz8LJhM515Hs5ter6OD4qSKViRhsEGkhmEvzXo+N3JBT2KX2qXeEDATFiH
MyRHNiWmtzQbCSxkiipBEgLvDs2JTCl4p8ba/YUr7+R0IpF2S98EIOxwSjnJS702
2QYr1awfBMk4WoDff3YyqLwFn/7ibqZPx1QsWEUiwanwQXGia58TXBFqYtuqZx5Y
J1Mjte2ynQ22NjYqqPJJYQnFJWwJplvZ6dpDYMS6MqHaFhTUuoD0uT1ctcqxwOU9
TBplhc6zTVpRY+Siha9+mZZX+GNCDoujPfyNndOqwUaAdcn/XsFwMyV/Qmwlef2Q
BYv7ykheqpk4BJG+DvogOeVG9UEw80En6lTRpYEPTCd9oychKzUqBx7Oy8zPSMcQ
wzo+XC/wSSdVU/oFcvzsYKWuJNda/vZQjOfTGrpnQ2gLfLIIeRPbAXif1y9H1i8h
/2POBnC7bk+5IF73mHoKoHK9x0HfcTKB/bILVA34ViLdN6Vy7e27jkMphAAhXKZP
m9Ph+ixdVw8k44tXTtVx7Xd4G+8y3rg3CsxDFYspR13lzLCObSf+K3iuMVbimFrS
CSU/GRMyP3IqE95wSo3vfovezfb+4JdpvTygHCulq+mv0G7mLZwwVvyyfPGj90X1
zKF4o33GKG2DdSYiA/Nk9/oiTSiefpAm5LAlgs8eL5JwuVGOEDn2ZEWQM3SXaZ+q
dS1MJFmclFE1wTUICRTUm8dURu+SMvej4ItFIOZ+KrqJUmJwZPxvTkIw6LOFFKu4
ndNiWhnTv3kU3G9IvjzGnAbcCpjASnOz64ZRo3CeAcSjaIrblcLr9HML95oTkwbF
NRWm2CwU3oair9XNCHarR/1l9tcZDOwRwQohFRqT3YIDrKevRJfMZz3FxbT9vtSa
fXNsP0J/cRTYwP7K1Ovv/FoeFwdI+VSWE/vfCSqY7wuhVlkMpCac6r9gLlPaH/5m
YcC+OVkbSbbJ8Lp4mpkr09uwzyKbS41nFf+kLToRBA6FILGnP7opp2E0+VtMiCno
lJp7+frQ4t/py4RsYE1hXea7UlbCBw9I+8MD5JYWSmMVdZxnGto2heUxuYR7XTc3
TFY4EgplSZtd+jGnQ+7EOw1rysS3XrMSycmmPz81mbsHvcat5BCiisxTPlUueJ/W
eit16unGpcAT3fVFqjVfaIgCysl7JHIiJmEnwt/CqQDN5zAtHkZ/jEutZhW4F01U
6S01sRlKAlPPIFFzTYAP8Kz2eqN5st8u2HUN0lTQw9ODdn4pGVfTXyjEkTgyCPin
KC8eK16S8QPgbMD8kBZsU2uPl7S0fBCWOMwWnwuw4HarKvUGXGEJ4tVMTGP04FXi
lOrCWs+AOt/8q4MvU9dRaidyobkCRLKP698Kp8WccC4M8ZjwOmhMoOoNOTrymLNj
a2WThmkUI3OXXw4qez7FW3GREhlKELrOfA+pQh60sW++I8Qk1mhxqpItgeSgZ4ju
omiohzvVGXsig1dgiTIhR8qlDK51LmcAwaYcrBD8BLW3ne/Y8We5OoIk+P0BoEsF
Od5JSw5iJDsUdVGd7uKxf6Bx/u7TUhHahjyV+CGg3yf+uXaz9ztgLG5LePtCc379
l++UUi+oA0Vuz9sThEU12hnDYdUvtUxIbzCq+5EtXucCGNqvUzX9OiemTqS7uVlJ
fwkken10gGRWTkzFH4aDTH7YIR4bSqrsEeCpdNAMgJ62UNT1fKwLRjww1jaxKDy8
3HEJC1hQJOczoUwFUyTW7YflWJiy9v0d+ttusx2bFQxwHDtyGQIUuuFw21gOQu1E
oU7+IwCgKQPWhtFikEgC3sfkDz36Z2ZzzdvPS3/G2PrTnMWc9VSEIzZgne9HYrN8
x6uVLml3Sr+KqiWAknKxL/HtPVkxjQBEkjZh+4Jzg/HF/hTPjqgSghNS07dPC/KG
HlaOb8IhosGKDX6iiLf7Z0cDzrsOWArRoLsWRVPHqGAa0GfWx+zV7AciAESMM5Rv
UfQY3HleE+Xt+GAZOPriq/rJlA8vXySGSCXc2j48Eu6Y69kSzMXOibfVQhEl0T1b
7n/DHHUxmsgAkgxAPDmABmvbNTsH7Q4krpIX2xlFPhnfOcaxeXCpmdYc0LmV32a6
KhRgvdjXMSshofi20+pBDr1bLe2IFZUnm9d9DW/6Bw9uFjrhdBH+j64RUPRjr6yp
sbA9bkN2CXNgWpT9uGhTGy3QwQEt9xQQ4FfvyccBMAnHXrAPPXAH1ZvmW9URO0g7
75HfUU+pUBMC4aFzPLkIUNq3gA6Zi4008ARWy5InC3mcbwbV8qx44KCVuGX4X1N1
ZPwWzC0NbbtYAyC4BAxeiub/UKbVCgIh/7MpPYpAYSR1PgNAnuASuBLxBG/2QnRc
Yblpl/lvvmduD660Z+0eM5WSv33r/TvKZHBRv9lBPj8a23853YRPW3cFR4WO6FBL
P/apT+54LGTgXISGnSZGjuLDDebkDooF/wvPeSTgDApMoqwryHRcaSYZJezBhpxe
5ASozA5UqfdqPDEPzhazWvPWMgbXpp6BXI+0blLHBQHJjyzRJ33H1jGH62XhVYmW
rEWI/EGwJuOjfScCbgMKJKyJIA1cM9wkZpt4WcslcetjpcpzE8z2oQpljRjsmJKk
odd+6mclBJrtdMNgICRZPm6Wef5JW3Vq5umSuRyKK/DKpvXAK9TqK7KSy3FCZd/D
bclKBeBV28ZyaIanFAoeNRa4JkvnkClzRp/Co+V9K4fxO74dHfiMbm0HrmvegEuS
3iYVHSpYNic9LdTWMgAzGPRcVOOz8zbT1FXrtY1Az0g9VZmZ+08j0EevxlFAUVGQ
yNzj5fclGyb+0mQQGbaUwdBzLIuZMzQoYjCUPBWvvEktldF+VOKHazIBpi76eNn8
W3URAeaUKbVDUH3N0oLVLW6N5q283a2rfNCk5e5uUEKrtTkKiMQoRLTWu1d2c3RV
xIimNM5YfjVfktbfEUjP7cWC4UMOsdprvmsmCZS6B8kdW5iDMpF63dlmJYG2Yxz5
eMgJ5i3af9/XKDILi5ih9NT1EiNTK1ZBMEbCAnCJ1o6jTCEAWOJQF3cAsROXYYpW
xR8eCkh2SCfEj7QxNUemLc4iwN2jgt71CuyLkRQdjFzb9q8Db2PGojPhEiybRvn+
FgaB62W2Q5Y4BI1iFXlXGiEQHlLxMdLvQnD5TWoMcWGDWfoFZydxyyB2L9B6LurC
f9j9v76K2+opfg01bVXF12CSytPpMuENZSPFDfwp/oNR7ka1Zm6+PIw5rfOsEmIo
QNh9KU4RSbK0+vB9vsfPZXoyZ//vjZ9KKWKHMgePc4s1UJn0yYyTXMR7P8rH6WeS
SXNz3KQyiPYocsAmVFsCdpHXlkq72IzkjgvcuF92d4NpQ4dLO6zUXnh5XnGTXG2P
DdYzmQbcwPRD9IkaXdXHZeY6PaMymeLckXmRbW2tyV9Mzh/0h1XWq3HdksMLxqEa
H9sWGlpUaxxX5TVGGfhIuyyERTkiXunRUTGU079QHCMpFPEwR3rdybUyQWtk8sbR
ZdPLBXYOX5JeYYCwrEK2oCrVePPRmeOZBHxJRaDpk1DvppUHquY3j9bitk8z8iE9
KaeveA6z93WQ05u/yyjEL15EPaJxo7UxyI/XHXG6MzewlKAhCY9NxuNpTXuwm27q
Js/NIEayM5YyZYIMvW3HOMHDhMTg9BdE7JCEzrf1izvf+Hhh0Lb7UnueXhHYXT/J
PxixbnkRSnpnAtzg7TasgINyTHuV4svH4D1UFRWzs+HXfWlzREL6El/Yr/jQyRC9
2kB+fV4cUS4X3ncHDZxYsDnV92lDwOSxIcL6SrP92GKvS0P2yb0mmi0/RmBqrdBQ
U3r5ULKtQSGcBK+dJn4LLmS9WYQ+Jk+xAewCl2hfH4T6QZThg2+0LCf2WG4jNQmU
yYnDiZm26MTTdHTEGRhAVLfFTd2gQtgJZ0o0M1RcWA3z7ZQ2bPjKJ24mgaVPXzGS
JB08ubFi34it88FACZ7VmygBM+e+th8H3c0qzgpOSgk3y/R0Sb0E8HTfxnCAXLH3
4DuS8aQ/oJnV2nGYRcRvVcCCRM9zmAP/DqJUPFar8usHeurzecdJ+G4Q6aZa3cPl
ZYM57U2ItKPC3bqsBtgLCftHGVqE3aXwFJGNnmvj0/6/LUIXAnPDKySdxk/MrCm/
XlNbkVMHiCHqd6/sCv3WyvrAxNXcbEMw9/QIjEOkEmDgFr8p13LOF2dMjDg3neFt
trGUvRrsZlhL2TaEjWO303c1NIVfAhp+e+uTCbV1LFTHKvYW0DdChw7S2xNse9cQ
Jp26nd43Na6pZTShgcqoTODHIUgz7Oa9tjDbMp7sa8E0Oao55VxVGiai4usx4n3u
9jPj13pckaLG4zIRKH/pj76w9h+XO98nEgz1FHLfjqbJKz7ixtq4LIawL6R/Ky00
oKIv9sjrqSY1bSXmTJI+52U1xZmiBmGo9JFhAnJtr+k0PulJwdzKChlTJ6DzGbTp
oY36z0toESCQJj7hrd8o6hZIMTmATlUFlNiCxwaifGGybpC8F0iBYU2P+QmA2Awu
j3J2Gi04/E0my5/DCJL0JrLwdOFr2WdrjiHG3fbhKOlwJ6UssEvXTp4eCO+SEZHa
hH7lfI3rcvp4+Lgovb01wQ0g5/8AqvmlGN7gnTdNwsu+sliK5uunzo2sy8qYwI/H
z1uzMdTadW2vstY23JjUYzYSvuzc1LAF3yTtc6hBGAirgtJhA1mexvD9mfj5Jg68
evcg3jXtxFRKprWq5plep5IkOcrioSXZa0JvB/7m95PYLFfslMyEWQUKkx4NF8mM
ps/rr6zenYS9VwsdN2HoEw3RB+tjHGuQTfIdnGE9oSfknFX4BklAgocCzjWsEbWF
qDA8EzbgrG1XeVqffyo2rQepP54Av0SLHsrcPq1hSJVvJdO0/xjmhUs4624U53uB
IF7XsNTshkjEA9m68eNlhTCcE3GDZqo7c7pQPauhhFMnMaUFmbvfdBQbyzRSewMQ
ZxFf0u2TGs4BnIkjIi5DaiIDNPgH04Z0CkAEiFsteAyB3Rn0S/Gf0B5RfcMw14hr
S1sTsJMnf84erymfG+lbtJ5faQRsbVaDx7HZDYeyFn6wZ4Wnls3BOS8wQUmegSJY
TFaJDlw7tOFDgKRg6qeOTJboxve/PXplqiXPIkntm9FPtucm1n37+GHO+5/iIp9B
Eju4py4FOb44UsW5ppX2vAR+LgQ/yRMdvzUEYiM8OahOpWN8V9u5He8ooE6X29NT
nAAX1nXJXPD6NGS+hSTyFHrbSpBQfhEZXEuv17fzCw66vRfaqVRZD5adCEXX9OcU
ro+qulnoVpaL0YX5SA8iADXQkRLOu/6/jEEYKTWREkPcEenPSnbywhMP0wDY4Iv9
knzHkC7eAK263JCQnBaLJ3YlISZCf0P81wf/Nrhh29To1CKyKSY31MqvXG/iJAW3
DTasiFrfR6V5L3ibiykwdxDtVXbTzmBfM64Kf7h+Ij4WtS/8qOPscmHPRgew57J8
vFtSXx1vk5x8E3jotN4SyoYAP+89cNvydVvD+6hlmAsmdEESTAq4P74tKg2eNEou
84y931WHH3f/C5krqCh72jWChvihAggXSlho52hb1sP/1TiCDzAYtTra53mGYcCo
Gzvz2V5gcXWqqGT3AFVKMPVnsvXbU2xCvUFhhev023le+fg3DkrOn+UndhUBQdS9
v/NKoZ9YTXjBJ3O2Oe0cc9SsOLiSrfkT87DIbZRIDt6oIb/kld1SRO8Yvo+o6wrm
MOmSgOow96q6uGV6M4beRlow3GuR/VQjYyK6/UX71blGtzTNKUnwKNNtO9w2D/5h
kDouAmuJDIDFPYtj5ezd+sqJl1PnvN6ob+oOJvA1k27Bt36hiz3Z0u6a4HD91HZJ
Fg6jSG5iQU4g8MJFjMUkuHOusHZM9i5R9+1oxWs5E/6hclq2oV/mFypKxtjgX5T1
mgmHrUvxw2IoiBBxDXVcmiE3xqv1fRBIFWuTqbc0TNwO1YF5J5SM97NveZGaT8Dz
A4FfOq3wbdO7uoDNQw9q3fyo7vahWI5MqfgEWKnGbucWg9DfMJVR+gf4vaTtF69O
aanBE8PNDbOVx9QEIsKJUXjJrxNgCWIqyUHdfbcWBeONiL001IVTp/QGtF6TwwGX
SUnfh5TZd88pXCuppsuGG0xG9vIKdonq55Wvmf2kMRo0BV9hl1daZjNXHFeVpm0P
/8tZeMLrGzIMDkvLDvNmDnWQvI6KE99N3DTuSrN7MTzRHkjolTdiyqrGhaxmt62O
8DYVtxlnMl8Il5drOA3QJEG3DcgtoT0Tvzq9yIfCcMxa9/eJWolafcli8E0mpnXZ
GxKIaZR0qzB9Qwqjf5KXX/4H8HHFjNXhPGJp77WMH4fuzBSNDdaMQb4iMFxh8CAG
f4ERJBlir6mMJaRaYJTmHnEgHpmA9IEr3MaOjVFm5W8Xu8RRzrBoDN0sHFMfjCYp
2ZMjJoztszh2ub2usDdcdqLDMf7xI2MyB7xLXm++dB4pmpJjnrQ4a3tpTtb+LU+Z
z8lFevZvN3l5LX+UuizEuUBROWmoZgxvJgYVA/P+uuY+B3DOFJFiW4hOye8OrnGz
xhjK9/W5g226faYH02HX2thxKIj4Vt75xXgik5/4+2lbPfUu/Zb3Gk4WoncfKT4g
OnSYlcIcBiWnF/ln2xsAcisuwcYd8HGwRdWjV80w19gy5jsWvrEuFdcZDNhDNnqY
KpD55btzQ0pvO47wN2+ACyR2JT6r14o4Zrz8n5L9HGsUjiuilWTodjaXpyLcYaOj
dw0uXP8oJIXlvflz71t0Mf1Ty4SNhk0XCpZmHWj2gOwz4NVe8p5+T6+2RrO6Pbco
cTHZEutrg1uAvW0paaGEJJnXI9NQnld4cLqk2qJKZulYNAKkeZbdJi7+H84Ykt5Q
2WO05iVMqra7C+vzu6fHoEqEq03lawRq2CsA/OqAFw6rmtXXbQKN0gwiE1k/gIXM
12P3U/HLJ560yoFQPKDgp+WyqG0FmRQsD5fJVGum4g55IfFSOBC//TvlKCxbHam5
nscGdQQpOWr96L1uOzPw/eRWJjtaZI5acGJF1t7IK+ZR8hKC8dFTCo+U1jRbzOls
TIq4YSZqlaX5tmlft88cAjymvye9arkg8bpbr2SlhSTe6APfAy597wMIhPNvyeD5
2NuRTGq3iGCgncDbWTV4k/meEWOHeBckG1fkkW4Y8Nm9grSeVhMGWZ5Mp2LAOVoF
eDeKJ4aZ651er710c3sIWDJqBn4MgkEfVKU2yQKJVD8YAUSwRXwnt7Vc+CvdCGq/
+mwhwYFOg3KZcCuBEUgQMO7j5C5S+vbaMh+zvtrNuNzcsMw9EVZGWlfXz714iUGs
NjCbtc2k1wqCO1uup0cPKaAXJzsKVGHN31W7hwnijDhGGihVK5EZ+X/UNK/M51q9
SW117JOYezdoeyGHbUMDw26KY3+kJP8akk8ulCA8awXI2ronbQ4C9hizzFsOh4tH
h4Pt4qb9mDe8TMzBphCqGhytcGd8qDfuXL8YWRN+9vvZzjQ5xfpfFENm4WfzYuhF
OZjtR2Xg2lcIjbnSRK8iLJfL0Qm+6KInGw5A6VfmZKwpo5f3pwWZQWAHgUMt6yFj
paoHqFf1H4vtwr1vLfcp7ac/G5RllNszVMvj5IE6bSUtlR3H46cyvGUjS8FYlKK8
pMqfAMc9W/L8G5Pi6rjl5q0hO7s1VqhL6cfdQW6ReWGub66N1UCnpvkLV6t2hFDk
RD4iE/hWhbaHXEUqcJtBnIUih1aeNwLAVG0QzWugQ/ILCXU42+OPppnv7scNySgp
Ga8cRpIDhk3w94tDUde1OStLNRwfxtJGBNbcEZuKeclojenaLnXt1RkxuOf133bq
ux/uJh1CF49Ds6MoekOPCPZ9HH+uVNDjibxLff5TN6cDfXIcmFKJPAFvzv91/D7n
A7/H83/L86uOD+rKPxjXB86wBoR2DaULUv+loYbuaHEmGdCLAc4gINJBL82amy8E
rPBcIXDBVl1s2GD65NYGWam7PDCJjLMlPuiIZgp+kT5vq3adayTfg0XelbfgqI5v
ETtpnMmCone0i+81Dp1XV3aBu0SYgL4sYAvPEEWWrcwKpHPB7eoyvS5Nfkh+E43J
2tWn8ydHwsZEJ+b4kihCpXpQ+87VtpXGMM6MYn8gPyLXYvXTLOUipHKAG+ACPigQ
w1CLSVfEc2T5n43kb+gFjKTQVZa6I4fgbKUAChIKJTvq/g1Wc6SYM5uVEGA0dzQH
VJGzHruQGHNdfxN/FgwjU5A9TmzMY2P05ZQHw8S3fYY/rKXZoX/usDdz3+lf69WQ
OsgY12H6C/BT/YogyqPN1ULye1QCwCLaNnidK09nOTvbx34LCbzXy+b048N3mfzH
z4jtIKi50FCNyjvBPr6bBatY+IBwBXFRBLiWfNEuBszS3K+oSp27PdCliNxJkOku
U3EfKYj7XC0/kDzPWe9eMWBI5C/o+DHtQJSoBjX8Rzx+s0kvP1vbdFQUBWrPdxkn
74VtKmqDh7PMjrwysnMIVhj3vk6evTNDEvqqNsEHcLz23/rFx2BDJrm9LI4ow+3w
Cmh+2NJXjCqL7/RSndZEhtL48nOOfe6dj72ePoXBVpBWpzy4zm4hzaF7FmP9rDLs
mrD/FmYmoLTzsEiA4GxaZe5icpWDGxJgwEJamJHaCKLNOAb2BTjyFJ94n36BWntp
lzN3yNmIcpilL6rJ5Uu5XP03j+e0Vqr0StOxxbXvRlk0OvHc3K6LIYWL/GTc0MHR
1FjGks8FJePP/tGw4IkOxuO2p92ede3UPBE6TYOjC99i4AO6Fv6CsTgGQZ6M3W5D
vN9lFtk1QlK1M/ppsfg64Ub3ESLUxgHQH7fPQbO55FFoOg9aQwruPdb+0HnkyGkh
gqL+dL83rr/MWIlIXpoeRwEzKGbbOmstFeJr+KeTI05aPlEuN5tvNFProvXfVjOw
Guvq5BlTJaCok8UCNrCz9b8J+BljdJMnhjm2KFi0WTe46hyRFMT8TViTT4NqE6pp
OUsIQ96vjnkah1Yc8YuKdL9Jov3nB2Rf5ZRstJgBrbjTPg9N/w5524E22aK+z6Tw
xxLvxsuDVPsqvDhFJXzQiBBOLQMQwkUGGtCxe1NvquOs9i7TEzs+OqlPqddLpxnW
VDTYI4Rb88hnxwraSF/gAkfl7dbEB7FXm/Cq/5StbIjr4DE4o1J7hOCP7ONgyfe3
muRA+kCW8KtyxmSx3tXulA/DlPh4MufqhTnU0GSHNxP5rWs74FY+N9t0KcZq1Ift
NXJL3lHtnTKp6BX2neTdERmyYfluXF4zdB14JLgkb2s0fc2HbAOCDN6pe3v3FkXa
wkdrta2x4rxUyJg/FeOmtr8+4vzH1glEGD4IJqtNfC1n79mhwA6bnsAGXg3oylZ1
5Zn17GW8dfoFPU+Lr2rh1iRqSBoY16ajU8ahp4m2/rI3TJQICNSgwGz3L3zOGzOj
1N5M5keAPx9rI/oXA4f07dINCcH6TgnYj3GLhw3Xq/74HvmQWsko/XgWCZHxImiv
062h+Fqx03hw9Dvb4Mrj+prTbpnEo1kdaYxqGi4U0Q+1eF9nTnQru4qBxmm6714t
yP9unbbKobyYJEL7ZK/rlqtTD/VWMm5bfjpqscP6Sn/ZU02t3we6Le4kRHe7QYx5
/Xw0FR7kmp/6I2/27m/nHZ+JV399tIQHEnHpZ8n8e+k19MKSI+caJnKiF7yM5CRM
C9Trw4aFNFB2rCUGovek3TljYiYhBn7LrFbc5577DuBsi1KY6iiq1zuPnzfpRkE3
tNWNAbVXwsrkpOW3hUB82R4S5iFoOt0X1is2sLSAIEVtXHkYoVRQ48sOHFRU26jk
jOAqUzsmnE7JJeBO8KQJSNRoPbqof5JALce1uVZcRuorbrs4YJmqC7vlCaE0XfiR
SgBHwg/6jhyBR/LwS9koK7qjL9k1YHc/l7U0YIWXytkUuwrTrrMtIFO1cIUY5/lv
fLsaLqGWDpBravVmhO6Xpl+PMrD3aAXO2unEyx1gqir8o/IVtk2wN992z4sn+YB6
9NUwf3kcPo13DsicbTXs8VsRV1ykaTzTiHCIy70vvqrh/HBqUH67ptilwHDfVvJH
E5A7QqCLwdnYQhoMFqg3ozptwbvy5qA1ZlaNh8sRfBIuC1p9xC6AFSCJJPfvE96f
UI7Aj+gKDgcWHz6s4pyjmWqH+KWkWeNR2PYIcnIelatJMurg/oMBgImjKTdP031H
embMuQkGpD6rUBWsTRIN1sURjBJ3j0O3+W1l9DjrsONpC0qrpxbKLiev1caYCPUX
aIqgq7CLWn4rzL5KH2vhJtJsukda/5q22NFmpSoOU+qZDxO38mJR0cxZLzyiOoBq
8mSIqnfQDUw3x8vC4i1SmwuqpoZX4VnfM5BjDMGH83UADYlTtnJEdgUXbatlyhcR
TqWI5FvrWboZvk1carcqnNmh+9T1h3z+iFTfPOeYGClZYmmF8Gv9T8Zv7hmLbTCI
5uPnyg3VPlhNNIdyGlJ7VEv7jSEXGUcmx15MM/hDc40LsYkrpekSzyvijpLhoxBY
aeCvSk4ywVLMezRtvKl/Smv21VpVp7e65Ol7O8pPhZ5cso7IniX+PF2hBXwHhaG7
wsIAnPZpdidDOz5jWZ+sXeQOoKJhgWUVJAkczjkjCiLEYZYaqXwRLEI2RZshwbYz
91UnZ2B7L1m2hqfargGlpIGauB1lNlfIsSvWCvyAHXxyaMUEYJQ9VIFbzD3kbI68
xWL1atAOZzrrj23VG8iSBI53NKWzFTTdON7Zg9uf2/GXPEqgvGCq4lGPVobKb5q5
7V4y+tMFkfEicRPHWpYYUGq81hhW65RdrGXP+/w9FzmAnJiI1YjW+T7xwdUJ+czh
koyw8NuXEUQ/PrfRTeiJbU3hAO0q6vZaFdklN1AnSSANqNdiW5v8Xjk18zJAjuVu
rd0ygCStrCwmDscKwIk0Ghd43p9PH8dBRIHyAnV8JNGnX6Zn61Vk6aaywipGh7/h
0+OcU0HmQ7mQKL0R5TSbWgX32sIh3bZm3ndV+DTlcSb7ZHxxCgW7AlXpkDNG+dJq
DLpIGYvfy2lVHwOxy8gdmU5rpskFDDWqOS1yY0LNOCLs4zXK+L4GSB3te1rS7V5f
pcw5Yhzm6fNxKDkon39xyvq70l7wZW5I6ANSOwMe+JjjwgPXpJ3Mhbly7ZdLCRnb
6tSY5F6QpGUk16i3ks5m6sO+oiiIQccW74+32UZ2e0f1W0YD9/tpcQs1w5HW62Wg
700EeF0Lm3kR1TFCgUrdnH+yY2PPzV4NGh36yPS2v3TDDyR/hqKrI2cBiTXa9Hh3
Jx9v3bff7wfSVEwv1UXhEDKY8i9K3RcqEbIwUNQyU/LndylqNtv/0qRD69rvIHuG
+seXH0glaAy7ZDSFFivUapHHQYpMmF9hbnXUfccp9KpGrZYBzdGeeyN7aHwu7ZYK
yGO8sw4S3o2uM/jmzC0jA6lGnMyYKvpB03DhDBIwnWuvQYYMSnkUe0m+5DJ1CWt1
jE0BLGSoy7UgNVhi8TOoe8NdoTs8O5xbpz70UiR7RDmAIsS4WvG7LJ9smArr61IH
q0uwv+LvzwZp+grtnRHT5yDt6Mnhd3LAa+OWC8xO24Tk56l3HwSLu5+yJ1GkQF7T
BKHMp6FDgkeofDPBFMzaRFeKm0+7syHI1gN1I2n8xRU8dhXludWGQH9Vou4tGVkv
sdp2wFsAtaRooPNGFe0KpksYdDDUSdv2NB3LzXyJHk56g5v3yKRbZsoRmpN4E/AR
frrlY7HKxeDarg3o0UMYvNHaQxbe9p78M10Rf1aFjelzoY9qvGekU2n/PqAZibWz
LyOXfcE34papGEmNXokDI/F2vIUpNrzBGI6JLc/dtC1BjGoItAV8DDNJB8lGHkGX
0hGh40biE3bAtLaJDcBnt8IR1/flHss3J1OXsLPCf2UUfs3txPvFoZhZTRIBgWaR
3KjlxZSs6kLrTxYwnt3WMv2f1hVQ8ZtXysjn60WDkyZvrgGSmXcyRrYkCy+9JucC
9vJVaITIJ678UjnhMymMq+TKN8GoD7HJ2mFA/QbybdZ5FJoH5YLcLvMG1rIuqD/r
evJQ0HyxWCX2oVH7cJaqVA5nMQYVyfX38VS+6D0O5ERfwCWK04Dx1BOQVM2ZjiMe
CVBFQs+fGOSu3gHDTG7M+Qn3DvkezjVQ4LK64YlaYjOeaSRLl0+KOCEioZaGC7+W
HhaSiOFY2EdB628pk1tFAFPMzhYas7PHJOGIa3d+pRBsyYzculRGIEIEUdIU9+5G
UO2PyroLlQCUqNLtkeddZ0iPOckMJZQBRI1RE+Iv2/JdsRwzwmPB88njOd14/0it
bdOk4ecA6fX6EHzDwDkTBfsLxXpOACmDFffWwsPwoxnKpUns5U9VUECwPmTuxkEK
MobAPYFaiNFmRxz/tOq0qfCSEqEBOfaU+OJu+Q82N9pcOwbPgICbMj9LGtuJgQ6u
FbGNxRfsmtKVeovPTh7YWvHMkWN6VpqgdHnEyqLgHF2RaNyWxLhkUn0uMXyzbBYL
DsywKf6CGP/emtO3HmyE7aSxYxNEwK/kJvZjuMnKlnhu8S+9HZIocgD2NP7RqD+7
tBrqtF49/h5rENBM8TMfIsDK7rAmbv7fgFrb7UT8lJu6Zx8P1MGhlch2zsmb7gQP
e8D5s+dOfGmOzoKUIPcpkhAc1HDydbCi2hq1Jz7rJi4X8/x2ED76WhIxdVK1TImI
qAEsp21dLchDXoG7uPST+M82KtYn1BUbhw2NP/iXiub1RWWm/IT52lbN3B6nJvf4
lZGRdv+9Gcd1nrf+yuqbKBxyGuwoUq1HrWyZN++7yQvHCAtmdthjENZGcxyo1FHR
fnRwL6TNFanfUgXbJ1V/6MAOFvXGDmUzEySuFVVWJN+ml1T/f1X1yrPSsjUVtLsp
7H/tydXE33OpvkJXrceRUU3yFSYSitxxSQg21UI6uMVRHB02QvpskH7MH2qCMfeA
I49o+dYJtTkcs3WvcH14BpMqxq89NjiiwgOmTqlPzJKSxMWg+zC+UEM7a51ajVpW
RrjaihKxv8wS+gyCQ4PQJzh62+Akd5CS5TfaDbhDkvMx+5b+tQs8fNMOB7Sn1/l/
fzdZ1LYZ47964JM8L+rVZx1oO9Ecs16ouQ6EGvZvzFJ8hZtY+Zhbmi5v3hPT39EH
4a53nU1SK88RlbX55tyJkfKlD3dAbb6dfzRfkmZ7cIugmOBsvGoh2/DbqnSM3b1s
k/N3jUZLm1d8IY2YNz0xuoImr6kImddQoX+PvhVFPf+rz7qa+FTKAq8mL37tYUPx
be6k0XXB7EBVWSz1WvCdHbUgOxxgm+0TMJI0cjvfBuhwxFKxsVCDRXolLOV2YvNj
BjjZ/kFy0IVqFDOJWsk9lGI7Z6HtzY9fQJBBlQ1HrWnmQWdVB8e2QyXUR4zN8p/+
PEWwn5KcTmGIkiIRdGbLtPD0Trqe51nqluPhteF2HK46BvAgDMOchVY6dIetKZsI
jCLMHSr/okRy9StUmp505P2zta+t9fh0hUg6P+Fs9dpcL3LbVdX0Jc+VlGQEg27j
W/4B2/Wj3uLcJhSngHV76KW5pC7prrNz4UyZhsq3TaHbKgZMAugmWTvWKJXocd+b
3j6HJinLz0CuRcPXRNScetmU+QjAYdGp/7xkZ4S8qCIq9zvAb9rq2b1JgZEvhkCK
QiPkKvkEuvd2lLP5h0EGJoc1LQrcITgI8ZagrLJ1+5QF/wT+kK09fTqen4AgDXCC
ocOne9GL7vCJb3Ejm72ss++vPCX4DylMQGIzF77DKzHWb0OR6yMb5qlWJgI8YTpS
18UAithwx+qU3MKqANw94n5V7vewEfX2G2DbwMMSIoc8pHrWKBWzLRwwrMN2V6Nq
gYH8xrnzF06yOcmJKB91wMXPVxh9CDfh4DZlOFa/tb6MaMRG0xPhyQzRTqAuL3uN
qrcjf1g5/+yOIst05nPFp1o/cJ2YZnBCvGwb2zLritPa8C8sYltoJfSQN1UkXAlg
nNE8si32va0tf9ieJsk5LAq5R5EcPkzjzCwDcOJGIcIX2z3vdfw8OyC6/Ku5mTBz
wb4kQgolkpEoKJ7HN+X1X4bTQXXAGXt1aTQpqPDDp3++Ob9zrZSBfInvfL1dl5O7
UylH2Kak6WKLBclcXhrLPalLlXVOf7Vu34RUdr2f6fR24jO5RpOlFab0Hzbi8ypm
rpcp/bsSk/GE2/+kaBzk046D6NrwmwEa8KW13POYTyeyNjvpXyezcn9L3icnZh7c
t7rez3sa5dPdaroRAhqeyH+kxNwtf7YgK4wl4iRsuSG5E0GxCdSLNywNhE35fJcr
wCWXsY0grR4LMI7jBRB7CtBU/zEzf9ZaHpQP+mE1TDEAe92O+MUIyGLfblmSnzgW
BJF49SrXRt9S90gmF7nPDU3DWfFRZiHHY265jeiqKzSuCbA5OeUy9lPMe2XCNuLS
0EWs3WE4ywatZfIhODgt/jDHSSOsJHrMsiyfyX8NerJJyNSwBb0N4wA+E8EeKKNs
53SWtasRjfZ4T1sJ/xJl6BIrwY8zNopQOMl5jGTTlGJIFR5hJcHbXvFE8XHWLAqH
hJ4ruyQfWyecKtVMoa+23Fs4ovGxtbKZYR3IIBaQmJMJ/WDKMb8QT+xsY2R7ccDP
g4U6VvpTX/y5TIu34vV0Mw0kBIUPcXgQ6EsriGWgDhgDVvPB68Li6tElaBgit+yH
s+oYBOR9/O6IxuihtYpHZECOpHEaCAKPBw741h3hei5eCIghoDDSYpnWc4fVbMrT
cv5FZFSC6Cz+O9bGree2HgIADOmVPAbZfvngVuAViYRoub/lFEQMBvqg+N9OMIC8
QTXp0GoNSgvOqdiBQxg9lAOhJt69FOJdTB4xxcuPag4JBeP2qLE3Ky0O1S+hU9YI
1BnyYzVQvmMS3OfClUfOg8QmLP6RgX0A5Eg4/bHldxay6w5KoLYBx9Q2f2brnSg1
ZsZf3fE9gBYd1TaKjbYfAQbc5O5ibXRvh52HHBCbOABiHEVTUvVGKt7UyF0sCEXe
5f90nWujXO4KwGz0vpSe253m0m+A3Ir4RxjCOjI4+onL0RIcuXUuHWPd5Za7x+/k
s/aJf1zvfnVN84yxlnBeEx7lEtkOUpR03J7Pl1YvA1v2EJce8uoa45C/YD+CQ62s
iSVp1y2qy7rsIdx8xiZaaq7NCRHcrXWoOVdTpAMWEITswx0gwlBUwO3yQYWwWwFv
xoOO/xl8ZE91WYznehRD/21O4269LQ4IMXrIUJSlJmJwIdJVWt1DxODt5jXUgkZa
m66+dAeo7rOlCZzeJ7NGbc3lihwvX64ZzsggUzkksch7MTvJY2RXAjad/hBK1pdH
5GReodLjRoD8Axk5qKCzO0zvBRUkfQ8ObbAx1fSrTp5je4bF/RayY27aiVpRyyq/
ww2gQ9GJEwOItCVxuViXZLXxk80Pxpkhkck0m9ORhdVj44erg2EjVRK9gAEsE/zc
XXjvziEHxudZl2029XM2p1xo9u+vpZpsiKCz0bGB1U6IQcNyqJJqIb7Xjnf3EbSV
wkldy58ZHqXMbqmyaioL2H2rgZ5yBEfftJ6tpSWllg5b3jPPbWvEHUXHCAR+IySK
MMU0utUK26yVEMqAg2iPsGZUUbEk2GSkZWQLN5KU6w/gAqSHKAZ45lc+/ETABdS6
g4tv8ZMBlciRI/CnUWVt3J3GDlN/VtZ9kzcU6UEIBML+hQvvlqIgFjCLPmw3OXrG
+nFYKPAbh9kPkHJ+OaxijUykV2X1WOCTfIgQ9MQDXj8YlgXL/s1a5TVEIHSnHPm1
p7QxNU6N7D52XCJLoJcPNCxZXRan1+LNbFT623YZzIg4wQ9JTdjeN6y8zrESsahr
raCGC2/NUZfOPk/Ps3Vn2NZDoPm4aDNBRg9bsEu4TJ2PGVRookz3OB3zizQhzrr0
2P0IJdkm7DD0yVnroSFGBHubDDfUq9qqdtH3lAXZdDlVW+8noMN406HlpEt1s4Ya
NSXRyjfdE8t5s59zgTj0n+QwftZw8NJYWfeJRCoXOZcRa/WD7A7kJFK0FmaTZEBb
ugmNuUx2rPDbpRm0LbI1aWk5Dy5OSMiMZAFShHww0qteX5kHWduGFVXzytgiJeKP
TiYaYadrH+MpwIu3GKIHqBWwMf+EpDDKcmwtCRcuA8Ktv+8CG1ggUs4NYYC58Avi
KJQA0lVxCJO4x9Xg4KptnOoD27HqvW4k8IEqtkna5229X6UdI0daHHSnlO23yDhY
8oK3JNXngbpLNLO6Jq7DX4qf28/JHtEnHl7247gmLixIHXrZ1UCnd6WmGeSzLJ69
LfCeB1nOsp46qHO4qWqEm/nuo/RoVaOKuqXC2EZNyMzjm20BBHp7GZqBwoWzJmUk
cx3qjudIyGP8IGGNgHcp2hMvoq4rD9vPT+GWzQ65Hdd8Czb2MCfqu70Lnc12kzsl
jVl7mBx76HLAXq2qboKpOI1Oae5WABmoEuF58sfGw9VsSrsH1DES7h53+WYvM4ua
A8t3p4sms0kHFOcdrJ4v1Il8/9uQ3KoNMOSeaVjADUxO4baoQLj3b024nWvDV115
7DMTr1f59/U2DQlinjuQcvKIwQ71WQv/yCmLfU8oENRaoN4z9h43iHEP2R6W67Xw
Ibowd7t7jpfaByMyR9KtLqhWoxFDmSgIyuHcuY8dBMy0/TCDiMdNVyz+61U1rnOJ
7Y3NFJ2pzl79J/CSeyUlhogB/fl75NV7+susdQRDr663XlAajfXS5OSux1bf82kS
JJ1+l8KX/aKoRTF0SFCgdUGu4LuFFqw9/wB3O08Rg+/V3jXEbclhVAZjm+b7ahMO
63bU2ExbYzP+g32H8yv9/59t5Mkor0nJBuxD39aLfa453wXqgfOpLZPpQJM6aobZ
mPXlMm4d5OqyQEJRxomylikvJCT9gF7y96tITXlVpkMWJFJOHxNESnuLjnjbv6Ul
FQExbwZC9VF7gMFPRkhj7+G753VLGqvpKJqbzXZcDUvonAwP9F88gNoWr1D1HPPD
pdulfa/0IaZS7jexu/NFeO8q6d0gbCIl0DXFITyDE5hCJKU/n3d7ACA0Z3/L/oZY
cr8r41fKtW9mWO6Rc4LgRIDXJjO6Af6OQdAhSdqCvLwQrjR0Fp5YvZC5ia/5HqiR
eXIcWKN38gtPUYDVIKCE2QqzKZXdGrrvFETPzuXQ2lrY+gWTsO83LbyHJ9uioqJl
BTI/z4yG0eGlmh8VMN2gxvDQvZCGrz1/+S9WWo1jb4431UL3PjJe9piwrw/GvKMc
wE00Dp3edqseySA6Mj1p7GXpO5SO2KHZN3utrHl/j6LxlWZktLWakCuqJBwLjzaT
NyDHSfFvAWvxT9xpd3iGQisp/YxoEYutVKloafkttJzGQta2bqeEformgKyBe1//
DjU+H7/BCrVWtYp3ILK4WlK9rN/ICHCtWipbk/9yTyx+9UHmM3MuoALOALYMoy3v
bc+juVMxErceZh7fHixZOck0xvMFqWdPnmxe4hshOp7c/rx/W2ksv3LeESXe7S2H
D1wE4sLoCZxULK/4GyxlbGc+UauHd5LUU+hbvXCSYvknBDnVIryYRTOqoSGfq3hi
ksRuPDc+geDg4AfEYwOB7RhKiyKD8QDPLnU9FZTxf6x66OQoo/PZTZiQ/S1LAyqY
1KpdQU7RkGQwwSO+wJEJZVVrugblBtHSBVpltpJTAbgXS+/p+vdhNRhgwpU32dXF
nEYBvXoz3Li23eNQsBoedc1ZRDkXNofyjiBEzfgR/HK3/t87KQUOxv9aud1tOde2
o4qmXZ4MpVW/ZnebG4PLE2UU456QXE7i/H7h0m5WkeCNtrEv1rO/1qAI+zoSegGb
uK4lJwBeIMjOyDWduS2LeetxRRHj6e8zash6W1RMVb/hbFNs9tWERVITaYhuSdjS
Wg54q5Xi8LuDpS8fljQPbZzYjnLGjo6BMr65ceE3XCMBaT7e370lRG87YJgTYtV3
5igFERqUAYmStMjEgm0HqsIw0RLIvwArMatG2NjlbDo46AX4tMYpLfaCTBI4KNFW
3WWoT8CG6yrICwehjlwSqJzHkWOS5dZIdbAxyRbJ6/3kfpTdmC66kwUn0XbNs8XW
icDvphkvzVwBD3aNtckmP45AaKawVYD9zq6x8+UKgsxtJNs3JSomkjBxJG0eId3U
L7cpeAYAvwwVu5vRjbc7Er6kVqmALbJPzSGBNJdRzZpFPwimbCaCRubJGcTdCFNH
GUIkE0NZsyE57YIszr2PVId8x3qaBVhQHWZoM4rYcbJT7CxgCCteuTXRj7CH4FIK
ADEs74+78PzcPyKzLWcnwHd27EFIf7AGOfmcMVL9pAbaDOPqMX1oXX2y0D4SFaCX
cc18J6fyDlMPuoy9LRIAveILIURPKfb1gpSq72lB6sxWAxRIBh3QGZ84u1F0dlro
vr/BdbXIk11aKwYbNS2ZRWcvDB9bx6a4Ucyekat+dqSlkr+qvTGdwPR57aN3eKQA
QvpKXksX2ROSSVUKMQNcLxPOjU2/fS/xwsWNYc8F+2Zx9gmB2YiKCr2vu27Qxt7y
3+5k5gu8tgKGCfwq5sO/HtSkiWwUxZPcpwidCSSQfrufnzJLuahj2YrqbOXAxBAf
t7MhCOZHvuN/agi3BcpRT/CJsYM3/ZanU8caXM/uHKgzlnBOWbdAEAuPb+ya7VRJ
ICeStCwz1z1lMZOnkPBs5i6RBhYYcZGEvz+TPsS1rk+dSaAkzEJE90xINkRn7Z1y
XsWL1kIi4Ai1xT7BA/7O5atHqy6FfpwrfzIfK8jmStLIrvRhbj/ozrvFnK32Io0S
wj5kzB62S6xUM0KqwyPmKoLQdkld04CAoL588KhaJ69LsURUcw5/9zWgRPdHYuEG
USx8AID2GCxiK28RLfAorE9cNkqwtL95fBhqBLP+Zq55AqlDb3nknAQbkBagWwLa
BT2No0mFwn0U6L4felWW21nQnOuhXTHyHCFkPN6ddge0zzNQv/JmqykJG56RdaRI
8CLQ9zdw1Bmvc0VIgVBuwqjjVEBN7osVa6AWvvxWGtekdH0YoZig2jH6iavJ2CcD
4HQWpHiwAeueFpYqBptdIoGXA5creMPVmqPbLeDKh58QHaCGTbLmmTN8umkp+RrH
6CopZjbQyKa5DmIH6U83HjtQkP4jpi9uTBMUO2DKam92uFU9Nb+jBDwseoGrrW8r
G6RDbeyto9rTsd+TvXcH1OZ7ogjte04RTiAWOUrYQZXymOzZl84xUwIT2QpRgOfh
SU6dtnSxrqI5Uxt6wR60N2MHHrMVmcGtIyRO35v7vR0RVTd7xKN+QHpdVATxX0Es
4UFY159cwOGO26Mg6nywuR9E0QZ6yms7guRaPi7QiLm8RPde7LyJ4kGMPDolB+S3
U+30nQezPWidXRuVH80n5tfjdE6gZ7/uP8UQmENDnlft9vJyVKId0pc8Il/e6obb
EeD0IGi7B+k4RMmvUZ1yULvw6bGzmMLqR6wmDcz/EJsr432YIKRBgALLKzFByoo2
45n31nxDkyAwYDxCR5HO21dFBcQtL4XT2Em1KCzP2PBP/pxDMZDiJ8I8cHe40+Ig
GESvitmygsFZZWg7lAzoJoNxZmS8EEyodvtpFTa2VKqJh/1TWKunHUWtJ9mY0g9q
7FuMejWkx+KRTLbUFkpbhrPrnazeD+HLnuLWQau9064uFLGgGg5/on4Og/Ab53Ep
9e9Vt0xDAwO397eviyasNlkt6C4NR1EHzx4sCRJxhU2vhvOTt12Pd1Pu+5lKav+Z
pr/TJZi+NoiL4UADKw65hl6zGSrY6dwYPuJUvf91zE5SJY5iNEEeHsPtQuc/ocxe
miQfP1Z9kGy7DZAQJjT1GsUiLLlWfgLeaD/4LPJDdqBKNMGkGFnGEP1BcRcEo+cn
LaYSIiCDUMIebqPCu4b8XwPtQQ083pnanrino70cDuyozRWa8/lHsrDb7JXukUPp
PwwIdP542MSFCB+1KQdTUxMrqWnU/Dx+7Y1I6R22ve4AbGUBAzXS5t5Du047nIvH
q4yc/kOOeEu2VhAyXrXX1CPd8F3Fuc8SI9jLdXO0cM2jsqB3dcH/u6Pn5bSYjfEW
fwfpNkyYMMPdnuq0OOGXoEpPckgCCpGD9Alh9Jl517Y4mxifJet9z0dqheuY2In2
F8SJ3i2ryPhCWR0wrfq16ySVHeMRekQjgoJzarzrrNzrYGxJY+C2PTNHL2qHwrjk
pCpmw9LmFKiSNdG0Beb+MCHZyYdPtMhJvgLsNtSeaCjJov3XoZ0b1PmFymyeg5y0
ekBm4O3FEPEgP+WpmbbVAUHGxZwXhflsTjZXPRMVmiRTraA94mhiAIhyt9HUWddb
jDc9gyKNyo6/5eY/9CKNbY2J+9cZ4M1My0P6XAC6Fa8Uw8ZBlA+iea3yWlevo7WD
jfLSfqKaJEDFCHM7VAvU0jNorUbYJ7q+b3oZXDasO4kJLfbMbeVnhnzCIK/lTQDO
E0NGcxvEKVVfPkeMR9u1b0wQqCyk6oxMlYY1VOf7MiV1QrygO1CUBX4ZxkGQN1Mt
NTg12WLEz6EOxfGppeXNdSd3PTBuT/aS5zl0Nt8cAUSRhJ4XtJGThXeR8gd+N2iF
YR3/KEdWtdS61NwTlAh/tKb9XzWszYgOnUFBqxMhMyZmKXtj97GllfKmYTLWIxzV
GY9BWLDOdXtRBhvQ/tanFg91O/IYyAi5FGdZsBcaLP3JcSmnlOG4JnKAj/yBvhCY
/lcZo7x5DYyi4ZclvxaVPiPPRIT41bci83v8SeoZK5lBMELP5xh5x5iNOakc/R0V
OI7yWtXTZpc6muQJdfGvbldxQBSg8k1LkUw7BIGVUQltp2dcQPiuoaTmSxuK9Dtl
iOtxxprBLvYMFTek3EbswywvQfSFgWawGMKmqqjZXudZf8VfdWZ64nBCB0Ll1dJG
DVBBO3oOmcpzFtE9t2WycwJU2GpSSavJB0RcCxEuc1hjkDzElYUj6eKZ4fJsxo7I
U2vh498gNNj+O97CaVTvfOoKCDk453RN3lIMsrO8vsFODwTh1/xB4a10ZLx0PqMA
/ivUFSMPnatkTaBh7rSou7mMLZZzF+LCgAlEFhSSTadUp8tGlDLKace3WpRVVIpH
VToFVsazC/PbJxCVOk20gmm8Db3fjsYWot+0BkFPXTCl2md/YjdUdcHCBC5ZJaI2
vQjYolloIHNUGWvGXK6p5Hv+WTwDLHcjXnY3HGDqZD0IwQiE2oYlmUKgqk89Vfm7
GREfBnXaha069pRinqcTbQHkPMAWBOpMlozpCnCIDHt5tblhBX4T7Q1EyCHORYJu
C76eoF5wWK7oc/psw32JfXGzbMcxJU8IN2U2FMxjjPLPDBUs50CsSUaF3ppgdcuH
DIDmRiAkxSv4Gv6U1oWkxR8A+HI1bIrnwt1961Nw551WMlZzOnegnRA291CbSEgl
vkHqen84AdiH/wntQCLm8V5bhjF8hh2iB8zyqsiuJCvyl0WlXT6zk8ttj6+kQTWl
ZbW7SrZ1kHyLRFX5CbTsgTk+dAzUHBX5sTA35bTBkleLICm4+UaYthhAyTbB61Ss
m2lplytvc2NNd7/JzQP2MePLxgIEPIcPwTXUFeDhhVT111y+DqTcIxhtz794z07E
lmYF6Yaet745trXjtpDo3ENoQYjIvh4BNbKfYwCl1P7IvfiUz5H6Wis6lZCHRej7
bCCK5m/kOiFyrbbxVOn1CEfMrKm/+ce5N/V4kWerjC+pdOZAQOAZtP0yD/t6UWFd
dFOHLCOMTAwsQgu1haK/U6TMDnU5aE3EunQ4ajJQuxEFWXyEMWJzxLLlc2GDBUSW
JZe67XYePqyqZL7j6CsdpNV+NszgbH5dPH+u5afwtveGa0cAvjdTO//RYEIUHcFZ
KU24x9Hn5slYmXx4XfZ8l9NHKV+kPdeuunmzFjLipyi8AdMrFC8cms8127dk480C
wKEXFNSSh61reHK5BsssrbjVDuz4nA5t5w33qFxSe9CODlQ5CoylYhzH9bnkbedQ
0PhpTny6DRISQ4G96GDS+pMogHK2dnPKBMlXxYTjGJu3z9EINtYrfvVSLk9B8SGd
10vznDlc58eY3xNMdjj6qc1BJh14bBkVQLuIa/+L4NxZitxnRrQRDqdFZTkfSVGt
V/l5VLk+deomluZ5SO4dMEVza239MJwujYIQwdyh0j8ySxSQU4nkodtg73URhteg
8prheesH5iYAOFW5V7ionCvP5kSg5gzioD90wIvJaycgNqS3//jPBJ7blgJC2+bL
cswH4XQxc1Sih/ZTrmlV+PyjoJzMaWdKeDcQHHFSVQd3UqeLIAN9Sb7Y1mmXCJe1
LIZmrTNDj64C+qXcMqanYOkXC03wCLs3C/Dd/z4u2nhkaoBO/5PmK1N6jWkKS7yx
OcaXy1VwWqN7cipYoVLpNoznZegACcoKt4cJLQpLrn5vb/6nbhRpDhmP7fRj8GQd
scl1Oe0VVcrQoQVE1qJoJJNePkl7Im5EpVwI63l4V1XOSAnVSD3sbJWJvKHCvTVv
TGsIg7Va3y54ifeR+QxUgLcYWOJr21vxpjHrFijJ1HZcv7bUqC1VtYwvEIzvJ/IX
ESw/blbUOJgDPfgGMCEC0pI10dCNePSAOoKuLUEr5hH0j2ZTtlDb9XIydu8WyB56
kpdW3vU1s2D/9p4bkIJt0Q461GpJjHAPnM25ZlLmVRGWelSQlWig2qF/0XsMBeLS
Le9Cba/0fnUGxJsxMe7GM65KFaqMr1N24pk7j/batHQIQQQcMB1by7jJuTMofoN2
6aUPrPDXu/ro6lGukFlwpYvNfPQYhezKbt5pnruMwdpSiUhRhzFSNclCIfrU2+2s
cy3mPEndHK6cnECUIcvWR4GviimZp8nof3t2jfEo9ku/yi8qQ+QSCm55sisNKHnl
57v3K7Ksbg2iKnkxT65czcZ2gsDLBdaT9TVEuD0OdeVRMJnMulS5z4YZ59e0aIEo
P9LTYBKJrPPhGzFKHEiNp7Hg38NwOZesQgBVRjLjXXPB03THrvyENivQqzOALXjk
jem9EY8H/6/t57GboA3hHQ9Ti0l3EevBlwHNqi68KtZhzymloigST4vH9J1skkNX
lENbBt4+o4LQgHs7KhfehxhY2NMFI0AFtZpwjzCMhnFQtODvYCDf2QDufOlbWXzJ
5/vuRc3Y4MwAZNVTbxnZqe7DrU/0IGLu3gywbLJIO56jqrOCWsKbHhQBs8XTu+wQ
grKX0X7pEIgef6FenqoZyLeoKMQygUj7sLnAqi5kPXizYJbXqvIkABPJdhJZnq8Z
xmCthHPdMBsW0A6nQL7BE0AcakN82lt6qMqFUyoD16mqFEGw4HsxcYJHgOFcV7jG
YoxylSPeMvpGJW0fpNWVb0ZSqHGPySqtHHEX7dPWLrgzMtpvoPIJ/QuUWhUFkZJf
w2Q5bZtVohl+UM/TogD6U7bUo/agWp+OtpTKPvtfMgbPGbWP32DMq9WCMUCGwo/h
9NQyoMDL9mdh0rL8l96H8J3evjFTTVGGBQ23b7tBtnub++rGXkC8+kURQ4BBCwl5
/1FjIjCJEJhZ+d2xGk5Cg1SD31uYDkSxPxKDOT6XUrZiHmy8jQ6BaLk2M2o0xcpn
QUlsvVM40B/yei8Qlg0r95G+U3nR3ab3FlQ9xWwFaTLWmqX6sjMxs68HPo4IxCBq
Uz8tAr+DksKYho+1kOBljlG68qikC0fO6BU7PEuzrzO8Osf2D/Efd8aGwEdruxsw
83XuBke+Zw8A0WL0LQpIVESHgujcBfqUd3sD9QqCrnikAR9bAA19BkWHVqva5GHF
xF4p9Zzcva7RsluGkI8S/d92ajjtq11QWzww1TNg33EdIi21K+fhTOdawtBOzC4/
D9jUzW4h5cvZYAqWp9dLvmp4YCo8JbGhhKkE1UJsVCXuBBH8w/4E7G40Abf3yT8E
rRhMFq08mIZkOls44KPnKyo9ox7T7d6eIRDYAkuGW+5XSHBn4NF/iglxWwszdqyy
IfGVg9S+6UD+JCgW5Kf1wxmnJw/P/SDpy7sprb+R7uIE6JTdRsCGE16BvMPO+Kog
NXfkThJ0J1SGNJFKSdU4o/iLhLHQ615V/RSaWOry9P85rs3eFftkDeSPGMbRVsgS
T/sBVPVFKn5eutOnIJhH9HMsTwZLBE4fTqFNpKfp+2dWzDoH13ODkMBIsCYIkpic
vRga17lfvBxJPwjPpojjnS8CaNp9XZYuxAJkppX2aaEIWmPbw2SWW3CdfVSbKWOr
c1vnhqeh4nsC3H9o4cj1Xs0+LnvdFyLBISqPFkjqEbPbf0DzI8SZ3qQZar+qircK
SA6ihseu4AMhUuP7ZahmxJF4JVEWnkh2a8ngeTe12LITSjeD+sUyHQUaSSqfmeUM
cR+K6hOgVYH5b48bSXZFqetAtq5qwAA7VYWQSTNWKIJwdolFHquRZW1KJJ6SoMx7
YprBPrd04xMxfjO/cB6T4rrIEMevrDe5JQM+VIUmTxmKIVziSeojodBDeXsT0jic
lADGwTWRKAN9oZ3oDZrdF+gQmUQKSHTXkuiJhsgxv6iteg4uMm5isvy3PPORr1Lk
sYq2Pwd0o3gLB1U2vKN7WmOEKr0rQK+uCib7ysCD/vHbflPmO9656lh+blO3NzD2
BmXwFOACdp4JZ68j4uit1kVKmNqAepm/KzHF62sQAOoPd/3Le2yhVCVVgvo6r5M0
F5ER12dlCh4b1GKc8OY8N8yrc2wlkW2r6xOayM/m95FHFjUzR7mImrMxdMvPIDI/
ilGfSbFy1wrlHO23sSeBFH/AIoarBlkYF+oR97mwhvKZBtNg2oNt8V1Vt8MK8i24
ps6zS7EZTqQIllxI+hkGmzcp4Af2rK7FncJe/pDgpvJGcsaa1jkj9DHKP0rQTf+C
UWpaDBYToFvb26uAX+WuWDIWUTA/0FgJdfcEozKProDZjjh/ZnEnWKPs4jNvW/vm
zK54WGOf88zYj7y2pa3KiA0QzIDmR16+QUUZgm8ewJXJUUPK0/zRlvlwcj31yXEP
fkT/sAMUvvOUBXV1XXCFXzTPtUYoVtQWuNZAzty0/HhB+BfJIxQg3m0b8S+n4cgH
+tH5p1TnclzluJtbRljb7zouzEcUuzf4XJG2yYwj1SD/Vr43w5w4ngJYx+n17FUt
ZAbGVbb1vzr9qgq0SOoym6pvOwQcE9/KFB8v+PqejweppVix086hY7iUwd8HQ9wl
09QWJ6HI901xfZJP4rQH6MPLO8K2IR6m1dEM8HooVb3Ve8VXqFdM+njwEDzfVsOC
qpKsmlk9jIxn3dtvxiiHxucMPt0sLrrvHrFzygzstpt3E3ZDBfPZO5qyBac+FD8Q
DA8wTVJ7sNG55v8TcBbLyW+3mxXFjVMgdTTRO5UYyMfWkXnNpxS0SQNOaXFoEHdz
eFU5byw71K8STjZXsRd6GxyHx8jW5OTmDcapT7rCUdPjFo+lAW5fOQDGr7WGlYq6
Fmk44TU0LxSe/LCrnjUm5PiwX5WWyPeLHesSaQ06tGL2yLylkQwkRpcr7tYWNhBa
XU4RPGNcVUlM/wJWWBv5lS9099P5RLYGMfEsn6hulSn52sNTM7dmwGM0mr18dNY/
KgGeRg2Q8tE23lSyKmXT8pSY41UO1phfiqdgWIs7VCvHnkvD2ukJBC8DIhmvfJvq
/4ND9OueMx4GCtix28OucT4ThwPqCwIdqYU3DsIBFor9loNhOI/VF3VUBH4AJ9gL
4V+TszAKHB32c/QMw0BiVzwcmJd4+rGETw1AbG3hhvQQJaYRkhq1G+XMBvj+xYfl
/Xr1CNV7a1iOjfgmSj1rjAspUSDKAGDKgCA0juD1HtAvUzS80ngA40NkIYNvTb3Z
B1e27THf1PKSLlTTFOwKWg+gZ5vK9j3aOc0ZY1N+3mposevwh+vjQs0yHACMlUD0
nnI+m77gOMg4dwKbueJlQ/vv90KorxuL+hfdPFVvlHFXb308ugLSW3OQ9Ct8VIAI
i4Az16ePvftjh7bZmQTi+mB6ivBGYfD7o27k3t7AcdRinFdKWI7xMqsqhw4uzQEE
1921An2wJBAQqn39oDVv2KQsV9yffVgBI6mjihM7G0xSjay364V/9j/tzhHAaqbU
aoK6/YNqCMvvS5A4eVR5YMDmVFNAGHrQtXI3rdgGTngglC+zD+sSdrnggsZSPrrD
G2IDJxZJBtUtMMog28cC0nPjeFImlnLqJrLEIVPeLuvgqQ3VymDQTegRxyDSYpvW
Jecfo59taXnr/EtEQbuT9vh6REP0NaC7MU4rPB3c5GAhkdlCe1TWCcfmVSvo0B/H
9w9IcdE45ewD3hrKQoqQ50uCf04n961HsDdEl6zxhtHTEWHY7ioPKKwSj5gzqhmX
9VKDqUMWe+oFVkC/pDXwaeGxJbZe+njijfhJVLsNG++4k99J72h7glx4XI/L+ohA
5FgV03vUAjfixqDWj9ZNiuJPFPCkOl+b7WwxGG3bm9YrHqFNBy2FcZNNBCRIGcCT
+950Yr/exhB62CBvEiXb+II1/PUniWRc29eGTsnJc64KejC6b5NupKAIpk1GzCwA
1rzCdPi5MyRcrN82OMwWSK7RBa/uxMI63Gtl+y3bn4iYzD/nVYnYdE8kkp2RsyTZ
xwrEeoatiHQnfq0lY04e/4l8Qq/o+Q3Bz5OfqnJTqMHylTzbOlvak5mnrM9DES6v
a9NFeWPfk2AknokBJJdzCYmaWlf4ZaXI46yLLpnv8hFUcrjLCFOIXYbehZ/6v5ae
ovcNTBborXhaBY2Nd3cEEAeOJtahhcLhdTkAZFBhW+q/Qrp0kenjmNkr9gTpcWlC
MhiiuEHptELpOgO3j7M0k8yBFFtlPPBV6an4Nm0ikSOjpmVynWdb8/aB1hrpS9cB
gJkzfpqL4QNHw0IjdT21Or4LVlZeNTMKSkSCYQhI2YyoI61EcYaB16QZigAboABt
r9b/ONZ3VSkUzWEjdBAtTC8jhWqAv7++MqoPo9ygSAp7ScAR/NIEufJSDMURYR2n
y+mtHzNek1sXknspyXK9ORoL8Hu9ODmBzfTAHwKpME0MfXUxrTt7xp096VhS22fr
sB3FGFNYF2r1k4uCs192KhO5CrA5/Kln8ODeX1zFN0sPAHH8iYW2l+0R9Igh3j0t
GrAcu5XJ0RfIs3si5lMsRYD/5eNGzFJpG9PiAxBxqrnvxm1ZQ4yJZmZmQIq8JApO
RQIG2uUml2TyuKjwYOdg/3IIir6JZIybWqcBiTyQf5djJOAcx9EujdD4b/rc5xEk
1bUE1U0C4OX3+BFClyEuZqgjJ4Hjo4+llfzHitomSOHPbw3LgZK75f7VtT7v2cEE
or2DPvqdtWMYuboNSr9n6Tjfk3vQSYgeP3QaM+GkX3RfGO6m0IFRu7KLQlXJVtfU
jDMrq5jg6Zc5yGv4AwdB/ki4vmf4U7XRZQc9pQmkbntYReNgP/qwz6prixadcimx
o8mvTMIvYobxn17N3h7JeAGFlHE71p8UJ1mar/l2A/aOdoMCx5RFjrHv+bALH8xt
RWtLS9Cav2bC9fwt2dUne0Yb7WRGTPaZI79V3Q2ysV1knFs+lAkiqyej1tE3ZtJc
7VtLOeW0Jet0oHcRGsKtbAu54SgQb7VtianD8+4Kkph6IUcAJmge7ukha4rZPUvT
tWecZovHDmh0ymHdOynBH7KnboYJ5Lpg8xRzbg9ANrUuq9Yt0WQtPr65kJU2KOe5
Eaio6roVZdowu+WjpBkPg5omsDT02SrK70aLzkOtKfctiYPEOrD38TfeUTVZ580C
EZYmXMQYbRG4bUEuuJ803lmjtTdhqrQuV5aGsOVs9PFOfj9CUr7F3g2wIfwZ4qgv
IKTAo2tzYzlIC8kZck/mOuBRLn1dlcy9nUT6r2M/EEH081Cnek9FWA31JqhpA9Xe
S+UZYqUCYxhnh654Dv+cTKPnHGL4SWAk0TV1/qgOiyNTfyGQy07ipZXzE2zmqANx
o4uK8jvS8GoxSRg99vPYlkMVEKqSa91QmkPk72BT98BwKpW+m6rUOrHqEM1pXBH8
1N2mWgZpU6GIbTeS1nhIL+1JN76rrQRJvN6jSJugh0qFfI2LimCBp4wGTPL3redR
jng+NO/lH+noz4VayUMvLiptIKQH8bZwvuG9G00ecIPtN90RX5i2cQ4pjKqsp6Pt
ewh/ko1/13v2Ub+oUXTuxFEBL4pBYJom1DQ/VJgDgX1npOAssPaw8TuBlMRuRgJb
9NxoouO4Ey8/eD1Kt8WraGw3Y4w0rQMW0c6312zbmnMCItx7qOtcH7Gx7OrP0Vbk
pcqK7pyKSw3JfB34Oor0+W+MbgDeRR5tfDCsmgLzw35GyN0rwGKy9SBiuhAmMbIz
qavV6d4vrnB2bB42R6XajIw6bR07C9tBypi7aciebRVtFeJHoiPiIYJ/qwu6vLbI
pJmI0igxNvn6KYQ47KIRw+dnv5eFBkxztRAYoIn1JVQTVb3IaDEt1Bp2uKEhvM4h
DAgmRB0nMXHFleehIhNhKGtjAlGDQwru187rzMjDTyCmhgB4WKz2Z11nufd76m3S
7dw44c9WNd5mmfxiFRH7LzfemwlTuk6OIosroizkixhNRlbcaJfo4eCqx6zxarST
4fCshHsOcGGYALj1nNRD5fF7lZ8uvJjYjtZBW+OIGFY997tMeF+vbkOF1istqO9i
yKB5gpYlMKxczWV9J+frAZuqgfVFt0zTZouc4VNjFTvk+SUTysNdgWRbsDrjJjpQ
meqLAoKckvpPU4Km+L8RNiv95Y33tGo3aWRW187zVUAFSdhWIJQ/tsyJz52TM02E
tydeZzn2FOGKxja+iPJCxTno4Vb9IVuA5ukdSahyE0/V9uuJ1niyy3XQ1kt1H1HR
+l8pvN4AuqlyKCIPdSwZjUJV2gjX2hAdV45ehvjvQSke6WZRLIaxNppGxfSguRSE
WKCn451+IfIzaVdFqLcSPf5YxNVa08gXLSMtleMT37jM/rrPdl5kRatxqHLpgGl/
fMZuU7r2UECm7Vgnkm0fyqfeqYHOlNhF88Infxjwl0SeZdnFM0hPx4uTpf3PGn8s
CkHAdKAntKVIF4hJIz+AzQ/Wwt5P7bZniSH70bf+ADKg1LG8ODfT/ArABHQtCS/k
rKMmYr0UnLOCqdmYh9TlLJEHGS4oJc6XIw3PkmGEewhDgvciaw2iMDfWK44ARXv3
sy28KQ3rQ7ldAhAwmWDHy8mR9guh/Uuuu+K3obgdeXpSESnkUSSVcmb6pw4hibLk
UnCqOFZzbMEHrSx4cbpsQftjJSt1axI1y9Uv404XsmXuR8diwsqSe6bbCfS/Q/ZY
EXe/6G9yR/RaSZBypRf9n5xNSAp9jVdrMdrzpLK/xycWr2w6qKQk8CNvK/89IJt6
EzseLf7PFqqLGpumUlY2L0GWQNMb9D+WcMB3RXBjJBbm6p16mzrtib6uJSj1RCtO
musiiqell6Hb+ybN+4CikSq2yn7O5jSrPNBnYo6YXqahVxB/hMvur5V5/kjNVR6q
4zXSeAUNdJlkywNAnUVCqY6BSp5AEHbL0KMd2HmtL0VcqNb+BcF+f+bmVPcqojcb
Z+WdxWgJxGuYYLCuPjFN/oWEYvOMT5XeKDuEOnPOKhSpKEGUW/os6KG99IaQL/iY
Mab5NZka7k54VgBH9TNctGTPoS3G8Siik3M3BaCFuRWSf6qc7zNewWX2CwQ/ZYKu
VokJizc1u2Kc+9CuZHFl6mH5L+ndtP9sn5wAJn/kw1LcL37gkcoV/+z7fLKPkyDZ
w40Ky/+HSdZ/9oKCbqUD8ho0RoIU+XdGz+y8fQOpL3SIl3dDhRkdy2UQAkbbqqiQ
NyO0VFH8LwyzU9+361qUmKIPim3vvbJTSTEWb+I9gkvRGJ/BuT5tldpfo8GEWQMT
3Lqa+BJLH52cvHqIdHEKEqsCrvD1lrivAx1pN60kg4aFbpR2TMmE9mRhUxrcZx6o
ke5ob4wV3g/h+J/vL90yjlPZqsi+5qdte4N4LNyFo4dd+kFsLWds3lLavGPizbh3
vJN6SORFLFOftyHFz5Y5gfx+0Z08l37gwxR716RtLXlFQQojNws96LnPZxAEa8ko
12JsiZ5HfIKJ8+kG1h0Xuu9O+Nfex7JkvfTq6xtpsojJ+/cjv12iYTpUk56RbAgt
r2fQMihClh/pg7o8BcSuhsFq2fGPMI6qTdN+5R5kNu0Yan/QON3lOx7W4Ycr99GB
zdc3/rrjrA420DVNuZnuJY3ol+jrpJH7hpN59Q3Qtoj1gi5AIKTQMHyZ3TvKM18j
iqg6M9p373TsJ1GthGnuN1/YN1wUe/8msRHgDCN0KDyKprYx2Fa0Aarw7lxa1rq7
UIdVqzbk/Sp008kSbtywhi0vTzqui0pscB91Vau4sDsmiyeyk1ZWLtlrbBFkkYIx
hA1Aw6W8+zNKrSrI+kA23CQ+Ie29lOFCaqr1XOEVVuFkyOFY4nA6LqbT/+Vb3ZvT
7gILrbLliiy7Sa72xBi3NZ6YFMxsArToqfSS7wG58YOxXdxc1g9njZ3lB3XEFCD7
RIqzcOwrZ3WkqvtndeEaCK4zRtmL4DWaPPuuuI5ad7hoF2DrL5qUlAmnNCRTcwzb
CTQ3d/N/ly2Hyvw/mDMMwqd0hQZsRBtTmNk0JBsRXSj9qjpCFr8vsNj0eQJbo7g4
MArNGe2wtlzsgzg5NwZ/Arzyg7+rPr7WgelPBYARmHJrHiXG+zdEH3DsANnvmVbN
g2GqIG6PKdcNpDO2KjVfWzVmTnWPavl/H7rFh2tPSjUO2L44wrakpS2dZvUeyJW4
T4hnuUIRm0Gg4JSkd6naZpEF7W5eb8WdSfvNwoG3Bg6n6nmSEcGCxZT+2Xztiwko
jORRgANq1ptY+a8wKzW0hHTYcWUlfSJGtMJoCpHSQUNp3JaJ04MNNR7Nc39+8if7
GfK1kATDUevPGcTRyUG8ORL1b1TAoUZEhLj5/AxUNYW+yirqXcAfTsgcrf7pW3rP
8TdwqSqKOhfwRrkIyDMSQ4uouCUzyudxWXgbvMLYPWDsca3OgDEo5ICmotBGMwUL
wzr83zGBAG8OYUsHBOYyl50HRXmk/1IM57WvWOKGWGkQKDvBV5GlvWe8Mh9U96l1
XZgTZL7IKfL4L7dpUg+EKUrabH13Z8XON0o/XPTbT82/b3JXvNhOY90gw8c+SUTM
Nnu0mzMvdeSo2311TkWUF7yw2hiRJXl7wrHKlffn4sc/6wGZRdcnO8bkdEM0dkDF
1hqXaper+qKVO/m5GcGNymr2zcPQ4sX8nJDp0x2MYddBzO5pZTZNFHkLRWjmGh4B
ZM0lo2k/ckaQqRXFTnD22NemwHXBe6A5zYWmHY3TfJ5gqbyUWbWbVl5qmjm2UDMg
Sw/CNzb8HKBzyW96BgeuueMlpYVsrPNaoIq8VGCXt+WI3HDxfgjlb8afr6kQhAA6
0enwMVxN8+Mrm/GEqklqsIdGtUUe/ykzdBT+5x/8vZPfEVYoZJ2wmyF7ieSgGr/N
1nCcLp/Q6VGzhg9GHyxG6ygl9OJh6DTxpj/Sosc6MfK2mGH5x+84X03aRmh27GJ/
JOFk3jf5d5D3fROVROazIGdVrycA5G9YkDKE9VYQtsxsJ6pvOjNco4GM1dMEKHw9
Hb74EvU9aBqu5UuFLrnOGJ0tf6fSsC0TVQWZLoSnBNB11NFqOhkCtzNFzmFkQnNT
fhA9vUQkFop/60H9GWQQHmMrXKkI1jziZokSn1n5fADowyKSFax856zlYhadL0jo
kbruFWGxYUCvJim4gIUTK8aO41UXkVa3sc4ogzh9MnuTtjZafQ0LutPBnbnKMx2t
WLi0sCoi/UT8tfScdM549eZ7MjEkyB1Raqf2Oue9XVD8gA6vS0y2/A1B1witxNgf
nazyfm69JKjBPhs9+vWF8O/iBa34BqX1r/tbwOOZT8YceOnm71ZLDT+IXybCQSlD
7ECcCPvLb3GFbQdBtcOA5dBI/fgphBVhJgJAtkg80ZUGsLjZ2lwcJtDN+p0t7CbI
SbDdq4dvsuVsm8MMyubZ8JihAA5MzCYGpeaauFFkQxOKZ3T6SC5pIdTyr2p+iSYt
PmPTr7h6oGyI7VI/c7N3dwB5zKcHaRgnQDiZXOTes8NJsuy4CU1hClJ5SjI8p9zU
bwfTrxJ6mVQnMhZV6g8hk0C2ZzwCX71aPan+fOcK+9Ocs4Ktet0UvBal3OiUUaOM
QQ6V/+sYaEsQodneb799SNIw0TvuVaHxWR0xlL0nWSuok+R57wcNcKs7N1ee+/xJ
sUYawXXtlajdZDADw4XZ2WChRUr6A0+5RC3xCHLegU3pw2aUHDrR+DqHx2EW0Pd+
yRNOF1KeQAnSaC8kFWs48YN4vum8bPbwTwbzfQfmlP4sS0TALnFfJhSLJxRcjSRJ
cPy9fuUmPuE0N2gncOiGRubKr+zI9vqpqsotFCmOEO7CdGL3bfYMa9IIsFhY/Eth
fhdmg2Z8psTLZJGRlFdFYCvQmxlovhLAeRBrY13yywFgAyqTxF1BCNLuaowsDlgQ
pCJiEh5fEUwaXXQg2Ey9cTquhtacCwh1EdeTxNPxxHN2A4UgO5tUMnuDyy0ucEIT
eNECmUqpMrjr+viy8Ug4YukKJ4p42ePbyUAvlYkSFpbJxO3g7evKYu71ZWdp66jw
3JxlEWfS3pgarsyehMlba8RbnCi2AE5hP2Yzs78mhiARCQMM3iOkH0BhUm7Wf3UJ
wEvmxDmwHBPfTdYU0uSbFpLR4CO6eXSS3AN3f++hJWV5cyFi70WW7KLKETzcZc0r
iV5MLRiS0aVgAAJZ1GpMHzaFsWZBCNmj966N62ftmF2H38K69h3pQSPQ40CSwr2M
E4eyVAcEZLIDcL1VeW8+Zz/rdiSNsJit9VzOxv5EmpXTpa3nA6ALU3f/gGjdR6W2
V86nDWs+/o6z+znzaQx+AeiiFTZTL/c/e7U7uEJbAVAJqzzvi3JHxWCXTe5TViJU
GDuwJHgfgv99i5sf8+eVbzXEoSo2uGhYoHqQX9M2Qso9PdeGC01DoY0QatLdM3N1
GhtQnF0od0T23uNBk6XbNQiROfIa3fx743q+4UtxcFMAsw6wzeoejsrVWDQH9Lnf
EYndiUFF6/stP1CSHavv/2X/IIVhQ8i+5qaKCtctxo5EHvBYYtKJ2ZlG1Zm5a3Sz
QC5si/cNHouHCepaD4DvhVVj8DcQfRGR304fmf2t+6VlpmmuIaX7j7ISfi/hFv4R
EOVGo5vVuUWK7OcdW8xm3IH6g1SY9/xtRe4xVtZSw5nJp1Kn8Wi7IlQkN4EbZO+5
0JU0BoJkCF1fvbhvOdNz8dNrZOWOCcdfr/u0cFc8pvJVLG5EKWktIjkXXml6vIBn
HnMs5ojvV0yC3CqCPEmh+JTJG4hLhnVNqHAIxAu50i2cO06e9qxRrGZZE/6UTxix
aId/0fSog60UBZbG01oD9qcX9KX96UXjhuFrf97o1gA8oJPT1wMyYaRVxUr+8GVs
urb95PWnMwL4A+SVYRT103R2SDcrJ2F9a7sfklBTlWlkD0SoAdSncf+xIRGN++RV
O64JDCAHTfIqu8owcv1RnBtKzAxr40ptUTG9nl0QzwQ0I/ja7ALcVKBq14JlY8ti
NEz4tvRdiogFe9KOIWhMjlC5v/ddHTP/BnZKtMX+bWi+a7XdX/Xf/oSEKy3HSPHP
ztifKtxLFLQj8Ub6oW+SMWDanCCqV5W5pebIAStNz2a0RTDcQ9aF2j9VYmrPGaDI
FjkWkT1jkvixb4VfLMc/GlpDJXaOyL4ZV4ufkackC3SkOl7pg2sdwzcPDBavNbpB
9iO6HwLyGPmxQN9b7X0XITel/Wcb1NtMQ74YSLQf6yvJPjdBQqIgrxALbxPaBQWf
UJ0BUWkQ4rHuk4OcYLX5CdDfoIYt8i8Ptf/LLm3A+huuASifvicKAXR4jGfvW4PP
zjwqlIlygFhjOiDupJfNuEs8bp3gSMuCwP3wYfzHYTP6ZQHen9Zmj5D0jiDv459e
yeKndqUIAyOKuUYGEgs5Xjgum21HqN3wm21QRhqrVi3hTMgRQxnMoJyQf6548DSS
hyxz2ZPp70OSWPPDYyVf53EDdDBDAh9rUq/eeeGa3CBwF+XhOjsD8+DFoglBITx3
u+T+//uCKkrIkvmKHVHejXvHsLMaRsehY259SFqMgs1JHQg0Ilnoy7FNYPMuZGQ/
h1l4kPzL6jZ7Zln3Mc8M7sGvb0DnnQ0zWBQkToWa4lAop0Dt4+lqkcX0iRnmtMAd
llT7Ti/nWxqVRj1PTd1AoJ7EWVotZpKeXA6Bu0y4xOyBK/ZX2x6fhLnFY/Y3KJZc
DINCt5uncz+o9GrnywQHpeSwV+RFkX36lG6u9RSSIlYyobMlO1fspOWel19rjgys
9WCiIuyJgZfWNbWgm5DVO6TKG7wh3trEcNREoHM0FxC3wFXrwRyxe6HulEbshBdo
WW696p8+F9GnNgvQM8jVSxOH18qhPJg4SeVoKvPIsI91rQASqmvcKyKFo8+kjyVu
TWI94/yO3nqNabKDifhr4aWmhNMO2MF2mC9Tepz5uXpawPwECkFa7ZgXFB+AInnJ
P0xMhZZZQhDlmQ/D93YNraUTvCcww7PzXB45ydkcXYoutGhtBNprNNui2NFUnMcZ
fctYltl96nR+pGJuhA1smPw0zdSoE33MGOgPD/KvUVqOAQkw2hzsAz68P+6hF3/7
pHaOF+4GHny2645GMoZsZSW4nUK6zxynjkjmCqAAcufkz3//aPmJnuBiiQDOhfos
B3O/m9/IdI5mDbhFKi99f8+jjVHVFfqYCrGAFyy8LVbASdcZfe5Z19sjapGfnZz2
72fXMdOHn8xav0Epb0Mr03VXXoDrEM28wrj8lEvX8cbPgCAv+SJDjuQOfau06hpl
f7JPJN3zUMQZdzCeXmyHA6kjp+QBbt8ZObZwWCQrROd3vqckdPpwaWll8DOFT8D6
dpSDT4pn/j5zPoMuH9qa23shTJTX+0lYjb92Chei/X6K9CiHuG7LeUnxl/OLSMQ5
lQMNqqEfl4jaNP6GQhNADG6sNx78sHU3SfSrjAYkLWZ9gLWTZ9d0x/MWrW+kNNkB
9bpGZh1bHMxuJOVrykRoy6OhaoV9XJDxNXEpDoY9EVrxfROWeqvcmD5qLUyZjlde
nt2Hn0EcznIvZ01feSmo18nB1OtV8ItPJ2hip2Vku+QSzgvLbsLo+IPb3Xui7fQf
7ouLHk58P2hJPIiABx3Kbaihcbbf1gA09CvIKCU99ZJCF7sDzoMrhO7XteQbAaq/
XYcDjYZyh/YfFAjrsM1yO+KlQ3gIA121AcWzm2yhUFTPSNR4VtyWKN8e7CfDAUjK
EFN5xqXXB6M18AabSVJcsElPVXWzgcNivxZWbYH9jr7/rRau1Dh1xvfl2FwKPBQh
9R1V+uFsU2teqo2SQ1ijhANOQXpDT3z7Zt2oKXmod0uAKIygjNkXz9z5fDwS4pnj
r53n8/QxEzLH962T5GndGQOSPbXcqhsG8tptMtqZHTbb62iPEAs+qD5ySfozE1HH
dY6z+N1IG0v29x2Pmq9LCuGkdwqHkqTU8d0vadU82fLdqPcXUIE5fd+ptvYDsWZA
8g2U+DCDetCocwyISeJdRX6qpOq4lXddTxSsvpf1/dkM1hFcrBx2WisIoZ6BYaU6
PbDj4qDv8ps9gWDJ5xK59domqarqBm3PiWdizsVisAzyfjzG9hjmdYV+kd4ns4qx
u1VHBtEBKSa3s5cEuYsgRG5i+GC/XOipE5lmx8ZCgn2+5Z5MY9d6VLOlp2DNA0Sq
23M5U6shE58xavPiHbbzCB63iCNQEerdpKR+z4bLOUw7mc2kGvTvJL4p8/g76KZ9
q4Fu/sMAwhFL1t0JXrkfPRqT4GsTBsfcwT3VfJVvl2tNAU6mpmawCRGIk4TY41oo
A0xh4Nz8FKBQon3a24dMw6lpwHRMQosgCaL1iJ9L/1qI9Iq5AzY4AHZgtCSeNzcV
6e7bsPt32eiyMjXCHIduOnAp8k20+av0SCAYP4SHjG37zaYjmyXjRCwLGrIqcixj
N4LB3hQI7sOCls3gGRWmbQLyu+Sf/rBujUTucLqsQn1b2CBqYS4rpAokheJohb5V
5/qWbhfjY5GMxbWbmYkJOspNUQaY1lPOyxPb0Y8gdKPJnX+M+aDwK/Q1/bjzfpVQ
MMPUdrpBCFveT3d7jp+BSuSQiEtU5/37nqDW5Odiq2GPAPp7sMia56xm6iChdMF1
tx0IpdiWD2s2U3zo6bN77LHM6Ye6T6RYja3QzcluE2iVCvZ+4WkAKEl4m8JepSCV
LAu12Eh85ZRFqyUBd8KoxbufgyKQB0Ii1UMnHq2kuAYJZe795cmMOx2FJ8ToCuPY
glSUHSdWhjI9kpewAEPX+fonOh48LdRFHkkuEWGlbuV/bomPhYFakY6UNVvRU3Qv
BxMJ2VYlYnrCpOGua/u8rJMQZOlAqqdQyY+PR0IP3lgZxiH1+uADWR6b5eLrcZDv
ztcDKkDwdpBrPshG2T8Q+5iUpSNVducUMFYaXM3Iqe/rC1m6SyTbtdaZ/ryWAm4S
9viGkmd3o4dPEKx6+lHfaeNWBpAyxrWw+CH/xLV60zuJLy5FbkTpcxHR6DYESi7T
hNLQlFcllwCEgHxC+5PpDNwoGf9Cq2m6Rv642lzCXU7fC0d0hoVcbBDBxfCAbYlD
3WKmQTLKKAU5ArbJlwaq/gcEYU0Zob6DMXEd2B16AotXuOPfvuRgJgkf8W8CiOSv
S5kowcZnwQw6LopSPWFLqtJsp0CPLkh0Ut9Gm1rOIQvzb2K/qfdWYVe19y7cCEEY
peAGJU6b8TifcUNk052LAr52fGfLthzgXx9cJnjKPR+mPS1oN6AaZXvxqED76k48
gLRhS603CZq8c/u9dz0Cv6XSITv4khjRZ+mw/3RXrgEfTeN2ZCdEG8OnFDEuAfIb
8ORTtxr96hW7uuflnYrfLTqsOwQrBePFezi9L5mLDSmrr+lomeUA0pVrYniPt+Iu
ndYK0NeEgUGL56X+DpJTH1pgK6xDj8eMpVJF57l/rCXwlwkzB2c6SObUF81+WN3M
tc8ex2cbPVvyBWFuNNnPSSnxH6zZZYHSUD0uB14Urts3zYaN2e7Ca0uwTV137c6C
GvdDO8bIZXs7wg3AZGgSolrauu1aXAguBM2XjCVKmsRlNM+IlTJJh61VemaLUhd1
bww0EFWtBdy6sPN808LuxnLFYmuCPavjw6MtF1WtM34Fn2JPycUKTg/aGXcj3yJy
Kb8jpyh9jNaqnxK59WWD2ClzzLun/9nsilf3jHDlB9CNDv0fKxMkbaAC6cJwDqw6
SLVQ3oLeZC09qgL+lyRAoXn1HOlbwinOC1oLPhiWGA2awb26W/rfV4MRqmw1RzyH
UNC2FJKjAG9MsmHx0YH0IyxznmtZAx4QSp0FZOv+Gev+cknny5KjQgftiZjE4OMv
4NnE784bDbwPBehUfFnwNgOqvfFfY3ZI4LCinCxgpNcklzfoemGOnzmbC/wSBlIf
VB3v1w3rDzbf6cJL4uMyi1yZ5ALJbaQ7frSX6VnAqsP5+nfwUZAHQXDKteTnsSmK
cMChV7RxNrzWX62OO+7B4L/4+ozVU0UiJbpXJRXsKjyAOF8vAayVVda3J6gsgTpX
8iV131nf4YV5kIdDyP3uXPI2JmdGgGCJR9Zm7gO7KSd2Wb6rUqegki+vVKxvl/yE
rsWN8I0cgEEuZ42dBLlviuRdiTXxcFjxflFT9BGzZXY1wagM6fx4FRo5j9qsQq4S
jRxo6Jk02KRhn4puGswwV/DcrWOX8aorGWtEoaAfMKZ3pgmcupGI7avQ+HNBE7/O
yny1fwzcUE/Xrul0aRrvsyI8SZsrmnzB5xl9aYgoVrrxFGxCslXejgrN7Jak0KbD
3OVGYqcp8no/SdOqRV9YjA2iigh2ynCadHFU5SAeUGxcGzVl3qY5jaM5ScJRrc2X
em5u/KfHm/zIRYUhlTUCpMcHYoeQsuR5dF8f1guExRZtyXNKQKq0lFlcs/VoLy8H
8fwxaOPdjJvvGWlvHQzqVUejSriPQScGrjyFNJ6ovKYlTdm/x5imjPOfX3WHKRS9
hizRNZAhvVpDFGrleHN56teXkCVZxl/13lFt/AGTKSD7JUqf1IoczbE4DVpxQK9n
JEWFVo5MPI46oiQ3A4bbKUcAp7fp9aRsZg5xVVZxEs0W1vRpE+yHFHRiTO2rUsul
JVc8BYU4PgyZzotAdqXwn426lYVysxx/meni1tn1G0jKFyaMoSeJLRq7QWycgGM5
D0ves59x152cb8w1hwFdv+8qabMf56WWwNwC79v3Hc70pgug2Qw0PzzQbWPqkD9A
kifbB0/ILYsoLogwFCjNjIfttqcWlLaxUBt5a/VdjMkuLxFs+hsJTFT1I48L7yGY
2AisqpCueX+rh0nM4Y+Wdvd34w9FTKCuNEklszTFT3CVHwyX9XlINa+mIdut+Npf
v5jXHSHszrHUclIX0uxUa4DA5P+Ufv+l8nAiffpRPz/b5FStz99XFhufKkwF2rmV
V3ahGZAJj94OjOcwTeiLJ6P1lGXfL0f2l4GAKpHrOKfw+WhkXOpMocjVcdexVZNp
O9zROTUJyPwUlDGNQ06IXdfhPSYFaDMzdONEvX1PDPKdjbbJHu2vbLbwST0t1Z9y
IWdLpBoIArAcF0KCQ9/8mrdvT5FDBO+gODMGrwl+nq9Qq3armb5X13U951bcG2Iz
UsbPzdRf8nv0MCO6FNTHyeyRXFxiuqRKKf+MxMhM/N0oAm947q7YwXoR1DsN33Hn
s+vtIRiMrRbzEow8v5Skb8z02ZvG8BjC79xmmwP8YxqVYEf+5O+sA+cLEVWxff37
yVN9qyF0zyY0aZOnwXlwof67Apzgzukk7D1ENkECasIrP7Uu3LORp8HnqiVK9NBH
mIYFemHqZnWrKpmkiBrA1pkBIch/Tq4N12RHZ+xp8+UishSLRYdwSWHfhDlzpnzt
xxJY8Thq3D45hZTRTLN4R6jWEt3HgL0DKxypMLqvNmd+rLugOM3j4TY7ehJbElGP
Br7CqbL7HYHkgT6wQY8xjXM88UuXkltqQuvodJqE/UrsTxVfhw7eq/EDeB2Ldhai
frAB43QlqyREJGUWEOIOYEBvwT/JM83L/BtxvbO4EfA5DxK3SAQbr1p7dhohwate
Ouxb9v3hfpmaZ1GI7/S/q8Zz+IxLuwRf/vMNqNxHCeW7bUazKcUyhA1U2vzlwDoU
9G3A/x2dnUKRXhEyIhD6v8Gg3+Z9LFm4qShGVvO6FDRM+3Y/PpFq+q8HvzW1Eg+y
nZdfPT5tkAtlEwHhy8lW/WQl60OvFimNI/gBwqq7KaQ52sQKp3RqfU6ddq1+bZ8n
EfLPW7PwK4P/hxqR50xayaZKaWgyVojOGg5LU4jUuAqIGjtV1MZdCyFKUXs5w/Ln
v7GmCKSz3FFnDLB6wutlbvLK5ixuttM+fRIryvd0Ke1Lk+ot6AaKXxmR0SIk1v4X
G4dUx9wvqgCq3Y4dyyFUVeFP6Pq7UhQXSImv5llbeHS//64cFCfsNmHChE1LHO+B
SPk+EgVrnZfb9vSV+aseSC9mJXdzdz77qFFt5fNXtRjN4D+hciqL+Lsq1cBuRSEP
XLpk1t5Khf+CfQnxBJneg5sSc2YX8r2iyHeRikLy3b9wgj1QAqQ3o7/XcaXT+U6E
r35q3CB/Rqya6CR34WX9DQaQYwkYH5icEdmRFmexBZrCmPLr5EDqiDmtftYFMppM
ecEu4m4/AWVJXvXKITH2Gr5frEDtvR1JvP2VrFR+IqQT1pypQ+uE+KA0mafZxbgs
dnKZZulouSePCyT82+tnD9FvUL9gpVunU4BlnM/P9C6oRfHo41dOGfHqRBbsuxOS
akcgnLTaYfnQYZpXZcI7o7fqyQZt7Uj7RE6BFQYrTgAEOjWoxARWJncysuIJ2E0g
RW2UEJWy4jhyxiSRJLunBQIt6cKrag53rif4ERX3na/oSZ5UamgJLjUajk9jBZVh
9LiI0lauCoEkiZCbqUh96eNmoDC1Kb4mckHxG1kxfzaglpWCYnNJIVPJF/+hkIhO
lXXAKst3OPTG/6uLJ2wHhG/KLgP2xmI+FJkzHzzXMPIy1W5dlUUzcKuzzCA14LyP
Ogw/NEFN7RmHNZ9blHgW/xBMe6s8FV6TMgCj6T5kBzPxulF4Ut0rEQ7T+QUwu5me
lEps30y+gBA2z41YWl4ZoVBL8PKr5Q/Om2LJTpOsrJH3jmeRz3mcjSJXmnktiT24
9GRqnKcfDabP72bG9Fh8YTzAV+Kc2lf4vApLnFxXvEG+p7kVyxO8TLpoxkkI7zGD
FxaEboHvyQECj0f7gUPNO1MDP1C5FHbOjHLRROmcoH8Nkoy6Bvkds+oqshqLd1SY
wNNXteehA+HhrkRLbfZzXIyXpcB/WG5WVZh61+5QTKzfl++nKq8eddpzlVhVMhCD
KYLhpdpmmXQfSlvtHlsQp31yELaLImC9LgWCqz2C6XDN2CfSMlzHqzXdp+5kMQrn
PMa1LKfR0u1vOGbvqYrBnhZydF6DJk4z9OGx0L3Oe53QkK8oZQFOD4GuwH9Ci6vC
y9+fwA+eO41aGyobi9Q78Nmhi6npRCOqoi8RtylyOMqycXVALpe2P2EbUbp1v0cx
8/XHgmPwuFSYGMCv5gjHbjFnZmn2oe3R69aYdfD+S5a+cvXTVt+LQzVDLxxtBdkg
`pragma protect end_protected
