`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IiUAhH+OTYxz9OzXBRT2jANybPEBVcXDHRU3+Sq7cR9zUwzwwcDp7+PIF9+YbAK6
ztotuLOVHTRcMR5Yr5xVtNGBfq7olpryWx7Pvqk8dFe4P/iOSUd5aRy4w9LSnU3F
MwGLXUsSvwoMWzoli/Yh84vicazIVzuTWKzO25qPW1I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
D11DKd8+uoEZoUWyDZYbjyE/NM5TV3z4RQObZUjyU3g+Hs4iCdiVzSH24xRIct53
Z/lHouKncEjPvUX7QNgwzhu37UAdR1WU1IXqzmbC2DDY4ft6+b7BGHjZLDsUbdgw
H6jbS3Ofj2Jt/fmYmHqY2vRzHh3eMCyOYcO9he4HsK966NcNKKkwLxPIS0fqS3h/
Ninqh6xwu55E8Surf5It/NsBehhjXZRQKuoy753JlnihzUq5mgpLMf3ws3VHcG7/
bZ1F6fXTQdulF2w0ZTET98TEC754pO0er2l87FsGc4mTq0VPVY/d+MTYO3WZ86QO
hSG1Gp4uSWmswMkd/rwOnD5xC6PFbgZxm9eHtfgFS2LT2RN/OhW8QsbjO9BRB65X
tCif1wt+HRm4Mo0IfBRSNG67rFUP5FcXgcnK9dIPTov9f3QsXpLPmO+QGc4Ec3BW
5EOKKWVizC1dg/ChvagRw5YUr769FC+EfLQWJTx5Dv2RPzpxKnme/cnKPk9K2x3t
C2yDGJ2JizaT9mq3QGUXNzgtfbYojZYBUT5jctxSMxbcrB9NHxiMN3Cw1MFUo0cY
NRSPM4oWpbgx6u2rMXWxVu8k2cUfZAUeR0xdbQ13JozrGQcNg2+PQ8X2iv3+wDJi
74q0seJNHOGeGc8sD9mr++vBx7zcEJTM6TLMO76JUuzKww1bkFyuao/VBsVJlsuA
mNzSEBgwhImQVfYAJLxovnGx+JX+/rXe9j5vL9+fv6+abgZvU1pXRtqZ7I18PS6i
BmQljArLhhwg7h43yj85n6UDY/OE2ywVvFqgNDb5A8nu/fxvU9NHSVAB1o+u/JwZ
hJc4EQ8/2AHKDo4xe4M0GJI2ApCSKghBkzOsVRbDildyVLgvHETRSRLTX/Jkdlc+
mMjxPOqIAVNcx8yNWXeNU4/KX4+tcdm41a29avKokJcyrsvqBzWfVoavPpJPKeNy
9qMZx3qYcn9CGFSJXaHkcG0Zo2SuLPEHjufgqOdXbYvbXPZU9qfiR2l/o+G8VQWu
/9B8JzEZ2TNTJtlMjtPsPJSx5po7vmCTGq15FQczSMRpBOXHL20rH0G8GFTsI3/u
/8972AZb2nJ0MuP6UxmP7OKJqzVWzhTc7yiSVVG+I5h4GdcIT/+ZVC8nxMoxa8g4
hxRVcE4m3SrGs28094xmqfvPb+Kc3AYNF9iZtJVVvZLP3VkSsN4Pd+13A9lnXe5y
zSh4xh9oqPbjHidB8viVwoVBdToiDh2338ADwB6f6R33n79tea34f2XUmNTdBEm4
s4uHJ2QQTDwznS40wDkZecUzvqajJ/t8uakPxFR5/Gt71vJXeGvuIOFpDpXNarbD
WSolPWFBzVH7+wgYtWUyImNlXr6g9/BNrvgMaj6deoDw986Mm0Zu6LJdfB+E+USS
OfDK835t886eVJDA2xrCY7XZ0MpXTdMinzc7aHfRIRHKXMkK2SGix5FBli4BY2dD
O1zqSv02NfpU4lIt9iZNdajkrUQX67NbaQFmZlGCds838Xv7swF1px0kiUJlAWHB
vsSMzBDpSmwQyA8cfQrFhLdGws979vYOecQMyzq3J080w/wkZBn4mNxz2OA98lQu
59lyfENFTeLQsSv3OfRMjQA+dX8H6sn/5exRVd0CEN+pWaonur9RCNI5N/8SUX9s
CgG4qf7IVD8tCmqnJik/T2R19yykO5GlCh2nP+MM+a+xZ1BFXcMCjzC/bktBTlXN
1pQpY5ZFg+nFSIgHhlBDn+uxoJQjbWCPuFGLQWLg2kilbLP5WA6H/58poNV0cCJI
AWDIWawKBODr9fF109lvykdBT90hDIt1MP8kjNuRs6WhYiLY0RPgUT9u0GA8KijH
RB9Qf4KrUtw6r5vaKGUhJMVKfdgpbFZbMVLSS9hD3yDU21d6/pCxipu3uA4Pcee0
RqCx4L7unq/3NIoXmmk+f4ejwa8FIgUmWNuB8sKKffqtDxJLnzDi3cxP9HMuJ1bL
6SiQ9SUmRci9lD7sRPhtE9brRwGowCqZy064SK8kX2aq+Bksz5Zgd1eHP9Qtlyd3
2YvBLp2kmEHcDIfRpbHRDEkl91amf2d7vBz2LmQ7tjpqPVl4N+Lmq7LdXsiH2frE
aC0EhrhWK3FSuGLyhuatuSKenBLCiigKsg1Va8svCMjojnNZ2tzIG+CEGeQn2+uL
MET+7FiVBJszd+aM+BHm8GSeQ3AlYawhxg81yQNwqdwaLtu0OrTjxbYsBytdMMYK
7m0nu9/UqWrDEdNSrwckaTtBfBLYBmdmFxT4SK94o70Lb9HXTx/s+in/AcOyfA8Q
cVrudrcAWMB0TGyhGY79KxdIecqORtLWnW16irTVo0XZIOSpWdyt+jtFeFDdXabQ
Dlqy/j/dyc5lpaO15lyrTP+7chWew4AiYdsrQqx6hOLnpR5nDVYW7cT7+PFcKeZQ
+nKp5d/pjNUxfU3KHeDdZzW0mMDj00g6EBm4HOOkE2mWruJLzkR5znSHFDfqvV/p
2tZvuhWOk5p1FR3uGe1q+o7pFOxQYEUYi9IAsCZcotyA94ptL3pmY3+MZvyZE4bJ
u/nHVdXzfuYgNtEzzHUcB2sXOTllDE7Fp0eCP+ToJlmljY/erM8QO4gFCTYlq+P1
OHGl6Q62ScfBofm1rYGxTYUnSCViPI/Itc/S/R6H9oszaviEnnd7Z/RvPUMi1L3c
WYzFPWQyDE2K4i7gLqunqUCCzqB2Y3KQteKooYVa9J836i9eu8kq4gMtUwuVHrqZ
iMiBrqIS9eSnUlMXfcInsdqX9Vg+lO/ZuijKaLng+S5vQBaB3sabY4iSElLt89HG
9f28aZ/EMHx1ZxGrwy0yG5G5loluywnTvWMZy2PpUaUfl7mjffQTUebsAtgn+qxk
WOsrLHTNijEPVlDPtbmfrmO1InUFlCuKb+XaQTKOhUUKLSdaMua2mkR0cxbsSZjO
5LOva04Lm3Q9Ixmp6Q+dISDNaPJODy0tkGWR2mJ0Ov/yGSoUmv+Kc4hISUWDiat/
AxK8+H1t7lB2tSg/7pXcD/SfMXj26GsQRfEPBCthznSbsKUY7bFjYscsTn9cV8CZ
/vVwCtzsSnQl7RTmbxcqQbsLJQODrrfHp54F79HwYRFmR3kxEBEF/q1bX7iU3cDG
Xl/jhXjBoohwkKxVB7zxBSrJfMoyuWd4svXMz/n+unQWeBAZEWIb9KmwVCCbMvra
mI5AjOOuc8yT6gP9ltBfmT0v1onJ0wR5vsRitl5jgAxlU2hxpOZtLVAGyfclyS7i
N4SAr/xhE06O8dT+uOLlMdU1UyakdqGWGyiNA9s85v+JXRvQwNaW1yJmuvZks9kO
hrOyl71wNct0k7mYus0Rc/wS/iIqZm6kpSChXtlJDrjTj3wfcXcYTThE4x7Spczv
NN4QDob8KPHeJCrpvLpaoRMHpoCHrZkzlmAK4I+vpPD/k6fRWWrwZ/LMCg1wFa2V
vZWb2XCMHaGnCmxe08BQPQ5hoEm0z/uZGEHoeA3Ly3ypGqLK1DarDzppZ9Id+wjJ
8ATyJ5EnonlTInbi7IgiJHr37+xuz0W5p9PS3Wdh5PvVRTss55AsbLY6Y407/oQr
kJbHCPm94VJ9ITbJPQU1uRbhYfDoUXnFqLuOfYrp2ZLgJTHYepM1P4uAOJeAwAvk
cEIVw/4veCf312KwJZjAVaTIDicAPLvCEC+TSpF6kA32KKZ8WxS4whNH9GEmQHFT
8Qft2DwepwBjR4hxx3rlDS6q529w1OHZlfTgQuamcekhgHA/33I6liME8ApkPK6a
hn4i4ra8mTqwXgBPfv0MjLai3khZ+bMk/sKwNGwAMEg2H/7pm3kou+E2pyEmaMDx
oIsm230vB2LpGqnE74jqsyaUA1VqxVdwo2KsgkAxLAJ4/lqN/2UVf66v/NBlf1wR
mxgnh2lFJu9yWfhD5cKn43bf2LYLY5OWIY55znfP9xVWBXIyH3ZTGtoRZXprRBGc
qNs0RLYje+2gTZckOF6lAkv4s2dtskj+E8+6LiCTFe89jsnnn5MnQ4+NT6eCSmrz
hg55ta8iBLZzSo9RF3ZtY2pxCLqYjN67OZa8pa3sfI+/CMjYAEwVD090oxavC658
bjqait/SEhNm1iv5tnG6HDJmnOd6s/usI5lnFcATTK0y59cfudG0eeGtN0nfs+NK
YQotXwIYswjwYlOewnc04gr9osvLe7cCX2OF+ZVXDHGEHZSgCWSoyVECcolxN0DU
hbMY+Qfl3Y0TxCxMf0mcCmn/KvrP3xawHbydZx0PyMXZJYIVpQge6tv8/oTpM0o/
yuwQyEHcpLSppQb3uwr9H8zi/OIc/WQJ+RtQDsdlV8XZbixS55C8IA+ihuJPGQLw
ZSWCBExq39KDTgXYrJIZgSGVzREvtYofY4PkwVOP0h5En2lJPo8jaPjXDS66xKAa
o5rHgA8ivBS4KYnvYc8gBUl5rPALuRUTKNNQBo6oS966TvR81hvtx5lPxvnFtLHR
cf+PnEIOITA+m+zNGzW8/4VlsPcdY+lShLVkyxdWcIPfNrD6rmtl8DH/JmCI1Ur9
IIuRTxX4acqxK7prkxDdzs8sAITSQG+GbsVpHdkJ0Xyh2sE1P81KmhkbsQaORY59
mRUAuooKtoPLcAtKjXI4trLREnCS9p4bVbfdbWRv8lvXFGRHUhq8/lOCQh89o8qJ
G6i2eGPM2LvaRV52I+zkaC0qZsBrSAzjOzjIQZsuEBK8UDT8ygS4QqUH/Wu2SpDd
bt+saxObV1FqtFg1Ux1dl/s1rWXEus95E8PMyv6WhfzoAgheWcO+W6bBPwXQ+Be1
bHivBGPM7r2IM88mEGHvNmiaopxM5PuZRu4xxqv1BkTlSAmePK3om+gvSXruWdcr
TgMiTiRnhiAPYbADRUT0SsGkgadY+AYgSd4FfJXTgdTEHHFzHDyCXpY1n30pheWM
1J2JpPVufW+fNK+7yP5tDaondqWz1hxjQx9YjTd1eRyWsmhhyObHl0k+jOUEeOKW
zQEsXJ8oQpA3KHawrMXe1j23D174PnQG8nCB1bZvzbm3l6CzbtGbas/zx2S8DhPc
ZFjlegI2piKseFu9gjfLAfr5/M7+lg98mrZgHi0JVptZhxxNHf4AZgrDX7Br9o1a
7pVafAVSrJqZKcXJOIcCsxMwjpkLQ/hIS31nqMC3Y3NeLYpK0Rp7176gS5Su8Qtd
Qy6ycH+4fdoXuLvjPBK/TOISgb3+OooOVKT92Fy0v+7y0P05XucLkglIZ3XUGE+A
X7cMaeCMjIbyc5tQ47V3Z9QMzsry7ej1eHq4jcOB5RsfabrUJ6nnWWJX118bkmbo
lrVlnv+B48ZNwgaUwzbhCm1C9+NF+VMZn0bptMmuQ/6Lb3yXy0FsYnTsgH/nYpnu
EYhcynaIT+yOrDrO92V3stsNaWFtC3/zuy6boR32SojdW9DBehvX8HLQ1UJghPto
GciRrW1G9H/2EbqMcOgCJAucpKQgfdPiKaFoaRT+iT1gKPZPFuNG2CpO8fkh2h4V
WTlSxOO1MSyODFO7wYt9GM18g/Srl4n4ClpEd0t8kcVHGRwiZhiEQD8jRyIQP/ga
Iyyk0sglNoIaoBg5xvh22vMSAZbFCgcnVQUXjimUht0S7me045psl9VeEZYSQqLv
Ii0P9FjIcusjOs+WvUWDfhpecuYffG8fogyExob8O95gJkQOgcLlOK60J0Xk/XH7
p3ULCLBPeqESyXP3l4xWcYbXQNGWvpDk3qoB0XvDuc/lLm8uWeTiK0wBrk34hXc3
qu5RwCKxV+L8/tzFf7T+aOKZzvRtbZtWYVaf+xJKl7Kshx939FJHR9eVaZ3P+CiH
iNDIO7jYMb8GPIoLDzgYTln1wDbzUJ6hR9RwFh5TRnI1BZQytPHW/6GxfkGZTanL
b+j3QtBCFbe7jlbkmbvwHmY0RLOkghxvPb3wW8RNYo2Y7aXcGa04/cz5LXSeQENL
zcAKfpgTesyclkLqVUQntPN1zWTNw4yKlctUCr+NEbDsHgnKGnI91atPazEBL3at
katjijAbdUxI1sdUA3mjJW6tr65GqWoBw6EhLaFvKPbTbnoTDRh/1u/n/i/zZjv9
HCy8HhrrZ9w9U2g2xm6KGFSGZfk5JR75lPe4nRGeYNGRAVyTECXitZjxJqCv3g2V
HScfeUqhd/HDvafs9U5s/SqMGFk61fXEnQTl+3UsFwSkjJwTI8Y0e9RuiTkH2Fnp
uTc+I07qtRhInTQjhwQw1KTKEkwUpoy4m/FBtViTCekUfuzOKh28FkGZM++YP8Zl
vKSPU1tQGWIwCn4erP+3oy7zPOyShM2UoqPxZPccADYiX6NLtl876+me0oSw5fQa
lMBZJ7HO+7JhUxCYaKYPp6Bu0/lmfRFhAa2AgPwsF3oHTJPSfJxPR8trsp2F2bAW
/CN+I2uIU5pezJBQqxIVYbeb/36bSmH0e7+vHq85FDhrRwQg8qO3w733ptgMM9zn
qj/u9v0EoqzNYhF2+eVjcCMX/E9SSsy/eCYWDWL+vvMZ11ksnbqjMsYoVTjMfTo3
Pw0nKh4XuCyG7B4V5VDpcKV3ue/gvArNSbOtAU2tzXsBo8Zxw63NiQuBGoEnCfPC
a0i86jSRsv+x4ZsTEIjXMvu0l0ZgqP45XFoEm6vMwq8PcDDG6fdZNfu9l2jpdYyf
veUXSE4ZEA/s2ZmwQDtfV7wPy8w/NDhqZ8sh1mwZJlAvj8wu7ZZqlHXiLuZIc9wP
E7CoL9I9dsp8Q+zxGLwzLOZ+PzUBqQfY1uuj1un4Wx3j5LzTj6vu6vOjs5MHU3sm
xCCQB0+k6c65b9MTtAVC+ZwwioB2TH6KInt5EcfSPcTbq7Kc18thWrqDWk6YahPq
Q6/Orti33jfN8EXNIK51NGFR94Lpjv7iWqrmeiBQgIsD/DvNi6hRHiHYzlt/uvZH
M3VbXyAEPt4Qm/5lxmap28aeEPAeKzL7BYtnYjA4QEiSHLcK8iemRvT3Dt6NUb9x
7Spob+6jfI9seVX+3WArlrzq7ZUWnVptT4suQVQUUuIuif/yHcxYjDDpu4mE58b2
HyP/nR05QG/Gyh+QAAwlRGCK3q0Hl9e0BZ8yze3X7tGfD4+iGuHcjI1sBhe4hcYA
F7/eP62f8Vsg3q3FbXIJ6iipKRJgLnRZOb1BuPtJjWvaLW2G+ihonA2FwyQKR1D6
flMSmkoROy4ul167eg3xATgDjgBXCtLvg+0xbBudxCTyGWmv7bU/ojtqf45qOaiG
nckKFJzYeAcbXyZI18nJUNvstyydo/f63OuzAOgBSnBFUesuu3dyBVqvyoLh0oSD
bcwSy0FsFm8jVNt8m7CfYvtW6glyLOhYn5H5bkLX47XWKaMc0DAXiqS0Y+lAKi2E
pl7/7dxye9BZf5D09g2ERRxkKw9qcNFhHapYpiLmA6GumEFJBDWo/ArKoKY8rfi0
zxmvaavyUv5EbXsNcERwrw==
`pragma protect end_protected
