`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jK7ISfnDTFfLKANZ8/bhaUk8bvCapAwrrfMXXeeMSK3raeOL4KzLpF4lzaftaZMz
FQRjTSIFZ8k37WxnDCdVH+jM2eZRtZEEfVueWcrURIp8bX7keQK90RZWEQ9oB1m9
CiF52yM58gQHJsBddAk7EhigqlWQ06JfkOSNW8Ihkt0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
XWiEO2WlZt77xOJ4pXSpab0cQSMSuAXl7DGNXx6aBw7krSz2sf0/E9KzuX6C8fcn
H0IJkBalBThm6Nt4ITPAH12d77irjVwNZoFmwdfXPIHIMRC3QHBozEp/beLMwQmx
MKTCv5Vxo2Hs/L/5vfjuObPC9vWf7T1Rg4hn3sIg8GZGC2TQc9C2oPAm/ABd+BtA
2xz0I87ishT1zalX4zq2V4HXM7kqhStMxfNdPLLgAV6JlVBjTJ+O+y36K/Bsbg6g
c20V1OyzwzhXSO0X0vtMaLgPMABgW9lNRpKkcMUCaF+6QQ+hXbKDWVyxaJtHU3TO
Hw5mjvx5UothTEwp6RlTaYSTbQRCk8AhBS4BF0i9SaayT8i5onO58m7sczV4Nu0H
Jpt5vi3KfpYF00G+zwORPUFnzMfL+xpXzXgWxthwjVw7NNr14lfphP08RQGqCeDb
ipUHnfmwwjMS4j86YstCNyJXWF+eluM44gM6gz1d4qZx74ZgBX7/3esez7uHAPcR
6DDBJDo7O2kgjQUdhDYgKRmCB9Bu1CtN/g+itYTkaaHxUocri763OwwH5VbMfBY8
sPJALiwTA5014AVDTwfH1XxkQ5YdB8W9Y16lhxoSY2WBexWUSbanKLc7WNQ0hUSP
1wno/18MaVpkZhbcp27qCLvH5vSWSkC5myFheDAKW9fXg8wetmSUC6DaEl9U+0C3
ee0r+fIWauSt4sRZ0Xqsgwhx2WbekGJo0EDcauxMZIUYSS93o5Pq9lX4UvhE5Gtl
YPzQhdRH22tpPrAqqaItyI2tdaJVY2TFHlZBE+gOFHKcQ2+ymo8U23pdjloaKDqZ
gud6sfmm8Fm+t7iEwgAn06CuD3w+waC8PxKiBXql1WmpHzvQ4Og0kJ8YbCO7fEd3
PjiFYU2bjjr9utEmoUsjvY8w7M7KQ1ZKLtM3HYHGJ8ddh5ap3SnSQsUZEZyVjumv
aEh8SzSxKOiNNGBRKLg/PCGSWwopQgXq8x4oCsoIiIqpnOiVEph+uZflVZ5+e5np
VytQcyjj3LJ14azdF7GaAMHFaFmoCHD+4a1l2yOK3ZP44IL5/TVrSxQTcYNWOOnr
okeR1WLYvyBTqWs2d8MG8K/c3GHVAnDayIW2EIvtOeOjSRnGXYPPTULLDYT7iNsf
dP+FRVFXROQ5Aajy/tk5rjyVS526X5ViFSTCv70ICCjAejsoc2ZeSSRWtDHhL2mD
ePReP7yU4XeN1oFFTtFKWlNZifWFqnTxgdkYxl+Z20+wGVTKyAj9gu6E+PDiUmuu
HZtqkfFuqdo5Ywm5SE6ZZDWVfihEae6BhozFXb77vWMIQ//o6dbCR/gh4U3GiCtU
FRLcbEgoZn3+iLTfgJ55Rj77yEul4VKEDZBaNQk8RPzwSrvP33K8ZJr5iufTnFrl
ZHQi2gSUfmPkzLV/BwuBtPOTxZhx3WX6njvcFTiGzGppEcJvxV2TnHV9Kl+g/3Ys
khbTqUsMTboUglnQvvwcQGY2yDDvVMEzoW237BVC20NJB2P2wyfpYt3ZE+c0Orfc
FIA9lS/mmB2midkhexVIJDlS8EOEVgHyM/CvmISd2Bsk7lInuKcCnqR5p1rzLN8K
lHvyrzjOrfkpCtKjE5a7Rhf4AjK6GDSK3cpHrvTLSRCDjMqK8zPb6i8OALlgYvnn
4JKNyDV8LKP7SHRbga1Kh419vJY54/aKGMvZmSDO5GxxWfstdwgxFMayw2DPAef2
wF3vV8JB8ElyfImgm6gebFEdH4EfXpFvmMPT0apb6YeUttXhXbIeS8pBH7haYpC1
aOchENI3XUOlB0vWxpElHAMcreveQt0ZjGRsvWx9N0U97olgvCfGKppkzMDxJxy6
vbS5qFnr9gh8mpQVvtgNuA6DniQEN6DQDdLRWhz+HekzfyoqDT7UQur3PKIqQUax
xtzpoRf6+cs2W1LnZVHjPLJqbvhBVY9D9eVdqS1atMe0UR2IblzY0LhGCXXyHED/
ooZhDgC7XSormu8p8IkPXPC3cbDh8LG1hNYANB07rko0TGVS86gGaufWSL5d5XaK
2TAXL+pUuCEL8jd4eWa2Lg7tcJqQmltU6QLL6NJK9nQAmnFeTHdiFovpNyxQP7gt
M+R8RGk6sXXiX7BIaNkA7lOJGw9gsUgOCmhLsSaPVyzKAbO/g85sK06t5JVo4MCq
u5Q5tmhtsmZ2b6ClVqNiO2MGW6vzYO/z4UBOj7LWFCRF/sL6M8V0hAF/IymXncon
AQiVb3xXRpoBy8BXZPSr7rGuZi8JNqcLq8Wi3BJSDvi2MwEFCZyvRD+8mQu6cQgk
c6i2xW1xpbPozb552neglIqQDLoytFRJprrNnEjefzxdoXDe0QHDjkp5/FC7y+x/
zI4L7+eJez/Pn1v9ERG+60vcrgcFwtRphRDPJamVr3DNqT5LY0lnWFPy1xHq1Zam
69N3bGyavFRvxoRxq6eGzGGZE3i9+UnSTyi8ImyG7wq3EVcSERvsysut2BSe8Ekl
oU9DePx6U6I5PJ5paTMSqoDwvehfeMGrhbhjocjLKPaNjSjO11E+8NHvJ0XMHiH/
5ZFklWO+qpQR8ZRGTKdRQDwZonqAvn+zNMkB8p9p7YDwTeoClOBt4r2UBtdq38oX
D/QwHmg04yx8OrG4amhr0HyulhgZWHWT3RXKa+oDBqwchaPlqNkLK/kXLnV8ZW1p
Fs3IMmeGoK4+PX6LIG9OEmOcDaRyE3mpAr+tDmYRweWwMOpK2ji0hPfoP6E2Egfy
BKt8U5YexWU4IpcBKdgS2KlM5otGL5hpiM/Y1AdXrmIC64Q7ppeCb5uAO1K4/42k
scFkxAEhhYo7xNgNNTWrLgWvveef3p08xjvekXzttfJk8fH5ooUVHYnuFW7x1U45
uREmzFSbRIkTPR1WhpDnNLWXWvGDccub+6eqc0j+fsFu4kZ3Yqu6tPfuWXEm8WVL
As9hoO5QKq5NBWKV5hVI4Csy8SIOO1QBfLQyIgFdEVLlZPC52lUwHGMV9SBqtWii
xx+gpEQ8RaMCpgdI+RhWlir4EsHGw+5lQ3QmXm1KdAEWvfsOPBrjxCWE+znJJqCH
GEueqTWa7MaVFnHBZo7S+sB1fZqYTzn5Ux9mbnRd8N0W+yLU/dtLkN63DVFp/xGa
imb+Tjb/ddeh4Cf0ejOWnHOhbGn3IRd717lQeNgsIxXqek43dIhrcjx825Mp/6Lp
+RhWRoWQt6ormHnyGnwAuQFtmL2aHQXIbhMlXc/JoqGFrozdBF7EIAr1rzO7UaHr
i9wce5UskDT2B25QWk2fu6Z8yfn28bDsxQDjUrTopsxNU8cH2CeQSo+zQDmHpyvI
NY4prSdZYMDUuD9248v5wRST0YRL0EpR4uLAydx6G0Q/ztpz6U3CfxkH+TjrDGja
fZD8aAtd7DpRItYAc0MLl/8xvtANrSVUHeYt46+sIIoKMJBccdiLwByh3QmmXSxr
t6vE1mrx36/TUdVgcljV4nECDpv+Ch1opAz/FNJoGKA2FIICmKIvm687SmQ42OqG
zjnlkpwyov40R+uRjjL0vxsUFCdicSU+x/pmf84rqe79vq/6EzRjsxCppRiY9mGk
uOC31J13IBApAHtZCSDwn0JkHQOhEG9ByClCMFKZwpXu31jsR60y58BrYtddq9Om
2bmo2FRIc7TRNjLLBSKdvpi9BpxWYaknzlb6n8c8rueY6Ex6foL/B+PAMhU4I0dq
j8ot4584/u+MoWrWfCWXK2/t8SezinkoqmnLRJro6YPFiMWozC2FUzL9oTG0zUiB
QTDcqGFauNnYi30Glk0KyzvWL+/6Lv0gX2PuYr1BGEpVzzMDc2L/kU89jKJZlDWQ
hXv4pqpLb041xn3ZJHhfQyaDIZJwiMRemWQD52bUi6QuA3NuiWWW15vr4vMZ8C0C
Qv1pzbVQbTaIYoYb5jnayo9/pWAzoh7gfE0TYj9UsnP/n641C61wFlQIZu7Q4Fat
3qvuY5cP06C+BgkHSYwS1Z8d+cRzGeXSQWZcGL0mf2DpLPR3WlIwaNzO1IVUgLC6
0tOFWxOU1k/X6l8l0l26IXp/gkeuFnepoPWCTZqxOftatjegXtSfVOWRKITdDV2W
ubqaRSBq6p2XVPImfVJUAd6DBxzYnkknVgi20KbCvFRd2sA247XCiHgo0tefmrSr
BcDF6BMmxLwD+up8btzSMd2QqY2rQghbBGK7ipqlvrnR7Be98riarmjn4HxjLqoD
1Lxw58yCbTXSPznQrz9as+vtw+mTbpDeLuZjpMHW0AdcVLQzUoGnXpVrEERrJDVp
6uyawAp9rJavrZzB2rPIB9RQzdIBXy5Z9OVM1oD4fZG6O9wX3mTeOL6ZgSEd94bl
pDYxTx6SzM2sJe1RqtvRThhtAOqHJjVKRkhURaEvZjADcvwT9LXqTByjxBbcF1wI
lwp0GE/TqO+SyEf/bqzfJtiQGSWj82kkJGRoffOwBnVapeNw3DZTTrnbnyERG0fi
VV5drICKkk5hurHrcXsuuS1DbyubFgO87VAUcv+pyZz9S2WGKwrk6mex24VSp+zq
lVQ4ak3e3ehcwhQmkZ8JSoYXuqPPus+yR1Uxnqa+WdNc2qxusdOLpD0DO+8hlHih
xW5Vo/btysoyL949lUNIKYfhz+k4B1jR1Mf4RE5cL/TxqhNuXrcCsAk0ZnHfZBwD
TU7ycRIs15xPsxXQpfr+EB5KH/9gLVUZKsgn4/HVjjIvWoysG/VbS88Pbg2DPgoa
jnoJr5xnlmO3EUDKBT9neRxb1BiW9N+vYh9yryFicjmcutrg4AlrLUzQ1dlAhL5R
CRgWEWQdy9gW0HNKfOFhZA0LvGii5YxBhFiVLsgf3DfZ/J0DBu5NtmIwQGnZwrcD
zeuY5I84kEKJxN6nJejiZ661+Rbv7G64oeY27VlMEhxt5US38d9lbBSM3Bw56SnW
zAKCFF8f+BKyT3g9nrANEYG+/LcnRWI0Dp2Bw2Aysib2NpKsbgS5U2I4qmwOGCBe
a7ejgtw0C+rST9bnlwv+3zkFRQPWj/jMukHBYFwxOEhGSFD1R3Df8BITGIYo7BDz
wkeyD3ImmNQRP2E1VMlBoN1rYqf5xKkm8BBakDvL6OnCVl0U74JmYxFfeZthveTi
Lo08rGh2Rm9BT27Hbbt8eOfQFzd0Yn41SPXmpIX05dnb65Gu5ieKrHUoET3ZUf8Z
1nVQntxl9bVZE3HrCUCrIIe1b9BMttWerRV69DBvRH3JHgdDiR7ZHoL9GKE+Kcxk
6Ozq4cG29lGJjUqwWx3wFEybeXYCa3QoUYI+r7FgdB6rZP5ndZoXzXJ9oFAEW+BJ
0qDwzR52Dhr/ZsM0lnWy8tAXei1IV+8ygzgqKDHcsHwBhpxXy24T2vpnVeZwiAab
3M66TojS8mW6ZCzFpATOQfs9CN2/Gu3JNzuX3hhueAuRavbkiZt+P5TFk+EKdKho
Yhb5LzUVEyqnfg/MQp3jVYpd+phRvCzp56eR0jBAlItzzisfPWj7RdkgkO+AB2oY
Z2H1nuwi1iM8WlNhclVBQ7ATBokzQtHOp+J1wThCoP2BwQxP1+UQX5fVDzdM7ZIK
6LTD0wiBUGhOpoY36gt+PwqQY3nJUDnA1kBjHiaY8FqAusbirPOdGYOXzALTYT4w
q3nPJhgmzDatR7opv+vKRDnEk+o4UVzx6CSc39orgk3GOM8Q499khV6FQ9xMgLXL
yPfYBgrZiXPcQJXVaHvbx+WzUvXQRI/IF1nrtsU5NAXK1WiWwE+wxeO2wWVaAIm5
ZdBhfyY7qyh1twk4KAwD13Nd0ccweFiOIHP1yD+Xsf7/5Qj3xz8D0U4Xw1fG3N7g
m031Jxf//mVw7RYx6dvkKfeRZWASVfAr4ajTNkEv1ROoRI2CnFr1l5l8kKahG6eD
kiV1W4sjo0+FKvN2K4jTk/4EkSYkduzrzN9gJjlL8QftLmLO2gHRN7JG4BEctYRz
M/7rUP7geZoecoUL+xec1941/UtaRY3Jq0zUhdzlTSlEM3ZHFPexCmPLi3E/ymaW
L75/RVGFFzrdN0ZjVdSpzD+bgrF5kwwRlY9pBVlKfdo48b7RNnyPUE33kpLP4bP2
jujkHWXI52IwMwLfvDui6wdY7CsPEra2p1HCRFmvRroE5cSG4uQgm1QGqEA/nwRD
44NDo+iuDVieCm9nKDjAGitmFQjoBU9gXTgm2noEomajxnt2iaet5Z8kdY6NxKFE
7MQ6U9qSCX/Ngq3Eqa3noFe9wQThyNlAYpAtsHkBIN39Fuob9QVy1deXGph/KLr3
9Wc84dNqqkUkO/oqovPetlri2lcBbFhBat82ZMZ6hpPcdTrVoBuHub3j7TmboyNE
yzaO/PP0OZEl6eR0oDQWKf3p5WM3zp4pGIUB4CBAfLYoQSA9S8YQ9omSDN4Bh/Ix
1seEMDd+uLGUVwB/56PCxEFx1MQItzILrH/xX4BLmvy75Rbir4FplOiFVesL4mK/
jvLASCak1/ohXlYF3EpWM0q1XTPJc8sV9hHGH81k38whlFuJBh9vdBZ2l0kSYpsQ
UTeZtASnV2lQYDbV72xA9YJPVIAzPsHELnDhkBLyIdcmTdR4q8++PKwy7012Jk6M
zFqyUT2dyy8IE/9RaXuEFESPMZVwEXu6k8brYkViWQgonGwAQPHkKN/f6e3mM2ce
gg2OLGPnZhqkeh9PzejdBGv27ghNs14I9G+ZZZL1e5a6EVF+lMGbDlzqS3M6I36S
jZBGDWSKxqQ2f485ioViphrGSjLQMWMllATAiqppDlAVFW9xmBxIcDgjuLYk4tx4
3WtzpBaDQXT0K6iY2dDAQnESODW0BzK/oyzIwisStIyo+o5LVGtlHRCY822CeKh5
eSprgp76ltiXezBiwd6QcnJSPYCrBheIMPrGGDYOI/BmE2Vvx8GDrNdrCZlDz2C3
u6Es81hzK0Jmi+luCtlHi7/n8xF2fgWqYpzXHlkWzljK4RhWIewIBnwuUOym8xsu
jlQGrO19dYAMw+HIP0tjwn20IZLTuqvv/UwVIUN40DQVkFwAnXKR0L/Cbn1uwyTw
l943N/4x6KXglkqoOI9xzEPkQIZArbd2XX2RKeMxGHWhCX1UaLhFw3PgZymf9mMI
vLsLRtWhjXL/8UwIBnXFUfCatxLVS4aH6I8tBZe9ui+DHLq2TjWrlko8Izz6NZla
cDj2zDbN3kF6EbenawK6t1gTONKKNZgBLk+okKr3fpvUNU6mfsAgVh5rCQcMftSi
8+3RmCPjAFAofZ1+Y32uOpdp1t/TIBhQWy/BDo+Q9b9N0dlRfylGUOcSa6jFl1Hm
+IBz9KpwfDjsF2YrKjyw6jS85MOZmU6NSq8YM43RnjeieH2a/98o3bbkFbVpLMbZ
sdnrClRABGpZ6bc0L4ld2c7v8ogalTUAtXe/gvL9M2jB6URDhmpEWXdvgroRt68h
90MPw2BTEnj8WPkXRZViE1SplrAeFqMSfB/GT8JZEvcl7bTZjNRfko3TUBvUjTZb
xV4yLOnVcrD7fMMuuDIXDTJeCJn6VAEQUYd2kjSwZbnrZseaZ95nwozLuAIuosSn
P87OcPXqmY0RN9fsnxs5ZvyEcHlBP25x0lmc/Mt/iNQFuG4fSV5XtXXDcT5jYNqK
RNmrO6RJ4U8+O4MJGb2ul9mW2nmRRt9nqHdKDlOj7Nnt6zBYe4aWzC2cFycnAojV
Z4w962wXkx5xPKVFb476vXy7WG59pbrt6t2JJvzhEaT/jG6AoYwS6AkdiSCt9MH7
38VQsfgTythUahUw1oEuss23L199fvFlc2OYi1tAMUHAyg26u8PT8D/LDefQuOUW
JCmTVmTAzfHZE7PLAXfs3eMafWABJxQn06UVIgICsybrcC7RP6sF+n0GRnvbHsXE
gHSneTFpf7rcI9CYtUWGVrz3FW5Se4qC1qgZW+L9KEKteo+CkQI2IQs7x6711NlR
4tMlMbJJxQzlC4uOdWpeOJBsMHNoZ4mBw66FMwBamIyUeVolNBg4OVRmsgzPhs8C
rmXLlRgbj0iX2p9OzuRUoQxEK+ocKYDinRpKhMtvpty1W9WWXsdprwAh/jxUk5aK
HnQv/jXxo14CgtDVNDPLqeucJa5uKJkJ5N+0q8TmS2zP4FBSkFNEM+A+qWNdCX/Q
KlDOR3ch22pTxH8y9kmkLZz5yoXz/b4apBDH1a1kagzky5KiFnTtuVhTln3xPu7e
jeJ4yA3LRnTVz8/PDAsheS63wXJ8xDDgWydIJDQhxuSmq6ncOEYjOLpbxhS/uGS5
MU++AD4MO4EHTHoXcAJ48Pq4DzuiA3vnN4weF2xT+7s3KAn3hFz+YASDxtpJ66Dj
yFNN2zHA9CdaRrmQ8u+NLbPptagrqGeAjCDW5v+1J64V6mMo+py7IJM4gGRFSNLO
z1v1qOuXG6UYdBQ+NqX0YorZ8MaKW+eDoIU8T5Z2TbMUtrjK538nBCiGOlamj+og
x4PmpcD+43ExGaKE0FuD3xuuz5roDKts6qD0HmhdmJvM2GUwzJqGqwCFmWyw4Lca
2Px0SAdPnWVpsyopyANQDm3/M8fOjMaGfI530Yl0E2QCx/T+4mjP7n8Utx3Yi0CU
Zv61KO/vOLy+YR4rWf/vaKby6wEKQfHFVhzYLM61Mo2ePVVkNm2a224Hy+5QHA5S
imryvav3DluZIN583zpDDNvfV69qyo+goK5h2nsnTRE2YP7JDky4OcBzcbiDGv45
/dgRuyxXUUPX8vioPK/oM7rVE4/L+Qh2NuF+NZBBSPOvjAhk2uTQZgro66bsQ6Jg
EH9xLH9yAa5x5C5Dx1OnyDZV41jNh84Mwb8lflZD0HiKtENnkV0dXNmwP5dhtSPF
MwdJ8Pd4ewb8N9hXvJysZsd4hHDTLHhvap5/xVhy5oIJeuNZs264jegfzOjZaBE8
lOP3VKRyAdLWfFnKNUjsTDfwqWiiZ6Y5DBX+lYugZHWxOeJplPpxhCIKXRUTTLjY
zSgpQOCs8jgf99Mi8VriyiWXRrjtLCWzlakYShKDKVTj44tQTcW5GQvOc7lsWujO
RR2tKwKiN2PpwNkMwwSCPg4GDyrwL4ugAbABJ8aPcoxPVtGVyDWWMBwwTUHGnU7I
3brfph+mOjAQOon1Go11C0HPrl9tBpitKJfc52hm4uI/1NKj0xXTqGxOcWSmlfnj
/mKtrD/eDH7Mtm0FyzRJjHPvOE6qOIvUWoVjX+nVsPTgD7mNUt5ohsO8u/ZRLk/W
ip6gNfGLGOE9aoEXr8sOF0ukUOp5MLIVgHE7AFuzUygyFvJ4xnIFu32Qxyv+yBXs
novGNJWidVJmgUtEnks80WWtPvv0XmcOT+WtTMYYStZ94TW0YttSTaOVen/aI5is
U+iPVGvwwS1K3Tkp6TRReT6ygLYVrExXJtHsnDdKvg+BPugDMLxmvkNFXnPHAjLG
J5hW7bragkZz7hyWhqAuEnYZ9QPNJiZftmpTc+d+CqUxZugJpQ/oUFeqz+IFLQet
36GYHKn8dwKy1pViKWBx8cuLmTqGTDJhvbSlfqUJhUdto/+wa7NlUsazsBnPLQ7i
jmIcsRwvwYNY/jZtXEldVF915c27cJ9KajUiKkz8Enq+1qfZSyNWCAahHDZSNiwY
3nXUrvZ8gPbs04QaOfZUofrFIxcfsuLLDOOW5YO+aCbGjHZYo/6H/eYwURTZ4nv5
dxUcxzvWyNweeCx1Nnt915GGWPqO9sHts127g9HtinVLGWAZm2Oz3YIL4MyY+MWM
a9SmNbCJcG9h5Xa/06MMe1t+A4XYa+EjpTFLgqLAAMaQPfJHx3EZXk1nOIyghx+J
K1HyoqfncRnf+XziSbpF5ZbaU6FUgw+ufFA1IVOg6VqP8kdqyL556B4FBG0oSMHB
SYWowplmniZMxct7S+t0d5Mqyc1veXYHh5qMtLFPV75tWm/uk0u0udd/aF5SUzTu
P3yIlk9TSChPVnfRMXlbUBeXDxaBFm3GnJG/qEvyfnNxKz/pacY+jhDf9sqnI0Mx
zsEkczYnO28jAAc99wz1J1z7ukC3iHIBi/TtARD0khx02LBs6PQC/rw6cTEhqqOB
K0/ePxi7ZAUhiwb+RjIsqvObNVubuC83Zn+42IquFjw=
`pragma protect end_protected
