`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
olXgIR+EAII7rTQbnJd2IrVFpx4KalcFg7m1cFiBxiwKqUBrms9aOkJEs4IKtTAa
n5l8DfzTUYisY4PKpdBE9fMHfOBOQp9bRnCJtzEFOgJdp5Por0yP2m8GmvvXcvnm
UkXXWx7DOS3MnHI3IiErqDqgJyrSCH9Kp5jwIV1/4kI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17360)
ytm5T1aZlDv9Jl8q/XwsFIbEifJSCp5MjOnCPQac8p0u5qUM8hct/BJ8HewLmxGI
ks5XBb3XoDA1+VHdTjZu8rX5zmn4glSr9MSWNWgpMqvfrD7smhx0EeE95prAoK55
4BNxhe29VLPxXgv06q70KNNOgaYqjrRAOyEDX06OvhJeVqOG4saGT+3jEr1h2yQW
xvUsNqychOm2xGdk5NJmdGpMKxd34RV8rpa5SYiCmZycYGgHzeAjZjZ9ggdymAJJ
k25AgBbfrZe8RX3ZecmO2CvlpevU87VZrk1a2wwUPVKkiCkesynRlMKJZJXzlXed
ITvsl/RrKs/VeF2sNrTDwTm4rc8iiEr0Tb4kI06u6xASOl8c0cgkc/5lrgxAGaAb
ibDbP+ewCkyzIblvGBXn1vt3BJWFrM+Yf/HmPMHMYY7B5qrR2FVAfFUx46h0qDMH
cl+RJ/K+vBU3H5hi8Oi9GAYQMumnUowcPwuouC6HXVwla4ECMxGVAN9K+PXzaO6i
0x6qJ4HJrsyVX6HWVl4vX5EeAIw4pCto1dNF+6eKgveOhfrbyrd+ZvvDzqgRVoKU
SgU81R2wYwSnlPTwsoB8PyACXjD4oEKNKjWV06EaGIMu6w+sSzobmiMvl6Wdif3r
5oMhoHK+xpozvHwpmv5rgwY4LvRdFiNitOd/Gbek2Rp0hrewQ2ZwXelLJNq1aQBQ
mbaxHZLkTmbdoeXo/5G/WnY4Z+rrZCAKqsYuacOocsTkE7Jg57is6Kd0d03hEX9U
4x5MqCATkK5JXaRLZIDxR1P3oaQcvhS83DwRo+1j5o0H3Gij/cqQrUD25db2IeRP
b0kWU76zt4VRJnh6qJOPd0NBaPw6iGX0zb6fI2lHnUw1hC/YDH6N/mPUsSWYrZDR
aGCfoxobdtR4uuBdylQx//1LlbGbHXd2kdIIZ3oHrq4ej2062mHV7ZUchoo6ya1u
bNpnyHPSpj7hb6M49P7AWT/8PHraaCktwWsSEbAMcBL7tQHuXorK7AQmfg7/g/yA
YcRlCkYO3iT4zv8Up2NGjJCAtQYc1YLhOo1aoFI4TacJfRbIvx5CABYg+vR4ahGC
MtDKZ1vb1rfyfUoD6G2EBCZATzQ/OIxie623heqzvK/aMGyjVSsq1Ck8arwKwNNH
gzbi/sgzPs14ip5SoCwxcWJkll8HiW+emYGckJsr9n/i6cTdme3So4p67Ktqyx6g
n32Malnvskt60reMfLx1yN9MAZ9B/0T7TOFsl66QPoReireWYHIypI0s01DOCyw4
iR1Dz2D7kRlhjI62Q9nIpgP5tlZY2egiMeEiCuh5tmlTK7BKgaPXTufa6hoYtC5a
vp0W6LeybOPu61kSOwZMEmfcPPDidOAqFGirzlcNXM4YUxVjuLCxyOZLfcHCCpEE
L+uBscUu4AbKT+gmvZ/30aqz8M+nSSzD5DeEKD3Lp4m4TtlJ1FiSkVc8qFniPcH7
z3TzM9LkX5ed7rfJwgNCveForq1VHaXPzFY5zgPif6bTL2jEY34kkvtXSFkrd2L5
NV5j8HUCJAV45aS05ZNZAx4AEWYm+v6o6ZKSlSnfXHQhZDPtjLaB8SUmcjnR2Mcg
ZMLAZwZjcKI4mTIuIBaLqCkCu8PBu+dbNludOeYZoMo36voX7coy9sud9e35s/7s
hp1WK3dtbLHKlYOBdwGxnL9G3orX/Xvc9mzU3iyc4jR1f1mw66i0Mlfdg+S0NP7J
ZYhjOhWBb2MUTdVRSsu3yLLk1dng5eVV7Pj8AWTPAtHVVWNowzBjTa/0sYTE0Y4I
MBqwTefborIVswFKuBC1vGfO7qZkQoGAT/Va8Zwz0KGb77Rfxw/4rXa/n9GVnNnW
R74ql4tNr6NXHlsC36Aha25O9HQF8CHXVlpYvh6dSoGU8n2p4PxrZBt3NF+H+eL/
d45r2J748yDpShmxQhocMZnOljB3HDbIPTHtMSBTdWtWorNFHeA8uN3O44ok80GN
/2LkZVycX4ShWrdxNv5veDg1yl84dKzGE5CZIYk3d6TO6tbOaTUXJkwiqS0kKf+W
QcflctTcs3f5r14nQDzEUJq0x2Cmel0cve30QROZWzuZqCfp/G/HWGtjuOUnm2LM
xKFgsfjBl4VpIT8HWeklUlEMjPZMcAJ1+IH6eoU8SKkrhKJvex8q70jaA34ktfa2
9eOcjQQIKhC3UdH8iUW+BeV4sR/dDq4xIYtEvsvvLYdwV3PqvBJexIDMnTGXrdNA
1Rb15L7cwRZrfMxQGGfyYfs+JsgpfQda0q1syhoNsT0d8web+guuBF/oez09rGHd
s/lutdJjaODzMmut3KIUCcdMLg/2wqSyqCTNPSpiKPigeNhHuj9AN7w9z43CtXi5
8AvOiG2boEZ48/7uEr/qQYmXcTPsP5I4BaAkn+U+xSX9qhUV4yKc3E3I1wAZqK6I
ej3PsrtV8RxU+LI4ftVdRhnOE4N0KMKVCaG5wNZtKWSQYFstBCg7h2mujecsDmnf
raN84VQJKRWZTJ4pyww6ZqSxgj0Frykrg1SakXLNNJ14BdElnSceba1DQZgFwlb5
/YHc6oWXyB54FP8QMy/+x+opyYxcgMcUfAHiySF+U+llbOkglb4GEaUq6lwDk8BX
iC7YbChDZYTcUmk56z+9VqNKgltunaHJ659gf9TwOalppcXuKDZRwD+b3J/QW2oB
th6SnbNKzqXKoAbK7KH58cQ0ZA1lrSEpt7zagOThNKUT7Z63rper73ShmwT0s/Pu
9fRzl8LTorrWE+H6D8UdDi1C8OtpEzpQTjbVlg1dBdbxXFNR2/CRT4D25mlYtPgk
PbiN46KGZqwX3yDRB6RvV9rBFs1cu19D795Rj+ITog2SbN101RAJu4Xibl+3I+8P
+BPI2RM039Q/upsBm30zuifC57zS4h1J8NkuP+o4QPv8Rfef6Cl9XCQibWRYs2a5
If+M7z9zLI/LjP9VaTJL+76gGx5lUYPU6FqKWr86KJNfk2lKdHko8DshVQCZxiph
5KwNRodZ4K159oaLEq3OnqUAUdygTb33kQOs9RnZ3eLqr/hxLqT8T9YrkOxBSfwG
8b4vQZ1aQDbU2RF1LJexhp2bQaEPbsTz4030SbvlA/IdTa7Q31owLW3+t8lUWx0L
vika+MpywgFJZMHA/xo1XIt99dMW4rx6wHJixpCYCJkebAN8Y7g0O8i/qcSXFWso
By8aQJ2NIUkDJpU3pduw9nigY2fCCjN0KrW1RC+41sj0byaS15AiW/RO9A5uIgr2
Hfvl11noPJ6vl+6TTMh7Nsg9SN1UyVTaxNWtRJ5B3DIabPikG2boMD6lsnQUZtoF
zFo6eUOZW1aCLfmGuwzauprgQsuU/nfO8biC6wDhEOfASbXIjFwxwSWJvFAnEYhr
PR9Wo0gllp0q5MVBP4k0OAZc2UdO3P/ms1DZm8tK2AiraJRoXGGeowabnMpiUw6P
/rAYwAY70B/UQXrSM5i/72Sn1m+xfycT8f8ilPic5OhQxgKomRtPgFEC4bHXYDLU
RJ750rb2HkFFPZZRiOWd4OSQtndxpB2rPvSe2MIKebNny4YavAnr3j7L3eKc4Tup
OfLWpNBHqoJevo+Og4Y0tMDLV6mBAoVwB0dffGLc1O0aNF/egIgcjVgWSS6hFVMn
4IQvD5RE+d7ibf8jEZo+LU33j5o1ssP8kA3BUY1q6XTB1dI3iEq5HIsIngQIhD8D
Heca5SjdYs7cMNXzawn9HEv3XQJ+C6j8scMst6JMfUzJZUSl+6Pi5tKSIPbGn8lM
lxj3Lhmain2xeVorifHUYlRQoJLBE980IzFedPqWd2OqFw3PcBwvWXPRgPd8Qc76
uT2M50oSyF5GQBNq8IljuAblXrpOWdI//EPZOG2o9EFKoGpuUTrVlpPvj8DyNLQ+
FB43qmeffbemIt21gUkbQ0IqC8i5zReO9NKn78wHrpNx9XZrijY125ut/n+1zpwX
A75uYICpGSR0Gxh0VsLWXqtWc09oF5xS+gnNQypJmJYxGuoN7V4aJx7jwYoAP2ap
Kl/RIFnl2dttJdwRXEZyDJ5eCzM2kGjtmkJ7RMHQ1jLrD8ZWGGDAGkQBRUQYjItr
fAR5a7c/OTiv2buBdRoikOSTtPfXn7ftb9Y00hC0ssEc/6V6giaqghznyYHv4L+t
59lY8c3kAaDXIshZdOeL84SI6AZ2CpcKe1mg8woTyiTYLVrDY+F25b5wyd+XdUKj
9CGsxOMm5IO+8b9qa4EyoeT2+612wSVAQgs0KyitfsCnszCLbymrdnfu5L3Tyl3s
OmVJRYucvKF4Wl1OuqixA900SVFtsah4u7fmtlyMb1dbFHdNF83GuvgwUay0B3/t
2XlZP9NvGVWWNfHSw8T6yffwNr8QuaIyGoJNe00K92yUKS0IWkwjBPU26FZD7qo5
nyqchabyFr9auqCxIK5zGSHRFPL/WYt6asxykKDo77n4MI4+VuvughwFgcubXpel
Xfi0lAUw6MKPt/jdKSRwtHmm3GdPdIvib0gEf5NXqc/Q47QI4ubY9O+zNfB+IqK9
uOcwPwdQDz63wMsXi+mjXWSBIHW3Uro9RKsk8kdqFhgv+cLF8X/Mq8nHr7q/F08m
C+Ayq5uxP1xygzGuw3P8pk9YV7Gn8bJ9ItV8mmM88yLeXicHt+0H6K99TNXUrEOT
Vp4ry47GzruaB+0CxDvP6IDhUBwQveYJJKzoHuPgmSEXArCdBt2lxL96Od92tJIl
+ofXKisBPXbUgPHh6w49nY/jEXQ5fNy0pRVdj3Py5AHSsAtw0GgiOWVuQq+eKBpC
zjQAklOg48BcXLkPOOhCTs15DhIs9/7yZTWNMYVeeQsI4IB9O1A+TAW091ZVUm7f
b8uomqkDWPHiFYyQ/OjvOr6FaWr7pvBqe0Xjz6DxV4u5SElUbF42iosPjW+RM2ie
hAH30fSkiBd70oPei24KpkS6/2D+ysQIuDR8AZMXCT96R1neb828gL9Pz1teXQ9t
d/Jx1w+RonrHLDzGshADp8wkZawgMDHD4ZtI6oIfXnQOcay8ce8jP2g1GQXdT2hI
cnZ1Mef8fcgo/L2I1yPVncp21YqYYREswDQg2pTidlyhX+ZlBeYUyguisrZxPA19
VcMS4uavVNyO+zy/Lq3M+ll8TlamFMJZ3SnLWPtNREEcLt3ZhpcOT3Ht5Tqp3wAS
25ZEioR7ipV6vvYSxv73zKU4DfXFDCX5BsKaKsy0QGUp2qSOv6qzk3R984zndKLM
Us+5CPHHzNS6S8Pn3AjGQ+W5V098hPhgrwBahy689h+POrRwg2+z00QedVJxeszC
ubOQ9MBA7e3J7f8aJ2HdThSSOfa81TST6bEXtlBatzv4ZnU2Ln+IKOtwp59h8K+S
5Wstlyqqfu9AALsPPf5lBnL93q4NAXPj1zf3gJYiQf3U7rLLivT2T6VWJjWAuFpO
FQA1dj2DW6KT1USA138v9wbywnOOKsvvCX5+Y/mVdFdt9yZ/ZROQAE4mFsdv1kGU
dLC663HjIvmnt30aCdjewJqTjzFAY1e0C1QsXx37BpS5bQ2jHgeJsXyNPyVmnRXZ
zDRoTm34Yb6a7v5VtQBxJMpzummASloD+jwIsPpBqKr8MDsl+BgYm6IbOAYgaHAF
mK89EFLwFcWw4jP8i6DIyQo3yHrBE67W8GAiPXWRv+hnRg7csdFZyf6ocvb6U8mP
o9+aErIm/u1/DG/iR98diGPnAVmrMwDiFtte2eYLJMjQYsCvhoGIlXE4DQBInNjs
JhCDLVuj/4hQ9vbe6XDMB3IWLz8E2W1HxJgRdW+Z0YGydOdR36sqPnn2KgtoYoeZ
WRFBlKZVM2dbnSX1UcxN3BfPBnbETH+WMvn7lAaLJ8W3QIZnj80Oht86KO+ikcoq
EYMOY0Rr2IeCYWZc5xR/WJLAvONAecLYRgIEHP1jabPeaNPGd6ndmdlGlIFVhgQR
oAKfPci5Tu+d57GQpUQLs8MRuKEYYRSPoR7oSrOrAcREU/1Y1l+q2xrj7C1pa8hT
5pFLeAA+WBnw6AhneRkwGvGdRfdvWpon2n/b5YcO6k7fdAtlBBgscY4TI0wbNp6P
nIWFn6oESF7WhqW1aJwrO9YFBDgy/CUR9VpTvF6v3JMVN2KKO1E18DUaeMAYcUM+
wr0LMU1DcqNznoQu2O9A55tE/Z/c5Hv42D2J8kxwreeS3ChqaaA/F9pSTsYD0usW
W71b/L/CSKLEIpE5NM9lphbl9A6NMF1wccBUaqnSRul/A75QUv7o+6vK96qmB6O6
udiZhqsnpCYzJYDxszMVeA8ySOw8INT5PqZ3jElkRgCugDUXuOwdcpXlEIcBz+ge
MHKeAoEU3aOCmSl1kR+owOnWuvf8IJ1/XApAEfiKyYAKnbja3QBvli2mUrXf41WT
yd93m300bD+jtS+ng0/plIkRGn9Lgc2QKs/Vwa4ttmzeuKAIU+kdxvSaXZ1JUjyX
puv48kx6FkGCU6F4PbLW/89Wgv1LWoxRqmJdCTSmIOfyfCdhR42QfsmioqO2+gd9
3zfEFg7n0NuSJyhMuxf5Y6rofs/3GyZIXKFk0HdcgjITNwW3Y8o6fi2lK1yQ/YGd
hfmTXj4P9mw66LOnhzSq9QoKtfSO0FSW+9lzxBWCV2NIqX0I9cVZFQR4EHL6uyp3
GeG1RcjGbL36iaWSrPUMmurlnwQiDgs10VzT50XNBs4Tw0OHXWScdTxwA7i+A+/4
vRfYFpOARAXmcNMfwI6lLKISYjmP3Yv6fa+0OAWjuskCGevmo/qPtjV4T4XLytWZ
AQpcS1dB3ZedfpJTd/lr+zBl0HFFi3Cbrp3egdP726ltFJhKloAkGPQj7J2S+Zvc
RSyJ/ajelQjJcUjivwvlSevMHxi6d3yt26frHLlC7bQ/vAi7x+tK16Kiga0H9BBX
UDRvuVce/x8dK8JW8EcC92IZkX45VZ5KzUGJWNWV5VSIEI0rZYXEtmcmp90s9Ksm
Od6UkchbhStGzNLUrto/leiTVUsgsEtjbsfHnU9JdVL+XYps28k7Pv+pLVjB0TZk
IwpD4QVCnn4RUhl3obclz/LkZwr7HJ9m6TA+2/M3ZV89LmPj5VP/ZVEj3klwqFsO
WjXs9LYifIDvHsexzg3sBkxVF7tuEj0Xfcp9aid8y742+UXxfy8frvAT2drILYVm
fSTJUnlCEOZbaGjp5saeMN64k07EStWp/6LhdL8tAbULSzagfTvvBDpZ4c4dsmPy
4f+DU6ic5ckiipx+X8zV2a99dwOYIEsOiz0vYZZeR8H1wVjtiB5Ci+7zbYwtV4/h
1OiQ/zobXX9nJjWI6U4njpQsd9t3EgRTdP8mhY/9EmLTo3RLYHhLRvQeznW1xPm9
QfXw61YcVR4FhDPIAAxbJ8wmRwTkneQwxpb5G+xMSXhGeIDG9CsmavHFqaD6dBTD
xmxBVH28vz6L0V/LGeLDlGqEgWzwU6m/RwrtoAKmMpbZStrsm9p6vY5lFv+sC1e1
NCxu6YtyBCaNrHBcc5WH4+dWZbBGfNz1jtK0KyBlODE030PxTfZH6mqDuQuFRArb
A/piID+A59WaZRuyKNJpzUSyDdK7s8FumYwdKm3fw1dWWpzVoMTVD/I0u0lIak8r
MfRNtSkGnqAZojzdP0vcFuur7srEaP2dREceBxz7shSO3p4JZMlaWxznodfy633P
I4q++JUA/FJHgSJEgT+Fn+MhAkBtSutW1rOFj9Cuc4M7cP665uD4FUCFajzB0nEZ
qydIF3FyxxSQgdqS/XvLe9+A2n2myDkDJITv1DKl+2EvwCMrsxLfGsKmH4iWp6Kt
UNKf7Tm7xUQnxxbzaZEsC6kNnncizV5yb/g8x1i2o/G+ShzHo85YTiMWm6ghlaeS
J9mW9gtAAj6jGMZPGNnkm+NKi+jrT6Ca9uLcmh39D5Ootvbrqy0u3QaQaCQIdL0D
H5v2u4Uv6KUdfDcUckFWQ/l/5vJ+0RaZXEkSxW2wVZwLBSpjRVxLCTqmrmX25SjS
NbjOICYTrBKlOrmLVzyxnrw7hrRKALqQu6Iwnor9fTjhmTiMHi0lDyI4O0qGQn1A
+mW6WAjdMFppH3tvcpYUiv4o72uoesmBgW0y5Og0hkRguelxgNe/wTAwSSdimqEo
5hTQYqrG0DNp7rOkxWH2zvL7rvuOe1+N5brY/cWf1reGTsWdJQrsaVNLmCLcP8uf
R0OU8CHyQeGyTwCdSluU9/jBBA+adUEc0dJT3YheUwzb/eosJLSBMXS+2YCtaUIt
jNSKFpJY0+oOSFhoalo6B4sN09jkyNbzeb0I5dW9aG4O4bQ/o+tZShbwhj068ERw
tSUWSOeUa8aozfgK/6pfQT9oKyX4WYl9DcPL5Tzh9j6tWGBA/ejJhKR/GkCZ2KyD
pfGwD66d4zlRYolgNHPTnXknT3vvhbKkegnxtxqc2AINmtn4AehIqAWI4wGhQEVC
jJ99kEgv167w9nYr2kyCsNp4SaAjzN4jz4noOJaAZxrMHgO6rfwbZwprkAdWUCU9
8+fzCQfUFGgLRJsOF0cRPmaJ3D0k6PFn5Sx3m4FyI/HhMPioXeQIhKZStlZnYs7U
mbbTnm4AQwga3aZMI1YLK5NE1aN/11cioBAdyrHGWyJrMcCk1ObyCqs5X9zkH2UM
iBm31R0RIGgBPn9d41k/xXIGvPOkE3HjrvfqaIl7YXN5PvmrfkOTEbzjJyXKazfr
6wCASEdNSULkHZL6hwzP8aSTetL4PvcFIOaPhLIOzldJNrGRRctwwVq6HVvpOfx3
f1jxuq15n7QHZLdtCsybb8VdYLEmTvKDDB4VQb37vI2+YBus/WpTEpfsnvzOQuYw
Va0W00lBk9A7qZztzMwaY+F4Sa0htRs2GWfsMEJicRHElRjHmfSZnzhMdhhi8Rak
9Rs8WA4tL0+WN1/Xv0EhvcaM1ldhOyTi90jZSKd/Itts/ly14Z+/OtP4EeYekpfo
XHBhXSV1Jhp8V9QNxKe458U4Kp6JdSly+i76bok+yxfSw88YgOdfpYjNjestlFRq
q8SlhmEmxIQdv9tgzjzgoIleZo+QhnsNr7Rxmaw6Te0r4iA0afUOr1TJPG1tgANx
CCjtLqiPHOdQuNWwnZT4semrhPaVIJUqw3nFqYS12UYI6Cv/7YooOGR6ooVy/9p4
T/V/Sm3687rCws3YRuUCmA2u4B8iqz5AQBK8WGjc7ILVslUoPhdB1hT8Ku1eU2lG
gnPMSEtAw9hX4Rm/nXWKZmnDzyUwHxNWbx3Zb4xSVCM/jPUZjKzz5a7G+yTZAnNJ
FojDXB7t1vKjvi7J2Ywo7AWoPhBJ4pEQHnmEhxEJdKsBkwEaG8y43cQmKJxv+x/c
97vgsrRxlb7nH2BbiG48ml22tu0kao1XpGMKoCubVTHlMY6OFrp/oHJf7fyuFVkk
LD/mugUa+aS5t6iNYcu03oq7j5CEHMPxPh/6jqqQgHp7+aiIvJebjX2j/A6gU7qx
fpzIfGWUGIfChB55+Hgn/XBI1B3cXwDQSK0FGPe1KCeBWfnYcaP969Y6edjDoy8q
xU2Y/Gp3Qs1NuLguWaEq+bI4Hlc220+gtCsZT9DsQHo9llcgacVTcyxyZlm27tpf
4CdiZsGZKa5MAezZwiORwFc6vDV4hN6L4D6GAZDe9qnhiBiIRrAG3tkNGIzgrm+T
pjF26P/3a62yiiXIA8G9lJmEZlGnf97pQ1lDiBjW1Yzv0QJanQQuYuZYrdH9rqCc
bGNPhyvyu8RuE3A5vqqBpa+HtNO7WjaDmq+ez+vgEZWxLqCVM9tF/cbOowD1a5rn
qRd9VqtAghfQb5U+hVbXbbzVrVoIQBmbqz4Ikh2mucnT8/wVtRWELnCoapID6yzr
nYFvX425WLgFakWc114QxSHF7+59oEE0/EkTgePUMGVMXNun2O3s5cL3kwHD6yl2
eAVjh9Jj28eevWfTvcmLGKmRzOlQBtqG4tX/o9ST8vBzpxv9Yg2FSGdp15YXHuxQ
9uSXc7Oux+4UlJsqEeQHcK7EwaTeozk9rrfr+TltX2KuNMPgrQ/AxI9gK0scZoGK
9vzM4+JXt9egLT3VkF9XPhgYsg8kNy8WkNv8rJpxUJ6YuUJY8RprA7VaEdPGkUTe
KNc8O1UkrCQ5FiNKlYTLVowzgx86shrtVMbjwB8ZoMMsnFnO2kgEi1r36RJSspkt
vcock3vAUfVQeViu/jBA+hNAoYpU+8NeVUh9b9bkBnnKc82qu4lDTogp0UXos60b
ekTWQBBZuBDjULX1OeKSm9+Ox+aQjKet8kIRcrVJeZiMlhf31sIICvPJvnE/D6T/
I7YfkfFqpnSXdS9P77OlfXbv7b4yJbVQm+YDeFQ8oLcJvnO1i1/aREuNgb7gPQKG
NTe5qqGskEpJ4RIaHN4bJ/njYygvQF5uojwbHMZxgD581WbpgpsvkvvTQHK5NXMk
hWEo5bSScK9AMDRwr7NocUCThwl+7BlRUV/Yz1tN0U8HAMD06q7eHEUgmBomAyji
qDSP7URYfVx8X7s6gaqmVVIw0OCktPJaIPTjMn8Hi0wiw8yrCJmlobAYvO0SuxED
6l2nUV5axGWwKLdzWpRzkutAgtZiAidlPArErOVBWh1JT+Ly6EMBKnA+hKy0O7Yf
i5BIMECCHe0LdGpm7Zwk7DnrVY24JLSw7Pg3YNzuC5jXxeyD74nAod1KCOe5YCAu
4jPu/p7OvE9gCtxBoyufc2zk05qRYuJPv0+LJJxoORjiEL6+SuGQ8H9rumX4k7ZK
GHrI2UpQP4LVE8iiaKk8H5+u5LjM10s67kEQTpwn8GEa4+NB1gEVPYfbmv7I0lB+
foEf91qkf34mVEKFhzomzOM7siqfPls8wkjJt+lWOkuL62RV/YF2PWa3uaRgfiBR
QcWlxTtXSOc/FwgL6CdKQaTGK0EkufFGlYct8LCAY3dbnfVS/qCbvKKydhif/BvY
6W0rBiew9BfoXMfsleiWW/x7iHuA81S4GJVENYWCabGgYGAKWKhqbOXep4gYbUa0
WOqqqHxVDFrqln8dm9BeX/GjjIivF2onGyzZIE4Fk1bdoMlln/pIclbx/Ou5ba9A
NB1EAOx50/DEcsbXgVPMSW3/3ip230smAfKDO8yZxepToSoNhU1fCm9UXtlhM47Z
aWPwlp5lLQNk/g6VLM1d+ZiKbMM3tC0jqMikvVr2D4K7k7GsO4TeKdZVIlD7PQP5
TmuJmv4auQP3Tl0e83SnZSFmiOqT18YuQNy1bSSodWwIeATDhLZqX7v4XBtPRS2V
1omQdY+vg6nt1Hw0ncbfXSVpYf4Gv8vPjdVcBdiRF5U5yljmUjHk4WNcxWIa4zHv
FgGeHZI7b/i+kU1tQJC5B8iJI1wrsFUCddKVY52DPs1CP0+YnaleUMyoU+Q8xaZm
L5Cph3N2G0lEvyDLGFpAjmfolOhC3cXQbJAKgZuLqJ9RgPKnkKqQ2toLQnUKgyjJ
+3JH4FOxcVmBSGvGOz9ayIAFtauqzMwyTo3lbAm2MVlpgGh+Z55UB+SSPgNKz6Ty
Eq/xJZWQYCHpvBylECrGBYdEf67wGHQv9J1lr2MWghpZv/90e6i7kFrg+b1jqq1Z
MSsGIY45rB/EECAP1Sdb+Vf5WEZTacX33QOZsfAO8Zy0Y2B8m71nlB2Qlup2uXK8
pjJihdEDl2Q+SDEyUwn/+UXdV/a9pa7wNYU/GhOMKiSxIZefbPVUHWge/jHyY0kq
zpQ0MJkIJ49ulpinu7FdILJsATmNL0y/YvYlXnUCN8OvebQK6Mtp7ZJPcqrKv2Bm
gwxizdFgPhsOLGG6dz4ipf6/1seuXQyB+oTSQcDZ40Omk1NF0USNNBDTNFs1vJZY
MlvU7P4r5cIxCyFY47W8eR7u+26IiVKZzHOz8NNQTQD8Xycosqs5su4WfsbzWsC8
um4uRZPu8mQtkk/GqprD7lOpBf5tuvoO3on+GDwE6e4dguHAHetUBkyhYHb0DYXR
a7rY+viLutq1uVhDRDS0lI+QtMMwjcuEDDw3RkDO4vgx8fHnxUKGkRqJqB+Hgih1
uevsPaf/4aQPxExjzLAB0oUXG2TgwQjMXxaLsBVdOErRhhMEs5j7i7sPj1CroXSD
rDBuOVRaUruVb6wbQIW/VLwjxg2ehsL5mo0B7dpHMWREMdeI5szNnFSrYA+FxHom
zJGfJOHcK8V+8fBh/9oWcjfnKasNSDiNaB+08UvcbNmAPFwxqPXK7NvM5tPfeLwk
XMhpOHcc+9ZkxslKGEDHC6zGm1dbaYNg2sV9YY0DGiZpOqmmGNrRHKahcZwBhNVQ
+HUIUKWb3p0K2UkKmXNZcSIBTVh9nn/cyqhbr2CrfhUvOsYHECJigQqOlKht/4o5
xOLuhATlgoLWqV2sM9kTC10vaVCVZNsVzqPWmk6ueD23RjWPinFDEbezohmNFiP6
GE3eydx7wsgQPiXaSbWaU+TtWuK6z/KzhBkNtRvr1Dx24G2K3FZ5/MStCzMmQP67
nToemqufnKjYjvDsSxu6ZznWUfvqQrTAQcuLi6jKl8reXfMQVsWY0z6DKq0W2Rat
V/XBnvqzXYEaaUbR0c66iC8GAZvxUudkE6rykWwBPDk0+9RkuDGyQxWB/Rx55wSF
57jsD9icuYwlAdjMijrbOOPjQECL8iXyxGguTpBiaYErKJN5eyACSCPXo6Pq1caN
nN3A0zIeCQefSHMfox3KPZmbwLb8DCKxXoRazeIX52Xnl0W4VCJLyqHNXCxZN4mC
9bd3hpGpXHXY3oqwvHlzEO6VPLC78PX4y2x3rV8JdvX1KhgVTiYaKho19qTGUhSL
iPhX99hZMW8H38dsHDz9TSe5aGbGxVUu5IJF7+pant2s5ikIcyXuI6EbevFH/a/3
CQvv/1DLXT5VaajHT2WRoMbm+vNmr9vIISDTUm58jz5jb8B+ljhPvG7+fI44Np2n
78bZGFUUBfpHZKg7D8fzeGpjZtXJOzfc0abSXfZG7GSxmurUVVicWEuuveglcoxx
BXWWxlHs84OSOeJWAo2ECrw2c2k92bRcUsUAWwtoVIzsewj5p+0yvmwnGR3EE4Ka
hxAzVtS8sLC2kiD6unqgGU/3KVvDO1UKLxacIa0JJKujlmGHNqc5Ir0G71LeC2el
vo5tTgg7jPV4zEt3Cjh/QkR+p8lmoaLDLBK7PiAe77mQNk1aUIV32NVPQ7R8Smce
RsIpoml73ur15huQ2sDtJ3XfZmeAej/R6nnkWlfkto7ZE8d9H/G9Ey9eK4ZQmdof
ki4XxXy4wn/3ObnZc9icdptsktQVXFmOnSjcSdQAlQROdeh5YurjgJoSCoIAxkRW
6ZV/3vn/StxrEE2w0rEGH4/M4HEEelNvA9XOBkL5bQ4nDNFfycrlA7nVFsikElaM
MAdZUwJHFRTq05XOXdxLoD8BVlwiyfHO1UUyze/S+Ijuguxsy1K2VkzAPNhG/qIw
vypCWPjQTDjEac+xtqQcLUTJa8O1ir9rjePhYpaScOpCteOtFjPO3c4yIe+4y9uL
VT+1I/tHUUklfCL3KepyiTEDfN5+0KjiJbxs+G0jaqyOVapjPpcxuQiJiH2TDKKv
GymoKWcCOMvBD71cHKhDG0wzpOCMj3pWmJOhLrB4/heHS9zxjz1GRhnTe9p25JnD
Bxu0GT1hNttqPO8ZIW2+8LDjh2H3hDghagQffr+yc0VVxo2dag9+wtIT3xvpId79
4MNx7BTBGEC5mwZZbhfNSDcMb+kBKYEbnafhbH32nj56T8cN/POzCBRuyb9YCsMm
swL31S3sekK2pgo4fN5TvI2bww3zJkob2OfmGG9yiwsx1BbbxfUjN2wvKvU0aJEw
tqIPDLy/bHgOsGC671tAT8xKlWPWtaafFJXfNIy82CLcDFZc0BuZgVSrsThvglZC
Bx0dKt2Vf5Q57cQk9Ua6rZ0eGwfFoxvrVWafHoCKO9QOQroVmulG0BeYpWbUGB4h
XBhKqcy8qRFU5HQ055Dsfr1xh1xAG4slw4fxc+RwCRW3KcRi4Zj/+xfQmtJ71qu0
j66jekodvs7ZrqBw8tKRc42xT7plISUs3D8+v/JtviQ/RJknqDVLiuwEOv+TZM+d
ZBez5c+oIZFW4ODetlzr8eZAFmwMrG+wMMsq9v65ZuvQ7nuaYAztS6u0kHEE9u9X
1Xf/mFoIRMbEw5gcnDlnnsaBvHUxsCmFB2p0i1eskZXPeel9Vce32lTQ2u3LbbtS
NkPasEpwM5lkQDRDS3EMKzCdW8bemOHn83F+aG7o1uBQ/yTaG4m7jkhIC5xvBlpO
+oh1+BZ1zKVx8jkyHziwgBzWQeRtrjP4a8szqt+uNWaA1RmLSAFhJdN308pRzGNj
8DLZyuU5Ulk/YY/9ATTaUXtADXYtyWMu4/ggyzfMmQ+tFny5ne80Z6mpBXwEZ0Co
yGPW4/g8nhGw7+1rxqQvH7E3mb0z8E5iZOcHje8T0GgvsVjK6L/I1pMrPm+9GbnG
ySI6sahX4KXhWWNX5KACRVWyaS5SlzlSQWwMhYRNQ+oFi1QhEhAn0Fjp5U7Iz0VJ
EEtKtN6I67LxM347aQfbf8OYwV5JmMCcg+k/yhlPX8WbjAopRTHB/aTdr1OXlQWv
DKJJuL2JbCT93aV+fHsK2T3g1vzcjpD3dRcO2ddqb6aRpzzoPjY3CbjlT7QZ8z23
ToGh345e3GawHjsNiZMTdqKxLVrMx7lQddLB+Ui6nUm6lVod1+sQJ6aiucxVpeSq
o5YKfb7dugyz5N02lV456JyqsYNOHPAZpzNSdBdoH2CtGrwG58fm8vcKIeZ4X8Yk
lgF0AdFnfr/c7a2+7cQeCT4De0LDWLjhMB/yTlVgWGhRmefBYPT3CYciZIfkAyO5
6C6dBxkhGeqEBEbPx5vkimxTFCg1DNrTl4Ws47FRKwzOcI2M9KfQ7FsOo/ndc+s8
vVOzaA7vkhxI+6RJsgXA8z/+zUOwLz0shOszExiqJLRZ55BhJUZEQx711tHTPrWl
gV7cTWkywZbXgcupid9EWhk7ZoksiQI9WkrTETiX3Qe67fQsl9hPuW4C6ILy1r6o
9HgjTThKPgO5vNq+CNAUl6UHnQihDBK+jMODh267VkI/uK02ghPjzvaz2LSZCzag
SiLBobV8uy9cOIteD+d8Li5k6LmtNVgaCp43i6SqHB0VdYy8S34rw/gYIfhpmzOV
U2nNvDlDhHVMcJ2T5nNrQDDl93W7P+lm31NTWopkn0F9srncRee3rUzJBiKDwAIf
ghs9EsaivpAbrmdVH20MSUColuzRlvCwZ+gEC9PhrTOv2PfaEDjUNnlAAhTrVOQY
uDovd1yx4kFR6u5i/UxXMZybo4zgqk2PD9di6c3WmuSngtnmUFPEs0gdV/q1wXoj
QfdID2UwwQAKGkjzKzy/A2q20lYMusTzwcZ1i266UijuZThT4wB3eEstG3p7nN80
FoZXtVxKKq2MKgKWd4zj54TypMtlsKyemBOzdhXdQWlMOnVtmDNe6BcYMRTQzn3x
oqYsAQjlCikME5oB6lJRaoLC71N/4wwUL+66tV1tZdjVjsprXMfZpxXhE5QwB2FD
2vuTz1mkyeTvQmvyIHxyxBxlnGqA6tpGNZWXzf1iQ3khc6XmIFP1Dfz1dLd6Se0M
5AjoG0+pHFK4caFTm6sjEqufzDRLgjScshDX+LBLw9lMFvVyjH5m+Q1hGTyfBPVo
kpW1fgPsLVYQSWl3NFd49SmxdJDV+90CzpdfxDfJQjAIw1cBzHB0IMQmTH7cMsYB
4Ct48m05ozaky+Q4UsESna6j+4Fdu1bGjPFFa3/KYr/laa4tZRdI+as8oUcHYhYI
V+nLfRtil/0tyfpKHGsOD67HB47Uf2e6uoR768U5/4VUHvUqaKCDDXQP5BL751m/
VgfxF5H96Lk+LM17i0znsx8nKG/KqYmMeTTdyJnm4H7hvvvw+ec7NVgyTyO8ihWR
6v7D7Ur21aqX1xyN3jpBdbQdWXPjgoZDY58Aa2MURsnj5nsm45T9wxU1FCGxLMZq
UfKSj3ZZGNhoCQwiKxdDtyR1yeU/XtOGBCekb35dt8sgIOwXLirrmX9dSqlPAS8e
Q81bA0uo5Tf0L+qTeKIOeV3PE/dt5nvguoE+xbP2AqaF3Upz/WPKHfxHeXABSx0/
BOMLibJZwoWJR0hpxnMA1EfYlwuPQlq3+W09ukO17xOyVVgZSAkH8J/D8ckKFSx6
OJ6EIO11GO5OdfaZBFv9TDtYvyDzKuYRdEl3ODNNcwH69UgiSkUnxuu0UsrVd1rP
vUDq/Si6zCiUeZL8mwRyT/u02+TMNTBJ7ZhcxdPNZD2vClMRlbbns8qnqB5+Ysxb
TKhnRa+xO4TyfRXRjIe2f1q0bpkvqqxTy5OgnPS5dS4AO3RZjg8QE7zpOHJVhDSq
jwC/B5dG0PvjNN8yi2g21/UnGOQxBZovN4h09igQvMvuDsTY0eriR3QcAkAcRqaV
LYlF6ZVeeHkMYAnimjptdPdmuBU9Uj99Wo/NBpGG3sbt7vm5IvdCoKFhwiCD0a/t
cNTszB2h1UdCNlNDs/Pl8Xhw/Y0aVtwPX0T35PNpPcLgEaAotLPHu2gEZbRYWIhM
3Fdt4ymG1titN7Efab7RRielfO2oBvcz0EgqPCiXYfbXKa7KNaMkBAxIP+fG9JC2
5xhmArhpl4tINXLNamCN6h+5Ps2f0JnWWEGzdo9H1nAR4Db9kP9wUZ0EOruoHwyl
PzOBfzX0XvKt1GgHyrvP1BPwxZWvdB0fO/gneZZKAMUUzq92W3nCjCefU/Wu2Quv
9J6ksYJFQpUezKiQxzV3S3tWsGrtGn/ArVIzU8d0vNVtGIE6J6NKGfRVo4o/jTyY
EhpgeiSNCCks0Jx/0XKRcObshLTsZICKOAhCkLd40KAuEYoNXFZPClNvkPn9LV2C
nmRWfwk+Tat5rhwTz/ka8pz4TDpFFCOZIH4DncWd9FydX2wj5tFjJvlvHAdnZBHm
X4NrkT6c7xZNESiQV6qZ15ozGkNVTDgd6+wByLH/Ia+FxzudTEk0hTrW2YAI0BAV
2BRhchx7Y5jx5MmCUj/xvtMgZDZ24u2gntZce07eukOXZPFLJ+u6R4AaSA/vnwC1
WCyaUYlviLi9nbjGqc3Ar3SCuq1B4OMBDobafz4lyTKRGhu/++RcUNkgQhVLE8Uh
emXHD22WC6hQwR24wlFNtJHKkbU1DAjhcgILR+vdLuZbM7FFDZ9mlKIBcYXVtoKS
aEhYpvZepEhNs27sYHsgFkwwsluHT45vEInOyI18CCr1JLG3AKiXd+LrLfQjol0o
K5EI6iePVinZ4h+8dY244cfySEATproxmekSO6wy6WCrEpSFvSxThNhw9E+R/p/b
XKac3m8Mxd7ARv/rKUGmoRyL4q5k2rYKOMY6ugbWucI05cDikqKSNC2ZGSv8AgaP
x5IDMj0sClI77fKuJR6elohwlZhbh3CqsrTe0EdDkggdtqiEwMl3pO3+yPoVjVn5
B/C34Uhpl02JS9TVVY2HRQxZbqGKSkgVzROlMYHysYSvHLJ9fvq9y3BWa9WwtUva
4YGlYzbcqrRUiU7UlIbyqBwXO3VlNCRK/FN27/x7swfjrBbY5/SaZ6yHvz0b4blO
m2eNlUz8UNftHtbuT+NwA04agveI0IfOQbv0hAtvB6L8RNPXxfP9ZOwsmZ0IA3x3
u1ZegRoFmsO3P+i4XxzTGFoEeZyIFzQN6sQoyMR71+SbcFlat1rGUVwMpo7coKNX
wspygjIxbBmFDgSZQJ7EH9rKxpGWYvDd42o7tAI6mw3D/adV1ULWSnyjiwWqxreZ
Zn31lF7QMNoj7aaKqvDrEqoCo5x3NLWtwRcFh5mr+3N9ZqfoEbrKO74MjUqcVRLt
FLa2R8OBG7LH6JiXgFhaup69sOxz3l0ryEzKD2FAmAv/E42SbckybD0j6/lMRVtn
H8jnTdFdaPG/OLpH2c4xcutW2lSbLc+M9zQUDl/qWbrwzzb+BN01vO1VRieJIzBu
Yi66oif7cidEzQErA+FHJ3LZWQCoL+9DqTFNhQi5xt+EckQ+AEq7yc4XVzsCi2dQ
9j5RxwkADJOcLg9DBXEXdNMSo5ymgWLvQ/50ClSbIJbxUSVFHq/f2Jz/N2CWhICP
jc/XUrwUD18z9bCbBiL+MRkXOTTLzBaAdk88wFnNZXjtdcds8FeJaU9cHmdjx6PY
HwWz+nMySOiY/E74nDHiF70RwdQwQoNCyTimlrYnImRB++qUr6zH7Ybdn7iA+poA
nesSAdEHTi7lsGRSIyvFJGUsg6b2Tq5HS2mQ24utjAnA3MJyyDRM6kAY2CTJqqdi
/Mo+7RbIW10J3/505MNXUw345fo7JZ6QtFJNoaBaeV7v72aXlMr0pTcKIGkGKMl9
JghYG6E4iS/JbT55XpGP7Ryyp1tLEAl9XWW0gukA0jfVlaO0+CZKnGh0LkQPlGXZ
T6xc6dkakDwY5JgxZ3ofS7YqE1RfZf2o/cVerNJ5E0qBYBRcwiHzbaXJwf72F2CQ
wyZdxSt1rMzRhxoHKHARWdDtAOOKtHsiUktgvAPvSLkjVL1z4dIt9hr+GY3QUeUv
Kn/JTP+pMr9V8s1WDZsgx9uC5Yg9rAutiJG8/3vNrvXpqx651HsGozV8rjMz3qll
AkA3pimaTgRSnTAbgaawk+DSZzI7F66zhjv/+BnCgpYJ541/G5cdxDc+1pgw9Gy7
fj6rYPVtGBG8nt80odayS8UNHxv5UBskoE4uIqM7iUSf8l952c6OZ2bMZJun8uQ0
3T66FHJWtADClyEwDfCqeBTV9QhX6y0FY34QuGo6EowzmPj1+xhiUbzBea+NpUeb
CPKSSI82M9y1slh1XVXlt+CHYikJmliS0EZGLgmKQlF2+tUXQelHp+gzNj1Yf3Ld
/BjroqbqolzPx2wD4zbnb2MW7ZahFBSOawZ2S2W3zskTvU2gnovAs+iF9+eMOSbS
IQIrBxd/x2UlLnelZjr27eppzpaeWd25lRA9HyDdtrAthj8sXBQJ1qeUzyhUMeqM
ajrcuLO8FDcl94sOV/uVF87hNiSBgALJ/5ZRVdRoYxhra8iiv/XCPDS5hYIidG2j
b5VoQU7UScRJRw4r7pIrWPmH6gUpwMs2Mob8LTVvyaKWwk1dnvHC+6DuyUSsxvxm
q8WPLe1PJwEVgdTK5v3WPSLdgZLNdIuutR04A9tiVVZIiH9Hh7jkG+UGjUmq8+kd
GVPA2Zo8Li5nn28FYKQEQXM1l74b+LA3r6T19Z/h+Ks4iJJJBE1IjyWtgqjx+y5Y
JpWCQuHcH9nWCH7BceHM1WhO8KbHlmCrMJwH5nsJCVhX1TXRZh7sPCQIkiN0IZ6e
g9IiNVvwZx731yFAEj4cHFtp7L4P66y+32Mgn1fJM+/GcxjUXTPJfizQdp92puDt
HxtmK0OgEUeDv6anq89Wuu3DMHkCD2UQpDpQ12ISUKDRP5UG5HF+h0y7SiG+Q58t
hz1IBfob8ZfSeppu9Rm7AGuiUL2L5AVmxD7Qsvg6R2ulpAXcdzQDEELuWCnJPAAP
vk9iHwpRMfpX/A78KoDiglQIQSEhlzxDAU65Iotf2WZuPOkqA+Q6vUmPRT2E5mo6
XSFPJ5tAJn9Z9++fzNjhT7yLA46VCiQ/v39Rht9PSsO+Qb+09g7ZxcrygaKhCAKC
8xKQiZ40EDEBsjyRuHeh3td9bUJYCu5ebJPWhyIFZRV5nZhp3KsqOkb4Jy9TmifD
WbaOTa/gAGXFNGWTDvOHhIUG25pYjwBsr+73peDGIRZHWFNmfCRTUfgIDCUr/XW7
SUvxcrsnpcBEpJ6OQ5WwMX9DYH9jlJ50y1rGMPoDtuv8FTgagRRPvkL+DtMFhdfv
XNI3Dd8jMa98HFmI7rEZ8htTTy8Z+w06ZAqqJfY9is9PU/Ou0AUEAN/ZtIIr8DIE
Anc9Ft4XSnHaUVvjPN0drMvJRbOown1FFBD3I3c42tmGuFTYFgR1AC1okS4vszfc
NqfWkAQvL7axjFwJ0sCOth2UcgSW1uFtSxTplFBfbMCd8h9jKbBrD9h88QN0abxl
guzXA3+WWti6UyNOdEeh43hlXXZIT+KI9Mh/hBWhtzfXuDvqivZNkH0uKwCrpGPM
Av6BAuKq8siDyBBNDzWNB56gSqIYNq6e/WUfgt1vBFGmsMgyeAgKJ8rfSLYb4Fhy
CjaXmF++y9pGAiWFvvvRw8up69+tkLd2TyIh4g8hXD8w/EQ9EEA4K+/NpRYsIfb1
9ejOOjs77Prv4shINZNtNVgUCPqKBFuPHfGgObpojHydFrgSVOBXue6x0p6wb44n
wT1jcxyGrNdLNdjAtDIN4WwVshFwZwb2XNWHTGbXEZn6msGXRwRir/zKOwiRn7yd
8Q57mwvMwDRO3T05uQE/Kbp+AvKHMbnrXtCTc2CE6S+hHFIHNsNINNTOY9mlWLuS
JTv7+zX72rp9LNbAxkEaWe+zhJxeA+fwU7Im5keQpavsQ5So4BFq4t9h9tcfjHLR
i/Gea/sxcwAPp/cF/8ShDKazN54Qmxa8WQtsSA5tYj3ONLme1N9pdV8Onv6MmIvM
bQhx6PhIAT8htYfPyabopeMgdm4ZaZ42XnoCIxWGLFp5ivXahe8miYRlepjdwHCn
dv/aZZMLJcnYO64GKGzWk6+cr5bdZTUbD7i/6oTkf9i59CDlB1y+VUL2n3AQ7eU7
9+/NEM8yAhzFyVMMMtOe+zUWzKL6tLB7BAIWz2L9tt1UUGkOD8D8XAzWPXh93/1o
FJTnbXe87OmeETrNseFqepk2xmTG7CgLqiqijMLp3YXhnQzt3hLYJlbcQnwdjp94
zTakYbPLid9yNMxCnKpcz0VG9nuLqVHuG0XQlCJDfba+/NGa+hnIrZrW8aTj0SAN
/anbhNo9eTTUepbxzAgdD8Smr1UKjy4wq6J6aFVPmtFBAHP3G6Z4spn32EYB8yGp
9vY6g3rI7IZFLEg1jg5TNSXa3nrwBla4TllQ2sNJ7QXQSEQDwjgHtu3vX4oourom
utJFEWE7+nUYuG94Q83kP8C7aOCsRoNOJsts0m8R5jegcHbND9ORakJvKi21iIAH
XStJa0YUt7hvXaPtin6EzFlihZ5tFnTu3fddlukv6VmpXwUdY1gEJdFIfhvb4NqN
D83bB9V0pWUB2x63YU/4r7AKlsVlIj/p+HjIivPiNtZ3JRnACTC45eRzrmlctwTH
r3h1I11RMK0PgDWU/HunIAW+xbHVYP++T7W3cktKG1AL/curKAqKdk7cnQ8T/LWA
kHll/P+vhCuZAvcsEaXLizBznjN6cG2UIiIFvLHIuGQyXVyXqwnGa6ipIeVE0p7L
BhaaLADqT+2uElTyKl1QjVPlrxw3q4Go77TAQoj1f5aYcWVgi+pZVUMwTrRRT016
VWLkOJ01pdxdyhQw9Hp+r+AmTLJvpRwUWQkazh/z6sVB2z94nLBaVmHfnCsClmZm
2dqxljIeW6lf4FUgtULoH5v+J1lJph0fviRMoXC39E7o9P2qsYyUwdEGkGpCa5yq
EU2B0kn/yOCKoWC5NXGoEXP4dG8CDL1W6VE/Rz/gSRrGmIhEPFkl1GgtOU4Zl374
GJTNeTwYTdwPK1IXhYUimzTE8OQdqPfLrE4/wsq8oHHIVE1N7lFjjFg4/DZEq4WX
ucN5qB1CWCVcdi//ScGv3OWQO40MpuO2OWSgDr9/Ap9oB/eJOZrC1pPqy+uaew8E
N8TlHO0wgcxVFEDJOHJKc6hkXMU7zS1bagtwCrEFwK5q3kEc/qs4djBgYWkA+toT
3/CWP5Wgq1M7vs/nDANhNeEVQg0vXud5S9d3OUCOGDxcB32x0Uqz90U2vqOi3AwU
YDKBKbMUMH2e1qXEuEvrtvOeEMsU1eGSaL1JuVc/QpgPzZPqsfH2yD0puJxuqgN/
4xEiV9tJ8ECscbIEy3aaoYM0Ffn4Z9fvPrBMLrfDoA0QGX6hnvc+VVCamzrfKvWY
2WUXDzZt232qWkPlC1A0UcbEO/Ng+pQ3MdwBaEUN1EDY9ZTvAA3d+p5mUhJ39rlZ
5KKL0kaej0tU1sNpu6EsOjr6yyF78HqdJ2twXO8KBK2cVTN/qqlnjcQhjl/wBfgz
BKCFsJ+bxiRBwhSkZ84OD7W4H6ZMaFTO2BL3o7Dt18IzYpOsgSO1NCJgO5DloSkc
BmRWjSDkXNz7TQnpR9hK2MFPg7D+zBpXsfg7Ity45HSdUgV0COAlGLjt3eqO1Yxd
2w71a5YodAeW/YXhyz+cpUqt8FNak1fAsGZjL1eWmXcg3igU3cHUTWE1l7KySDp0
3saqaq0ZE7SwV4VKHmKtS2YPOQp8WRLmpHFcXqE8haCyUhJgV5keLsVHdtb48GUw
6VRkSTV8BYkjLcINOqAccttX/Dk2pClmeMZBaP49OjDHhF3tSKsGMJzvDUgWCB+5
oKBRlSrxuEBmhnaOWotvsB1qBqz6t83bI0gLdWYWewWUygD933KIk/JZZNIU1wLc
jvWz1iXUfw2jUmH2K6U3HRQlzHCNCyD6v2h3RVqgnxWpzIcJ/WRC9GoEert25ne5
7tNkS4nbK5zIzpsJOFaQbVxciwgVS0S0coHcNtoA8ns/68p8D4xt4ozyUqoIFbJt
rVpOrQxJtIUZY+zieb7ZGKWCegcB8ULYOnuhMoZt3ae92Njg6npJK0yxL2AYbh85
35I1myspW3igkoHq9YmDeKU0hrPfoIgZkG58kLv1+dTUMysndT6ZMUV+nQjdwMyh
7Alz3Y/CmoHLfKEP5DtnV8aUK24hDjpCuzJZCeF429PuN8r4oJg6o0JroBXLxtsO
2WPC24pyYLbFOKRh3oQ4ZI3TZl3kWisnFP36vbbMH6ysrMpZX85lnVmITxWXMwAM
A/Y6lzEjLUIK83PkH0kdrfB+PwM4g02ofyoGZt8qAa9y/CvCLfqZr+k/Q+FD2kEz
noLOMZzUXg/gOqPLT0rULEoigFIuEE5Ht05u5aaNZEbozXSK3dzIfnWkD5/HXuB8
ZEQ5K3GSXc2xpN7/EqXZaIq+HK6ArzEXQKlqG7VdQSdz6LXxd8Bj/bTDrDafSC0q
4dATQHx+zUe4AiTkCshzpv2LDxQXNkLPdjflxWlD9iBpUV+0e1nKXxJH2naZxIb5
4Sfkk6f16TNYggEB4a0NlyEFyboqpYOkBd9kf6HVXEc=
`pragma protect end_protected
