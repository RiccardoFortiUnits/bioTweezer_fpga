// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
dlZooWXSz6hYpYVgP4T8gOvJWk1t61czugwBgsJg+VR6FgsBB9tiy4P9JM9lV+h4VoJgsmmUp29I
CxJTgcR9VHDOr99fgixweA/xIevvM2hF8B+KO27oc3F69VtkWb8p82gDLUDrVdjG0eeueJw0f4FG
uIPDmkl649ajKtIKG7F+6CtZkoizRVPvmzGF3GPZUpA6WUD1WDoMGPX+y2o+eFcfZBW+3NHE+/hz
gce24Sh2YwI/T2tCysDhmCv0i35oKtnPMMDngI6slx4tBguaM6Q41OSiyzCzebAewTriIeTQ5And
9rIK7PXYj9wSqprvNsCiJ3ET54KfBion1HOeqg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17280)
VU2nP8nlv0uYHy6RfoG4KVW6nsOyOQuVZIc6o7gpM3DBO6TQxCaVj6/+Su05RCIs8+acDCbwgaI4
KrFgelC3F3vqyERmAsya5ZATjflvQ6okU6O7FJfpiwN1YGoxc5UHwAYCK4H9z0jteQ1PFA1aGppg
13EHByNUBeDc8eI0Wztsn+Uzpss3JxxzSB3spPPXvNrqhFQYwIZ9IPApJN0L/C15gQXmqeV70D9Y
8aXUMCbTdxMLtZmnS2s7+e6dJ70Z97jgKeTIiGHEL6278jGkl/xoDE88dUMAbJBIfkzA7fq5TXUp
2MCI48pQ3wf6O3KXDxCaJI+/oypP8sozPicjeGCgU5mrQgglSS+XjbKOSl8sLA5ctZkzUpqTNsth
efOJ+m/TTe4t2MMQUmJafzpmkfTVhktuYIkshojwDWj78LxZ9pBIJtgNv/L/z9bvONRy8AJJel59
eyEdVTIMizeFy0m2gQYCrZW3UZOFW39KImtmUwkLltgi75BmUw/7ytYkDMcXxMTcSC4FPqB28Y2A
aBHEKqaP7Bmr28UmL6uMf7/VFkPtswDxoo6ZdTjlTHUOuWNIe0lYlvXmlvTiWD2UPQ+TG43Z7ZQE
6intJvUpqlET/ZTEY4/RbujGbMfZTKLHLpQ7wdQikXA9i4SOHvkXeYKKyLsZ2Th/2V72IjuVhmHM
UIHdoo4OdfIsA3zgEeiw6ENIXsJlvC0GIHtE6s/c55k2o1cFphP6WcRXB8bGAt4D3ggU0M/44ngJ
0tktT1LZFtqkOHW1g1eLul/crksBS51GayjKh7JIb4yMyC+TZ1pRyODXOhNGEB/0GMBj/jnC0DSG
1hVAOOXltNCmMLw7PJiR659ZXe6nlPSzR6vb00gQbPYvIrCmGdJVDN/DRKRD8wDtJzHSU7tt6skk
pJcLwKs0N1KfsLbtbvvlg52Zu7cJXoQnI8/UAHR85WKCauJNeXpXMieXBjVvvZS7zcWBZ372fbJ/
Y6kJwlGD2DM42Sd3HSwqcAJzcQmDLEYB+C0A+TDErxxpRQyz8npaMibUTFsJatS5cs+vU8ZBZkVJ
8qGHu1ux8Kt5wJ/eivguvQh3miidSgqO6fPvf3lKO5jCO2EudQJTAC7IFh+aG2kWlE4/XF5HwJYf
NXYExqhaB/pSzHP2RJVTV9lQmsxXwf4LP3tSs7bF0Ide8MMmOXTeGY4usYrULLarmJwlTvHnLjGz
nvweiXvtIYQO/V3GbtuXM49GwuaBLa9yDj7uW+ky7XXLbrkM+HccQaJ8/JhYWc9BcwC/GZ7LFY97
3+MMhQ7tkZw3G+ICHmgGv2Sed+fIU2DlG3NCGdGwF9tRuabpI7HhdEsgv0nEH71IAT9RZWHMR6CV
CxmuNlTW5SRzTTBb70lL4794HuigB+n8IGukZ9Fyit4qy3X2vk3x3yhy60DUzJW5GAr0EW18My4Q
bsrs0KQtEIuSYIAo+3bZvNL1qOIA3B5OWbI8qUmHUhYUb9PUsoQEYVU/Cl5gTAH+RlFz3fdZeU/3
ApFPBoM1ZB+e58PYb8+b1Qmi2ft0uEPNKzf6QmvSV3rkPgjmLgw8zDR3BD/2q0Rt72Zn/Lrmhtcf
IjzZpZREo6EPjBzVOs1a61NTgNN1FVHNXYmfgjAUZcy1tGgfLylrEedwv9YSKxzaLJc5cpvysR1P
tFzi2ipAjXlNQUJrxm50VjN3+q/pckHfjqHou/QSrvHQKDA+TTUJABEtivAwN9oNwVYM5+OjASTu
4yqPh9jqmIL6YsM5KPXfhn0T9ga0x06xGhkSXDlKNpbrt9O5WG+7MZKiWeioAv1f6Vx1TXhzqdqN
2E4NsCRptpRSq6rWxYOjb/x7PAHFIXvg4iH3d/x1RXVE8rUx69B2Q1ASnCQTe4ygfQhcJDh3s5El
3LDi1zHL6l1FSHnpI/FgmnE1vAQXxr51EwGBG0a7vun1QapnoXU1Anxz3MuM/tSSpQ/Qv/ecRgcy
I18aiWx9MrmYLl6RIX3Wyl6Qfnh1sk7UxHkLk37htGRPVYhHAnTCthH4HcJlXbkQXdVhD0dIb9mU
jYVkDRPPUEIf6tNHioLiaaSMeMuGiCd2Y2SbS/GF2kEtevdeJulMOHZAVb06N1siA7yY04fd3ct2
zmP9iwmbCdAvYmh6eK1YdLiwF51OlrmnW32I7nF73CkNnYpWwNEIu7VNkbhLEJ2fPcoizlzNnikk
NpwFr0rzLuYfkEkjINZUx4kboRo9tiQ9qYosJqv1yz3zFXWWI+f/5Aaoa3mS1SPkjrLyyStmqUfj
H/0yLqAM31kbt67wqJTcaBNe3D68UjPBmX6CY4fK5fjB9pMge1KXkClldphGtuCIvci5WABXiaUJ
9eALkPmDvnDl1DLL3DcP7jZxKGM7rfN4mCXm6z13HoVw6JZx4mjzw097W9A+nErBKEaRyJDxzo2H
Onhj/3apbopEJLY2623AEkncrtSqC3gFJSIIao0UC1l8jFhLq+eOz3UvaD/d35GhD/6EyKQv0BuE
KCcTDWCE1TNyMGcN2iqBCj8oQ46mZ/jRHFo8sSXswzTI9kbQkxPkfUmg3hhixt48iqqeRXDsDvDW
9NH6TLxPXjTg0OAM4Rp+z+HgpblUcZZdxN1J0u13Eg9mfEfU1JRMRhDqs5yFcPCzntaVtypQDMDx
XLvqajDeoHZVBtKqke5xr9i6+aQwnFRy1C5t/ycipa7HwpksS5DjVGSKAynCeucpSOIGQR706d2T
8DgSaFBe23ezLgTLT9qY1hzpg2SDe3U3jwmSlE9tdlGKF/aJ3L4wfUuqhTmhJWhlf3IU0p7K8doq
WUrGs/5y2tgkaErRM7qVF5MZh7gcReAVJ1AZbf/9RVzCUD7lThp233hHguW61OXaeiUFd27P7/ns
FF68wIscx41gibakbkup/2PxxXIaVmJo+CCFS7eVn3W4kO35Uf8FAD/yYbVOEyyCd391VYzjxa56
/qT7ZyubAewgiXanptOUzC39JT8dsKI82FvmELmLFJITMLOtWRoSR63TfSqe2UCIs8jeMc2vTyvX
9XeIIKVkAoG7T1tHTHxVNurrjk6yOIgh1DajiDOMPDuRpUbBGOrrDhzTax4iVXb/Q9MJ5w2LuUGa
sutNeeYqj/fPsoST+FQ53ISOGOBtdT2U5srYs8KSPw0CZymj0QmKr9eqP/6L9TOR0FsqPWWueinC
QgIzugkSBXrtBfIzhwlgyLJH7FKR2jXX6BW2EhpF7jSxPkR921bfUEEL+xXMSX1PrC/QJOVvmH7w
QYmqwwLTzyXOeSd9+l49x4KT50GgKScepJJmOZ+455pln0H0L1zTkAOmAM9T3tETgPVxVvh8O6DB
ShmWow6W0yWm1onx9trpTzuHVSnwWXTQTsqYvW+ZwbfMqfXv9oavsXe3gyE7VlXOAnrTZTvtZobN
b1ey2w47IWw/NBexiyoWE6foyYh0qwBwUy0fbxQWzAZwriPyfQ/WyGE0ksrru9e5EyJRjqN1DkSq
n6rcYmv6bDnF8cmo17rRbTgkEq4ZzYJKB5Ew4VyK2F5WU3ccaFiUe+fYJ/lQ1WociBaaOSyM5hVl
Q4Hwqg4jVhXf4sH6MnbeP92WywTF0FZRrL4r3cEM7QgjxSpmCrKa2NPdXBJwOex4AxdOMCtsm1aO
pE2KoOWsMmQZ6GAMYPA1BnSLSfnB6rK7DE5DvBm0k4TJ/EvqZgD2YxqzCvEFRsMpwu3wZb7L+UPI
Wj2anMpYuCeacscl5DrUC8JGTYXwSbecWu7qJuIjXnEC0OAEqPFQifGGxqhmbnj4bTcMrzif8Y9a
nX+QfjV4E6KfIO9CW0YiUUYgfVNgQTvyGLs4Mlcb049pkFhsP5CIk7vZTbao8401eR0SuKAF7zEf
Xp5+gah6JJx14aMvD7O1jhjkkQ9ZhWKqa6e1A5V3EqDQ0SvQ4D5bbmS4DsD+/WQNKOT0xj26mPgt
YQVZ2/RIf3jzddL+tUR4n9zAgdlTo/5vHYgwYiCxqayDaecqced7CmOFgJxCTJiddUbNg3zq7E/T
lxdnKbIH/gAB4mxaD7FOuaRveAu3BLu5PwCdFlPwV4BJ5o8P63/GCh8WjfnR20JClyEzFQ/1Qx/o
tXwu4rtx9udnNnKBoKlTU1uXNVyJKYfpDiDIRSBVzczieFKVxE/c519JCEvNDBthrsB0OLQ9ykiw
/m56nR+Y1EH0ncg/07wTbm26L4BgLi4pzV8BPfNrKhMhTCq3t+meC9DJEVABeYReJ2GaH3a/P6yA
y0Yx9PCtPh02fEBLYBb8drkNLEY3KMIT2hhjahjmpBwr+oUlSP1JUHt8JrF1UqMHM6vSdQjsqJps
vtoWjbnTWc25EiX95OCmkw5/F+ny81Akv7but7Uw0tLtrSrVYxl5s92nxcCeTjklRK/TIKe47Fna
3t2MFqWaFVPR+npxkOXDPHChZBv5ibFSjT47GT/viKdspkI77wqnEAuCkDtsZyTDkiq6kqtVcxTE
TYgLK3UcErUmMKonLxZcgT+kBXCGKI0IXT15TT8lMfK+RFO3WuXyBg2E6fD7SrfZRy7HtHO5PSt8
wjhX1eDxJclvAa1Se9ZMoa87kEWXiEu5PGYPO4oPsC0YC8qV598QeusBWW/V0s45gkSVF+B9DhfM
w3mO+C7LNxsAiHFCssaIEEUtn6dhyD2D/6XD74n7sS1zJAcdlrsgCU81388LcgmoPz8CBNYO15PP
s+BE/AeOLyH83pCMo6cSO1DXmd8wqYBMR/ByIsA9XfQgfnaGV6tR9KdiLkyzzBKM4MjM16aFCFvp
/I/BszqHGPJYlNLh3/612hN1isuXm8/xVqiC6EQF6U7E3+oqBN2pwkaYN/aceDYAhrbmEUPgyaYA
pgkPbqWs7JeiqHp3YqfK8SB+ULPXbh5slWORZOM8oemaSlFECPlspfg6YSxmhZjAu/h7dxMdbNID
U80ja74+LUnjECZT9GY/4C0dDcaPUeDvljwFUPPQvfusp2lUF5dwST0FdCryU/KtdYOGLzX2gOwa
c6eHfk39iQ6tPrpnEDDnP3ebs3YA6Sr8xSB6o1pmKUpMPt0TaxxA1FPftD18VAKUNXsIUw4y0Hqq
EToy29mgweeGxjeoufinZfjAnpAmJ2KNbAm2khCLTduMmkOt8bz2i4Go4VJboBlyqnXzKKkQEbX8
qKeMdOW/nPRgirapdYximUW8HnWbrZ0Na+E9ooBZG6kNxKgm3EofBKdd1R6EeK/JfOiHTmPu0gNh
pBCWjV96LZ5Rt6fjDICR6AIQF5JreFV68fNiWbxnVvU712c3AeBkcijgz+2kb27oRq7tURwffjJJ
TAjOl91ZgbDZr+/XZ2DWMspQ8UMdiy9LCoRIcp/iYdQI7OxOFmDxP5/5alCYOpgTL8tqon7PaO7/
YcWbS0WuHALY/tVXaVZMuFKVydxYVVM0ZUt6TIxCDjRKdzX+pdNmMyUbTIn/T8WmgkMhD2dG8kXt
lEGAKBR0olJGXUh+STab4xRAZHUVN6jy3MR81hb2Cqe7sIuJLq/vsqiWZhNIJ0ho1ttGOb8+jwo1
ARmlALOy5ojntYdf3REaUPPhUyu257vZe2LTMya4Xjcef5NBBPBgHmT0K36gGsPNioj6G0F98907
Pw/SocQblcPdr3UYArn5vHmYTdbleJMm7fUaSLPrRJdhvOlmLRlPfWfkj/Oc95NTau8c3IPuWFJv
FE++FiFady6EVPgRFgetV9vLa9BOGWm21+zzIMFOH2/8435CUGCDcwjfYe/ReKwQVhxN74VTuslh
qfeizsAWMeKR6yq9MWmKTvEwb1RWid3YVwSXqu3G4HJSaujPFFannb9GZoWMGs/6L1jaNxJdPsQ1
9/+jk6lwS6oDfuq6H6iZgaGmKklF7HiNRhpdyUmPRVAjqYMpBVK2uMUkYqTlrC9J/5tzisH2/TVe
nbGGLLM0ih+p0CRQtAybcxrQd4Ze6nhHNGLYSYAhI5FigS+pYU6iq4dp9xjUnSwxmxlA3Dc7mjPl
138kr/3gPsj3jkCanPXmKd0LKnXlO+IA6C2eiE+FEtVMeLqpWw/qRwxDRKTF2uNvrg09ijxXjlgk
0/JAWYuxE9uHjSfbcs+mFcnQhVhsa3MokklJlwnYpqySaoKkWi3rV/jHn2De2O8EgjjH/PksSm3P
54J9/KArjtsGYIjLr3vmW1Rh0xNaux89Z6I+dhSgdxMshh8I59Gj/rEJMGb9jkWwkxjyWqwDF9Sp
unM9emxdVzCZOFP0HKYA8bp5gSL2uu6/5wLt7CmEu8J+68KqyrJP6thag+BwNtle+nyMEk3M04un
o0VlJqdz6tdOQaldFGOOmWu1W907mdHpsJW4KppU5SXJndpZOhv1mOVUvT5O9bMfulDPq2+T/A2S
TgcM7gyLZ+oWTATUeDFtcNqwYE565HQ1/15DAiGd487Csy6xozWVg7B5PNAImjeSOpdUGNO6ifWb
JVKwRso4t/t8sLP5asegfRX8lPJW+dCf0NRVPM4zR4QISyMS3JEvmu+J4WTyrg98Pv3zRV9j6fYZ
xwmTByC5V8/ieI7f+EHjLdtRoOLv5LQr6VHyZlGv5Em0P8hGNkKQxEUxyIWtVwvEc+fROkL/NIbX
n/hniOkuudaNXqznqZKRmFRw/g2cXUsO6FPheSnXtsKwWXPUGKRQjfc/AnZMT3TxqXf6Pi4TBwnX
oVM5/tCib1+LmlU1dq58ygGQE589M1NSIYNA/x/jiiCT1kXIU9ZgdbyFHvrtWTI6/xP4P6H9IfAu
mluYGP7Xk3kdxgJyIhmExy4ZJuKOAR5bYKzTtLU9vO/5VO7LkHql8N+9jrIgHC7YYuCPracuQFU5
6+xbc86hTfnUDIU4qeEp00YcBFhfJLeKMLyiTdg5wGov1VnrXRcnMlvwSSurebQ0J3qZCNN1a+FT
EJRBpMmVno8TS8KaYaomlDAYXXy788Xqc2E1iUNepzK7K83D5Sr7rWW9ilrVkAK90esvJwmZ64Im
KIXecN0hbqslu4jVzLHiuP34e48JkfcwchCaIOnRIYyIVS24FU12EmsFajipVPY4N+emIG75G5DB
w8gBlPBLn0u5DY62On7sSjey/kQ0l2etv8IJQZxYrIxqE/43iR7+HR/PB4b0xxjPWdIej0PWDmdV
s9hG2M6iIHlnC0tKK8nIvgUUD1HIyeVRs+SwLmQv7alpCaQTaFVw/xxiPTjQjzmJmsWDrGHX2X4F
Abx66ENunJD4L9c0EBieNn7nGdN9XxeUWgFQ6TlOeFL0eN4Ty06SDh7AY6kEIN1iOEOH5JDEOzpY
XfPGc1WROcF0cIJYbrGYvDPyXYlsFdzidV0G9OsY5MxAhBNr13bW0RcpmiW3G4QfCD3xnYXAsIgF
bAli3Ll9TS8LyYlQQKbX2NmWd60UcFHW5dTir4pz7nGBZxme6lCduDi6eZpWggzyMAEVd9fhWQJw
OGZ/yDSwmG4o+GBB9iN/uAZUYXhw+Y80gHTsDI1iFV2OSc0GOv1ranpOUApoHeQtg6hl1x4xzjWZ
T2FjxkUamQvyGZyaJjahfj4Fz1XlUq7IkmboIEq0+loweSreDwCRwc7gVhc6C2ihpi9Sj8h3NT6K
Vamogm74sDouAeY/+XfNasEj46TwYh7ikpGKO3TpwX4kzgvc1+AhrmT7RKemlSHK7vlxRkJQj+az
la+vlmN/12n7AwlLGVoehvw5R3gC0A1KvzXwh7WWkKwRC8ZmnCwNyof6VjBaRHtiGdkcu9ifNtnv
jq8na9Z5uqYHxshJf9L5FY3SlIe4YCByBaH9WH5DWms++AhSg6CQsK5UPBpsOeb0P9OanuSBPAx6
WuksND6DkmfU4hvNlBz3SxWpJQU5LdKYSXVJMoYFJ0cyIfj+7q6wajd6sPA9OkUSA458mDkrPxq/
SW00AjAux4bDf5eEjOMw6IRqgKLhfD205qr5p/HZ6YFbrJAxv7YqIaf1mN5Pu0h4s9uzBdrAYhNY
FnigRDQII4xZSi/T/uxkjW5y0x0NcFz0UpVJq2sFjTcValVLpp20jGghnL8agxxTbFwlUvZFdGa+
OpkCg7FBZATjTXsx6yId1UPU2LjOrH6PWRsSd80PtLxJ8v/no7XerFqRrVpaSMQ3KlDK+C530umT
mEdzeZwrGvmlaTbb4sJWLgu3m+wLJBNoVgHfyoyDQ7UTQ1P0nA8cgeRMYFaXgX9Sj8FY2MSklvrO
r51kRmH6aV8JcEvp6ZLzSbHz6jgqeJreWvsmKhEliH+aNy5a87PynX1JXNmkB9OEeZ0/64Wqjgvx
VTK23jYKjI61P0VgXhV4x5BAIMMRPQzrH8lu0naw36rdus2uiRMonJcX8fYd3EBErx0pW0AB6kqF
/+KIpQlJziC2O+ReneLDvhkx3O6RQnGD7+uv02Lq9l0ncO/dpz6Tk4jdUiMUVdWvSqVN217PK98z
Do/LvD4VeZG9VoYGMdnGFyTJwJaT7Js9qVhlxxfYtRXORRlYCpC0NK/z+kLUSlChC0KoSBgC5EPA
dS+qhNL25TnzqJlPwkocny4U8MWd9Ht8qkfrM07I4l6FsUNW7/IaA/XL3+89RZ5bKEB4i9GemgNc
wbykhXfiJGnRuGBco/f3JBCDU/sy6d/h5yRR/nTn2Sq3cq9+PsNia8rR0l5A1alVzBGyEPF7UjMf
AxViqII5RC8lrGQdRhWa/noMTolKzmjRANLmTvatjRTxbg2EQoPLH6BOtGGQEGcoyxchxyVmt1wV
4qufgQlUR7dOzYKfNYWn981w9MUTqPnuHGNCA0sHO1aX9xaloZ3loMGKj/NuRpwnY2OvOyDrJQ4A
n6h7RPWNiMhcZ/bt3zRrLEz6vswWQLSWTikZ5KC9P0gibQ7/Zn3LSfz1PQwvLhuhhcV3x1l8pBIu
oo49VPKJfYwkSfm3AhLoX/xeGt2CUSXQkx/6mbYwC3nPTsJnXQISDT5/dijevVzMVzZX6qHBRvPD
Mlq+vdB3bTT1LzOqxNCvyzoLxTHFH0ZakYS75fWRveM9OZBmXGib8FrYacFoTp1RctHxc1c4S0Rs
e5f8I4bVv2cdSFnn6RiIrj3IJYfRL4uleFJLYhoBY12n+RAfnUrU9xy/ELJEX3PvwwmfhPSffrwD
bC4CnbPKDpgsNKPMctNaqypTfu4ueCK12lfWeOaL9MlbvLJz+5n5cR1C4GE6uPb/+OOlhHLSIkog
y7oFhhcjtAz1yKDN/B3w/EPJD9CsYjEH0PNsJsOkmhcJiEOxbvg+UzCVRUwhmmTPHo+SMMTaymMT
VNyou0fU7duvAe3m6moWDj70snRbeKo+ZtZ6QlixIlpuifcbS2x3wbhlfrFDg7+Ce70fGZ0HJo9D
7647pxKDN+Q/nvY5zZekUkmZFmpgu8tUkA4BKl1Ay4XpuRgEWhCZj/mhGQuIg7jGScFEQoFlrxww
woXnx7B1sfdQsY7Lph5JD3pp58ECbMVvzpV7YNsErW4tRpNRcuZ5fMeiUj+U7r4fL5cuACOZBc95
NhUmsToLLE59kuS2cA78qsrlbc/8bG5ywrJqQb+1uleyxt2rjG4pDxOHmOVBRGQIh7g49MTM4fya
njvRK/N1twKDFrIvwp+/B1XMCea78/SnSLIZboVzzWF0o+nSExbvSoaJeUn0EdxFFC2WroZQPLDP
1ssrLTq4NfOjHq+h9tpckuRFMONyFJu+fqaUFVznENwg1sHwi5iQTKxz+vFYqCEi4V5k9urEEPaT
6kAWZvN4xBpw5i56lZzPR7Eqe2tnjM7ezCfyeXV+NG4SEa/G6WxIk3EUp3MQl0MljbrbfxbyfLGT
WOUDja4cBDu5ol2o2OMo5mTEiQzUR4JbcKSHPJLTUsezF1j8t74r3K6Np8chkro6OsBebFSlFIy9
nKwtCKKzRlepgk1QZ4OYFoXoikvYKKaV9ONtNjrI0Njmmup1r0zn+nxiXTuWafnYdJW+45XZMeSX
dqDjBfBoH9E3B3pke+3veLFluQnLW9yoDChGbXMnkddTfJLYcPx53vuwmfGedOMjEKOrAtE33ond
hD7oTlaYb1pQ3loZ861XsWv/L99gMM+tKLnqALEHfA/VC4soNYN/lNvw9rtyEC+f4SSHNK5wxvLR
jO43ykvT0b5KVZJTPLotl/qm9o4+VQ14sl3gngiPki/AoQjZCKwKih32JBWRuyfWSGi/dQ4zLFPU
zbFpvaimtHxfn9Dv8IGvml+e8uHccwdsk5zyMQaphqza3XtAMhfYS21sEpMF6FDG49iiTNtIDXTd
Cc8wql9s46l9WO1fJYEFvp3tld3Kt77QFbtZbdJ+mhzqnrOrrM4cuvgeFSTaT6UHj7kbDbPllJuK
wAjsmK1eIUA5EZam5GdC/4g3+58X7lUvpdNwk+8qhAO6db5kWPxpW5enoJsEC5seTfFVKl3YLRZB
rMWWkiqzvTVC/oT0EZGrR/8CbLYHFcAlAgJSJvtWuq0grotzNLVvG1IXA1g3viQR8oHMJkbxy+vj
VdABNmQUFB6uI/5b83ZtcnF3X3NLmvyJa82c3D6i866ExbgAv/o1/s5Eiub8zKtCrMWr0jOsgtoh
WyFVadaXmr7vxJnQMhiPk7VQFarFr77FnYXvkanwUqbiTcfKCEdOOLDxSqu7X7esJnrVDxZJqxSv
q2y6wljErXbtYkYRx3rFN3uE1biMryzJlR4F55IFE+cQaJCduNBbKYveZvB9nwyF2PVBJu0kvN7A
HeImkbHwiqbQaTSDPjdwEuVc1dp57QWgVcarOYiFp2TnyG9PQyDneeJAIrrWyYSBHa35MVSnsk1x
0fu3UVoEKM3Z2WMLfwm1aGqo+6mRaH1hnJWYCXAtIWtyB5wMEtQC3OG/sak0vV+naG+oMri1Cra4
8RZ511fEAAuCxSq/mph9qLh+TtxiQ/Vs9ibJ3rF+Yq14EDtL388dN43KRO79ybquIIA84NL9NVFZ
jTygnbk4K9w/Jb0otlU16wfNwj5ywfPDbjDY/oKdBAG5ARBXt+GrWZN44suyWf7khrutXoEO9TbJ
DjsYtnyaW8XtSifYCYJY1ZOVhcFSMjOE+Ld3QPWXRbtueuvho+yF86DDKfue5tuatTM7sLxNwc+O
v7CDK4Z4+KTeOvtIKbwOHo/nBSOr/4z1YRzJSYT5CE4vIhaaan2ZkrTf95Jk+nU/GSQOT9AkQZ2I
RH1sXg7Wt+Yhdpw8Vv+rGQqy7hQ1ka8d0FDRVC0H4YdBcdE5dg/cHEUtmDA3F54/F/Q9QxMlGrrR
PH7Blm/T3YiNRJj//elRqVSzJqdBBj6Dc19qUfvlhv0wfhjC4o4beBJDPa9c1ipaX+ZNkeepN5SP
XUuzVTKHTULBWQrBL5KugphGKbGcLosecvxTEKH3GOasV18Ygj3QLp7yDz3MWzWO+o0+VPM6bWog
wo5jHxnTl1OU95YMEJxrO0e3neodQ7DtvgeQmfyqR2BwHw7wogWbE7RCFDAulZ8jIvC9cRhDSOIC
+hsax8xX7yoCvhkAmiVZe99YLx56Fa9RJvxK+rJIdORUz0P14PrfCaaPEjakt5ezhOtE7SKXbROg
blWbwMR8E6OYxh4UrCzOjMRKwC08UBK0CtQ/MmZ5UaJjY1UE6lBsa2U6nmwcxdInSg0jwe+1Dr0/
5jfrKcmxTtRD+8mfyGNglLULJuvs92gQZ2k0uXy7TsHsXRfBlpEDTVMCQ8YDWIvLcznwlK5QocpB
IpwZUhmzlJjg+ia2iheAGiFKBu/OYheG1tLgGVb9n9x382hPzDmVB/p/mBo6oTVtWPOGJDwZ2cpe
c1M2+O3Yi++ozGMHmKBBqFexIenOzNp8O6mj9ACx45cGiNRo6sH5ASBPKBxNx3GBS8AYGYiEwzqu
3YqtnskdZCB3I0Hae3Ln8DFa3xVs3G5buzHnJxV2hLUtYWE98CltG6YwnGj7lhSWsySLYZF2sMKy
FtvJW0BHBL6LFru3EphRFnKlWVHsfs+bRcAmdAmFOnW9TUsBODp74vxChRP5zouMJA7Ju5N+aOQR
kjXp5lpE2tl+lYUUKQi6lfabNv2uy5CD/ssBAvgR8SKwKVxIP54PluhYw5sK4dolTI0uZkGhhLM4
ugDR0Df4P1ARjXJ46xOvDdHUDMvA7TqvLsuzc9kTM2moAoz5alNOki//0bjCf9RkrM4czQLHAZSY
kRcVT5FlxLJednNIelk/aG5MlJPAcW6XdQu83Y6w48yfxkoF2f4J0NXNsUW0NQin3Zj/pQ4qBhDx
qQOLk3Ro38V8l2nWHUI8qOB4HSOl4rMZ8wz7M5KGuZoI89prl23iYeWMG/jGky6Odw8KsLVyn+gp
zIUmGgUUq8SYgqaPUcRFDIyocjgNOv9m1gOIH9QcdEt23wKG0jZz/JqnqKgiviHieA1xa3fwvqO2
EcN1xF+zrmWNzmXJ998aq57JQyLMdSPrKsNyfR3kRriKNQaQINTg7utfJVrk9NunI3QRYo96Zg/u
OH8vA2rCCw92O/jYGFjTkKVboSJzP59IhV/wMIsSFABwMq6tcPW39Vem7GN4C/my8odalhEqfmA6
pGo1sVAPrwkINwk1PhltMyOFC26SvZx7pmmaa2ElOQ7hiHzJew269WI0IeorOFeibrhnxfevG+73
cBEY8Fz27SK51FFF1h9ovmu24IHFJ4pG0Ty24ZIEfq4cYq0zmzzcZDg+zJUwKeY6OBcCBC1n1vAz
VdHq+QzzKxfDQemmAXN0W2nLYxmBvNasYmamm5KULglqNdWc7V6F/J/o8ilo3d0iBsJ1vpMoEtic
mQJXmPUPO/DipVCFiWhywKrf1qeurKPuJWf1aqQmvZUQqa3cJQRQQKOAVkbT/tjEtN6FIX0UlPpl
dlwbHC33TPVWJSgC3xmQStsQjiFUCvVDKH5wt0ykCe+nS+/o6i8NpR9By6tc4NCB+IjwnP80Hi+l
RK8KhEtQ+9JN8bZ5QsMBfCICFKfDBEsuGm4dMq/OTVImxa1P9Ms5HZrWliYYnMZ1tBLvIgew9d/x
TSfnf8WKzQ1/M0JpHk5VBCxRNVo+3LU76eBNqTENDKfELGwuYDuKq+PcfBSFD+W9dDH5oQ2wLaY9
9iGCSnCwqPB2NbYXtGh1aGljEVICmDSx3jbFli9DpyvDZnAkKwAw9DKNzgl5lWs/GJNvVUvQnsod
KWrKA3VRskPV2ewWewQJWSWdp0qNq6zceJlz0sNWtPVPBTx7OGfO3Y0bT90yaJl118fdQYaE6by8
V4sCEImh8UGYHr30+XDBbKahu1J3SPmr1dtIS3QJfGnA+11abCZc3Tbn7t7pZT/m4fVKAr6fTrvR
3Pvtmk2dJmljMa5M9EckeQWYF7dYaQyqRAh+0xvmJ/129le81GX2sIQEMtS/pFeBHsGQpPJseOG+
+XCbAejo4vKLZfXOsC1qhaEFDC6D+rgnIedOByN5OjbeKvWX4I+69DydnTyU77eoWyW3nVzVfS8g
1Bki/lXmW2Pyi2XZMNs4EDKa/nYkfOq5yCfltn2HSnuSvBc6K4SNqpOOn465pRUCzAQ/E/1q3Lpo
7EX54N7P+1hsV6ELJpIJxWHMSMyaeRUCHSzdY8bYopYsJ3CVbcEJ6lFhruKLE+OzKsoKsQitfVfu
y0DFTDnwrtzDnftzru/sKYUJCKgWvxetkC6s0ha3hpMWoKOfuGh59eY881iY54mea58TNFSqP+6s
LBIbOvdGRj70931FgbshhOuTjNoX/c1c8nw+ZYetdpv0fNl88BjLqeO/vCmKAOfiRO3IklsjsdKP
2ZqT605ERA1BdYNXZNDhcUhr8BJoOtnVNA2YoErvggIye0S/YVKd1rah0S1Qz1xdRfwO68QfnNFW
n2/lxDwD9Wl6R/ES6RcYfWqracUh+mlk7It1m3beTS99j3ZRX9rwNvQjJsxMxyyW2a4ItIizP1yv
J4TT8VKkErZf+yxKJfcPZZGRhdhrjf/tYTD3N9WyX3vJxJUv+tGDJehLMofpR0EmFrrTEhqPjCni
eY2Mo5hsPjxpA7iKYqG4h7Ta58Jp1VOeqaY5FFb7cjaWsEiYb66mhV6C3uLIFJRnB8yGQmaGym/W
mEVD1LiUurJAUB4Kfh+Fe7GVUIt+E1eIcbSQNu/u99/QkYZ7+kDraxwpFAR34BftPpwr4pudvSVd
iqWBf7mnoO8VD28VBS+yhpdXclW4cofZmMnlglP4q46jU4oDC5ll5f4QdkHQRoco86Acff3lauGo
3l6E9yDiuWqYGvFxtG9tqkeABbJf82Ee9CFjichaN3PdjqgXsRT/xGJELgvrXXfztDOwq63CZP87
n0YJgiseIxSbQQECG8y8ysJgDSfeJYNCtc4qGML55+y9ncSHYbSzAvJmHpHVYRGHN0fpxhGONHOj
ipofSCO7QoxvIC48oJhVwgBP1KBbAQ/nIDV9/aewtTANvktuB9uC/0TXcRqxmOuK/liFFSTEvkH0
NArV6tDaWqpmlA940wf2paYtfMnfZS46S9yaNmSKBYcdJsecl/H3DYVQuEGZnk7/sfPols65eoti
qJ6ne1xBfna0PAKGP/onaCiwMQwfB6Xbby7yTtLOoG8z+oCtAzbgY4xGZWnOq43ZtmCzEc+7X4pY
dq9qSDmwfhZ+w1s4hDTJfaqQh+5OQXtK4au91gLHiLenFGbXj1K5XSbZWWsH+CFFPGAP6m7JplLh
PkR3VpX7ZfAtht3qEDhlMgPpJi5lq4Bxsu2mCfgZhRNTrQ7m1GqdtwAbSUB3SjpvdyA6R9SDBr7M
MjFiiI7ujlewd6iAxzfUUfaNWcSmcW0S6kKlLvhVMq5W27e9IhF7cX5gZVG5BXQBpnd9sBm8si3u
NVUxjZdAak78LKRjpY/z35Kagrr0vjsnD6xMyZ2bRhNgpa2jPblAE81/hT3XMuq4Bw4awCG0eV+o
pR7360/tSjEjXHUXUra1Tsww7P+jeIkTjzrCHOcQXFsIz5DBhpWY/95aX+VPsrltsChyK0einp4r
eroQgCKogZ1VZQRRjNkrui0x8xwI2K6sDvI4lKAfKqGLdvzkxgq1ACsG48HQSP4xpZJphZcYLPGm
edhjygfI6VxkXrOiq6UdEWOJdICFOT77hDz2KJlqy6rb7KXaSdKWTeKh/2//bR0LZxxnOsCHyrTF
mMvLYbJtt45vA9+ue1WI0fYn0/QMpDAPTI863A6/0Wwjfj30YPQlRlwQ2TQzdlwtMmtKbkd0rvR1
3GIZG9+KG6lE8YQiE2K7vdodfnRmL6SLOXXVC8hqbHDWt6L6U7X1nueQjdP2iUJDcq3IBM513Bwf
8P2WIv6BHnrOx2w7WBmYOAuUWTn7WZbGSaIxNNCDWRnM6fq8VY8/cVDl4dKdJZ3Ab+XnS9uJfpYI
7wJoRNakY1y9BL76lIh3chvbl2qJs6N65eOnkObd55Ir3hiJGunz198EkC+zyiQGi+/EoDNgW3RL
iA9U3Pqltw3Abu6qVNdeeo8SyaD+07AzXAUX3RoxW33OeWL9Z9BzWTdi0uzAALSV4pptV7v2uZyd
J6o8wAAgf7YBNU9ZL+XsErwvOJT4P5ge/qC1Un4gUBN13DTrI1R47dJQbgeWsLHdMZc0K7WlWVio
xSbRYE2eYJqT19aSh6VQSoxmJ8yefzWRLf0gsguPInoEey1OKjLXcU1xytT1Y/3pZmz7ex8VSXKn
Ez5y7utucWW4Mw9pZiQKrs5U7cr+zGCzLo+KNIFvJVjz+wvrzwp2wFr2C/fLQYBCF3Uo9yn+zGbi
9Oun7Wz4NxBni4+C3Qag+uz0uxBDdJNHeGCNyXzdeblW9ZvT7BWDe3rcoueS2LP6XDhCtNLPuabU
NXd9Gufg8SFwcTPbnTv4cwqO9ezoXhyXPkbaQGYNiKVWKMDKNbEaRIwGlRSvp/u2tFEKBNSztVrQ
x8NQO50HULA1ZOwS8ZK3wc/2AIw6ZifEHQLzz+FMVaFfYCahuW1igORl3ZkrUxKTyrzobeEy5eGt
UYDyXGIOSviwmdvin4VyNQ1/8yTWvZkUXR9QBJoOKFrU6haZDSdFWa3VMbrcFDHuxktiWj1CZtu3
muq9yBLAPv+Zdt/DlOpBMI4GppudFhO8134bGmvFRHyWpm/LMslDQGNyzU5pUSftPHBMVSF4U42L
B4pd9sAA3QhM+fPV8Yf6ik4gmgCZcMjrpeL/aO5V1guNXleHhanoRwT5YPi3AQ6lshRGCOhvFkPV
rIgm12gv7vCWeR27921I79q20XUVZ1ZMrFQP55lfT5PFTzEpnTH/xNZYgNDNcj2D5u/1XYQNKzWn
SHOJiCvZ7B2SgGKziaF2KYZCFTgytpGK4l6X3N1MqwFUFxSjp3l9yLKyz1AfLRpwP57uvyOqeKxa
+fNN74b87w2LM4KXSzGqUZzW8iEvxwsCJCJ+4X1u02WA2Vv+JfCeSD7m7CB7lloeCZbs3yI3OI/G
VMv33MJQHSOpfuG+ArbD2KcGYLJghHlie5oZvhnU0bftiW2zXYJ5nHrYuTJb1fmLeZOcojH3zs38
w+kqA1KZqdXYwEIcDgbCr9EDN3nbQuwDvYrZTkSrIUwMCF8n8ma+Va3rySzqCVe5EAyEJbmyHDyd
CTDP1EpwBuAUmtZlyy8K47OcqKiG2qxxZxH7krXUAKjD1oJLHMbcHzTg2GB4ETIDizxY4558FMOH
Y0ThJEWxlwf+DQQUhS6UyrHfEyPjm1Xo8FhZDrAbiIeik5WMaIhnIme0367moik5gyFOJExIYIKY
mNmUXOcfyhKerjEGnXVT0UjpiUQvbdtavnH4NifxHivAlopqGkcJg9P2emtZ2KwiNbN2SKh1s0Qu
14Fogm0lWxWzuPfI+A1AFJeLLV1zWFMp+2auPZ4PvK5vQhx+VJ9LT27QeEbpGeOM7UaK070kfa2H
w2FfYgpY4Y6QN3EWkqrofFcf1Q8mOglRetljbzk/GxlZtwf3nB8dJ9whmDFfqoFp5OTmgUdyeBcd
oeVuY5fmYiiR9mbIY0iQEpkNFi/J/2alBNQPgtwS0LvBfluYbcPFVp1O1moSVHDFo8nqm8PHbU3J
qxkfxOqf88+yHy1Run4FchoKvvmTsj3BheagvB36GHOCwrG809PVHIuMdLv4CVoJwcd17H++Z7Iu
9uiJQCZ4nZvPVjjns9nFqqfyHJi58OpirfJMb+kGP+1VC1sxD023fhJCQ52zoVOnfIh+9L3jslJ3
PmU+HhslQU+MDL+5tzu/fklpiO3Sr6zbCogii5WHY5hcD0L//PNvYWhivnJZG7pUZXEBHhFU6roe
aIUmtCQ5/BQUR9j5kyUmhoAzPq9TwL/pcUzncR87UezDvYNgYJkz7BY2JsKT0SCcPgOhpVXIJRqF
1p/O8M7w3Ye+n+2ZuOJZAPBgA5lRy912t7R/wN7SVTo60fPhUlIyS1xMon1ZELff59WARMLM7LQb
pWdOkVsSmFt1JgE9tySJgeVLBT0nSu2sFen+WYUR1Df3VF6+gmDtav/3JxCXRCjuF+wOREo5C9Lf
WRtuevPo2jvJ49kIDXW0uw7RB2AyLCFub3g7My5eSi/GHaPQ1kAPggQTGNJn9TZz9qlXspJjwkeE
+SRROkbvIKNToiONxqM582ZaNccIZqFXJBAi9sOm1lqZBgx2ouFMHCnsQyGuMKWSrFOUYiE4QHx9
Q+t/XWafeepzXveNA0SLAfVSMBi+yDYTDd3nU8cUNLZNGd+9AhRqXNyxyWAEaS19Pw09YlCM1Uyg
Bm3zU5oszlxNvrvStglx7Z3WDMIN5tCw9yR2G5PGU3pEZTgNEbBHf0h5QbWhFDzxq+BgkSxKs3Lk
ot8MQKzMcBdivpV1jRi7uIdCKq1qoynIVyiiBvnHQjJw17TldbJ+lSZseP6/gwZNFS9iuVdylI93
KHgxhTiuLjg5ZTMm5IBV8G7rGwAfZfDO1pELctZGOvJBqNEd+YpABCfjDcNWQCQ6f8j/R8vAZswr
2gCrHguB2XFoFONlnW9OU7U4hN/Hj3HDZJ5ONcs9FkaaQHtyGnyitEvEng/+8NWmvJrex52mypd6
ZuCnQ+pRj3aMfbGLg0E4EPCXLcK2Q8x2i3wXIbP8Rbrv6nPSFJgkY2GiPhYyXYUbz/uUc5zXYVwD
2MLF135bGAy5YoOJzurjaP3Q/Bu3EV6oeAN1+UYJau5wA/dU//tc17WeBjp+OR5mOmCRA1mTlbWc
btjISBleG+7qIXFjXX+BM3XrIkxiXbwvRcVzDBtPB7LDrVJ/narAFVVFnLJ7aTWxGm66mXP7EEVs
ctIhwH0p394Sfq0JYDUWBnvpCRzlrW/eW0x+coX82hD1P11NCHoisfC1tANo70PXfajisbgNpo+O
691uMIDRRGSQ9sEjhWhlWIOTRlKPRrNhRnkaLBuJ7QW8KgtgLSutDLtlFcQomuHAEKWvQaDQ98Vv
z1ZvTzQecSm3Y0aagz1Q2QTdQ/OUTSUoIb4RFoWnQmwAYfOQWHNm+MkfKNEmXCki8Ed2AWYk1uk0
lf8oJX40AIuK5HL3KKQdQ/DQ7spYH+LaHMinTMiB1fVhpMVbaNCAWgt53iUZxavTO0aoYqrkZd7i
/lHvNIBmU3Og798qenvtWDFL3+3VDDQJZogX4WRwQXww6eUMh6R5CWb31v/m61Q2P2NXJMfhIn9Y
UNgcfWv6ArXs4BKR7CZUWLqW3E6IhtM7sirnd//gbAh+xptTliw0MN4CrpXrydgihj5Zpv5Tu6Hp
+lop0f+d2CnVPUPdxZ3ed2G+WQnCWDvv4UzXFomV5AMboAw1Br1xnrqo3Nw/B9aQN98hbB2ZOUhd
Z0BuOOOCjctIoDUD+JGIzAu9+/csteKlZBd4ekAhhQz7VJNqTWI2rxELEP0p74kQ32AHzJBOz+ci
v7cU/3Xl1WD9SqCT35DmNDNGtxoFSBik+9Irt1yox2QsU0+3n2Rmr+y/c3dYMbdGaF1mpV3L8OWV
2CywufcL8cvm97eIDB9IQzKNFmbJ/bjy7MlY+d6UvFBfdGdG+8SIbHRtDsaLQrdOS9itDtpXdmuR
0gXQtzEf+wNUM/enkHG6GX5iV2l6keli9qwx9zX1SJBeE/Sn2crq6DQ1UYKz4oHigZKLu+mPDx6z
IWhJNHbNYZ1BruINQU4td71TjKUFswoqhaLIcpWqtwtMFvP7AO9ABpMqK0fQI8i60RF+WktKjwnc
Onw+wgMgO5WT28EQ734kEcq7/ZhT/v6eL8e7Dlmv0fZnXUt8hzZiuIMBe1GQ82daHFzX2cPHGiC3
dzd4WilxVagCycv2gJ4/oFA2MZbDPT/pfXoWEPquLWhKJTCPL+sS3spDEvVrYvgOXiUfVK9ka8j1
2Te0hM0eCQr+gpB9+kE6D3tIJ5yMXedCskG+/FhV0MaiKCVDmJUE3i4HOlUiN0b/Wnknb37dDaBi
n7HYS9Bc9JC7ho3zsPgz8IxxORRHQlConnQxG6IzM4abiO4COtOJu40JVE1tgmzu45Z4uA0qYpH1
0msTkXrmmoVcHy1Bhy8LsimU5AGYbsRHGjrw8U6hO99WjXJoT0YFtuALrLlEPITMZf2ue7ErRa+K
C7Xizf3Iw12fxEDP0RodNKP+j2uSsmzhSYblfKcF4gGfc90DyPyB4Se1xAphbMK3bi3xlN7YJVYx
Hz1DAW+YgQXXFqhkBQ6sXWkAyNbygqkoowest0u+LNqY8cdyW3roHtGDRuV61qWgt61vR3iSYIN+
+HgkCuQNeLZ8WiEk+XInysvYWTLcgKDkfxD3JAHqskTI5cKkb51uzT+y+PPyJ1Ep2cTBsmiPnB/v
D0oGZpx+zd2fw3ncK/1JroY7fDM2zyp0dEPElD+o9MwtMU91qIirlaBVtSTKzoMo+abYIkl+cvmg
Z6OV+vTJtd4wJOUO/xmYOtL3bLoYsf3T16tfIhhTphYnsljUXFzFsNxqqN7lbVei40hmL3Hs9KRf
rEZdpz8s2MGTKItDfeGmChvBfT0C2O2XfEqkK1VHH9JHP3PuGu8I6m/CVY+ElMLEWoYKQAHvWck0
BNspWVNLKEyJ81Bq0wyCd5IGWJkFSGEIZnOzKXdle0KFQmzGL2zxdCdMv/P69a1P/suAGiWSfUFx
nFtfiw/qjBUyAp7q3cBDvqAygxZAasZPtj9F8gdSIdINGABSCfj3kE3aXPQY6sXSyuU+HX5M6W+0
1aDJg4FNzqFmfyk2pyLH6nfAl5qQLD13EvxIrj3ymtbgDtpWsPskhPkwdnf6R/TWIJIg/DsxlT30
bCB9SvKRw1vKkTYMTIauGvdOLnYYmh5m+W+yW9ydWDElZBtKd5s701ouTfqh26uPhXDlxaRel+dW
RuPFd4sZnZqqAV3ctweNzqDQGHJVAZtjx5oVOugaTpHnhndnQKFqZX4PQKaMT6SWIJUVwW7Jw81y
PGPSvlAdel1AnKYiKwMcPaLgRZOzsHq7ELoefSdIlfncL8KIY1DwWWJ8rac4c14VKjoiD/Mp2KXT
89HXn1HTMgtOTAVkMU9BLpYckEq2RUv4aNO2NCDOPkfO4JkgCq/gqbpYsTlxHwayVTzcIjC7SvJs
IQFZytKvnSyRj1PRnf15b8vkbpTUtupb8oE67SWg4ADJN/Cyk9dKOBgT/CiDPYm6M+cunBU5kYgB
Fiv5NRxG3yTh3ftJRBvH1n+2SP/BX0FXwcAon+C8JwuEA5Y1CCT0fujS473ILjNbUdqbRUCjVTfx
f57gmv+nR/sC4x8kB/9W8XIu1+tKMddk7NY2Bc69/iPsZibQu/rgGnZMtE8V0eLZ/f9UxZzfEgrV
/MGATzNnQaoqpGZkonbJQNts4XcjTtiSW3vCiyjoCRhxcVvOPx/eMallAtGJLPtqSCyfQAY0Test
lC/Can1SzKpoCIulduyN+PW3VIocsJFvuY00mGorqZs87R2CLcWAb+f1wlm0kZ3ARLFNuFLF2gKL
vMelbOC/Ble16JfBJfmI80etr5hop6CBky2FWYjkiJaNM50w9NI3Fz5IFS21ep/GR6LxNfoyuuOI
HFRjrm3h1PiPcp5b5iy6G2JX2gfHmkaO1pUaM5pwOYN3/Lac6fh7j0JyiAJ2S5wZjUOJMnZ1KbCj
qwuz68nIRmIDzgU6ogpxRu/W53TrssAmQKSLOhiaiAm83urc5Et8Ez7CbR1YGM+ibGrXF47ypTX1
Rm/yFJRuvuj3Umzvb/JtOgaaCEC7IxpJivrVNB0S7NpcpoKOrxNBwsrsYM0LjCB/+p2vVR54LeLf
b//Lr668DenUXNKGFx4oTrYkp1ZqYI9RJzqlwvFPC/At7nXGuE6LVQwbhzvN6ixfTvX55gLAQWxx
dh/LCzzIv8z1rF5cOSnxUjq8Rsj+TS722U67mMms24Cw2VdrPiL2kyz7BEXJDTm9dQ11JVTCECuO
baOJqsuleo0R7bQyrEv025oCSuU5r3UCbnFrKx9Fh8BOItVXJ2CvfObWDkwg9Fx5hVft6fv0vLC0
uDaVgRAezONgiAa4dCyPVQlHcWxc7tqjgkKhuGVq0oYEnM9nR0ZvgCZR6fC0OT1k4Pe4ELuQWynt
AGznGqRNfQP3EvvhKqXBTnD9Iqk1fpdZcCnhcG7hQ23Nj+jBhpj5cqbVvEPAKN9mEqeAEz0abhNy
S7G8ZMOF4ZHLqt/OjmBqMqF76GvyzxWZPhAnJRgcNTHWo70cR5PuKvPYxtc3umq+dgbObJtHBHDM
tovUr9pvvlJdSijXkTORFZuc6Zw+I9vKJux/Lno5gQSVLYaAFiCrEb58iSlLoO8evv21JpNp58iP
N2KPijREDfuB5GkHRwIrEunyJ00zRT355ojZHuVh6Mo9t/AzogEUshJu9UbzsKeWMCJJZZbrwn6E
HlTfzibI+CnQ/l1Oq980qeYk9fUXJbuwCtJ7/+mhJkbW9yiwoIbjiqD5mvG+QEdpMPyDVdwSsckG
G2shTI6Ek4WsL14zlwknFViNpIfuAn3oVwnjdY2kY5No9fWIsg56OOJPkvp1VCHjJsU8OBvSEjrx
uZ0FqtlVfm8KrhZ9X6WHGdup8rrg3axy1ojske20hjVQXUAuNN0qrLEAIQWnCgZ5rtYWVSexrJgP
bZ1Cts8Zwld9hAK7CNCTjtv/MGWGN1I/lxP0iNcNpQqyNgJqtc+aqRodnPwdTJ7AvHaAfB5bXS+K
qXEOXbuNc1PgGu3ycQjVzDMI3PDq2emN6rjskNvspV7AGPON0uCZLagAOo5P4/OqPWXbTTu9vzDa
rthICDndrBRZXf1NmwIbL7Zz5ZzDhkSh4xJxk6uWN+nG/aNwWoXSo0ZQLfaVLLePyD9m6aLcCoPD
AVQaqun79SAyZDMYLZcBZJcOprOau8l0REDvvAuWZ/806WHi2azERSSYaURjcoA2zgJMhxhLu4F4
o0bF81jy03haqcg37WbL7Wcmif0V9SGNMloDLjDa9VKoKVDo6tEh9fSsmFKNASv9TkP0TsDSgp7G
DRDhZh9IOA937EGQO4LIspTkKGHtI3IMrybYMjuPA1pW+W5RNcIt0d1kTXNYS7Pc3P3banJsdlBI
ARga4YGx0opgjG4grHtr3u10Oyv33oM+m0qVcAIwR69lGSq7UnhNLOu1gGjgcwRyr9GMFZO8ps8c
v7z8fHCMn9iU1xUCA4G+Va6CVSxjHJJygPMx7qcl/YbDJshJhtbtkWEJcL0hzD6L9WlBg95slgDw
DtgYhOh/CZW5GuWSJNSX8s9Un0UpLfdKqgUPS/zrq+iM2lqHKwqy+BPIAdgxSk2FusY7mhfyHIXW
jzxGK11F6Xd5H4VxcYFp6K3WGCffT/6l8dI8QHo6WCH30xg7HujeY5RDXN0d+x2sE7MsN5tJg0br
bg8JLacM7TWeDkgDNIBity/lONjonhhrvkBHyrI4wWjbGTKgyFFMLxT/HAAg26GSX/5BzYpNyb6F
pMSJr78YAnHLYt+0BX7eVSUxfwtmIZwQjPy80yIKfvwkzI9jDf+WDqREEsURDg5Ai9xhH/4Ghb/k
FPYnAzPKa6wujc1tb30vZKUh3FFVO1DdQWqzdjAXHQzKwS5+y/SkbhhdbT24SDARJR3I1fL6LVMQ
RQEyivClvy7W
`pragma protect end_protected
