`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NnoqlrXQschQ4a2eh+9Tm425YrIX9azJ5mNNlDnw9rtbK7gA5rXH1QNdty6c1yl5
amCau3m/VNgfdC0VuKcFzp3r08qVKZG3naxiAxtwAld/4XXt1bXuz2sUV97MTCyu
eA0DpcExdpoTkUJuYlPV6kve6wAg+qt9znwm56vnuAI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18352)
SY7O7jVQdXRo777SEw28uiUKKGaFHen5nUxQyFK+66GYsJtge6UCVCV7/zFJhnue
j8XYpwbS7+KcWkCQ7i+xvev5pEZOk3G8jacAiHIpljO04oJUS3J27mnH+N+xDPvf
wZzLH9tBo3DqxsflrqOmpeMcLraw57x+dCVUnC9HhUruNucFEulA3U/oEWGQem3i
me4TCE1WKbwhLmMIFj2SrKhjK1SoFdSNFtgUoQcVCelVlkLrc9hWVcn4Y41egUvD
OplvspQx5FHXQbhsB4A237vHXKbme/iChzF4mRxb6JPir9gurU3ZSGlfyuBz1Rj0
bNP2KIMibm1UBgoqZ23m03wNIKYaV/edcwE1YgfMEBRGRmi4hdY0JEQcuR38Yx/w
bvDz0BD1zLSWsXb3GI506Lvfq0aoYwzBQ1OOcOayxSzyMP+Qr1J9Pj8GJbVg7kBM
cQ9MTuZKghw4guqngAoI/KtOQuuOeWPqp3sM3So4yAt41WrobklfmJdxku3c2QmT
v2oZMe1csJo12+Lig9RTzgbh/CaGshZAtGOfVJLaX09hYt5TEWhimHy0zEL7f1fU
egUHWPUA2F7Z3WZCLTMu3t7fD1qDh0WzUX9w9+JgsM/2RjL4z7duJoCSI2RXpFPY
x7grfmZR6FDj7qAuRJID15u+GgPXF9T35HYebWPszbNnsSLyudGzP6uxhcE/Um8n
E5J1vE2lNeyN5NYjhHX44mb1pCT92fPOJK6dim+3spCXgsHhI1V29E67N5xrmnt0
wXaE+BGtxhlbmrwitsUm+Vjet3K0jmvmkB8dcpPJQsTHCzPJXhkEBrgpyEn1mHsT
oPz2dZrA+CupSXVNQ89r029mVADRVL+nlV4cryYnNXecXYoTTtyLj2yxZ0EjVV5t
/yZ1b2QipHqnA7QHDr2W5RV5Y07QeXzBngT3h2zNZbETrAjOrn5joO1bCKMV4tQH
Jvg7MlmEZpW7BYWNi3RTfNIGCTppx7Zz4eFNWI72lABgUiL5ss3x7G8K2x9CdJ2c
0zjTjQe+73zNH827/+WeqX/TmZo16Cl7QWwsD2e5DE6+z+ZD10f1MnFGiBI6IRoT
OfFN96c6DXSYQEJ169w6I3kQc/lgAOhsFkay5wGvKZNW3Ay06oYJkQ+PUkZSD3OW
I3ghmGQzUdtf403wJNssld/CgU4bkNVJaxoRJ6QJjFtPra4KOdz54JCnYWJkhkDq
wrAJ8IMtwTIQbtkBU6Q4YaNWkiE7ZQ1HToqqRkAbjS/m6tYkbu3HP5M0Qg8at63G
WBTzUyTuR/zVVTP07rPS8Z5UGx1PPowRwge3Bcvsr8dlPlliNYIPRg16LU2SNe8I
/XX89b6MEaJ7A2CEEQDRozukQPmI5nZWeSspXQjpjozwiK582tHq1LDoKjtIXiNA
kR7LldGVeAr9aK6SiroZ9ePondNm8qHyhHUz5udVK3D69UdbNyjsY/3WQ76LMC3g
lJvdUnoPvXEY5TZKArj5HVa7z29ooaehivfEIcxN5qZaxhO9pKZRU88+t/RDN0XH
j09v4GfLwHoNKotBgYNbkSE6RPbtF6LDLEZdfDzjxY5UZuGOjXEVqND/6J2PJRPA
NasliWlJq/kOTWNf2RjwOcRFiKIomu8RpzpUnPAGorHpV2YFqdNfWGAdjfcfbfVA
MmPFxLTDANVv+ZLsl9CxSzCeZ2zC7XIoqNxMNkfliEQd4A1eOc5uMlKsT0lGFh3i
nGZaY+4sU0EqQ4XtyGCsevvUjQdAAQLEjwrdQDHKI5qiJu8A31s0qhGWPQbl180d
fhg39sY7dJwdLW/pom2mN89zl3ienVJkMXVFnukFiW/WxGWQRwuiEFBQyURIDduH
UhuhDhjHJUnuM9mMV3IoRBisVirqZABeCWkzzqBdOUcGgKa/GTU2knM3icecpRAD
cxdDTuaL4sE5LXn97B5/npgaCBGS/09FpYa9JxF6df8zulA928RKC5Jnbyb27aSc
wVF1hK0yUZy5G0duelXrgNDqRfnh5LoPhSoygD6hO2EQRLSul6F8vZxn07h6uugC
o+Y3f3p5VD7gX4yckMJVDHxX0wg72s3d+gQbUOU7agctNMOXn9vmsf/4VTTNUJVz
Q6NN/mAwmLjt7IoHUR59afJkeEE0udDjcCDkywYNJvUiERzRxrhGrqb8bP3dfHaE
84rgfeM6/eEiTm1y23U2bnug0VgDPf8DVjcXOhhlCBUKBCLBuVh+EO3StlSISJOc
64R6cnIwURCRgwfGVKx5BEc66pq9Y+mAB1FMgnAlSwUS74+KDNEFwyhpgoDEHD2P
oinR48j/fP0xHLBMcgeJxY2JMm5kgO9EIoAvfOPMEPJWCzp2ececmAiMsGRTeSd4
nmaB5Hs1dpLntO50YXf2j11B8YAfrv3Wxzls3fjSZu94GEIPw64uWQ65sTmcIRZX
frizIF8Xk6R9k7Uw1STkt/2BHO6mZrOUHt8TQ5NMpG6ozGkFpQRmcxFrKCRovjtB
Oos9eyRDTWB/9OzkMhg0863qvIZ+WZXxbXgQMmJNtsvrmozT13Oxus1gbWmKUfOf
VeceLBtSj9RZKbtlaBIXChC6ShkCjvXy1U7q6ItTECG6jESlx7RqufmBJPtsyBSg
iYVUtBPsZCRU1TnjcrfFG24xhaH8dh15itCO+J3n4pv1aDnwMcMRTtZnzss44V+v
FmSTTpK0+OHLkx+vaOvLsRJd30CLhwyfb1wTBWjQ4DIPhgonn7WcFJcoNmTESDPv
s2mJPoXHWYP1wnYiXrEeOV4+vqEs2f8AliH9bCCznn5TYtiy56PthP83jrDXqh6J
nziXgHumPsBMCRQzQyiHwXm0nwRo6COi+yr8Zao5cBlbG/fcnAHkex52vK2z5k/u
LSfB3ZontIRJ2N1AmGM285JPJZTXFXwFxYG6TXJo4H+2gPMN6lcAtijDNCM9q9nF
6dImFxFHUVzJtXU5W9yaXjgEQCOmgDRH0ZtdsCX64odgRmR3/9kBHt1aIr8GjEZH
O8+mWeUgJFqZB0bhAxBI5s0Gc/Bf6kvXCDbszRWusq/L/NEk74cQKB2wbnrsDOTm
Egn5JctzKZ+n4LTodyvmpEWPwSt0hX78Fc8Dxkds9Z8WzUlxqolZ5IurTDYmdxVm
N+Bl55uvaoO33omx5z77KtSaPwCG3nmPks61s4RNnyHoeOAvrRsmPATBDXReaFAj
7YyZO3U30kvyrzi4Rq8JTMFwnmLRHRRuU5P4mhmP7ix+Tlacb45T+FNaqt5//esN
hL+qdLhOZfiDHX7Qqxm0fsnCYif8Cym7Rkn0hOaN3HQooqnCAhdrDmq3iS3kg8Mi
dKpcAySqDJykxtkL10zMDCtCG0gcysiHyXXk1PhYaeM7kH8kdyld9g9Rj5avdAFb
ep1HnqMXSacgsXonU0r86FN0ufY7mStW2rrdrAgSdyiBVfHS/3KTrplApnsBRmMQ
xDRUZbrOcRH3AvrfHV0MgBzbC0PFbxJAUllQJb5NkHn/PAdTT+JohXWLMzbcYd/a
dQc8v0wQNq88NoNJ6kfECfSfjG94/zv7CwYzf3chc6iZ4745O0Kic1yIAg5XqSZ/
kveji8h+IRVupichm1l/YSRdJSQfc8LbhaXyZozRERd+G4vG3tDrJ36Zh7f3zDv4
y2JDV8GSOz5KPJTCAFBTEDpEFdJ6RZxMVKrSMLU9WU2vgGlZVW22qh3zNdUN0LUS
kvhRBQe8oMpVUr92IC2YKmchvWyDsbo0C/bI05aSPd8bGxtOWzn3PkVw0jDaHxFv
2iWaAvU0iXQC7wxCdvsZRoLdp/r7YIXPiXOhD9f1DFvPFhGUC+MGUK0LWQjPDahP
F1m+B4BYnCmCjzDoODlc+1nRBpLTDMsaGUVGCdAHPJqeFnp2Ho/k/4Tdi6EWb+8B
vTZt0dH3wbF7eBCayetQ7+/UjlD7FigFrAmVqJ9dvPb7mVdUO/EpH4IXCV8NMA6B
uY+neeB6Sk5tpwXmIVhEV0GBrjPB/vwx7ezN/qoUCDjSD7n5s7vBbyu2GVCfPEkO
y1Ll9pEWnCMTDABkD3tB0R6Sqwr7cD1zh18nU8fGTfGx4Ofnh0i6cNKMSsyu5oT0
nSQLiTBI/Ckk8DjnCTmeVywyvbSMgGib1/Wx/bRwRwysrjm0N2GTlxWN85CAcyyD
DXrVX8x9lG2maQjlqmChv4+jq3iytjTvWauEH30l2hgd/M5pYRO9VCAYD63maDeg
4QQ/Ilrh4HujDS1WzFmrUHWkP2qDw93AW469SMtOy6yYeAPv3xC3SCoMPB5Q7R3K
KoYpTd1AmFMtYroWRQmdfKClpihDaOP9UHHaIyt78O249iXaGkAj5p6xQYFm+iqT
lfEA14rNYS3scXRDo9E04v6UWS6iePbJzatlsAGLcGqqN10BcHEsPGfFHSdgqwdg
V8mGQ2IK972xIJp+q6Lfqpi16tdzajXXcNsia+HZxApcCSkp7wEBultVZymAkBCC
apHjuNrKdh/hfcAPJYSHpGUVocOUuxDTJci1nx810zTrL/R4r1jmqkHKIThNxRpe
NtsNhEcXEbez5WIwj4LhzCA9Iy6jCw8vShU1RpRl6unS0I185hzXAzIz4XTTce2y
B7wwwtS8Ur+AQoHKsnkaW66f+o2LwBKxpVlYXJr8d1HpkIjIyGYmSgZjS5oAYLCH
XA3u7l7s1ykbsfUDWHh0Oj701ObEuHQkUdiV90QNduE79YzaSCeDskyIAVRQfCA2
dLmF+vF+rV6QTlN85xXH7wWD4uYKkNZDrlH3R4B3VS6noexoUPzDtY4GXZecfOam
4vuSv+Xjnq3uHXG7/CdXLNXGi2ps5PTRsEvPOnGPo57x+HifoXwXMPWSQ969H4ST
dmFevF5UZDoCbHSsnffP1nI0sY/LKc/5vpK8AMHZwc+N9cBMUAL97qfnq8TYEQlA
U2nSafOwh6rFnSTr58J/zstW7+bWzDvmNxVxdnA0v87quIUGLLkUAZ12ZDe8qVhJ
Ga7jm7qh03lohGQWEjrkQLK4UiTXehl3yAEELtfmkUlv/Myt/m5+Sf7tbn4argUc
DJ4scXiQ3k+XwK/K9/2Te97ILg47ZNOAUueAZvoD6RCX/Nt74+eNPhEQyuJT5Ioz
3MfBYn1uKwa1v6yt1aBWvnAwmc5gJ12kgcJBRrT3H0mxDzUQWPFJvZCAurJx5JGX
VAxYAMmE7z4crjZFlX9EPzUGOHEw5gbNVP3qgKjG7n0QHls3G0VfW2yNCaxF1dSH
wYEa1LTYhdpt7V3o+ad4Mx5yZGapxflfksDSTNyspLRZvBHsL7ASyWxTecS5KN2c
y6CBBCMeIyQsz3te3AqA3TiVekH7/ekgSoOg2IkfVIQEk8YGZ5LlsXX4v3kFHE23
7QExFLjDvICf+2WVv4vdxllw6cKhl/6OBKFGr3g9O5CyIxguFDYqC3egnjD4G7qX
7GsebN1YIRWZk8Qo9N5ccXl+wvOE0ySxpss7GThzh8MsCVw4gP+TM/DjcIUz6bK7
J3kg6/j0qCJKjVTawCgJdtYGGgngb8+o1NPmnABx3HuefKlEhNVFCTZeW5r69lWN
kQqv/O6rncMB5XP0z+x9nc4HReqe/iUtxDkmcoeXqWrZsVwWCBLTKRpo2Ps0+yKL
r2QTVkdIDVVZwlnJ+xKPuoGPGJpZJCqZzIWiP3qkx+axQ19fTYJb/lnZxxUSJYht
d9/Gls0ClbGb4+fPCmNbc2t8ssaT1SnHy5Ihc0mibxRXAu75wF+Kr1ZnAAOCDnWL
PMfQEkDNAyFpsbJDKMKmGFZxFyxBcEMvangi7b8zcsOP4iPfXI41BUCWsE3ggNsD
XUr4lM4OHQoahybR0hdyZqsT/39oKKtCX/t3Y0FTyDiCT2Ia7QIKs1ByY1HewfHW
uSZZs6h6K89Yf9aFyvy9M8N+KgnzZIjRfXVIrL9eCjiQC0CC5gYlQfbZSs9QuwUX
nLxoWO7M3HJL9OvMAT8o65211qT4mQLfnKgz/IA4+Aed+NMlHZbHp+lZaPzfynv2
A2MwoNe4QjRyjZE13pJQaO0HJVpZYrFszR2nzCAhUiCmpnNE01/yIiM/tLIJaYU/
/535YJ49H4hbXQiGEZW2B17eDEpHIiKoB/amzQUPVuXl2vywGo+kOYzZiE2BavCl
JuB2w/YtFvIcwiRXPrlY951chIHK9MXWiq3y5AxHJF9ZCa+fivpKeO1c/7lAj+ZO
LEYOZEgDw0dJHPpD1lkgNR9zsu9mqC9Q3pMnQa0FaGYwnaJKny4erbCR5hE3t/Md
BWN+9jR03ycCfbI6oOOYENW486njhdukRdqf1pMm3FBSdK+fiZ7osjjVZ5P6V9w7
Q0WTQE2KteAJiThd5LHVaHzc6vnVIKtLbcV/WcYXs1YrxsLAe02h3odwxHQypTZC
r5310ubRQQKRtkTcMaA3yn7wBxYcBlekOlxrG7UHf7evfMQLFiB40pHGRvfzNJiD
nHvoMZGgvzhvA9z/DQIAY84drL4OQ2RdyJSfTtmYMaKbRjg7DuzRRWfbdAPe+421
KLyAPFXigDVTqxS9kiSX3spBWwd39ivkkb/+z9a8DpZbhv3hUxu09Keg70Mms2/L
mdBtFWK13fMiEsQXPPr4jKSnUIB8xwbUeaNSMjMrD8diuhxtlqGDDRSjz9pAY26l
TqWlCS6MHk8ORKOmn5/ZytXovNkF0vr+ztUVu3n96gVYLslpoS/soIB7vpL8gY5j
p2A6I1KmJqFXTrQD33x6PbZYKPxEcrYpxVu8UbswxUCuvybKpsAqF5P8ODLAwgjG
jmZoX1LOz0MRKbh9qWXyBiE3DiY79xXVzpD1tpjmzB6Gy+0k8wlZ+VCSMDzNk1sJ
EmK4vN88O2pXyl8mV+QTIVWS/gFmF8Ji3yTzy1BG9ZGBCJeCA1FFerwm2Tw2F02h
A+VHeKdev9n+l93pMEQgtP/iQLt8MZGIwfEONDwfulhim/yg0AHcF5/qMxMCXnn0
LmHIsZoDkU9ntzwYYtFfthXN6AX1aOJIOeekQ1Z/ezLchc9fIRS+vCrF30R5+Ibm
K8B+bPiJVYscMjUDoS9ZlWd7nwhr2wOh60/hZBhtIceUXQaQnM8tJonokoIovlzr
WfI7YN+ebGNaFmj4jm8wKIZBUaqKlxk5hNYKSkJ1ZKSGwW8X0Tw4KRb0q8dkN8/4
YofMsv1QfVZhwBZsr4IomU6J2l2UgF9WTBmG3stu8Ku3GKHxfZP1lM9tGFUFzMJ0
zTwV6r2t4pAwuE/oWDCaED6t63u7VqN7Bngj/bdcVU4fzChtFZ79qmhZvvPqn9UJ
TsaNJowqkP1IoyOFKYR10hBHieixZN711Joy7A1Lg4WJWiU01IcARadeRlPNI93h
ECsGaqAssBO+jaPDuJNRJQN9S9KsFhi9rhVYWrmzm2maRxRTKNHp4lGbIusz6rw6
5WDclLSyC2jlybXxor1xN+7TrGpH0800E1JofQGxT77MAlwficF2P/P1zUfQvgDH
DnpyWxtR1Q7Yi5PZJx/DlButQTMegiJ+x3vFINqCNOiWnuVpEui8SyoI8FvZTms0
82tOTGzWsfkwa33yAXplCm6jVOmUKe3zWiHl8vg8WZLzakSFOehMWiJjBMhesQej
ZqZrQGsJWA4ARM7igPGTlPS16kJ8Wz8Spe+GF0H0cc5wr2jPuZxVfcpOkMgXF1A0
TQlvMiBYPHs8j4sKBpOQrHhuPCC/1vHQIlJ4lm+u54f37txC4xaMK/xlijwjjbpo
9EaSiHoP8R02yepLABlHqp1Zxe2eY3cgObw6aOk2qdZ6MfhYyLtzWubCgEHDeWgw
SCzE/eqHrt8LVOrmYPgau2M4H3lcyy0k3KHReV0vP64Azopjr83GtF3N7kpD8V86
BjG3uE3YiALkHC5ySJ7gEFUgN96YMSNf0G/CHUq7PLPLw1MbjNcr7Jn2Er4/MixK
yJ5OsXmYj/N8CJiiIX7+cEKc1zHc3wDq7VhM1kEX7eJxS1Tr58sg5CVxApwbBXMU
BnaxlIp0lL8W0LsUnK5v4Uf/PjU+AkIXFokv/lqblaTwFPN3Qie5Qb70hnWvVpz0
BHBes3taNrZ7sSkrhAsVHYkj8PRS/8/7DJNOgFKwId9xSodB6EizJhqfjJmT6n2E
5DgTP1ZEiDzCeqHYVc6YWZkKlriMV68aqI9T3CDV/XDPj2UKrfKCXA8CvVjDMRGo
kHfHTRy2YHXzh4w7k50OKePJg0CRSsPfGj4JnJqwnmIYhglqxomz7kWGIUB12YEP
crRd5ib9qy2eSvdF9GO/p2jKoXsRibrOFKl/bQX7OVwlGd7WSISdDGO0tOwI5cn9
AT8wVkmSbVg6+UF6P0rVVUIMa2w+oUvw19IGGyUmF+oW8ivWAhP9cha0mbmXE41l
qiTXZ9uKTlmRbXzb/w0kwoV0i/a8eKJh1B+YeYGS1sOHO29vgcsMtzsjATkfOfg4
mrzP2jFeacG0+ViSPmFN4vLcYI7IKGL7WJU6+xKKf4GFfo8nR+IkqKP8HEyhvJqf
R8sY+ocGMgKsG8msdh36znodvPI8zAEvZjpVaTaNClNkBDxqaVkPfDffLQDL4zMd
Ie1towh4eEaocvNWzuQOoJ9NOqh+1KdXATg+8/QfaR0hi8wDKxwLqCxfa54/SAcA
vH/olEB2gkVJ6/osxo/XTT/OSBKEb9zprq6bs5GbrbxSw634zXKamS54ps2hJRa2
bS292YEmsVL72IF7nOOoCCN744yRVNespp0LyiiElmbRvKQT/PA2DjL1B6rX2414
oAOqntWlvdVlBw6mNkYFzYPr6tyaygOZHGaNjPcaPUP63ZebLaDaReJy0pGi0jam
dP9rSvHPlqYu/sqgWVCSO1Y9PRGZztes8uSoTsu0JapLDoiqsKbj/znx2dXvcsAu
ciDajhnFAXRuLT3Xi4aULJICznHNS5Z77DQNJ+igLeYstNUlgxuzw7JCQ/SEwY3+
KOK8dmg5Avvh57vLMlHb9hpIT2JjEatwxvyz3E2fIZTu+XtSW6/bGpGxRlsgK8me
pvptKLLbx1WJUpXIu6W8jkdjh78tboZNwVygmBQtOy+sF4y5rpUU32gZ9NMwBUsQ
RnbAkum3GhaZfuVhfeMPI2H9dj0/P+L3AJCcKzlCr/OI9pIM6wJ5bpSNOt1Wo/Gb
1lk+2+DsgglBPUd+RJyTUyWbbsJOIt5G02u1tcZWkh1B828OzlQwE8ll/LG+rmDX
rnU/Y6NScFQubrJmncXFnrH6ljO1lM7+AJ8P67lwl43ASFslbFGGhNJiIpUF6vdf
TmJWEJgHvx1GXg3p18YTgE0C8cgK/Ms67aBXjAIlTnVYIoZPjU/cpj17bWKILhYf
l3X4nnjgSVfSLeT5y9qoR1md3FxHrLbrNZ+jXlbV4DvM+FW5lVh00eTb6LiYv6uP
VJSyVlVY1I3gSDLheG94HyE/Jp1Fa+f7K8Tgq2zje4IOTWY68d2NYcdaUr33Drmq
hoKKbSrN1eAJaFPEZ1nBDkWzKQEPXGxUIl8bGhYYSyWTSlfe9oWfWqLcbegMi/S5
3mWveh0oxUqeTwUzHCSrchzItx//HlhlaXJyN/Wl/pUAvKiSYUG6vmXElMdeziOh
mgCNelRp/qZOXvBOqbJFRttfKSzTAIVDvD4uN/3gWAXiCREGcfrciW8wXOPc9Xew
thWehgZcbJY3XcdRul1u1WMHIj19a392o9ud82dnyuhyYINmpeF4Hc5HYRbRAxtP
8F3yM/z/XXe1zXoD20LVi9ZLCh6iw0qByMY2r6lCWMWJBJO2IJUEZ8fYsfK+BrFD
2LiKaJqdnp35YpSUInGQvrTtNR2IXNPayDSK8b+brRB9jmTXvdzi8lI7HDSOQne0
kkcg+mEMQOUbDo/DhELOaKHL18ht47584vgYMwAIfCPO5Z+Xl8BSyWeRFP2afqjJ
bAoi5qeRxMpkwXI2PNItYN8EhLzai3GG+KF6+zoPqE2fQwr80eVB9eOIH47XiOgA
gXMwzdlTUJEx2QobOmYxcShAKiApkjoTMo/UhsW/8Ii/3rd2rEc1deVKjqHiHWaW
juu5omP2QWRuylVRaV2LK7R+DesEjlg7oSV/lGZvj1MPxdM33CvCCaTS5bW4Ymaz
rFv59valNFySv4bkzs5UsTiHRQ37a5ugIyyuTLyc5FDscwavwLIaRVgBRLRUCovM
H4pO3R+KWsrZExBI6ahiJV0W7PGLgOkS23ZyAeE8IzMRl5zANq+vN2vSpgiwyPUQ
14C6FU620oHKUu1VKRhCVw/AfivLeo8Re3njzfQ9uc+QZO23dm/dfOGqAl2fhs2h
SCyzTszErKKF2QvoZX1f14xa8jYsV86lMYOu0eMRNjv8hR9hQR6GQtAvzyRgNXfL
4aBfcSHsD0b1AIiMVcmAAGvWBlUvCFCQY33yRhcrkKSV/JCpYeizrlj0G9MiRVkA
LCsFYPjJcemb8OyuycLbgP4ujPFmraJLT59mLQm60plum0cvt6sCynwpABBKTa0r
XsO2g8VkqyJAXpmJZuiu55EIFONh4ZterOwortdNULKbuSD7lfsX1GzagYQhphRe
p9gumbwqXkkDz+clW6osCvnHIhgq77hg8X3p9l1D+EMpu5pRE5+VuHnhuouUTXkG
hiCnH8osaf5JsP1Li+xRVdijGsRsNHmsJWakwXxWRpn+TumOOdDYf0moeokch7Yu
vQ+DNdsT3KWWcl8UsUlrI0f548mGlw2zl42sjIFe8cRjd0Z7jzjKFcJsx2wKyHt9
TrvOupmmhScyMt68SdfyKTrnHL12JdHagiKxIq3j0SuiNb/lHJMh8M8uSTy52owP
AI0tAJSOc+Ovp0biFwgbu1V03R4+RvFGwbOK3IvEajb05lxyDtJ72DwwtWCJX3hf
ugRXkHkcIsfZU6hfscHGIsgeDrMYwh6rn49QTGvAacXl8ckF5XofSAmxCYyO4oXs
yU3LKw7wgtXep0qfvdFxSb8EjdI4dEi3IjlWwKoJrZU9qwXXO86NtUqAA/CQFtgq
ffz0DRq2glSMa7hVOq8gf2Ny/qfnnxQUpPB4vKdeZRHOzFw2XCcbGlCwCYHSaE/D
dnjmZo9EsrrVCl3kEMLNgEhVn8drBPc/WSuT331aVv30AupOu0smFdcFbFHXZed4
05bdcR3tjVj/mSMi5P3dWMAPbHJ7QcIEohbzY2f5HnfBvP28YtLfC3T6VPPE7/n4
/EhWq75rCpa5oEqOm5Xowew+cKed/cicMnxGG9SXNt45RjN2oa4NVWXa6gQV/ktZ
Aqgvd9sbeUS+15H1FBcrU6Lc9ObZVAeKUkbtqibjkkrzkGuEEICDVVt6iD3ESeDq
0A6xBKwfLQsSkEOCXjLyJNHmOfoaGSOwnQxlAVzn9u+d0lM6pBkSZnwDpk5mXWLp
A5eev4/Ta5iCifZtTM/zTgzP1uw0q28fpIbaMYnuGA+APr3jC0kG+iAakKz30n5e
RS/Cq7/D6qxNNxA8Oz6ttrIaXNf5P7eHn4lvWQRJAaJnxBsp98AIaSyH4zmCYvPI
wLEI50pbKiGWNAdUYEP06sgDHxAyqWL4r2u2MU+sVAwN4yrrT6W46DDx9/aZGpBo
HDLJX6z1cc/OKE/moZE35UeQZYmMY1apAb/J65Wm33htyNSy5KvAY1tC9jCvns15
vZK3eO54muj8o/kVnI334jLLnnSZPi4xDUZR4rq0D7IB+hU6Q8CP3JXIO1dkIJ0B
uZxqgLu/QSYhCKsK33IMw9guk3r09sncsad50boIT+Tb9B2ADG3KnjTTdjNFjFAR
bDpElnfEX2PB8QpiVAQgatFlToROzI8lDr+emGqP9NOUY+JU/bZYFiNa/JIutpd3
f76m7UiB/23Ab2IYxPZpo5hG0XvqRDz/yD5K0TMJGJZRM7FgIuv8b9Yd/BA7Vf4q
8zcAHAUQGK1S9fJnxw0mKY7Z4I3BRMOBWSx6PcDHzibGfOko0sl9h6P7aFEeXxRy
qunZts+KOX3rZLDcfSoG2RkLKuic1/81KW7n/EcUXdYGtl4B73zlXX6vtUBO36xy
BiFVrxq55mcWJTvwYI7Hp0WQ7sk1YxaTP95wlAIesLC+Gbfqt0nmKeU3SQ67NMht
Pl1urph0umhjXbhU6XR+5fenb5IhDUP9YAyg9ykha9cBaWp6yWthLLao/ySvvsmr
ONiyNwF/DkcarquDVHt/fO2i3YeaVT7qsQSky94dehVQcgHbOLaVEi66lt2O6sCo
cNbb5PNZUTUl56Q3zFB+6FLilEOrtJl82027Cf/9Xubc/sijpKntNmh+XQrrPq+V
KcsyyBduDM53Xlk3ZnSmBXc2uaibEvzRziVCU1Sai/PEnumqt7kzxWSy5des2/93
Qznfmm+WNry0G48hF9IFaVrzbEQb89/T6c77ugfG0Swxc0Fj4XbHIU14+MiKFYQ6
YyNY8QTMgOuauRxa8Smu9bgnPwdyla1aZvU5CDu80IAQrHx/naPwIorKpK26jDmi
zcASsYXQGHWCtAfQN30QA8xWW0QcGH7Z+AQTUDec4O/lJVhWm0VNr9rIdwrI95N9
QMIX0RcK60V04Vi2NhJC0ILSVPCEce0aNrB/qnpYA6cwWInmpqcXFAx5HLzs/veD
sVuCo2Ipp4/A8dtx/mLm4k0j1iXiQS6CPqbwCc2TsrhhwDkosIFtWNraq2CcyywX
0D9MArAgAeOhvTvN2IiehBtMJZN5GLhmEPcTxaiiqJMloemMkxxPmIycpPQNoZL4
2S0Om35OC9X4RI5V/yfRG3npR+iQog7vByT8iR4/Q0PK9u5kVaB5xa6KMiYYVxcR
PzFyiGQ49gNA/O37JXwTRPyfE2IqIz0JjIcbqWd1+knF6v2B330IibMun2yvPltL
g1iDx4TksjGFd2kxCWT49kE8YhLO4bUNpQkdjVSPdb+EuHjVBZ0Htf0y1VxZ2G7h
A2yUPQloJI5SnawvSrFupIcY71JaaZy5A+F3k+Jl2J+vDA9I+bjoz2tvNPY42sXl
XGFQRLsSxJXsl22gU60N4vBpPvZWzLniQuMuwIMJ4RUMyaVE/8XYt8qeVhpPX25E
ltSGAydgdGptF7KXQd8lq5o6XJJSTrAlEHRHAkA3CMzGQos3xkf0J/F48mDL1fp5
9+OeMQtQgOE7qIHIFZAOYMBvuRxqc8YAb8fTY787IK9GZISU4X7Z39GceUTZlIHc
MhMAiDXHlyYAlmhz5x4mDM/tiQcQMbrxqVX/Jl7DQBGx1U0I0zf9mBNN6GupDJaB
ahlAOm2w4pxkXw+2W70SMxjCFxgx8Q9oLJ0Z44oqF/HqPu/VXix8fwtJzrJrFgTf
mQpxzOny/ArNbbsXjyM6dIP49SsH2ABoz6bmyrILncsxLV7OYU6THlvUHjh+hhvj
9GCdQZ0DdchSMoBwJQXZ5YKf8gPIjrTM1PA+tiNPvkEcnDIA0JlpVPt5B7gOcUbZ
Z8pmcaX5GF+IME4h+ivztrqX2xtgQJ+LA1rQB4PMj9z4zDk29B7T4Lk0wR6OPlz7
L/IUJ0ginZ1Upvaywk2uUYb+huxKLqSZvZMe9CLixdln+Lf4xxSL1hKRDzN4wuam
HQBMO7Nat0Ujc1+pXZfwDJhBKtZCjcvcPyITcvPUejVhJeP58O+E2OhoSP6UF3oZ
Pz5/soDpTt5sVHMYZo0EopXDPFxL4g6+ZUmpsbwqkkI18yzWOUVFEwOHDnbt5IzF
0Bz7dW2V8wlmn9s2TyhqzjwcSa3eZRNVP7z6Ya6ApMdQ2HrUqfO7vikPdidy2/kP
tSr4bjhdmKOe1BNYbXzFV99/WiH26YJ3H0uv6/PhVKQhEuSs8MHjpNoBx1FhtCg3
aSPzMFoiN0wO8S2eC/WuG5KLUqBpvm0JyYvtioBi2qjrgtLEO5DY8dwYHVIsIYTd
/vbvIM/yApOyR+8uKk7CtlFdNFOl84d//3IeOtUpgHsk9gTTsB5jDk0YRlq7SgdO
d7TvghPjpyNqXM9nQ0eAjKZIzO12lmax/xSEO/0QfZJq9QxKMLHpTg2xjyg6koDf
F96gSUeClYkpduSZaXuHwym2YKaDNYnkkfwUHjstulZbA6zwn5Yd66qLvTx1adcs
jAVscZlwxEjrE2S1BdGbCa68tDf+kXqq+t8Hjae7EkU6hHh70gtQxCSt73ik09I/
bUqXKY1B4jeytujf7fy/M1z6FzXGn1wumR65jwJbhza1wm9c2Vb/YeLW3WhnQqFr
pydHaSP830TNR3IqmJUhHh1pKoo7uJYw8FfY6UGhxhFx8TbDqfWSiDJ533oUZ0gJ
80ufp+8n3XpjQhZTZpj1bk0x6VJtOJF6JPzuW9d0hS++8J/FCwtJWZlpCni+oJsx
AMSXiw2fFT39gyrkCdEfqxj5oJwtuBy1abhcG3KmnkzrMSyuC9gAXIzmSwZcrxUC
TCoJ4XzwAG/F9uXEUljtTL4z4AaEKGaBw1u/nyZe7mVAbKsSBkaQJQgiCR6wxjDQ
ORqzs6Cnd1Cck77z8IdFkItxFqbKUSm18hf305x77ZsXYJQzpg1EQU0WR3zCMk5g
UaOmAoKZBDKOt2nTwqvLgHivyvyjtsHFTspirmXoWxa7usEpVc0Xdn80hHeG0PnI
E9SbjQ6FKwaXCk4FMzDvmHLrZ9ti/1j6VR3hvFWkeWbN3ND7K35CIiaHPMb/BoBb
MMRJaEzDseasjc+kECvln31XWLd5CfVhIIQbFhRRO05nQ9/GRbfV755hnXWPcC2p
3AgjEWfTNvkLmaZVmuFh3X6aHs/nWUTGMji0KVj5DxNKcc8KV/NDpSzFkqIHcYLu
R/6kjp69YWosyBkJJ/mwZrxiSyt7Qj5sJsW8epzjpeI6WQ8h2+KWqU6NjWoUI+kX
uPQq8WFpDiJs33zpF3eXTVIvQxdz4o0LyL8gs9H4Xwj/eefihdOx1P+so4oq9zZR
iV+66GdA2n02vz5O6NPY2ZSWCK5WODcby+O8C5UK+F314Ck/2HTzKhm79R9X309n
a4rJZ3ZcSLkMdjntW+Pj9czWdoFi7AWhGWC3Vph0W+mEBbuzY2if/qOk+tTWakx6
Vi8M3be6VdJBXrjvrhfwx641Aexd/uYEHHFyZ2wwtEF4dm/5VbcPTTse3FXRr6mo
TcsgtFX5nQHZo+Bv0fHuMYQgBnlpnF62ecsBH9a9CL9gq67jWBQnTznsxRXC5FUt
Ggk6Kq1cGsQGi2qnrYrYokjV3brjSaliK9tfJjpXoo0/7I+lg7xoiEblS8umSXgU
uYHumoaD0cX5O1fz+QaVC+eH9jIhYGe9NXkHPbm75jGSOtoEJUIzYlsbkKM2tPD6
GQ2w8UBNS/1dE/4c4gBeI6iegzjaTJlTLaaNBTtuevwVyOKM83NihB9K0VrHnn+7
CY8MlG1uDv7jRsJRu6xQ11vWSMCgQEpte9spvfaxVy5q3hk2glyuOj98FOc88Io9
JVBbvbs2qIVcyfa6wJ28qAXa9zAHfFX41aNcWFRvr+r5w0ZEy5a/GYZw864w7dII
Y5Lch7KAt4HBEu/H/21Gbl44SZIovu0ARkbj0GgAtZ+dQ1vQbGp71C00SGAgGfhE
9obn7ZNXz4OPpaE4nN6x0s57CzG28qxxxhQeGRSgPdnsDtOEYbT/PWOQb+0pl9Jk
2azwrLl1nLonLoV3pS/z1jyDDa/14zLhNVzW4rWsc17Xx4EbQ+OkDbXbkre6C4wp
5Hd4Z8dMAV2qEiLgQmPQnwazlULQkmBE+JmqeV5sERc1fmYI3n7CUWv52mPRsIp2
X+g7fVkzEkP0D0o+dqQPe5Gj3aM/IrX1kNUEz4jwocgsQfRaPhOmUaGQiIDL3Fvl
FrgzG59y1iVvQDe3jpnsNrikyl2joNuWofmwg6SQ+FYHBlCCXF2mDDAFE1X8XqCv
Wec4U6mfW4a11TIi23JCMaUVjxG2jjHwlmCUwyGXCQUJsRCq2QRhUL+rMFPzEGgt
NaNAXETbbTx/L19WFRh0oAhZQM561wm2ex1etbfsFO0iw1epN/sqf2pJrCqAGKbR
qSM4T9EkChzQkuwBJjefLQ3J37rqcvKhmF3RVns9oCs9IkXkOOst9llDFSOzfDvo
01msNViYso+O305swYylZx92KJv9uIhYzSU8oiBlYh/fU8WkTXNVQwKbbBzPsNBR
8HS/0Y1YCQ6J6MADLsIpJkgxSeEMzTnpEEdofCMajQzEQfEQ60gS0MDvhjq722tD
kQqyMLvXYQ94yTJX9cz/cO+yypF6FPqbhsWdl2tn17SiZ7/eLzcy6PTQK4YUBpjT
hjMU/fmIWg+xqQpBuz3NRZPwblSwJWCPGehkGSh13Cy8kzQ85P4IIe9WuKiBIy88
jltJvOcoj0YHqJU8HFYPLdX0G8qUTNtf1xtPQIsteCk4HSHq3uw+lJsFgYOjGyuZ
4p/RndiiC4Qr1A4Wjp6TDPmInXhbslSFLTakMZT/FUKMm2Equ+TYd9CDiAzWzVKn
CeH3KJ6Aaff/7sP8+psZZFWEhsz9UtcNp7ZU/EI1eIREC5IyTLj3C3xzCXs1KdSI
AwWro+ZpDkWH/NfADooUzqoTlekbzxf8nw1dXOQjFr0ryQUOIOuVB+K+5IvnLVuo
2zn0F6kcUXbpFDN5ZiA2VHJ1Rb0ryXlwxFYSGzfcaESUbMAgncUXn6eTcS26KZ+f
ALaKAKRQkvCdwwnR2pZONo985K3qqIBHzk6oVD31AzYOl1FzLOJvb48GGo3uHvBw
l9chcSch6y27Uyk/+q20iIAnbCtzKVLTmhDFqMbH6kuOKy/W3FdT2VWQ3B9dEM4A
6COUUOS6ozcLLUkT/oh5q8hFHofWlCF/7K5M4z9VwJq0QGQiLL/pUPMEo5Dbnex9
GuT6yPRXbhCQDzjQ8UJ1yojjlH2PjFcwLG4JDecEqotqJU2VNFHrGZ0edDf8p3SQ
PddZQIBRVgnIMFlT1h5HPIdYNfRl18/XQYlL2rFDT+lqStjgzs7breTiReE7nYBs
t6iLzjNoIWpSPKeDVkW//50ZzJT1EWDKUPBFUs6KyXHP6ge+m3eDjey9w07Hy4Lh
Pti9nkmrmC9nWfefUZCzZ1KiUnbh6SaqjlRAuWlht/IxnQiFDaSQuppk3BPUNlII
mVdTsHDQlWZo2pybsdP9XGTuKBH7A0XtQF1AXAe13tViYBwHHkBayfcpZ7c/SVuM
hYu31w5AFFcPKJQHriuX26ecPKzn1wY6Yk45c+4FzAgtBS/XnregZ4anNleYNvd9
F7WZEKmgCC/20L4SoYIKwjsCpp+WGzfRbbhJNqCUFhLQvlNZFBzTnNSsBPVsfo6g
HcTA9xOGwxKl9uRLLiIGdXFO3oJC3JYtXmE5QlMCnX+Ccpu9LCPDI1xiaNW3AVCc
Ah8IL2FmMp8QjTXW2EdY5rpEIP4vDCgzUvCfQiDqkYCEukHRuim80s74wwseEgDI
DC0x0LXDzV8VB+11/ejze0aiIKb2hQZe2MEapY+OZC93yAnWSILdo5Zj8LWylTDH
o92DcJgK6mWsBNEuUbn0y/qizwTcb77mJxvl+KfwQ0jzQ+YN/UVOBdnraFVFjhFy
eeBsJg3dCmm7hKZCIIhubHAoGkAOgdjw2zJoTz9d+zY102zluDjIaHB3DfJGdKaL
hMPD3W8A9tI5ZETMRTp0SgZ8RblbrQLYZ4u936z8516OlKlBXKTs/yYLZ8zjk3P/
suL2DB3n/ZBmuMzG24JuY7HphhtmxHBvy1EVfGALZ5vLO8rTIaV8CqNjaHIr8Nbj
Ojv+2jvO2Nn+GBLSa3ZHA1MlbAULFEMgj4LNE/4AQILptqlcG/EevBm+V6omuaZD
A2LcHoTqUiNctpi9XniTwmhXtEolBomVa/Il1D5aJEq5JpaDnkdsOAcAqcxCakpG
el7Akz0CfE/bi7bhE6PYVMPf/BwkXcPXtL3I1i9Za0dwfcdaQQjpT8Bm1BFe8snF
ywUGR0lhMCQyZtz8iD+hw+4ylZeNgyKiLdPUViwMH2gQPKL0v2DwX4q734YySXY8
o36ty699zxK4LFWDqflUpP4/alg2B+yG/kjaEUjJ/R7vtYz8QwP+/o8vKsnhe5RO
VL5/JaAF5SAyP8GAjOA0+Wnve6IkvOQvXxPP3ONjO0RkV7fXu/x/KxSgpJ3472QK
a+YpY1QKMc5zvYXFWQKtFiRmK47w3GNsYGpkvowwoyCQ4YlAv5M6rs8R0RCmr2Wd
5BTCwXcuMclYQgh2F/bayIxL+WLsGb5n1pCz4+OOj+Eh+9CkBUv5IlM6ppETGat8
NR5QPcM2oByZH7ucXSkCqYuXX0Xg1yLoMb0macxbvvibCUZ95LkIS1Kj4x8bZCTh
MRMdS06TCNWBlxYWNU5Xnds+s4B+jCOSzh2Y/pN8tuJwyFqU37Ur31NZ3i9Bk18x
ljG2FxFw0MojMpH4arLtOdEcy5pvluSvxuYDc0KSAXfZdvuFIPXZxYpCmTg3Este
bZ+RuzOkF3XNX69fLyLMTD+gyDi/4rkUu5vhVoBVln6EgQgeeEHIgWuUX+nYW2Gy
T9AYzmsPdqsJWT0BzXPHL+4V0wD7iV22/OPXiZIs5kK1b5JmXvXrwV7HwZcVk945
AFmk1PbFrFpX5PjicSSiGNTGU6qqwhtHQXwc40LpHKXv8gULpu4wtXcy8CXau8CM
M00Go5QxjFcphiDXirXaX2Uqb0ekJkJ7rWLqfIex0okZh1Is83ba7NJpuEcTkCxA
Ef9YyJU5AtagGisD0z7p4Q3SJH2bCS55DdWc/T3Z5LhteQ+T3bNgq6yKl2hc027c
2xinmSBLUV36IZraLOpF96mzdsP6K8lnUOxuPGkZvOwHxyBk1ighx7VfNXNDkyu3
+mA+Xf75mrHE4iQSY7jaZjeNS5feoB/w7JTRHLPXiiC1tGS7j2SyjXX76uOJ9IuT
os/DTniS5OvU1cPgBtvuV0fQ70PpUEP1HnNuiSTvsc69+qmbeJvtInNlERO/qkZT
YcaaBHsSUdlWbc+HHTXyPA5g8HZaCC7tXuF7sagnXQ1LSNxoz+UcQ2u2r+xZz7v1
DnGfoUOpeZEi+bH8BCx/tEG3h3rI5AoEEH4zP4CQXHIw8LAeZTv4OsaqR2ein6kY
HNyeK2GTzcHYBTmwi46Hkln6A28xHBUqXMMfL03iwCirXbHb9r689INCXBQGQOBr
Ac8ob7B8Y88GwH3icVVDTrhTkPSVWxApP4Ef3I22WiKyaWQTCqVbcG7B3y/bEWTn
uwHwe5Ot9ayeMAQ+283oHxe2M9CBUdDBkw4Af3MBbpfi9gUC84ifVm/guLjRbTtt
LSsmUhJiPahdRA93Iac1ofqwoRWXsHuqrG7ogyNPbK+aElwAyg8eRpGAMlw+pJiU
euXzpixvQyFyNSdbpbURioMPv04L0MpV46TaLXarPWbDktThPXsLCric1UMMy18m
dzaAuRzEX8rl+BaPR6biAk5Jh9I15fgojNtpRMqnU1priZrhKdJr8NRR2n2zRA3k
StmTTNQnS6hugMMGAgN0WEQHfiz628n5e2yYl2DMJ6cYVo0KT5XPT3SenFYsBkun
31DQ/5Gk3IPi3SXUHdCxCsdbyCy/ysByt3EZAmb/f8SztVjRL0ZxrFv9aRA92/ON
sYbtjPXFw7ZsQEaI7/VUxMTrD8oIpebosCGL5vT5AXWeacsN5E6pvyXATmUJOiPq
uEL7zvNRVf7FLfPduvoUc8MrOTaAfljeFU6VaHG1tje7vaUtY+OAnbOUow10z9cG
+Iz+09xjqtmS3C6zp5SeDTQ+nw2mDKi6E2qCL2O75s8723XqFcRPDgaYXvU2tHUq
kMO5N3MeyQ6Ua6zRw8zglhVyZ4yhtRWYiJ/2JIxJ56xFEEUTQb/fCHLCxk0P9xxJ
dCh+sZkx55ft35WDZM7+nmVnYYzKMsKEwXyxA3ggsB3EJfSYtVDnLqbk6azFwUNN
Ld3EZIovBLBPAl2mCHaI4A86KPiYQdZC1Gv8GrlGtWVdRqg/NYEAbZj6/4ccJbBN
31C8mSkIR5y4I+dDM4M+IIASKZBt+IR9i4QVITOOB6AoEUNlRxsFlxFN1oFyoS+2
c8IWzflXsgJwOt1z3pOwivToOlDLmEoxuIYA+OAJMD/fzkP/uLjtCsUTt02+k1QU
JTofr/2K5qhdj/jy+kpzo4W62lkuiXmI+CSJS+MnZgAYOOJQ5gxTBLGNBXMg8N7F
DpyeKPmfSFw4Z8NCIicLM7QNagmCIW0hzAfaIJtvMKij16doUGGVGgAIWpnyIS5n
xZntz9F0aH8MCoWXY1FOX3SXXp4hsfN8QD2DVc20W+2pYP+Z18l6Ld0ClGunCYho
HZHm5DsbFmSV92l1zxVhb2nFbPqzUoEhoAt5mvg8utU6Me5OuYt5/kARuIys/Hk2
Cd8/GZ0dmbTBo77yrOjn354T57ZVsR3p8fYQu1m7lfPrFKXSiAqBsYqbggMF/pUP
5y6aWyqG2ttFhyH4scD3TlZKBlAPqh6/DSvQWcgLX55vAVYAk08tbKFx8zuxUuDp
zuupAJDDosytxAwlNJw1vSB4ZtEE4iOv9mA1OscDSekv/NjzqY13yZUM/jhYhpio
DSoiam36/nOAXtOApDyTqOiJVhPnh74wQanb1rsX3AhgujVopjd6zsHQGUynIf0y
YOKiPJG1MyHJDwqwSZlsf4xfgOCLdP3vi5+qvGyLZ5wreR+Wgo4V7xLU0xKUTHAB
BTQ6ouxyjZIwpS+BxsBlV0Pme/oFmYDx6VnIB4xINqIg9P7lHsKufkt6CUyoomlP
3fagmLO6ireITlUrl4KBaOtTPa+zUNaG4CQxeOdsi7Xz9/lcjILPl5DGrd5tHmZ+
l1hymm1O2Kjg2ExTkJYZdMLUVpvFXU7r4yK0Lf8Wt7KygvDB5Peh5H8RaZkpyITY
23Ty5bdJorWVdU+QW5fFKpPthgvVX5ZWKi8iSaqyQMLnOaQgp6nBDwVmh1u8LGL2
6nDtUUsVhfP0F9Udks9SzzYTZWr5s0XgIoOiippjzsPhJ4JJ4rAapnu3c56XGfgc
ef54FdQFEn3/+W1vqRXJ2GukHp1zU4ZmBSPogp4EF345QdFTF3D5Zbty5uymYkhv
qto+eEFXJjwWQm9baH3P7HgJz5CHUM4OzH7U+naf2Q6KQT6Pe0YB96ZSdKnNMwDV
HRoZQTLnsJzAhyvB1/q1H3QaRup+xiwfzM860Df/yzqDVeDKkkzX3Qm8vmwGuwvc
OkHonQvcwkUUXAvhOGee+FV+sk4ExTOdMqAMtg7fSlEJkXFpHk8jLnbG3lVmElkE
hBPTLrJgy0MA2oqBesMjB+fh8zUiB9pocxG2r/WXkQ66L7me/oDstDt/gz6STFdN
OrBlC99QgQc6vsE6+afCNID+3oqdUET2L1sN6L+9JjUmhJOHyJCN6PXNh2yaZXYm
YJGDNGmS6T/gmpy78+Riy+Hnqd40x42L3sJ6rrMIUQE6nBcu9DKEBG0RLXMLQ6Ek
Ll1SqVik6P8L68Sh5nXOuoArh4kFYLdS9j/eXJf10iK5iwS27+aaqdlTxSyVWZcd
n68yYqKfdqS9Y23HCC0ak8siIUxM9tGYVFZ3DfOijVrYee9hLEZGf8KrkrQ1nCGX
q2mk6Nr6R2NcbYFimvQntueLJbE4I1b5PsRWf0/yvAgJ9OvEbjxPiFXKKl5yaMdL
/bHyslyzG61ZzEht//VG4hD9KToTaPArhs/vIayR2OfQ7gY+jDRgIFmt86wcXWgG
vtgOKADzqmjVksql0qV3BWK6WrIlCiX6WpZ+5+AOvX9OciRaa8igl7qrK0MxvKDd
w+CB2NrmYGjJimdDDOXDtpXcq4hG+pYcESyHesPQ9ClHFgqJX59n63w3QMKthX6S
XbeNaabmQULU6VBQ6LK7b38NFy/sjurVquY4y70bOD8XtEiyuExD2f32y9yQ7xJ6
NckjfK8B5EYoHG8bmHqXF8OsmLHKL2DVYVr5C/Vt1ZOlSDT+ctoaUDA+ni8OVW+z
d0CzTgEg36iwIxKb0vjB5ekqjsyOmjxgTWaKARAXCdcqUUn9eCDHUYMeJz4XWlrf
KJIfMjYcJDVvvTDUWT0Ql9iRBsouFOVwb3zR6ZmNJiOheQ0gO9TwpUwAmQ8x7Ku9
rblUM+plmcRviK+GRnA1IGDmvLeR5e789ynj8gS1jMOVHYVaEgYzpqb22/Vt66An
V0NbxgjIINVbm5S7G1dFVudWSeTqzlXDRpXK6wUHdwrA6UJGAQHo4n7beODKUkBD
UKh+XC+lFgZJ/YAE6rtwx1jmn57BJxkR9hV6vwMTc/NfpO9lNhpJzmsqaj4aevQY
T3qnN/B1I2x0KBe2ejH5r83JEgVOWuvSafjBq0X7Xs26koiecG/reN/zwJGcmZhG
Nqrfqpf7G1HY4K1HeJFciqVK6Y5yH5RaVqOCbwQNyRPclPE7/x28FsdKtC+Cc336
AqqV98c/43tbvPLH5LbxHpyZF8bPIGZb5CPWqkvSCL67ZDlF7pC0VwVt30rgPl1d
IGGSBWCX4hw5s5J3tmrsJ3+NYWd6voj1jX3Y5J9LftB+G/mpeKPHftdfeZ+4PsoX
CUePEkfjxfUodJOM0WITY5VSys/vSnCl1jN8cvrpdIxWAMGEL+xL9OHde4fAVUKD
ErK34UqqesxO/H+6rh1WFkheEGh4SRLAtVKb0QQ7c7evkoGTFSC/gpwL6Q5XdQhz
aalzgnul4Fwust3x5NHDjR8kIJ7jdcDg68MpX7Q4BJ4NcPq7ntKWeJ2P11GXV0QS
IWNz2TqdSYh7qjJ5CNgSnV58PWSASL6AG/EM8wniuHDZDRHYIr0tKopL2ycvSNLs
WkVz3dDqj03Rk6RgASPOSpG89014yi8J/SPy6iCzu+cZbrCvJYBrmPqfvMeJ/Xi/
fpYCZPEmPrcTWenJwub0qIjUuw+8FynHBrP9XTef9LcA3rEZkac6EIsOOPD6ccq6
Q8h1+hDHcWhiME1wq1UQG4f6um7wJzdBeUhf5+Bat71piIoWmeYpPfwOUArAyoMr
bZv1MSve3YydLSBia3tkc8RNCKsqzimdvywvCCaMKaJeGwrZtkr6/lt02w6f4hcc
Ai1fhIgvAMYer8g1Kk+jddrb8jOYdffN73mDO1kaQAcOhKLFSZWEzE4LesfpS2Gj
RCSB6EHAJirCB+XMh7aM9T+V3JRKF2amclj3kxfVM1hIuoU8kC1cYpMZr70wSUhZ
OaL6EyxI5j/OdfgQE6pdj5zV5GxaggbF9zHQt+0CdLGX1HVk5aAPjRioui7kk5FY
OVYOGSFnnUDA9kju6IJVL/7jE5MyWuVF2wYTg0kOXnereCq7slWGdi0saF5JdpTz
PNKpmMawolUcQU33Pb0g0DdHIIBr0j/vsZeWU7M+LBu+Cjc6GZIMXSAC1N+4lLv6
HHPy3OfEs/eB7T804cp+Gynp+nh2d0bhNqhokyj5B3WaIcRAVD/nPaW+A+HW7owV
Z2QxQPP4K3hJ1e4WZirzZkR2xd4V/bN3Dupq7lbupkxhqS7+67ga5j8aG/+VNazb
bE9q9XcJUGV6Z3ZOO51suVLb+clqQxoOvCwsFWNU4G55Rad4fmzH1fmJ5gIhfv+k
py2sGjaqsC//HotaAIep1zykRcok/8W7bq9PyWlhNgFsSDju4u5NdHwHnQweBt+4
q2eEnSoKSObfHjYvHcd8i3QYCiOrBO/HRtda00Kj99Eh+VK64DO3u6habGwPr/oC
Ds1YEjTGz0gPpO2OZxJ0B1Ro83/K+sxsQzyIbd63qLh00mjRS9Y84fK59SZH+eDF
30dm9rH2OL4VkU1yarAGlFr1O5soXvFzxT4BIMBR9BA1D0o6IjH041GM1NEJwUZi
A/MgXvtmJqJNMarZQAA6pGtPA+nNAIHx/XQh+heyMQKTvr84R+zHPnRd2yPy9dn/
U8IffmSdFwdFtGIYqNtlKdmXYHAnM2Pjp3GeNaZYqX0FeEJeqh3a5IckoQ9jM4LW
+Q2mgWOeInWK+TO0KKTpw+R8zJeFGDEEVEZ0lvpuVfNBOaYue2ljFkIyKio9uYFs
jf/IPkYoFgY+14Qn7f59zxOPHnaNsv0C1sy6863AdNeAMmMPIPMhnGOCjs1M7Fvs
1oUEpCrqoAvXmsPL8EK8Y3CKNuP/ZVtyOH2LUyBIr0tgGXeXzoSl5/B637STPH2x
TT5uOzkaq0V7qlJfkm/qnRsyxa8JSl/uVX9K1tW1GZ64az8pACqrQFyA8CC0ESpS
cNEV41rP1/hYJbylBdDQd2OcT92PfdhOu0NBjvd2IzHBjF/ZQ76cNV3uhk3ImWRY
+j8hSLLgvTLAL4FzcZilr54NuHghi4aP+rbwExUow8iPjpfMs5BleS2NzZ2HXjir
TYvwAqptp9K9LcMHC2HFTOtn0TwJAVnTAXAoU5ghzhVavEXd+Z2uyLnaFoakiMtd
RceeRJouJzXH4Ofi4SnRiPCTW7CFzO6hRCJRUrJcyt/cMwPQv6NkIevk/CAdXcTz
vrNc0DZdMvZKcfnqyXGWpw==
`pragma protect end_protected
