-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ajBjboq4uNrVx/Xhycb0aUGdEmbSzOS1zM10BK7L0a6GQRE+1rIOBGrfna8byN6mE6gygbYgzXqg
WclrfKaErAErhC+xc/0PddRUoKQtNkmtEjXUySSY3jt9mGPM4GtmS7WQQAtoXwl2Bd8ZUFk4c0ev
JH3dzBGL00AqfZfiPVILLQxo1E/Y31nFFlw5ZGIvqT7K9eDl0ADll5vsZOkUORQXOY8IXOIUhYwo
hTkFcjHXz8Nrtzkhy4+D25XgAsRgKCsnpncKLeXQPMm3tkG6Fia5MypPvDT7bxGig13xXBnOv4Dd
Qvai9EZoLJbZuFj1qE8dRLDJz6Jo3ZKMubGRjA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5744)
`protect data_block
EcFxF3k4U/2Uhm9e762GgaXJ0iCRTsueACnkCNKmhzPY/MblVTNyK70Ut6APgiaeW5TOXPRi7P3m
R90BqZBX4vNqVtiucifrH9b6Xs6wT1jUBQZmbQpbQZPzIjftnKq3KElssSFiZmXgMGma+GTTM/X9
7dHLvvoVIGmPipQcyzOausHAAgbS3lIuVpiMuD33csrk0qxaSIXOTUSFSwBPelN09u2ZLHE9o96V
geSyGIWOf2faKKTL5I/agIZc6VKa5GeNScxTSCGT5zZmn8dJSfwIfMFGqOsNh8AvohyRe249GShy
dcJcJRvVLCHXHKEEoALu0UudPsnSdQ3zeHU9xyVCyndjlnEe3mw2ctDPYYgJ1E8c/W05kTm43FYB
uqYwuQsgNkcmntmUFqglDhBUnxaalF2xmqBpOo0/0sfy2/vX5RDeH6xzEVqxIiGwmlIgZdXuCRr7
x1vTr3PhBvIhaShhq2E41+p3FDzTR2RIYhbyfYB3Tevbr7bF5meveK1VPCxGF8d2//c8cVAz2IMj
2duQgy133+vFXW9Yy4QBhM1M2JVsE9xS+cyAKLkP8c2/fULaBpxoMbSM4zQ3v/3sIAhgKJNBdC5T
J7NRaYyj4ycmtslYpQ7v8p9rOlYKNoD9aLaYrbTvLhoK68eLIScvNVXiNVQ1uavBabx1Y239X5W+
jfcUvGuPrObGigU7dKyktlGo5nf2Bv3AMbCVL5hcwQTwcfY4CicdFY4+TEAvPoFFVB4w1B0pm8Qm
y4z4BDPZEAyHgLwCrmf+o2biOxgx6Yr/MyuznyK166WwKG2bXcfWkp0wxis303PjXce0FCYRSwui
VhVNRJ4xfZfWudSArZxQeSdgGEjiJqKW5dy3WQaobyQwttbCWP5OSgiDdDa/FsEQrNu0n66UW+9K
2pM8N5IKVO7A2+jLYdQMSR97nApByc1pyLD6EXedqWSn5fPddb1qWxjF2LITqP4OwxQy5hFRNKh8
xBt/6aHPIaTAJWVKqLXHD3L2pKY2o2enHRiPjruBXEHfeifcYdxdFs55f5RE3VS4Z4szcatZiFvH
p/R6G9Reb94G/oaCSbwhIBeKdDUh3Mdo2fbehq9/edWBsO0wkmdP/kv3K3vgyN+fABc/H0AUSCsi
L0IJi4M1AvDZGF2yH+EnVECx5zUd1FPdp8K7R0b6v4v9JjMZkvmYRTQPQVJe00Y7MYe+MeTKGlSa
A22I1YNByf8DF0XIdImKvbCVbF6Ht9KbQwVyYSrVvkJq+hUMtnxSpYzLFsBKHbbhuRIv1B9XEqfE
UOZMBWdQ8+cQ+Wpi7k7YHJVOTkLSSXKLrXMYgedml9pTZhGAjk8n5MoOhmRDa4FazstuusUOWn/D
vQwu/4hSyMkULc9zF3WTxNZYTGM11RLIJRCB9F6TUAFKKrKUpHaIBZ8CxkacrGdNJOYj0lX5Zdcc
8hnDQaflpUsR8dkMkIxNCzPH6vhYlUCLufGGqQ76VG8XKAVT6afgepPMLL2y3Mq2joSrNLzsArL6
CMaZiRLtYk5UzuS8HmJ8ZwmPcLroyw6EN9Wu9+l4PivUpp5b1lNkxOeB/Dw3tGWaHGf7vjoCHENq
oF1C1obQ8MuuetWnpUpcPxK9lMsH2RqnQkeoN25JazRI93pYYxWNpBbtY1n7OKVwk9YaXAuoCOit
vR3V10Ur4rIDrv8qdkJCZrO6s3aUS0R7VV1224nL1cdizDPldjAVevNeD7ySAqathxN4Jc59sVOH
c/ZgZDHQeVXFpSYkXFV0C0JsPtcymBmHjj7ntr3ZeHiHquyNvehGLiUSso7N8yoPLUjp0m4DWZpa
ESm/tGM+h/LpBqGrz4VEprvajgquZhur1gkG3dFx1X/j+krDRM8dMuzA9nrRbS2R/aM+uqIieHgo
wsn+2FMiCiRxElvpryE35wxAIlsKjRlg8XnAkRswZXhzGwB31qX1w2w8sj/DGy+5ZDupPsOmC0Dn
VWJP5vJytuwaMw3fRsWL5+iWsgwIAvwU5oRt0bsPzZUQuYGQNpI9IyaE49JblCu4sXzR7P1fRAoT
+85VM1EANeqW6oF2tGaFaON7j1wR176lwrjyYJhY1B67CVkgeWFXa8C+94KCtNEQQrpugFrfFPC8
JM47MRzVCKfV6X1zGNn0KLCKU+kP4Hubrek3aqR9CHfnX0rtHZZrw8dCRGB9YK+M6vYcYecD0/7V
5XgC/1KEMm7k6HyvWffP3+n8qtOiDHgeKgAFenMeX/AOBzacxPLu7+shBfJgNUdkYZMS1lijvWy/
rNKWab+uNpYNftBxl44ONs/2QUCm2X7WR6uVqJyLcCgQCqUyEBys7+7eRlqdFtRrSYfECLfrJ1ug
nXhFFnQaybBzhXu7TIWjytx0ouv6ucxI6fxaGzSRyneotLKx7cN1mnT0b0eDqsqxxCSK295M7+WE
8yAo+ZpXwwX+kqMQrnAiEh3LLzEZoc/LmKElDeger8RYdTg0wSP45up24kADgT41y0YU+50PK6gG
YxiQAFAbzKu8qNZLMRpd8KK8SJczGAzFyW3psKm6eaanrx+95xvZa77piDTmDsIQVizifmnt9rP5
tPVye1FNPve+XRNbUerZgCJizJXpDYZnTSCHqH9f8KNh9e+BLQrL5/F/I4Q+AqM9KVYYkgM8S6ce
7ETDOSDVzsgV7b+glxUyd7QNziiXRtv3KbAcGKC+h85tohW21r9A28htLJ1an9cvrFSLr2d+hJ4e
RH7QPGvUSMEyU5kHvnjegMTgmuGHOHlJUKDnS7aN/zjkjb0SCEJ0PfY3CasyNyIZdCPs8u/Cm3Dy
HOk/Xlj+lhRNyg73/MUHTmGJ3ShxT40IYVk7oGB9OVugl3fCM9zhWYdL+nxezX1xAU+7uHK9shzK
MmVV8npQGzcMOkNNwfgS8T3xL/eWkad95cc9rOtDAZG78lGvlRL5rMldAiZymOv/f8VgFSdKx/7b
+WQLzIYf0PL/1ypwbeW9o8fKkzy79gxHl5wUX8pI5K/KQ+dl70wqpylnzp3H+z71zwqXeKgNw9/g
mNVfTjOrjBE0/utCGmCxdY6NPsZRcRq65Qtzf8mrj94JBiBFy2w+j7b3X74BtDBtaecN2L1rkXVO
ZvpG3xXnYwaEktdVRcC4WDx39aZIurIXYvBgO01gZFO6qquTXewU7f/OPY393RSOauzAIKtQ8I4U
IJBzrwnN3yumeq4m/GzmTAbYLvp9S/+0IFevuAyMLfRO1JXKh2c7o0W83Xv+jZKI318MuLIe16HV
S45slGhSuD85ZFOlTlH61b2av0HLOvBoNirl7bsB5QwiObj/hDDAwLd544N9YZrpe3FVbbzEOryC
0pfyWl4iX+y+inNEAVnvKhYiqcISlGSyxU9pRPl2CxWpDcbhwDjPI7IFz2GmKoWY4WHY8oLHJ94t
Mgp4+Lfpb39Mpx+sKC1dFUTUmmMPNdmQ30gDDG0/bJkoS1PJYIZ/MaQwKA+uM4ANjhj7CWnyVII5
3PWxhw/77EEJTig9r8b9s/VQbatpEv/Vap8WReljfLSt1WC2l5k1TVWZ3jGN3HkTKarRvh/qASmq
arPILP6hTGF1eHpMaZJDAxgIe/cv3a2HGMFQQm3ggau1EfGsNjVdJJlcZ6ty+Xk0PobACg3L+eeg
Gl4eIPLuGRQbtC2zgKdwytzRYHzygj1e1QVBo70eIvuRWKSITzzrbhUT17o5Z1VVsGLRlAE2wW8m
yZNA1BTY7F0r4UKhWvrI10q7g4lVfIDWW/1A2fjvDIIz/F30LaPTeasoGd9ZoBBUKspww/fu4b93
YBCJvVieApKHFA9gjlRGO+purKdTP9snO2jUYvhMsBT7fntVPEdzgmHt7/yAGwquzlTJT3lmeeL7
7GaDW4GcESrJ3+lhjvZcNzTPGofrXtk2PZqYs/ri5vPVk0CMphoKyAS6EKduWj7zTN9hMEr3siJ4
4QiqrlHNyF5Xk85bVPiHITKl8yeiewj+sbFgpsu2sD86W66hOcqUnTXthXx8lick9MlUbqqfYu6R
e6oYtZI5IqasbT6c3JwRp8tgNZpdxh8Oi1gTKBif0mdQDwEa3XKGGRYh4HwxmlgI/11CMf7rWAfp
Os1N49IMwQhDH3MAuYDP8DZXj/DQvLAFKY9LPi94EdvVAa1FIHJ/cUPPcrO1jhXUTm55onaSf6EI
247btBnl8zo44Li6/+sW3AXiHpiaYmdXQOfSJUV12nxKXhvIX5MAcyvNSEAW3KrV1yCHCykBc1pA
HbvIpdnoUFX/0ZoeFO7PwnmgvpEV94iZmKfGJ4XzoSQIEIGxAK7lArI6LoWm/9YB1GQwbJZTYl53
HpnwungHHZCbc7fnRG9wC9tgdmVwaweCJTgG+mEcb9P/QpRUfRU51BitJyUgipQaqke7nlzCWEQG
jcvDBHFJyw/rZJ/fayTKqqfjgsC3/OMZkM5FUn4sTWTyvE5TDvmQ7JnfuRcnGZZTiBIB8C2/Go20
A9t5X1P8lJIgzBWsx1iDLjOvwfYq64YXUS6QHhL5oaUdqhMtMpJUyrkxs8/szNXNtOh0icYYjzjD
WruhkuWPNbRulmLIvzFXhe6OI+LRKVGyvGLV3I6aXtoMc+MeYkROF/8JB837Gox/IJX9VR7jkxc7
/QuUQbTQtuOXQQdu4fTLopJyJHfS+CPtz3nZrgIT9jH9KDS45s3+8kXU/XXBUIlwdK2qQ1LODL8/
38XJxYDG87fPaBP67xr2RDW6UJgnNaymUS1ErAwNbbCDLw4liJDf5w6zor+tnSqrYmTGmG6AmBGA
U5SDfuLh/2cEDT22jAPVJn6JoP9pkdeQRQcJYONpor8Ka1M1fivkQifduR6jYM4VM/szTi0/GoC+
YEhOsxiAO86ifmr+I7/Mgu/WW/os8Sjn+Dx8ROZWTHHTkiTyzy5CJ0TLpnfEDxfDFVNdDasjTvtZ
WPUCPesr9UsJvINEh/Q00kpXo6cUeXl1WQiy2n1I5RtuEni1s4/H2m2+Kuh4nS4QMF5uPaUiaopN
kxdmtWsS4NpjH/+pqO5KFSqt3RonBtnaR6nrM32L/35V9mD8D+IgOwBc/BziVA6+TTDBQ78YRM8S
Bwr/0X1dxWMMHhPOvL078h4NUM2YFOHjCfWDd0prCCCZ6GJM+jkAg8mHajruQt3BZLEhkcfZWAow
+DJxETAW5Hg1rIY72guYBlcz7Z9S1W+SsZc+KZyFh24GeWqJsmTKSutYYXndPh4JjfyA/BTM8Yek
JiF/jIMJiQa5gt0wDceTgcaz1P3POxIBc9Vup/TuQuXvtZ5t6yJ06a8BENXTiG/CEKNPyiD7L0Ge
E3j/tAAQMqrno/CoaeIivAwHIl06U4YkfxkQLhvdlgGgyt/TXRPNKKf57ZfkLVjXtLhfKd0jcupV
e6gneCxUCwxoiaTp55iENs8EInaP3CtRIilU6PN3+jOYj+J2edHXxKndrGqUGc1o+UaGhYneaOWz
pvF1pgg3J/36RvFqLnbBXk1GmeSxY+Zhg0JQif+HkJKF8VPyIbSh/toi8ubqmQCdwS0oWQTyWfLX
zdx1EV/ir0Cpog3wMsfHwk1SWTbHUVg13cuhoPnPBYKDjCwEvgfd28wYEy81a2cLJeJRwI3149+1
UIn9HD/n6KdwD1l3BmCHs00YTtrs5DPe00Ib8dScgZ2iSKURnVemPViY18UvcTNpSrY8b8OVc3in
CKeDcWDvt/S/seWLcry6q9GVTlzcuSOqdcCM2FA3OaSZU1HdKxyjoqxDruTyN6Ju+tPnVBWThrwq
cQ1T/R5SOW+bBaXTaFJENMMOSd1oTjanSazkbwmHOEyIZdXHtoE7pU0gbk6vfs/ruTWah/daeonM
ClAkrShm3Kva+q899GZXfYPtZv/d7/WdTGbtS8kH52BslSZNF6C/V1Ef53GwxjmCjRq7mULNneu/
cja2J96Rcdf0+s+o/hxllu1I7jAqVLbtrtk1Xm99UTSMoUwaz2X4r0Ed0SLYSJMHV8n04ZUHNKXG
By/Fd0Iu275gmLi/MTYt1Jd4TTvYm6mdeDFXdDP9jef3GBintFqOGJDf8UoaPJXsCbLjYnu+B23v
/W6oxRseNt1YU7NQQx5Bf1R/dD9avD3WzLlHwit3h6EzeCwLQDrkVmYmz3Tyyku8ME+XuYs3FR/8
pe6R5z4irL1TwGgHib1/WuNonA8mR7P48rV31bfR+PHr+uaXrM6HKxkBwepvTpIK0Ac6PbPlOtmZ
qyLsLO89lF8+AVNuV2Ancn2spq/fqKvBL/b4qQ8kGfwtqn+kyOnkgfYc7xs+pmfvvU3WzMu7cByV
7UUrgFkyZoaA3hFSI0MlJo5SOWdsu0MB0KOslweSD+ClVfMk4FxEqcXivm/OyY1yKBHPx/IOf++1
KGmnXGq0Dg61BJsNmjDQ1nRl8Ts0urzD6O3cX/sOAp5meSMKTOasBxFzRsn2zaUr7UPaw/9Gb9yb
etsGPHa3mLB7bMIVIHTcz4aPi4ZiseWCTQmPOZSk8+UHXUqZS90NtS05TwlBsAGusAocX6DJrisU
UKeGQ18ZJ4GMluqDmZ0J9iHIXsCi7PH5pfvWYUX+C37Vnbh3mkX3o/5Efub2vCeSmeioIMsSf77t
q3L05Sg1+DEsTid72AhAVkwyZaynkvfAYvLtF5gPNq/vaKdUBWV0aKLA9avTbIxnqH+YhzV7Zveo
zPTcvptOWLwff78jYhk3tk3iig/UvM46MkrUMEri4CELjSdZhyA7bDhEhaRKPZBhzMhAnGYQDc6z
PircGH6rZqiDW8KURpXIaOXR3t0GVZYMEV5rx5mKTMy62AUwrMpvIjm7tAIalpQw9IoejlxIc4X2
h8sKYJtn1HIpUIz3XOCHmz9HZ2zJnB9YuHZQA5YDAUlriN36NunltksVT2tIuvS2JKQkA+7JGXty
A/m4ShfEGutHRIppjWKzt09PEGcHnAj9O6pxm6zF9KIMmM8ejy2M1IlHGH4l/V+jArxbyNn1r0HB
1TMbgGYKY1B3JBSfUPtn3Q9BiGiNxZELWODMFHiUp9oycsxKdJqDog+KSaL/Lwr+996RoE3DdHG/
z3g+VcSEKfQxvSQhrRkRMmx5j8jyHhzAQbSXqK/vbzE/EUPc4kc6XqcrygdWsbL6aHDvx2yd2gZS
Jv/qWtP2FDcpBY5Ztyo/VH6OkqEknX0J25Q6AswqWKOnU0jH/SK4q3e1B5bRNUIEOTFidmHICraj
E2v55IGc0otbU7as9o5KdQkotsBkNWOm+8WBGIJRQbJpjq/WJqGJJiQHl/PW6c//kuFRsUh6XFQf
uvyvwZDIsVrhS+0yvdkaDSt+X1z1NWGXlWSZmS+9SvwcpwYhb2/ikv2353m1LV7DtFSeKUk5hjpF
1TQbx972ePiIKrX35hCdfgyon7QyyTZ0reILJLfUMyMZ0mfWKu7/8DiKR8EFnSCyQ+fFJARzo34y
ORreiN4/4VCNcnn/7719hpErKGpYDBPvmYIYZnm2lncbVyCp5hAhLNfle3r1FmZ+zvw17D4/AeZu
NROwjddkyhLB1QVviUuk+GVl3F2cDFx1uGJQXkxeGTBX7QwzRI+DDy6cFNUL+Dp7uEwPuO0ERdnR
3hkhBtSnhnsIFMIYYhF35RGg1Lk1A9bGc1OF4jORjzxdpfpjqMMYzcK7VwU=
`protect end_protected
