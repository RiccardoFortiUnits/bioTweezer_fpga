`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QQb/gBYQ3YQkSgsexF5i103CMr/suyOhtjGEnhfk6NnGHoFPDMbquIiGBEyz5PTa
0AsdyYkph81wl5oJRyoGmUQVP8jEg9HCAye+mzkFU1SMSPID11+4gcDGrsV2wFdZ
q2gO9yINI5tCNo8GsK3kXRKcljinEEsh4s5jMsr/01c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14080)
kX97QlEX23tGr+fvOxRbJq+I6gjTWYOT3GHDK+nU5ihNR7iaXgQe4jFvx+KLmdkQ
ShZrfnefkOUJd3CINJA4UypyhIxBmXBZ/DXxY4uELM1gk8yVpXTRMe1w4CvTCgx1
7ecMsCjkPPk3Qv+0EBxfeh3PzoRZ41M/wo3KNSwKS6VxJxWGzX8zS2rjLVFCEA0R
ipiYFjD1OVK9wdQhwkf824+gIkkCDINeucr29hMPagMf/mmmNvZA7LLIjB3n/iM4
xNGyH3Y8/YQKhddeA7V4Zxa2glp4KEIsvXBhxxy0yJkdph45rpoIIfK3meNh55Jl
XvRsrReM/VEB32nCc/2E/B4rF3M3AjY32MgTaty+RysQzIArfyK3xqN6qw8dd3Rs
wkG+JDeTw6Gn2PqGN3sYXKIuvrh0YAa2d+w6ymcHUchMZ14Hz9nE11HIy2dllgzL
ZM7qlqR5TtOYw/guSMRby5MCKM/JRnubiow7+UBgjO+DbYeZmdBwMmqwG0M0WXkQ
wBzBnuyz0yeNuRjwyKCa7+G83ftSE/oqddf5bm350DNum5GPv0xrBlPUdVq3DdDp
BHyuaWoeNOE8mLhl9u1et49Do5XEBgpmNul+N2ypv8U0T0CUd2NL6JmwO+Akr6M0
Hsjvkv0JzTLBM6gQH5ppzXrj/9QgSNX8KLpjwctIYdaC2I8V+Jvnzucn9vs2P0i0
0KrLNbvrqWPeTH8ox7Wbd8opFSCdrPH8BWJcNEOXIANCQkyc+3Jd3ZXcGTsTWz9v
NdmwexGkgZlqkbRdAW6ezlRK0qbdImvbaCk4iLEn81ugWdMdrbR+Ulyz4FNU/rJ/
VfZbIkFucXknXc/K26cRqeAlmkmigocz9Pe59SHHs8WTZF6AzHAQnR/64vajhxkr
Ey1USxW4Lgu5vBBzK2I4wMj74tBvNnK7AEnzUAG+6J83iiSJ2nO0sGHw0P1RKiST
XnrZWWd86RxjJA74sVV1F2sKUJpzUBSZ7WyiMri5l4wJXseI891znk/jHh4JaDxC
ESURqZnlA5W5cZTyqU4LVQy+Re+1fCeSKs9igZGMU4RzLqyCUk145+jhjlC1lWLh
RCn0qpyDKo6yN3pIAmvhFYFSwoGPHDeFkwqPjZA2+8JAU540doBu/Hh5/+TY2P51
Gmc4fJBYCeTqzQUbOGobqe7sQoxy8C4KTNy4JIRiSEbTG9Oex93ZLHCvuLqFFVqD
bOLDm0wpli/s4PT1X4qP+z9aC65/YAW2wSRqTahWn58e7jMwZXY1cK1MhOjyFxFO
J8uSGqcz7JeEqH5RFMu56FKRsfXUu7HiKqPHBkSzNVitNaP092383Up1DgflAbKW
/XMBFvYZkMZkRHV7c8qF3h548PH5tDFyW6BUnY1qh68lIB+qXvArdHUS/UIv1rn9
Jhf0B929k+99pvVLcHVcICrpICMOOJrrbaPihEm1lXa2YelV5EiAbxPU3G/tHXfB
5Fk1C6FLZP2Opy46SIjrDPvphJfdYK8vZY2JfwM+TAjAsrnAHKG9CEDsjkK1my0H
69xl3Hk7BMez67GaEqkgv7e2qJ76WsiDDDea5ofCt7Di7dOxYtg9Eyhq8+vLAKa7
5Ln7vXBorkbPmTLdJb791nGUvUE3rsg0xxkGntRKuMAfBzbnK9UdzvT3I+O7r8K0
wMfnrKvPKexMf8KgpM7qDQVj/XP1ijQ9eKWSp6GhBGeZkxNHT7T+Q7QRRToOCm8s
1TkWz5DeexiQg5JHV3MIEJQCumhJ24FL3vO1Xhm9k61rKMTdzyyhZwKzkksgR5Rk
eoxranlrsMfYtTiAsY/sNcGqpFhGWP+TgTBW1N5ZWi966SXiV/1xmeoKwoWMoqOb
+UWS7yRRBwEJwEOKuImFzN/fwlqkJJtsHTklKqgnJyW+Pne+JZIckailW/x11q9l
vhvNZeNQPNpxBakjyHqPFWQKy/ETB1Equm/hPLB6zwo0AYoxIrkvA5bkkDlgEWwR
B9xFjvBlVFThsFAtSIe/zaA3KvFhPyVZld8ohtbHMWdB+Tbmi3DCBOKIPfTXS/8C
MOIurpzZ7/+Ohid5WtrBXXbnqcBbp68GWBRNCW+UmbluZ7SJ/QMxF9D0NZn1JZDU
ONDldkVi8h1xNhH55nmUeQItoyfEjqEJOPbEIZFit8b63eRQAndX8qZBiyiDddL7
wlMRx6bdAhizNy5PQxKyBOtDFzc1/ShtAOjVCoXFuy0M1PXrMETZbmeiUWUQ0K1P
SHw8+5c8YjkkzR2ZO2oNmDzbXrrB5geHvjxAc1agc4NvasMH1BBaFIToCw8bC3/z
Gema1Ot4pCx7OVjaRub/xrkBZWTgWVF2VTh1WMp4CUoJR24jOJBZE2yoMaTE/qKg
P1Eq92UbfZY86iF02k8o78jiIbWWzFZk5MILE8wdv4pU8X8euh9KvwTnDsJ2qSco
/Ni/glyK4eZFsX3V7CS/vuPE7Kn4fla7lGzGEdb5MgOUzLFC1+1ozmZFNSTmdix3
FxfxiboMTWJa2w5pWSUtL+BlWSGAbsTGtfOnNhLATTF8I93JzE02NRJQcltIyYdz
btcQe5UpB7JZUimSYs7iLzgpU1lAZG3r4hJTqYxVtWJwBIqazq2flPFwnwXyoF71
waDph56PnJo1nwqWzf72ZmaWAUbrOp1d1s4kw2F6W2uraDFzX80LQZgiMlDYDLx3
hexat5AIciQOOki1eVDOIoWpL2740J5zAPhKNEgs2Jm2NmLQNsUMV99cN1KIx2s3
kyrab4ap1aitJS/WZrQ2MH9rNOvspCBfXsNotVX491KzMRFHckCgYvrNAbhB5X78
OWz+bB2JZ+wbHvQcZ04n25Fvr/eJI3W+pV7njBLHYurs10DdW3Nm4DM8BjlcDtf7
dQiE0vuA3WLFiYOiSk6A4FCJsgEhXKoDNcHUsUgQrl7B4ILdKz15pHwJLYjkNw0q
Q9jzef5wd8oubFNC0F0/jCU5kvLP7LlV0W1uFZBxDyLza0f9SAUB6DG4/F05S7iT
34Dvpk6jDOSC27F5vp9hI1ZGTYeuKM8M10j6KDfXOXlQD4qrOwU/v7gvT5PhE3eb
Whv0rorTdCIwW7t6cuseLHGIPUHJ9nhNEjduqe2y2cSzm0c8qMUvsd+yfdvJ4TP/
PMIGD4sTKR4vAcUGDuKULgnMHnWfY2Nxw7CFBcCT1Yfim/Ca4Im9J4yhBVJjm1e/
+Pg0pnx7qSYsvIm2595jUvkmTtyjuSbjmdXGiETGN6qaTrnLWjI/SHtoGfg0MHBY
Oc9BKMnkO6Fk7+T2f+wwi0tVLuL397y9DAyeBj3vyU1c+aNzZnqtiHQ2Hijyj+pS
vUaoxNcFXqTF6ZvIvtA0OsErPBRtQTMa4eovgV6KLLK18yoL5o/Fytx2hydRQwSP
OP4jMKChBFgwwEVjgSD7YIpOM8IGNQhIzvyTSW5c7rHNCOxa/0cUaQRrNoavAwWC
K9bgntEs5MJ8733cSaoYmtfddl6G2EnRZUphwUSOjuaZ+mjR2mkXKIPOqyW38x+c
YQxwRVUpM+2LIddvfmdamPnw4WyssbWIdV+Y9vGEIAI89IHbzSwVGrJuAZX6NSp5
Kh9R3asLBLd/eCuZ4hr8K/HJc6rvBO9TQ4wE+v3Qh+sG9gLsP5hgBBnRYyL2SvHH
/J5nJs3IgmK4sJI+in0h6M4sRjUjx67+NIF3XfeUVP8HjzSUoXxldVHbjU0tW4OH
OiSSaRBON1bXKckajbzxUBvW8/uZL1TsHEuLemPxfckEsptleN62N7VguWhjVgi0
7k287/t2g/1Gf0FlfUMHVouQOVgi8fVSLCFgeJie9mrKDec1gPWRCva3cg7gdMDL
7Vy0CpPdtJTAkbPOBpwAIyBMMq7/BOl0zMaVS5n15U+XmekrWRBQMdYsTsm/je2L
B+x6cXCkNbY1WpU4f4WN1C9kX+gSPdCtEOvkEciroMGIa2zbKhMLbTWXfwzD026+
chwDVQfXWj4ixBAiPDYHKvV6BzM78KcNbVAWGSG+P1Ezt1hTkxbvCXDZO5zYmytE
Ues7es38s6CeqWwF0yn597LhNJ+nq3ZeilmTDXnLw/rtyPGS1pFpqgBG1M32U5XA
tjrBqd44j9/FiBbci78kjvfra1lZ9Ejvvo2nfYo9ktFfWMAv7Kra11eDUkslD+Z/
ONzIxzhngrqgKD1XOUdKB01H4MIYlZF86EKWOUAHEZGhYE8OjbcPI7SeF44dLb9D
Dh4lYd9XEsWhsXbQBevB5CrJip70zx94ZK8pMRVPdX/ThuMY16f5R+JSkM3kVlt4
XJyOiVJ+YDuEBoHimx2tswsXjYPUfYHrzixJoN8jmJApTS4wDweEwzMUV++rDMvE
65Ru2UknhYUnScFgDSwZssqcudVYIAGQWHzijRlpnleztgtHWILMs8W071zI/OqV
0mL5obpZgwA1WQeWNqmeIwu0+VVIUqvRVEqgQhbaKUtaPTzr0S5Kbba58SPfDze6
mfT5lv59ecKEJ44nw4LbRkSaH/Jy+wdtlrpVXjcvBLldoUUTnaUrq6+qLTcrtuzp
MhVkpDUaTwjAMccrlYbqsBy1ESoA/jnpCaxiSaNtxxBzuv2JLAxYzlFo2Zd8WoAB
ogRciDzx0/PKOWcP1tvyiB2UgVReNacE4krk1hWtp8WXVMEKd6+LAUnL1x/3EUIX
dfFaa/D/k8OtsxLYMStlcP/Wi9rlm/2R7Ea8NrachO9bbZc3GuaUDScgZHhtUuOD
p097ZHCg9QniKWnGiKhtPAIgN6pC2Wlv6ga1jqWHrtU8tFj4evRDnrnQsqveoBhY
Q5G8sfQt0FvWlu1kjWfuTbUyDR19m8et2qDe33LBTBEboFo3TOYQqPa9wDMChCcv
eF/wTcXejJd4e/D3pmQpLaG3N6nw84PggTx4Nhbn65ZehZFES1MxdSfAf1qagO5l
oSc850xn+0Hy9gc3IE7vvMyj5EfPkF08NCXPV7rZEcmBOQeXFXbookN3Fdgnp2Ug
+B1LfQLFqWPaZoVkJ2akGx0V/2FuviOriLpx11FFi1J0jqKPd7dsFF+rorUE9pGY
sxwqIJFTiEqVD/I4JKFQEi2I+rdEdj/5RAsQ47AR+/siu6xEjwtya8QEwDvPZlUt
NAS7sHAovL87MDCdJyvvOM1hXEhvXx3MS2FTm0gwboZXviaUm4JRTYPdyrG95Gmm
2xH5pZhEwwPu60txSby46O9TS1FJDTIl0TjutYe2p1HZbG5I9l8YsamAj3fZ8nUP
Wppo8AgjcmcMgnEhCYwBI36bIN11kv2typjm2t2OIijvmsXqJfw8PDGPmfzpE1bg
U83/OMMidnGDieEHy/O0Lj1cQ0e6n8NzUNml/0uu0YqVZ0DmKI8wk+vdWGIK79co
37KL1v6HnUnUYrEPsPGHm1Ao3ICu2a3kyHcMhJQq90wgQ92yoZdPS8hLqZUWvKQa
Zwmr1rbLTsnyIp/wrQBcRd893hgiLOhHzlzEOJSthZvezYuRdoX6RB2SR89nsK5A
KRP0bzuBR9U4nB3FLhKi6EQ4+pbfhdJkahLlwkx25Zhlta7g+aJNC3AT9/2g5hWe
UmtiClPLrr5QhvDowyaPwdKEwiI/v4NvZkj+S/gTtypwuU76g1A9dfw5pCMC7Z5a
YBtJTSFwxBivfTWOioT6unnXPLomXVcvfc9rNyCzvsAFycunnIGBC//iC9U0Qt2A
kL/I74CZOOuM2owDUS+MMc4nKGddEN3z018XVTcyIIuhr0l+NHp6p97O5MV8kaNN
9X2abpdfItVy/ZwHnQ6j5PqFSOiKw7X9Vp/JHXREfq0MddD5+wayKYmrIKi27hHL
GGuWqWgXh+XmVBCtaFh/UGY7i/f07NsbFxAUeim9zTdHSzeYQbDFgvXyrLbC6gyh
a30iwXEFH+m7T5QDHAx8VuDylYG5wely7XB17giR9ZRiyFEsUJmt7tLSzQ561QLJ
D1utsw3OZGSCAX0H2wYMBlWUQpeMUvl3U9VA8d1ieQzxyjk/z5kFZ2sz7CPeeHS+
YHFzCZwTrdSRBKoWykRq5PT4Om2MFXZUve73xuNtQfc+cM4W5IrAgf488sm9/A0W
wuqI2uLzACJ7dEfb0Ylwd0SaANR9i6+iP2lq9x0rlzO3VFjIjVIVm6SEfyI+a5/a
YRfjfAyc50xNHv4Qi+yNv+WIjqKhSR3nd5lXUtDUNcyFodR5WR8OtF0hyxkmvdzr
WJOqo0KSLzLf3Cov1inR3+26U02y8Qv/tJX4+FevZrXNAFWCEccJlb3Twek5HIMS
Jv6MCi/V3NtMPbCduUzdjjJcWjFDKmChkWghWOt5Plbo4vPDs+vkSSIzdi7ovykT
9ufNy3YWcoQDqnIJM/cO2Bk/3ctkVME0iGzR/AuCEmKO4xXvFygI6wYu7JrXsRjK
iCzGjOo5Bg7x1n9VqWAKGDKkvtaBqz52WWNz8oax8q5nIqtX5PSYx0mqogGbKJ/W
kl+Ei9pCS0Iif31XJPEz2Pfb8NLsvMUt9/H8ACcqCaEyFKMDwdEF0XlzuagfVVZx
qyT5wCMwv2QZti2loTVnTX73s8jeKhZLDQ8VYPTF1b01FDUXaoISGAFCos0/5wwp
FG5ZSYQA1a13R15uIRGinfZ0UOxvN7Y49nMA2fQUn15fdQIGRrqdlVHZOyPW5Okk
F9XWbbr0vncTnZOTWadYCg41cOLpScUqUbSXYO5qWxzFexBljZZpqvtXupwP1zqE
CBsCsmoL0m3mYKBYGJ99dB32cKTVIYm1tFuKv7k8Pdt/n/HUaLC74ESkjPCTSFxh
H/Z+zVaD55kHdzt3pjGaT/pOKbQ86cXfc6FDDRAxt4wWg1AnsVUyTCGwuF5hmNXB
AylxYeqCcQGG5Aovh+KpvHOEiq/hoSFFefH1w52h9/9reVfEeRT/NWgQeaAxVn2B
Wazt8t9t80kZTIArjVR4CccmPx3HmK3j/yzPNinOR2j5u81766g/k69RVROn56pk
gIIQcEhAY2fcdCYNb2DqvqvbTdjpnc9Xyn3FpuX8FjrVwP61B2+QPEcmkzMGsTtS
IH/SVZCTqEfU3BPdv7LM7kVhwsaUOMx0ziZ18CRjnRWhq/nwItA+laPyEf31bkQt
v0uo/XCRxMC7SmD4sLUIJv5eMFCH1g+PU2JxdAPQ1LYv65/lgkCU5CGt9uEaxasr
1SoOPdBGc7xQrHvnayNjV7K7sHgp9U0VWZsKDvoF5KKn85JGevdtDRlyzj/XwELf
NkUr0YGNmkotphcE8mSsjBwOxMZ24nM8y7BXuXIFvUBuNvEwZi9v2EJ4aS6TzitN
tjzo6QAZYZuY61zh+h2iLsyMEbinJ3NLXe+G+vdcHJjUxSoUXOU6FRMr7gOh1eUE
/y7dplEDzu5+SZUpHsYw2Vz9ohBLWpmj5smU0ljludf1DVOfCLB2yCqgp/rmeMdh
82OT1v5rSnpkwrN4bd7ZAl6YUt4Rrb9y+neXg62zLJmZQwuKkTvmXDKatS9a5Y8l
71oLRKDl2H2ioTfmc/RarWGSB98g0TjE254ROo8f+Yy3wonUnDgMgdw8rOsypmuL
Y33uXhajXsgzjWsmCH3ppaLprR45JMckm/c5CwcZRHhRLieySjCywhtNnYq1TZRl
4Du2mLxduxH7/26CWawZEyQfXw3Gh3nPK5hfDjhTI67j1884DvToFMYkvmpB1d5d
9LymLXk0PAR7aZmRTBpUlz57LpyMfPq5tjdA4qMJg/2+SkmrcCeAnyQOTEYj831z
T+1CHlUJQCHTqlka3nsASV9F6F91CbBdFqYMlPor91UlB50xlV4zoqGlK5LbXd+A
1F8luh/s1K7kai0aV73Sb+4+HwdpPgchmakb6Z2qVlXldoAhItzhBQB9mOlNBrdv
nz47NInEQR3E75bdwikhz+mBGqAldSNVTJgtKG+91XNFJdaOccR6JmK7lccCow8s
sUfmrYT2RgE5oy/BFR6vFlYAFViVgYuzPMPy/IIYad+ICOudCNmuFwUZwkhCuJ73
RHqAWN16r/VSItwWKsD81AJzsY5sCNPWK+sWbEXUBo6lLwDa1R9HD0RwqmSjs998
ISc1ob8H0UOEl4eGdsME1NQh2PywWjLOB3LNaXHWvWxh63yYmYBHnPYTtj4nBBtU
/R6jtc0PbLH6TqBuDGJOcZexWsbU5D3/FI43WHeYykkoKrqhDEuR7Pgj8T7QzblU
GaKxZ/t2+kahRreXzyVk3uOQXD+cQbHdkFeDRWHkOsPjdE1q5Fu7dAuB8w3ItxkE
P2zP4mIxf2IZlfuKHXuyCv01pDAFg6YVb8INjbmh+4ZhE7ZISqsx0SiXLfHhwCY0
SAB+qQ6Mp2GADF9S3Miaf555I0Vf7GbO3cB0gIfkk0qumRt3LRNHaR2akBaMT8hK
bCTTKTzZX+dtEy8DWYgBNsP9y6zbaIH91xTxBAGSGFqh4sWAd43ccmkFsJ/EvSms
lCjpu51eKN1EIfBH4yqx2U1yFUYBnODA1UMtGHy57IWwyintimh2+TD6IP+m7m8m
J8ZEG+wREquzyZmmBs4+bqGOQzbIIERofbdynj1pyqnGUnTrQCTinYgIZ5ZWIUpy
7dwtDR8ENYcV6Kb8n91LrO2jK8mCgQF/TCu4sWT5suYKSExbtXOWucBs+ntfITmx
a2no+GPYsWN7pdQdwrikFFK7UnGdDfW+RlGKOmDUrgMT9ku01xl/Cn1SJOp5hOin
xlE0zpmiB0xo3w2g8H4uNs/yHXNMlLiNpZvuBh4QFOX5j5/gzSIx6lRinnvdww9d
xc4Cki9R/Gzt0SMic6kZDw1ZA0XvUV14AViolYcJ6KEIBQwQmtcuO3SjZGwbDwRY
kp5YYCqGqLuKmKokL90ykIZbPRDOG9ClNOy4SSNNutWSlXpCFbllCQ27g/d3EkRh
KnWHO68kl5AzEitVvZciEguwp7i5akNfIpx1KzQ/sFTbiMhTBgxRo2s9bZz3bozh
YPJ0vTs4HxMUMaG9U8L1SwKyDlB/hu997SgbBiTj/G1HoFDc54X98ZbgYjG/EP+R
jhY2OuGLBXEpdhOQpcXIYXEsq7pEyqBlbqM08DDzgMXbNUwCjH5r03Pirpm+B6PK
dGPkg1JNP90yCUKmQVUC9KmQlcG/H65OMEy+2JpXirmy8yE7mPxLt+T5eMbOzCPT
PYZOtJb/PC+Sla96Pwx892dvH3+GbRIMVg9xWBLwsRU9GIVg0oOaZqPAu7mJiUY3
txOgObfvwy73gZvV/FM2BIy8modL3jvJHmpKSJJMdTBHlQ2VRB4YVZ6EgoiQ+vPI
ebFLSNI06iljDYWdQFJzBBzyuLuMAw54tzSY/t6Ay81zzyuFjqKVHiLefqRPY1xT
aLWx6gpmBjgtSk87tO9Sj8Z9V7hWMj7fViqx9/caXYIncy+xsmQN2a9RewIjxbMj
fMrRgz2c7MEmJHb/rkWlaQEg4VnciS7+6O/74xjKzfi3DZv1KYB2iwq/4p30HRrd
55mOkiWltjocQfC2pIruohdQsXGpP1Z28QrRh3H8GGzuNQw1esMC7ahtL7zrHzOx
c3LvSBWKJ7iO1ldgxAaTFU0nUkeE569LzBIA9rHndw9BTmFTidvwX/olz2XF7kew
M+rvCviL7Fk4KTIguPmBt+8VRJkzF2JeSGq8LknDQ3qai2dGlfWkCPNYkYBCw5e2
Tvo1wJ5r+3RSUhIeTCG6ykJch3nNA1u9xB62aLnuusfoPvDIp5CMNOeRCVg/vJ3C
mQ3TUhm2eCH1Nuq9fK2UnfWGbLr0FhsiLqQ7/fnRUDb2zTRsXIvCqK4IfQXD+K8g
4zTKb23crMpLpB16QgiYbF+VTbDESXOEcV+8xgGEW0AJpqe7vVB45/E/KxPJ9McV
0RxgxoUcG3sNwR9y0wnaWJf3GyD13acMqyfxBdJRi3pX3NDwn09P/TXg27PI6eoc
MWZcvoB2i0hO7z+jDaoywAsft41UogqYwaiwEiRadYSEeBJAVfxMH7YIlk6pGPmi
4vAevBafp/JACwJ5xohEsBTeK050OF1HFpacsJUMBrGv5LqIrwRZ3K99hfTbKsZC
trHtPIbxabnGn7m/paLP89O6XrXq7VmHL+BRCyvcWpfX16KyCzAF8OASmv+qMXjz
6Wf9QGmo7BX1WHwxVmfyG8jYHsl9DeyS+Y9oYA01IG1yc97bDhk85tMeAHQJYu0s
E+Ku9j/DZw4+hDUlV9TKFpXA9yT3Afz0e/vqiY1se/6EGC2PSzYBpmF7+B4HJLME
dpnwEMbimm3rPj00H/qD1nHn6g06Uo1m1N8De3WipC/uTLLGsmQewKAzqky7coxj
7gC3p40gK2ZDVsns/fMpz8+bOG6Ph/0oChLvoRWlx7ilN3nAsZ7AlDyXZ0hbn/Dz
PCW3u87AlT5K8fd2Uz+j7xMo/Jm/TOgwKuwe+45SMi3qYxxoFaKs1XBFuOh5FQ58
UD6StRPhUznrMxFYO0LnpJap/58rpYFphDa3oUV7KjaUHWbrTNzzVLVwn+JzWdAW
6Uww5fmWkgayRXaY9hCBkWpKy3VlCacZwFAnfrdgkvXA1/3Kwg0So1UK0lkxf1VP
1WxgA1Vp/PmNh7iSDov5GelF+Jxq0rf9mK9svfVBRn9dY7M/ICqHz1ZQltLnwCjw
af+qQy/D1ux4A958jAG2H2iywZJ3yYNhR7rpBQcGpVpzVOPox+V5em+QWxed9n5S
MS0V1b0drcUOgPkbtzc4evJgn25mZytlMeHwQWBsSPG3GcVPLss5sJU8hAvvvjWv
RrxeZKXMXzZOHTCA2hM5h2MeNw4OEOwIJEydNE5NAJpyFP6TNa77uqenFeNxXSTF
oNi74k6Stikhe+0YTYI8V10fyK69JitUVy8KbTusuTDdEm+Z26VbOqnQqnlgjZaK
sQhP7AyaDBCaOISFuSTRKkkuFqZeZ3pgfs7lLj9xOnkkhnl0pMPQIfi3R+7imVLe
1Kk2a93SefK21NivXBdIQzlU/A1ECrvFShhHyN+tokNwr6NE4801sJ3eH/n0gA9w
ZVQWTPDf70mKOYRBjHlWUJA/0VCn+ge4fXdKnk67Gfth+/AJwNR9mr76/MlHSkld
co2RTSfgdXIs/G52cnPZH4UWdpJAvYc7LIwsBBPYyZ7KcbkwvqRVLak8dpeixTl2
t+FvG1QpdUKdeTM5ZKh3SPgQNuoGgsNXuSZjtMo7O/6XdgwKtg9eoftNizt5eNBB
92m24XcJoijNPm/oRfOEHP9kialKi9NOqbSB+90HVGWPwqG/8vVdKQBnqzRXc/7G
yiiGOSjpdgfRCbXceg0Cuy6eddznIeEEPv9TV7dHyUY5qKfAvUVklyMD5NkFoxVi
CqC6ZN+OIZpKqH8+d+u/F35D6Lrl+f+5oHFW8IzPHGjWjnMdtnqu270LRAmhoR1a
NHg78z0RQarcHwYyBEupOtZSBuuYPVMgLmhYdpvMP3ew+KWNVYWHKJo2b1begwKH
HGi38kjwWy7T4ObikTxrJrRY+1kvUPG4zP8avqK+Te6cg4k1O/JssypSiFAjhukp
Pf1RpvQ9wa9arN+WyhTVzIUaBaqw0qK/JKA0SRj+noJv0b4Hmqgw4bKUJXa/9aJL
COmMAcer7GiW79/RcTA0DDpwVpGBFC9QylDbwkZiKcBhksCLKjF+rYo/SQo7/vXo
KkPHxWD5M7k0i1a4cCnSD4XdZ7LFua7oA65UQfto2jVxZPRtSnX4eYjMjW5WtuRJ
fxe0R+4pvGdfKvi3akZppaJTddgEtuxW3Pbbe1lBUiDTu9yuAeME2TgkWEQ0g20L
OiCV1vEwzwDrr86GrVPGNkNKuIC9hNtZRQ4ZSrht0tkDN+yCg6HKJ8GkLpbOoNEX
d8I3rxnYtBh4YxTO36hwCR8OhQHvlipbihvC4VPjeDZI+w9LtqiG12jdggq3+INw
jhuVUwy6RXnDsM1hRCZuoUrF5oxp5n0CbA18MBy3ZkwPnQ/oXd7QeH8tL2ifhuTi
NRiDp5Cu8P26MDgUVHQ/fvqEozfe+3aY+Bl8NxmT47BwucCkPXaLgldkHOlRjcu8
VMdULnzIswJQqUe1A6KqJnxcLBCSz8apuT13u/btYzu75kuF85GYoJ+0L/1Fy2nr
B2blFO1JmyPSjOPPWYur/jHhXInGJC6KwzYkhU9vXwl4NDJ1rjzw02O7mKkhauWj
jQlG51YyQB+dHbHccl4uu4Td1rPHz3d35BhfW+83KnLqk8D/wK2wgnGUzSAywf9g
i+KHFQgc5udQDnLnemeQ6Pp87w/xnBQKiC4dOEA3IA+SPKfPhXItbqkLKmMBmzU9
W01vQHUh/W+uQvWW1+SB4SnahexeMv9/IumtYhYOTiHFLHqUYGvVhzRyW4t3yQht
wOIvgf8PhVaMttf+B6A4WpBW6JG210ugmBgh+q63JHCniBr4ot0kBGs3Nn3GTlrI
cVGju+XMdrh3DoahpmsdPGebmbDUv9dvYMvd+G6NsFgO64aEIs0fY+r/uT54F1GF
5HoalQLLdI84ycyF5t0NOYEcw5a83AfzpSzk8RcRnWC+36lgafmpd0kxK60/dsm0
T8Hvk3/PzJmvPXl71iRq1m0nkmp5dh4kWJmngErIkW/0weLej9Qg5bzIOp+F1012
xHkqZMVuEohE9Y4t9burOVFkFcOAwRXEMI1T3v8txS7eWRt3lQ2sWEYKPQdOYAb/
aRHw4siVBbBcI56aahQJYCbAgUWDM4B20bh2z6Ped+7gP8ktobRJTXRXKEQAMBSf
UcAyV0+y4RyPzBazjgN2WNqDPL4dZ2vOp1MQ496N2pHCpwUH8iYI0wKuErWwBdO4
/JbmJZqCBkrukZt3FdXEjuo4X9vSUn9BgJu7qXLtH5jw5/Dz8XdE3SSqoSdtXEcC
ryoFbrqXO6PslF2S+M29Vzvm8RgwpDOQ5CCa9v97EQNJKeIunDyRejgk32jPB70j
TDv+qxdV/hfE0cAxUJj0cdTR01TQCQ/g88bzqHZDVdk98m5AL7+XYKOidexqQ2BM
VBOAkLAlwAoX53QvIPooUW29v+7zIQUZeWu/cXv/x2CHqVUyXnk2J4ZlY7b36TY3
K0uqC3KtJbC/BEo10AUjof8N+bfsPooBJi5loSYCKF1mR2ofond+G/leK8kmpI1f
7fgHbqqXkn1dkKs1RFV66DCdQVLfXbEFZS/1izTGK+ULNg2I9CYEkdDEJ17RaD4m
FNifRL6ajPUw68AGmYeDPBPO3GKD/xG3jIGSZPBX+7Tsro0iZcoEKVq68zuzJCBI
uU6SZPLBCNh+oOm7A3yVKGCwSRVgFWCDmVMIHFhhu87ajl2g/TA+kCGSu/e8XpmJ
jeNKPS7ABmiZtLSM/x+CRaSlnwZCsDv8UfP+F2vISDzeylWu81ReooAORyclgSni
4TymiqUajBXRmT45n58rbLZPqnF5toMG0FNB2RA7LyaIUDSwvVz/zXaqcyA0Z4dI
i5oOvz22PHP91LppAWWZT8VZ6U20t0JjHGsCrX3XIi4HE+Ekf7KtgAmEXD7pH142
/noCISuHO9v8Ur18CyWpIompxQilhjYzhUJn8I0c6mbbEzrxyRmAqdmvCGEubWmw
4wcEOmtVNv93Dj91YeTbSrg2G8Wv2r+Dj6Rv1yAkj6tPXC1M31UANXnRKiQ70fHX
fxdMgaNGiGkhjShW/ALQsEgIWu/7WBCQ3IBtQVgkOEtWiHjXi1xhEGkOY6AmBQM2
/iQ0XKrv2m+CrLXEZxShexxVgHB8rAri7UKAYXWvv3dZJJsNYr/MM2q0UCg8p/PO
iq76G2N6vsq+r6mkbSJXidh0p6FIoVYZiS0G70U3ISu5mjWPXJDJp4sxOeSQKrOt
8VMRUutCttSe70VQuqZ22kXbGscgevc33RNAId6yQTwWysrF/Oa6W4+ykHO93Ery
O7f6SJEQq2iPhCZ91Nx4TsrVgIddv3DmD7Fad8NC0xsIEXyOC+6LzacJzmd1xJ8r
l7ZbgZNZKJX98/QknGQtPRPDVujw9huD+a3NIaw6BBejxmzXxXhtoolcWUC+aOjk
7zpvFsPxUwYP5+t1G7L9C206UWfUupxS+OcLN9c2Aaq0ldIikBrKuHzem4ZYPhgU
b46F9AmFeoVhwJQuLQjpRrBUzNCE03BwFN19okwz7nwTYnlFgA4QvvCfKvwUbkg3
adzMBPI2U1DEhX+GfdNUZ4dO+gJC8+JEh+1shOKX3t92ZUw3uyhzzBAQVJY1musF
w39XytmuUPniItVmVXowdFhmgvvCr1t1Oz9te/w+GocPyUUKwLMlxT9RrLHUuo27
k7puFxyoJsM3/yJsFuOjb/eDh0LYuyGP+u5sJlUWbijMKtttBU55wf/AqyT+DVNB
RCQgbx0fhIjRULe8mj8//CHetG7YcZj3gliTJegzKb+N7EhF0lmAA5siczdo/cs0
qWuAh5wYQk9g/4hq1ASnL3tPpzP0I3fefX2u2d3YvQDGoIq7J4agTQh9Qi+KfDYZ
yqRrRgaCzmDsWLGjHAm7i6m2lG9kLx3Egl2FJ5pnEy+CvQPvtMQGZ0+1nFPlwYM9
sPn/B0t+Ls30zftCbSslchc5w3Y9TsweG86iHHY+nUHCbe9X0y7d97+asLHDlrdz
MDQbNNgnlzPMcnzWUBkv3vzVDEbpFL7Ow/k2JNXO1Ylr8KbrCemjV4JWk0w//0cg
mP2J2VLjm9IF+gXGcSodmmKw2k1IJWzOQCcben6vavIL3xDLSTBE7lNwm2WdMUkI
VIHWWV/KU/hoi5254YeNyx0IWD3+NQ60mXGLJxjOKH6aOING5z5IQ0eE5rZ3z8dK
zS9cltqAN1UayNO1osnCJJ2qXYksoffZTEkSWpd+8sMWhwZKiiKl45a/RPbRuY1z
8Ljvjw46vnG6YXKVOMNY+jaR0Nsa5fopoAw+NsGKeNOiT8uh3NIv7s7SczO6I9jh
LUjN40PHNOThI3IH/vsLqGkThdbnvS4LXVCxLKwurYXBgzjYdcPaYpIrQamCDHcC
WnFpgqFzClaBNrB6i2II4KsQuyhoN/JmYiqWaFHTZamFKW0pZ1guDfaJia83tpj1
OP5+GGijyae/Ga2swco91m+m5t4mIN0TdlVHHl0mCY958VzELNPb5+75Hebd7AsL
rWAuyxrZetCsfUFEYQWjna37yjOaWwXutd7miHiBG1iwLnWUlAFfpXyxPYn2fOfc
hnGpilozGb21+MmYo3hdYbWAvqJhZrNkaO5FnjBgv0kwbfg2A0dEhzc30oM7ZTsJ
wWMiOXaoKkVujmyg+eDiHXToK0b8MBszwKGPfvuZM1i3U8FcgMrBi6//BjDgdcpN
a1NiSkogvR6kWqTEJPBSvLxudxOLnQJBBJ7abs5HNESJj9p9H2xiDbw2NLLejAsu
LCoFyifVBI2oj/wOlH/+Lrm7hXEHVqSs5jat2sh4ZA2F4PgCTjmLK77hky5hLI4B
ZuF6+PpM6/73o7+QMLq8DpPs1nrhCfRM+bJUPP1Ntox3XZ8HAG0UxaTqVpEIDWOb
1x06XcjTsqe42a/fumxOWduUn+DfSQyoO1jAiG78MCtrLfPmV9ryjIwN3tllwrbn
GwCub45a9ahl2DYuGIZIepqMJrBkT2/6tQ5AUIV6ZOyHPZTZiywVxDFYL+eMJ2HU
Q3w/wstD0E6Q26RpFxk0aOnJunjrroYi7XZy6nCWaUdIyLHnqLbKs37XCFsyezcZ
xGPvaFBm4tzquf1ozi8WeSeg38lkaTebcJhvRYUqG6E2jkYgVOT9pGZPbZ+3xXPv
jCS+FoLy34I0xcS/61ooDfkSnpt80gxNlb/H1loZYXJmjk6BSfgTmyt8ocvufTgC
AO06igabQmtxTXIr7Bf3w+qnaUgFdIqc7yHnojTnzeT1Hzi91s6WZVzdxAAQLX82
SPo7RefSlGeRb5SWNIPRiCv4egURijapJv0Mr79tQ4XSPPwUs2m5PnFJWIZjY5oX
/Eg1fn5HrKNsIqa1CDY/IDI8WvrI2TYu1whSHeYvFs+zDIDxiAfSmzaq2BR27xDe
LhJ23g9TpmP1f1eM2GpHIUSF9nocXzkMCrxSOu2/l5Q0gdxQKxTmxSDrd+tu8Rl8
Mienc7LKJ1L5cWgon1BLDV/A757Eqf5QpqLv8szZg30QiAdTczOGeslR1YUN1T1O
CkaOBDGhT/bDCcZyb/Q9YzFpP/aceF7PE69oQlMqMsuOKKzeSM9ROVb5AIRWsa+W
LVOixtu78Vu1FNEmMqKopQeJsmKzFv1EfWoxNu3athQmM2AEYGFTZVXT6WCCbIkX
llHp+ZprVGTb3sIJPemHK1ZSlP+j8tqXDxyUpqTMJSYrmpOL2A+9Spee9yC9ij18
XTJAvdbaRsfP/6lxCVDAzkBY5Jz8CnjQhqxIuc8rSSlO+vun4raMM8yzBZKb6uQ+
brHvhu0VUhRUePJJzh56MkjRpgQSTpqmVsnU7swwwEEgvFiaUl/u1omdv8Ebzi1+
POcIV7f0L14FT8c5gL7GS2yi7ZfGtsdItqUe9mYqqbZLUORCROwG8apdZFTFu170
TkQhCC0FmJhNOXb7+w7wMOLk7RKL7AMJO0XWrv6iH6r9TnkSH55eIe0k0nFCRbcN
sYxzgqKOIV8Gcz/9UFBO3bzm/SdWiDu7DkXeOXUC7ycimCwY/rijbQVp+vMNUeNL
JmWxCARIHXdCwA1gei+GrgIGxd/hj/ysoJ0LaQ3TFfav5LLQGty/2ESFoRspPE67
K+zdxjmY2t07Am4PPurVYO/eNd313z5yslzUnG7yMdnac2WHEJc1KVD7QxvyocK+
tknxBQr5caQSy5wnmZSe6p+gqwg7SbNF6xpaal/dokp0jyWNZdDuqXJ31V2VaabB
attdTP6blGe9qMtNTEGMyX2RAfK/mXHA6eFVRhU7RtEdvTADFY95Nk71fXEKm25W
/XeInX46AUpLB2I0LZHq9baCZuy8t6dKAaBLQ+jsPw3uhPqbR3Elh2EL/6Iqfho9
Hq0PsZzP4wW9Wtj2Vta7G4mWoOMN6erprIj5X+YP6VnKYN1zQj4ie9o8toMqUedY
TgNvHCXijoBc7u52wQ+7pF4Y7OcszD+sbjVcJGTTys/08gCJV10N+U3rMPfeTdgv
aX4cGjnYa85LywvvdieA9UEobCgUwErzF5SM9LSKeNAcsEcAlVIrRPNAGRMvIhNn
Nwud51PxMA23ROFinn7YJoNOC+fpzros8gfLUJVKWx54kSSy5Q4mj+YRXZfS2wEH
+FctQ0hTnb9/il3DFkXpdHGDcILa1ujkcG0P5riE5FpH1hXgKtRovhNrBRYK9y8v
w32XS51nAWqiJZoD49OqYAjb7eQHT3RrW4v6FBtQLtJkNFGGsc7dlCTX+NGt11Tj
mkoOZEnXwlugiCQuoqZ3lBwQ/vPlEMTG+dKfzF2ogJgD7fzgJltFTBMWZsgGB/Qs
EqQx/PadSTxFYxiiOtygVFaFQsHdV4GIBfWtSPJosVmDFAtM64wCc+ZHoYG2xpqj
PVQ/xf1UAWwJCovaVnLGrKbXu62x4iNi/CJqz9Dhqasujm2ixC1Ep9KyLG6MqC9F
nqXMv9lMgFONxeGfNC2SEKia+tRoCusXcpWHx7rvqbllGm6vqcfqZQFwnnddKETp
ii6h1J+mNhgHmzJGMl1luSr3JPQljZDcnyiYtPOh72roUmuXWwMGatGQRlc1ihTP
iVFHj0LG7JOvCVCz0lg/J5EMxerfAZ/SD1IWSwoxt1lkecpQhYg44b/3BAIiSj0t
iQ/3+2WU30cCx0RLUVb3HAmyLb/kew4zKkI20MkUxgdnjoaZjyXuydw3HvNksT4N
8JWPj27AKqayQBaETuA9vIpQqWA6bvXrshkeiudKd9BxwA1YrEyY94YtfnWm2Z5b
VotzR+g5FvqDAS6QS2dqxZTmxCtNuoR++tJecDC0evmDNIylQyjyieP50GUp9gPa
YJiLc3kZlHH+eyfe4cr/55EhxdQHkn7G48C1/TJ9m0LkxGmzHruayoLMY8TYQ9QC
wNn5LlySofloA666sm6jDgYjbD2AP/ijxeiYVq832QebS+MX+50HL5LHjvf5k/vh
+43WWsas76RP3VkgRp/4kFQTvPz90J2KuvT7exJO3Aa/tqkhLqqDW+0XQVV/N7mb
l3W3T5/MUrWhQ9iBXbzPskldUAOrhZJRoEWsxYhr4+iGL7LfSKzHQc6HA8b+KZlh
vNrW0wlhdkAxp3F9RoEkEZQQ/AwNQpjPfIKVee5fLZWVt9x4lVb/HIZ6zLoVT3U0
8CYhojqgprlAVbhTbHIFfHcULUL9vJShZxl6Coi/la4VnYXvFaAmB5+soOE1wevy
yyaTM9Fej/Goo4MTXosH/SHN3fhoSoPO902bXa/NoXWVf+XHPyeSU7rnBKm31K6P
J5XcRo6TPyj/CGzGyJLLtcNiyiEIizzpcek1LeHCfd4WY4NGfUjiO0RohH9bVVZz
dsOC/I0b32WrUqQAjQTpblanKBBHugW5A4V4jB7yvgebImJm0XV9CCWo1qGWakWU
mVFP2e8bL25s0qAPYqZRd4AVqxpDyFmfqWLBrIQXwXUXVJz89DpuZr8VAlRlNMKY
c7WZEHNZeGVZR8ol0B+fG7ddMuU8jKdyK3uXXji//hbgkj5lMzE5bVlflWtOSY3p
E/cGSGBCHAPMKoPJT2985Htyd+2PS+iH7rAk07HNVVogOM5A/8iR8wcedOuVO8KP
ieNEMRGLhja0GI9Bkd4d8R9WITbVo3KvfDIWzuII9cUzC3b+l+BQ/kqweqRjuKgc
Pl7EgXl/ejyqh2Fa3TJqog==
`pragma protect end_protected
