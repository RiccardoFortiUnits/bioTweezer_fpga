`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h5ozjL1B2VgFPsQerW3n3MgJ1Mg9r6NNfQBr0YvMs2QDYJXKe5i7WnhXaReyJPA5
lGoj7sMIy69OFROKi7fKVMoLB5QPDPBXN5JWAQxz/1NcxvzhHuGd62RvBkg6Fg69
2yH4L4nDb+C+6b+9XrVyCuQEmXHqGxYP4pOPWUo79pA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71088)
7nkYesZlFwOQ4YfFyoxb+hZDQZYe6zlJy6D8SKEMnesjf4psgyxNJZ1EHpOuYMX0
rKWlZbWNSRaGqNd7QrzrXqQ7lceiErbXn9Q7ZJWpeWO2SLJs79sP991zpZL3iP6d
rzAIbUJzYQJitn29gXy9G1w6tORHFXgKOPXmXfoxUEszUP5Q3Z5fK9LVS6ewnFPv
JCE3a0/o5r4aH+Oc8VC6BkKvTMSf+o/9cVYvnIkREa5V1sotBy/tj92o+kIi/Zo5
s79vEIVmqqIbTOGXKLlqt+ZgSnXp3m4FGPBdrx9YhXKxKtCk7GLpdIOqWgNIfrl/
C3kJ7Q4hvHTPFriuH3RmnxCEgQEQ6XyNIgUCuuZfGQbu6ms5YvyJgq6lVuY9NNau
ukbBVkJIaWZ9pwPQpBA3A6MFQYYUiTHIe6zEVFO+dZ3qlyQOdNbVA4sDOSDgT575
wnbW58eDtaY9A+Ab0DsADq0btNB/gOhR/eGr8Lr5kNNxgDzmRddFbVypHd9Lh1vY
gkKX1y+PZwdObruWMPLgRjH/k3bWb9lEMTW9tBFUZdPEQHzduiUlnqm1SnGDs5Sp
kOuMO0CoXXTBuLQL8C51KYKLNMOu93ZpcmA3xRiV3mokfkDe/Jv+wDywsOMvY9iM
h3bQ7pqOZUHAvbdQPIF9TIZYQt+jb38TRG3xrW2tMrWMQr6rkgHrthJP2tbpESur
fmJh03a1P5lJNJBpYvRgYZqqGgPdzvaPcTywjKqhJyc1pJWuu6GKxNHCFV9ezC9X
oe/0Q7Z9MGdGL++VeU+RWoHodv7cdASnRt+S9a3zwK117UtcZdDOxVBhn+e9zP77
Ff9j409RU/txANej6vJju02EHUlYFD+vlQ9U98wz+DQXaqU6H83kbjjQZtF7ECvk
LNcgD/hwK10yGTKwPN+aCriD/COyTjTho2YZLDUrpID3z5+XXVcVGp9vJX0uEzQp
75QDdF0Uaw8HjQh4I8NvR+E9BJH0zi6iTAlBiNdH5rr0S30xT4QrDzoYndVOsBso
Nnyi2E2k6AFpJaTD2jcVf/kXl5kwdJ+Pv3Kn91QLUhQ6M3gRRnh5bWH3DW6f5083
XDiXkEOlc8TtLMUi94oHs7O/j8Y26ps1bqkjWY/73AztoHH7SHNTbNdkMCFXxPn1
Ao/4/gUxUBtg0qaIhlA99j4hgj6h4cFhgulX78IOFOyi7cWu3GLy0j2U7ZHCgPZt
O3GeBiSqF+ZPQ36UZHCNH2sQkRwgENnwLSLHXmg0UEIOie+55+foWxdJDKqK/jXn
r1/1B9TIZTzbg0WlwdSPW5YZ+e2VH0hSXocxpjqHTP999sWYGEU8hKBHI6sZobtq
kxP1ycpAydwV/IKGEO3dB/ZZzG/ct+DCqYyQVcMBUeMEP+FkR7z3MVTGhsC6AA4A
IJmPW0ByqRjh8Dq5210nIMH8HNlTdWSuR76W6p8/pq2HNMyCD+ktcUm2DdmEfduG
ifvlLJwir7eF48CEsld075vWMhgJiy8ZzWCVYsAg4WFQbXggOVtkNbYWJRYFcJ1W
9tY28iNde2JO8oa8xIhMaM6AM5u+IuxX/NauWNO/mrEAOAFaMhn+ZX18hFCbqX4X
8SnI/oVIslFobXjM50W8uikY3bOGhLL6Q1q74Df9AadHQXWPe7FOys09Hu6bu07I
Wc7qskaK6pZUHcJf/aH/GWo+QAgG7eK85UPRFBjbJnY9eylTvd9/84csBQSrgC1a
Szl1haNII9COhdV+iatBQsP0DTdmHYtoiVgkLL5+TqgOygK4byLlffuTIzCEZybn
qM4N5TVzfU+9K6Ah+53KDluyZ7seO3ggdA92znAYDgCEa/02ggoAE2DpuNE0gU3+
lkmlhd8VgPBf8NAol7mHYAxFwSMfd1S6r8sxPcmlDNtmMxV5CRIDxQ3/oQh8/uqw
f4s3uOb0FpwDv2s7u36sykZOUiHNBhozM4rNginQTbjSm/LpHJqSFiRHr8DiMjNe
rzKfnx+Nywe0I+e4VfDGGw6qiEb/jsxklM63tiFv60sz9hbz/s0EkljOQ9/xC4Hu
/hDHEhuFpmsYzgHu3SX+DKWAe3j18IPmvc4wF5MSOYyNnh3X8zXhBC9iTxpRPUrZ
IeyYi+K7ipdOZzfJ+aQBb+j3ZRaiiMQCuQj67HwiZfj7JMdvfQAI0TG3lDorsbEk
EMIZ58Fvh3YleHWkh13qfstbIM7CS8U5i9TIrEBJAS+aMWf3czcegiqKcaikdQBX
8hOp5pzNkh3rEk9rggkfPO3jjt0KulY1R21pIKWrtOXu6A2k8bmS9PR/f8NX/3Il
VueOGE7VxFaf8IEXUdQa6VT43+ziHYGKu14nnXBGylX3vehPf40W+GMLyO53Bxz5
lhA0j6K3XMOMiO4YvN/BCLOnOv96EgZu1Hq6GplGi8qqPUO6tWHLvSb1P/dXzE0j
XIc9ow2zdoGy1VzbLcrFK+DvlSUdwBQ+hEgeNvCGFDc5cEhfW6V66jyZIUEZjbmi
TQxhDcJX8GwM+6mogtbNcrszPlbEGTIRPo7aDZPK8QO6k/DiztZ6H2LzOPUG7rnm
OtdnOPVmDxDBeBGLm75Xf6vK7Le/nuIppkYttTmg3FHv8Qdbsv2CE++fySz4Kg9z
EOL5982PdcoTuhlrEf+xfHIKMhjCYnbLiYQGZv4eQiqqAIqkB9Iqva2rpy9m8MkA
GZ9F39dmdBJxKc47w/klNUZYWuJApUkEQeg88y06jQ8FOKDOKqt1neYMJOhAXnSW
PvZIbKKBQxZlfq2C/lBTzjnBOI6lPevzRuTnRCBlj4OvWIsjXtG2ktGx1e3cXMw5
VmNiLPmbLKFl2TGLYPFJhlhesXEA7n2FFhyHf5LUhJ/vs+Q3BUttI14mBki1jjoU
X2TgrNdktZafNF/CjSbGlgdBDLKkuh4JNCK7QrihgSgQicnXCQWYoGadc8gwYy5I
4oorJ94hKbAbtm4KxDheJWf8s2tizwgJxDQiPZVQnNFJ6PiT75Pgc4Bsh9MSEAiG
VjeE9Ujl/qaJz4a9pVA7CYvbBJZflqTDwi4+nJOYJp1x9ojhgCjYJJgX0ca0OzJA
hdE6DsWVx/hPsQJDk1sUlQ0+jiS+10EoW3pTqGGnOtzkuY8IsFpiojYBSOIwUZu7
qfHN4S+0+CP5yYhmLOaHVh0ZAkhyAPDVRTXeHvzcvF7QnDtocpozEDFUPUF4jgfM
fwKFvUeBOHdUv+7O4mhw8+sv70GE9PuugJ/W2hCtRNsip9nUHcqk1RL8NCyqU50A
LeSQr13miBk1P+mXSydhlCctVLETpFkEvBYRfARuYFT5F7Q4ku1Z18HMCMfZ2ddA
AEuKkUg8vAfKsuLNik6FomqpH7oFW3GwwofeOw4BVqmtw+/u+phDHX89R1umQRyp
JfAplv7BwyDyMgrmjzoMVynKjSMSSuKrmovO/vkQ13vjMb6BIAzMX/29KDM5YYrZ
nfLarSPRtOky1lb9JuObawluu1e0dMQDs5XNWaHt3CNO3OmGeIyzhbGIo2Qa05je
lz/psso5E9lfD7kxuBx2hm/qsQAM2bK/U+PzwCjApHw6fqaN9HycUrgtzWfaqqcg
5huNtcJjmX0miRXZWR+HkPfTO5AJnX8l2JXEane3KX2IGrY7lmg8mHPfbLJCq/7y
kOaV8gKn05nS9LGOQMF9HvmaHv+H0P0+Ymqox+W/XCH6PwDRp1ujpN77Y+wPKccf
fHrnaXwLUfeVL+Gag21VbaKsy7f7ryVReYxh4zdr8mv1wpc8RBx5czIj6p3FaHUr
fuHiHLBsToq4PwFishNOwCxEBk2qdFF6GIM2wXdqLjUm+W5AYzphnlpf2WMz9agm
I6g6cP+yIrrXGMfSLVXdUr86JICJ8dQudrjKDtBS7ZaBkE606amcU0RS/cYaSbCM
H86kSPaK7zfCnA+icaDoJl56L4oA0DswFmblNYEReG8st3rwY0JLKQG/49QRl5cM
MyTOWqhhROSMiMdc4cy43Mn+LYKERyHTQBobs5GKZ2O93JiOzwo7u0EVX9WgVxLG
YzhonXjkEssV8OIsE2b65+XYqyv9DVJc99RU5QJtS7s5q5YX9SOEoB6m2hpso6iS
0u8OFMU1nWdMg60/5C3qSRa/cy3tlG8BsQw5mSNbOOpl9tFInfv7N+OYgStGtN91
hk9lZ5cpf1YLpezisBo816KNH742/fSWa5PybIr4bAs43vVR9kZMmIziDPSOPUH9
9QbFaLdkYrT9IfhsnPy7dutVdq4AQq1RMoR/cNc+xGO80U3eV5U6/Umvs10ZSkOW
MgVhKCCh0wF799cTmZrL5Yao/9HQkabZ/N0GTXZF8C2xfP3nRxyXaQ/AcY/95XwQ
wGaAYIeFi8uelTCpMuRcjd7enF3nzhyDm5ZwLXc0KD6wr6pevHiG8r72m3DMGJvI
tBKPcma/CLu8Cl5QrfBiX4Q78zfKzko9QJ2rgrIdVhp09En97TZK95f7r1IdllEA
Wkad4i17BFDf1uHOP98toSXEnb2egACcTxedRZP7cPPoSShfGRVf4E8n9/dBFfP+
1CYxc4gcXosR3mFT8LpNQUH1q7XE0J9ZzQGOWxeEH9/jbsI2dGDaDnAtF1Q7qH6d
QO9vBXr5kIC9iZJR5p+z4MQRdMQKToMdm5UpVbLaADkOoc3OTDpjSrasawnjre5k
kLv0taZEahXIklp/Q0Mgeej+CohgOTiLYc+fR8Gp0BfiZ3Y5MTSmXub6ntw7GgDe
FeJC7VJxq8uq75F/yJFYknAaIGD12mgZbKgD7RDX2bXd9mUOW4FGiIw5zyBECjRU
TDKSoBbdul5PE/Ik9Vi1P2hM+OjF6VExqD6Hbb/LHbAMdOEvTAZvI+xULt6ogkgp
IQ+aepU9uHCRFSJyhOBSS6FQFYMJ3tXz6tKqhTik9yGtClKyaurZvILIuvclymro
jQcLYhGaBvbULqWC/6uPGQrPUjPqgC8beiNM+KClJnjjqFtGSErjN/Tcn0gFcgKE
0IO8ftUs+/jdMA8ZI2Z8Z2X1jjUGZjZ4D0cMISyRci9oHqbudbhZ79h6eI4N5VtE
qgbKbG4T3vnR1x1XnIKVai2nqHlgbqZvFWHpZOnRStbnuVIN7Ebu0sp/4nrAfqBU
r9e56tUxgfAcq7MU9+7qmuvI3GEsozMXXquhL5ol5l0qm2P/6Ei/e1e87kQlk4M9
prCDqGmWAIqPV7fXnrM91O0WvuR6aP5+jBb0wsjKVCqHoqamQEtXgpQsdJtEpBd7
tVVBaev+XsK8FZiRH9NSKhluj8lxWPl/kbxEZDa1JBaS7QyunVoLb/b0BtDeSFI8
j3HgUhOuiyg8b9FX6ApZlEaa//V6hnbNaCfQG6yq3R6rednYzvLsIUcSI9DT0M6C
LTp7+CPkbPY/zNVAl99BZ4g2ViLYLosZlSUGw5CxvxZJv0dIn/rptiBjcrcZrEVr
0lJB8HmYyI4jZAaxu39ihrL3ZZ48aoALIuhkdViIcg9XhLUvmw0CGAbCqVRk/ToB
/JqeWT+tYp05h+6p42dap2LyXkcg3bQAQoX1dpFzOIdXytq2D6o5W3NFueLPQF5X
8xPZACBqvYqnM9WWvZCIyc9SbcAq3PpUReQyWGv7UZ+e5WhF4Gdy+RwHqbX1RXcx
x83GyYt3qmI61/Q0ez6j1lq3obqW/lawaF7drYA7BD2qcTcPUFDnm4s79Xn3PM0u
50yX6+kVMpyn9qFFhnHavFMZjNrF18VacoRnowtxqFYH9ddoMfjSf58wu9H7QOZN
gQ7b5zWdUEkxLQtjZtB0T3labcvj5GUeHak9llj3/SeCg9aoDo1Oc7wCNOVV/iXp
Mcd6BRYXPM+khHVrh73zj+H47ypOWcN7lDkAzMXz/8Jdv4kdfXK18hPuhs6b7V/Q
N7zYGbfCTDE3nZT2uKfZT6T4NqNalMX6AVLYsdd2tOdybDasQg9B7KcJ8DWh54Yz
wjq/hieKWV+xLfntDR2w7oUJseWIU2Tt2n+3oj4N4mVVDWU9swxeXyK6A0fju0ms
Ssc9Kag/Ro9bsY0WdzClHUgn5U6TeD6IuDnWQ7VKn4OpqSus1X3BLz79ld5qzTfS
JVHqFEJALyetP20V3CtOvuA+jNGV5140kuCbp8X0vlvY3hGzgoFxAnW/WgGvB1qN
XIPHf6krfPJjewtJUZ+76Papg0sSPvDANYzK7PoK1Gkfq2MhiFYodw1oE8HbOPJ7
3omOHxo/aVYI5yQWBQ760juREsuu2K1056iDpLDtAMiiuxiKswlo5bHUqx2p7eEv
uqd+jNLP6ioUNH0zazDma4T444hvORziOK7EMLgBJF1Nj1z/V9/rCVv8Z/5d7yBP
Gt8Dov9qnC2Y1n/I7eBdl2fxZWhBFeoQnfyrSDw9GGs6DUOQhPxs761j5mq3aUuy
Zqk7O8tK99ieaIuHNB20kIaV4LQolHiCh2Q65ij1rI23se5iYRSfjZSXXdABai2a
5VvzDuyyjc6wNUrqeYOxkm7D+hWHitI4S/L4dvSTl/uEvyseCzS62c61yb7MyCS2
Cfs1FiVMb/jSNwk9UHV6669JmnGmWa9k/m0ZU/jX+Uosv/1AVxm6k3RmAEMHicwQ
mh8JzyZKqKx1ePt7tIUG96+1nLQBojXsZIsR12vmGdW8wBaFhHlqdOHELlEMmff6
10biVxrsnx5TBpcIwXKZs272d9fM4jq9HeYgLaCmgUtI9bit/p2WHypT75BgwrR5
6Qyi+o3GjPbD4ik5DOFyJANaSGyPOd/1vyStSujrpWNfXGcOozV5fzSPby21RgbD
57N7i1VEMs39vrIuxO5EbYyEOnryM3715XRz6d5StpCedmP1UcLJLTBmkFjm8NkR
jXiGOERHcOtDKL/nn2YCK0jqwFK36DVM2L0vCA6f6/H2wV/sbFlNq0m6Xg/a6SR7
rgMzKIEYZly6M4IKE8vP1y6pjfhNPiLv/Br8kq1dej338+WBL2mcOjm4XP0Xm4l4
hHo6wUoGBl9kRTzAk4tZjEn5y4Lcn8zoGlUiB+qOtnhXFk2CNYH7R10QqBqN0f8e
66yTYoI7r1H+S+cKFd8klvjoY0b+dIgh9IEusz+G5xNey8KawhuyhyNvqQgo0AIG
eYtaw0TOruetYvAbDhOwKmp6AJigRvxqfx46ZODpMRFk5imsY0MLgpU+6f3WXguZ
fYKqEJxHh3zn51WePql0YiabHRFgYh4Y9z2QwRLhqJVl6QoowwWCwKQFsaKGcK8/
tluKlIsBoCNhaGtgd5WFTvK/8gj3K7Djcpu2vJ655odD223ilByWEVwTsVI95ZmP
2Ddm5QZYTpLd52ay68eCoAmHBzWOmQG7e3UDa0FJ6cdtnpKh3LstxmFBt6Bn7PNG
eCvGDvN/GxHSDGsp0STuu9vMR+VV6J4+AQcaQCF2jDf7TsyigG8++4KlayR+nthR
Yrth3yW2YoCutfWNIitYakGeFomh13Y5xQnGxxLLFLbcjev0kA/cLb0U5totzlfD
avupCIIRKJxbDsvnpd++hk7s25bs6hGqce9w56xi5lHp8ZHLC7BrI1qrVOQZL1gL
o/WvQBxTHiUmZJD3J5p5gTZ0dwuAgKN+PUA6YhWqyclomyHHYz9pRjvMR8pMJkCp
V5nHrSI2V3bBiJ9i30Cd9TYb4nnR1UfJ/yizEKiPCv/BI71BoOb1YlllqyFZOoF9
H652J6T2IzoldV9Vu5d34S5r5TFcfAfBlyCfaNqId431x4zHJ38a6uQy0lOcWMXU
HiVo5XbxpLkH37+OcL0hiOKj2xis0HPxk1Cp90FIv6VLsTfT4eEfIIs4eFucMvah
9dD9cn5sIk1T359ecG2gc+Oa+Dlk3SzfaNUiOTbn62wdq2PzhxwVD2Khcipgi1Jk
r2M/0RIWtegzZBsGKsMUiA8fOVH0zOGrorTvO9kWi2aD7iRz6LjvfR1LRIYKhTsx
ngi7SHZ1dCkfpBMASV73xO/JY5fRzaaXyLr7nNAV3KdOPaOxOM5E55UaTKOYUxpk
Hwz9M8Dal+wDrZ4HZfFPogL3xXk+MMLrzgN0946qV6nlO2kczKHe8WkaLIlCSx+v
qONXKAi/hLKsraoy2XsL12cGuqhWpaYo4rhsCXaAAnjvXSU2yRSEBSTIBZPqy+Ij
4iueDbQF2GNk4yxlXvxXIy6dSSlXAH0eqpP624JdwBG8Dav0NKTUOG3rRpd/zxCP
QaIb4HzxJIqVSE92ROiO3vXbFdUdV9NW42aIlJNJEHBpHRe5To5xLxxr3mF/8GB3
XLM5bKtAyLmmOEXAJfhUWmGM7cPudNxMM2RIED45dKifdPV0aoznKDhXlPXQeA4V
Cu98DQ7TuHgc4VnXWESx2dIPE8HWTodidTJf00nRGjOAPn6DN7S4oONIWRDPD5ZO
oEGZBWWhobcwkOf8EzsLuSLUhfrE3cotJNnkJaxF5hU/5IBzU/VlD4Jr3XDeuWqE
GHA1icWkoO+ymic1UsMFNnplNIvG1bJgVSkcdj+qMhbhViufh7xeIVYSAaSqjxyn
IykmmS2uzYCPKOI4XFUakTZvpbTwBrwBKepirPtFIKFdSbK+Ch/nCuhqALS+MCCX
xLvRMnF/YsI0jIDRpdIhf8Il8wjWbJ6EmOa0KA5hKP2ShsAMf/hSDlmcKHoXAyec
jjuFAaHS0avoJAB4Jf/BTdIeo9dzeu+7lPdwSXrthFW+2uQmlJCxVhoCfNlYD5QT
EkTdfVOvyKYxz1SOz7qM9AE52nt3/QQIMLll7l8gypeNAQTwHFurTNpaSDHtnnoL
OOhqnc6aFN362McabdpJOASbjs6185hZxsXwsjNVngI1tfuDraFc779qBd2FQNWf
g9ZKyx1WZDUa3/LrN3slA0OxwQUIh880DQpC+1E+UTDrKG8MzoQ44/bckUw0nG8O
lpRSCKgcmZVFetM3gY4oZzIMvxQZMgBs5gdMJAZME+zt+SmAvGGDmbU9xlKZEvxD
orPMAQq9ervFhmB8hFN4QF1ppJm7dAi48yarPDywuAX4MS7dZH1Jk5KZBiaMG6YQ
Gfjhxhv7jUpHr0fMH6iArqQnksQBOyC7YObSp+X1vP03054mQxfRQ6R/fDsOtcEh
Bm242gaGqoShlq1KOeDDovnPUGFVqgfwteZUbMAxkEkRXuGR4o5oOFo92T6TdEdU
qjiyPfMJDie8Knq/p1vxz7ZgFEExae9mhdDOIr61D9JHuaCGLYutmGrFObMp34q0
JYkXYi91WjOUn0IkDLMaaCX3QWg6DlD2PdowczwbYV0Q7BcdkkB47v4THCG+Ldxh
MKXb+/BgmacG8wg2trkX6zH0pu0jp/X2SrjmxPgZ9eJkBOHcMk3Xy2vRkjlRqgnq
N3dwLvko8MIPZA43DE3bWj12C+lKBp1VDAedkDxRfM+0oklBVvHbIO/EdQGtSC3l
Jv8/VfsPBVNUfTTt6PVPEcbE84YB5LFJ/pj91wy+wqEdwiOOl3f1erLfU+pF2+tC
yMiZ6CouevmU+ysJgxKNXpg2a1S1oG5Jop+1B7FewRkY6d3Z8CEabuQGNvJ2N9et
HC9RL91KNRJ5QShkSyYtf4PYdEuVOimKqksixQ7gfwTrCNTyUxZGpiKnmtS2Yoiy
Q6RUP5IDAyG5lM/pn5GPT+vP5heeO+0Tr9G/4HntmxuH44ptYGL0qFSrk+4ZKoG9
tH/K8gnbVfenuYIzRzveNa1CuT0700lZHaqJCP7DSdsFUdp3aYzo0jB/LiMnMocX
oscsbR8KP+/5k+y1LU1PcEbrpZz4iMif1ImODkox1gnnD+UEG6TmqynbKR3/S9ex
+Qd8gn2J/j7RXsH962qYmIj0ygUOPw3z1JgLG8LcokC+grW2gou2vx5ceaulPQF0
IUyGCF1nPyKM9VDaFQkLBNzfcHfPIqfAnjunzy0bXmZDDkiEc5j1K0Yu0wn5zCfh
udt/udPtfPwRRfJp1m+T9Uc4g35LgiMujTGTnyaytcd9JTBPUPT0y61BX/l4OBAv
gJUr3ZE1wEY2xMC4QzNpb2PnMLnGbtCGzrRRQUCBzvDIc+8u6umGZVbkLvHLhNh9
nuEuor/PWQPIXwGTm+vIrgJKfkDG9yrLqdF72jGtf4tcEYc1woqTv+dLtOtIxcry
xkDlD0LKyJ3oYq3eJoFTnrKipJrk26LLANEMK3d6Mh6loc2gLtezJl+lg1tbx+jV
ISC8MAZxBUvC7jx+SSUs7wXBA6PiZNa/wq0Mexqnj6DLSOZV75hkI1NWqk3V8n88
PHRAKtXMl4Q4UND56g0JRl4Ep/74+6hzuGwlVDPJkrlvYw2W0DHcVraCwLC+G5XP
3v/D1wLK8hMuW0JPdDEQp0BriLedIIEGBcsYqYo2zCNcTk+GOSbksV+Tn72u+M/a
N70E/e4qsXz0cAo/3lPQwSW2bqYZKPDroW/rJ0j0tlY83B1f9/ZIkubTbVc9mDWC
3z3wajpW1EftY1KhF5dJCGKzY3199WYBgjmG4Pax2e5dXf+JOZKRjvCSjEB1BOqn
OSQ5+Jmq+T6TNy7CDROlnGpeMBggw9JUIHTlc4h8w0faWakmjiZzGC+0bdtAEfjP
d0RxApUNa48U1YjOmkCMcY9UzG8v7urdyeE9s/Oiq5LvLOe3pqeAHQn4TkZYUW6n
QxWQVyOdNl5eNWEgyD3pqNUCGCp/sNbIPa8KIaW23IEb7CtY3HaI+xgquJfW84nu
2mUMbY4AAdTvFDc6vDSu7UVeTqmm2+ITnHMd5MmMk8QP8QxMmGL2gWbQwG3G7wUD
5Q6ia8euuJnepL6emsrWhvG4Ib/DFtJUtX0bJxwgzY2jeYL+OoByoYCwyHouS2P4
NLWONvo3/lgItjqMtGh/GVmhCgjiA301IwLgzHXbk2UKS45MIUNwhTAk/cw9N3Kx
QBeYCbzWJE1BLkTE0p7FAziGwBt9qd3jAY+zRh0LDBNeOmBzjCPXGWZ5FgjI41C3
mGblZU71KARX6We8B8q1LNObbrvmGFfafhUKaVnT3PJ7i0uVRJhE8ONEFh1z0BER
K3vItmvxkt66UvntvpFjH287rVAPnSSHj3T2E52tMlnE3ZT69kmtoCUldMeoNvPL
gKjVpvGBi6A74xBKWnbLd+oE8Id+mCiF3J3Wz73IEG1MIUR8NZwioRKfqzA25DdL
644NKETdHPzxP1MBCEoqCBQugkf1zw6sb7wIEzW3xrwuo18TvPt2vhJzJBy6wrYl
WeT1L7666JiIplkYrKiPUN5Noz0+6NnMBaWT0T/5NTL7+i2CC7yCcmtJs8WY5df4
W/q45SpQ+mUOdIqYswZAvyC7XtzTD5N20Pd3445Kp+NM8xTZrZS0Pi0AGJJBn9W7
v/noOl7az/UaPPWCcLuUiHVN8Vet2iAQdVQwqzwJSLhaT4E+ZDb1YtznRQv1TVTY
LGbwEoCooBOqLzHMjZIZeN73vy3eeHF8MeAK6cAFm/hhHVy/sWWLolaMO2opcPxF
P/3VPJEe+Ky1xUqE1AWiEfdlYdo44XR6aoYmZaYi82WcZFN/Dx3u0WymBd+py8GS
UjSctxo0L32D5NE6jeLlXFmQu+eZlXeqXOGMNivScf4i/gt74zCP9iSIMbOGmHYN
Y8UFWyyX4/Zs+i8Lk5TIgqilH1Nw2Y9BQj6ZnKrxcECfuYfHE141sTP9bqNODFMx
yl6vGa1K39xFVUoQ7gfMYE6pDROXcGkNNJ7+qc/4xE0Ak+wsPOFwYaEGHouxArk4
xdX/H1xYW9XXeZM21W4OTxCyi269f1sO7C7kmd5w8ZZ16QDyvj/peLWMHHwROVhE
nyPJoRZsWp+WSImC8H4n0/7/QAf2gJtus3b2w+j6FHyPQ9ecjBV+09e0u4oQWyxr
x8vzRTwqcZdBzoEelqP5QQCNmKaZa8QdVq3bGFtZp3wqJ6thbe4/pih2nCJwcnoQ
LC2KsV3WULOApZClrw0mSLqzVaI9UjIKLiA53sPzZEPHu8yeFOqooqGPzVqhVRpS
cRy7JL01R4fhTgKh7QYl4tNvRphAr/blPOM2cmY6aiZSkY36mOl49rt34kZHPeRh
eldGdCwio9sQYRM+2sDWY5ArOncaWhQnXi5Y6k2cRnVKe0aERnkYcSnQeqaHUQlu
iD3UYTdHhyIwB79meVcyfj7KYWDWrn9hklnIpiBJDq2MSTFdRUTsbR+meDYqXPfi
eU54x1YeI6OYN8tjQDSG8XaRNmfYmjSzKq91cwE4vyeaEOvd+v/TawpcFKs0AScR
KJ2w9cOwBucBbf+YxFGP6x0le4PpoLnHC54VJV1CoDzQ+WBrSyAfmZBrFAHpmexZ
9SWy87pNYA+jTkVGL0gcphroozk1NKHXDYYbuE1dGXS20twcKCc4OmFwfxLVkHHQ
ON57io88+A8+q+0im+Ti0dxGD4yXbITbAQ650jzNNez4e/xce/nXNHJnqfBGRHZt
XBB8KqiXqeC2j+TpRSSe7D7aehjDg6/JqNRtQ12j7+961oHTti56BX7IdYiRprA6
ZxwtadKa7tOCmlzf7eWOjLcpmEJ4IKJiBQYUo/KoCbJwQp/oakMipm5o+Uw45IYH
SxQLD9bs7IqX0pn4rfeIcxZNQxJs/F/3F3MNovD3Lz+H/0QWpbwZXN3L9DSUWC8p
G0psQ+Jc4SqmSuifTNgTkJGHe5GZyuQXvj8mOX6c8t1o6WnMsix6XBVgJ+xbrHCM
W975OU13v/20askqnx4ffo9yw9We33lQ5Br3HzX6rBDQumnHv763Ms9uaTdUKCKW
uncDcnUZHqFrkNADvJ39ovfhEoiGcMi5NfEBPjUqjavjzuHUQge4NACIiPZNYkHP
jrCrgv90Lz9E++YbcHPaIc0v+9AzNOVJEgh5BVP022W9798lKkM3YfSInqsK4kB5
czai8tvwCZCWIADKFQPg9IYdKhJfIZN+QYdjb3xRc8HQpb2mqlDGWz9HVRSR8H1T
RTf620cGL6SYfS85B8SB5xwXdf5kXzsUBmkpCakqgAahuSTwz0VdbHME+wKXzuvU
b251WYbaT4bO9Irowa+wCI3GKNAt6WLrMhvZUQNeVJ3ZJAWj5AwAzAGssh0wm7zA
GRMEPp+uh9z7VPB8s3vAxZ+DnxEruYwhtB9SM1Mb1f43xjtlSwsYFKI4nvqwSk5q
ujQ7V0Haj+TQjuNDspQ1UPY00CjK+jflaHIqnTam4+2b3bS3xesc8+OZIxYQoUhb
XkAPEWVILAtHJujVf9M4jhn2ekSTnrW5LFeFFJQcA3xjE/HHD0jijuMSpHl5a+ch
xmq190NczaldqwqhacHEo3Kx/XLwONQwmOzDhIohs1555xol9bqouX7b1ioHdd1K
0omRvaMzAipH6QbH6+8pJeR3XmauJarDQtpo5n5BRO4pqd00B8N00ss1we7n9W51
JhU4jwUHQltGIHzBl0jvwn9NF7VUzB1QtR44UR5ZruCYjxdr27ZVO9i+vD0sbwh6
ARDd8PbpXnLYRtwkw8P//jNaREhaoPVtjKWLo3zrxGY4eK4zTClMY8OUHnMyh/XY
EHr7HqSkUAI9DXD2YlPTwwmKIr3qafpnpNAFJ+QCSwkCrNuoBoLin8IreROnkCF5
d9WpZ+deK2VZhyQyobNcQnHRUS6ArlrHdhozP0VEgIfZcZfolZ+Tbew9qoBEHTRE
CWlFurqTji2JQNcCk0XRx+gGpOBlJ573M8y30PsI+xrRb/5PXMDpl6N0YMrTuvBg
wrBvRqGWOwCejAbpITr4ajbqnles7ZPU83vjNrS8mitazAAVO9htHmJRkfCwKE1X
AsI/F2yqV9KPK5KZK2P320CTyUgCeQNblt4QLfkQMii+IyIjJX/E6RtC7HZIgiMl
hAUa2e3su/DDX0RkWmV5kWHO5qZdRM0A92IZLkCUFBqKkDQsa+LPsZA+4m9SQl1Q
+MUXMV++EMBCPSSxxeSg8RH7AxXWX8nCeViPQlafen9mhS3zPy7HxUGAa/Hvj1C4
8JTypmotyeg5GcNE7xECn40QHKqjGFVpoTDFvmtJhVreoanALEenyKg6PBtzpmeL
U/3xSs1HRlHPiEb427d0zgx4pXHjSpZjir3trounMumnAeQqd4Unyxt7LxBZigG8
SRvw9dlFe/bI3PG6A4TSSWLc3kJidVnPlCN4oGAeg1BoJcDvUFfC8enP9OYDzZum
knt2jZhh/IRerG0dMe43ot43cfYqpI0o5T4iLnuLXb1dPRcVfW194vuQRnwz8H70
cc2p+EQD7MDjzi+7Ldgbj7zBEsuv/hoW3V5RxFR2U6hs15+vG7OKw1oCugzmC5Qz
4rJx/W0ZPv15aU0LkQK9CD2h9dg0FPbsCST5ThRAaMjY430ki/HyKpx7mr9mi1gd
Ulrr70+GDgx4WR4NR8b2TteYBGxiQbI5PvIeQoekv5t9jA0w7LNIko5GQ5DjOplK
QaKAvftEXL+mX8f/CqBU+8DvKUlb9YACEZ+AOv/3H2ay8K+Sp0eUZ0MWAyEMna6i
5gEYhhJ0iq0qVplpf+Frpd/bbVa82RWn/5ZnsEDLjL/DiZPZcoSw0YzjAh9Xzl6b
12K3idFpuiyaS1NUSA+EcUqdCHsBWjONOULBiK+qVg4Yf3EF4xfJttlaA7Gcnc+l
RbUtSJKTVmSuDrt5D4lkrxFb0JQJMbvILVtqu98Mdk8V9G78Umvppov2kUJYmxhK
k2tuL/C5mNL1soQiIA+3GWVNzgxZT+rGDmaObNQ4jNOjD6bI/qj//rTp+sUQw5H4
z3oT7/8U49DBP90r13zWXpFq7xxQiFYBwrk5Wqypk4fYyNAveqCGooEqgcDTXCNS
FLYZojnfdwSoymqy88wgbPFCT6e7PKLy8OmHrVI6tv1QpQke3tI4mgSr9W/W2mdq
FxHBzstd6i0il4X2wypxPLHyY3+xqd+tLOzXsSjbyHxWsB+4gFG1wFOF+ka5O3fv
dZt/h31tJQN0um76R9r+vYxVBNMHFD5PA0SSP6aP5RZ7cHo9y0LIs+/MLke+Enna
aK49Am8dfHpgf3TUlZG9XPIzHlp0sdyLi+e9GGbp1ALsr0S+RIMwXp7Fwww0EhaZ
fbuROdJTMk83XyCw6xVmyDFNUGjSafZprB/EY7aCdEAlpymEFK99LPpmPFmJxJEo
CyUaVwknEUTHG+YuXwoTFlUNZpgrcW33fSKe+1lm/maO/vRaYVuc2Dc68JWsFD6J
pAwkP03kfjjSXZZ53H6X0nzbG/PQCm01lOKODlSQP7Y36ZQbYkRvwyCAQfjgIgr/
+qxV5SXPxHakUTiFzZ1va7wGFlGlaKAbvSnslvRc/gvhx7oLl646xqioa3BqGMoK
g2res1BkeMx8srIEamNYUfdKT1/vqyDPvfRc1meDbTPNTjsqUYXBb872hWCLRFLS
9mmfrW9HRBjV195WvxHG9ZWlbiYY0Dd/MmhrdNT7S51SCfLC9pj22kkUEcXH8NC6
etcgqDb2EfWTSXpTBVDHlD4EZW6bL6bfIIAStVE29mzavFbtbPIgony0F259W4Zi
OVCbpjsuLkhECGNB1fgb7C7F02XHiAmrbAXbJpiDc8ZHfUmU3vv4AValgKfc1q+T
iZt25dZKNgSk81gAEzZLBSsjiFu+xJSXDJoVdgvMo140IoRBoSHGrc37/BUWt8Cn
2/O7JrV08qZwGZreouDmZz+Sw+VTPU4GW+iUwRCzZ4cCbOL+RrhkzMOy8QIf7pUy
taxBs+79iy/8xLFQm3g9yAQkjfOa2i3HZsAgMfjXhpV8iOdW/OwZR5zx1ozAHAUM
DrlAQzYtnO/DXMx4Mfg3J15jFgZ3J0g2Wgda1tJWHudc+RTDESCqNhcFv6CcQDmm
cJ7Pg4m8KJLIhGUAvTi49tTcy6wbxWlwRyE8mCapV3bxtjp7h659ELg3HmA5CZv2
Y4dvQXhyVKPQ+dPNgk1+oJF3m7a9fETINGQxm0rujpsmBOJBnH4DHK8AVckvo+jK
McYUJZJzcTRKgtAHJcwIN8tAufL/4ddadkFU+Io7lRzkEII8BRBij8ZC2yOjO/4Q
Voy/Ky3Bna49OgB1XVo16ggC4hoU1YE24LSoSNtAJQw0uzzpkrNZgAmufai2hfQr
D+u4UuTe/SHIR1LOR+VZQuIKGDulVe4KD2GKgCL0NJ2sMrIeOrKNZXxVSc5mCcSN
d9FonyVkwGwGfeLqreL0oYHKWWfDol3SzMqmb3zKND6IXnvfz1j5kkzkUp9lNix+
1Ie0PQljsF3KtZAi2loUiq0lFl3iHjAFxMTorJHC16Jxobz743qdxzNCqqwIRYeB
f36PdGA0knsqTdmSiAkFJUvQhPzkfMVbw/PkBMvOcTZV2yoHW3c6v3pVwmYcf+v6
XOsumvsZzhBg9IMpGrZYZPzKHSlAK6FeIGoinh13q8ig4JhIKY42mYRo7e2hXXsU
9eActyVHJ8bZJBn5YFPyMOgCgPAKQdrt0FwOCmXC9n1I7kreX7OCAjr6mqYlrQm/
VCzUbFxDqWwn6OTe1X1Tv2vJY1IUbkRdpaJrBVVFJLzurOEzmQ2OZQ0QgEtlzNZ6
mOMj6NhZjD7A3wBepB2IHXBPaT9/+72PdUGWR+kwlX6bXfymn30LNUkDkLmJ4Iaf
znzazFTTfmcWxDnY37z0WH4c43ewLiBzxFNCg9Ehz62qjt0yVTaM7YJ4B7F+v8Yi
mH1iP/pVx0tGRnfBaAaV2C0KKEYe/Dn+qqAsdyLF+qUFDzZur1qHF8OwALQlEalv
QxdDwWkKC48u3PbHcmKPZsi/Au2YTgRcQOyJw4SCDV53F28dUSbJ4JcJFOB5leq8
Sqx+Mah4ZItgUY4T9qC5EL5qq0LIv/6qN2Zub+tvVQXFRCULu8cmfgUthZxH754g
d7orJ29jkjxPSLGa1VJcVXESsGBBYXpX/HUhmm7R6vBz2xiXSEWZlG7nKXwR8jGM
QYwcpd3RZiyt52TJUJSIEfHz4PoV9SyU1v9j5+mAQbaEvTQzr6olyK29UG+g9fHr
RB6MlFN10PQbB4vTpp7nplSpGu0l3eT9zU9JWVl1H0a7GTjavieDPTwHtYaHC7/G
WEQNATminz/bx8JE6OCmvmPjB3hYPsWKhlc3w2apZQzLyBX1xT2Wf/XbMGjrhyDv
/LdToXoNf1XMHXozOX/lCD9zLPl9xqoF91pQwid4nSyIsdVm0wQKPR2ehPvSQESx
6uXmnetjr45CfeximeUMdLm9U4B+hCdQVqtj0yp2g12y/hJYe2JQuLOmu2SXM6IT
7dVie6Iwg8P4QvNCTH+QyCmjJwsJfEaDrHkEhLtgAXWAgqoY5f15c3Kaon9Xnifi
nWIktPA+5nh6HlfebBEQSd0LbrmyFIPLB3CDhEAFrjeIH8KivxHunqHL2WTCfbYe
SJNm/au6GInVWllx9bUGg80/Ky7pTKXLE88EmssUHM3rlgxiSy+ghzeeJxUgkWdQ
2u3HdwerhK48yNaqsoxr/H/xgkwlnfIkBlK2fLpfPS3PfcelT4Ei2jKp/xGik79K
CR9h+y8xoU/W5elSu7a+et0tWo495IDyoV7uPVH4kLoDEEkLMd+JyD8lRh6qa832
6vGk2bvohgbOveVpdU0gx+fC/k7UbMoOJH8iUP/UcPEw9AnfwHbF24KiWna7FoW+
2b0J5CyKrqSJ5IxfGRIf0g1tj3Bh9oDagRSEIxNvhhyw2l3lQohg2jS1+GgRGbgZ
8AyOurcYiu7B6u3xYI/S5cJzhYHF8qnNAnYJUC+MdaudCTkcHVAO3bSiit/FXomW
FI3J2VBeGXTG65QqBz3pR2IiUG0SRktfrXkhk67XGol6+AcBBRSdKRuGZ2kHaRUE
mFspPTOFejNvRwpqJpHOXVDyQUZLZYmlh7hM+C+D976qOwVcvPoVI9v4VT+14Pt+
t8xbmuRf7ayTjndR84AzYHQIriANjeAl2R9XGrZ6CUHxt25EZ/icgkykcMcS9uRD
wEwXQI/04ee0A2ZRSN7e/o8B7IqppDTd+OpAFV5ByESCR/lwMa4TCkZosPaWldOW
/oVjo4ZlkIqyJWrhaQhvN1j0uoTdfIICuuoQPngkWeSu87XQrFUTuR47xAsvJsjF
3vzMFC6cuqXV6Nmc2LEmiAx36TxuTWBIanhd85a+lA9y/MYC7+yTmWZPRlIpE5mb
PmiX6bBbaFvOgJf9JYCFQ9Y9K7QNMZDNTqSIodq6vhYuUc4Fro7YSoFPJulM7nsu
+6L3j+5eupJMFA5m4jyHgSnhlHlKdNJGx4b+RqXN7RQc/fSrmD36RiC5cHSnnjYz
Ye7N5L3qzRyS1I0jsZhiXSAqT2njRWwdZ6lnN8ly12oMdRt1tG7gEAWpT7rBDk/E
KpuAUtACoMePH5mN4tsDJv4HRq6CWZuZzlBWIIC6rRexirS6CiCbgt35Aa69Rzqr
JKzrFoJyKZQFwjdegETfL2srqR2l7wNi1zQHqO0XoJsLkLmQ2XAmgaEi0xVBGWsV
k4R9zr0/j01YqInGULHPwADjPLvMFDZWutpyvHxCSXYRzejSwTqMvcNBEHtup18e
7o9q7nfu3PDFbESYy90h4pEnXCF3YvFce7ODx312V4EeVjcD6HgM93vCdH2+YzHY
TMR9ziVthdxwSXQSejLDeZXeevt3dzKnMmJC7LL0D2spn0MGxXtHVuQELYG4sZc8
hJanj/jAtpdX7SeU69RFvPTG+mfTE+TsU67MKoezRB12DV8xyqjTgqZmm6apXbtx
wQTuS+3rFS1r+Acx34vNPKQ9/Q3ZQUcuxK6kv0yW22OUJ5WahliQmzwYRWmqPq/o
qQsr0D3/eYCdDYHzcTqUJZi+mzPnIx4MwUI32LnJ3UbIozOr/PJ8TV0qkEfLHe5w
SNWAkVmGeeoUHGovVzZuYNTisD5sUSZpPse9HFxpRFLLsFXxtfCsSgQLen3PjNmp
b1qtv4fYjkC5pOZD+LOlVAVzB5G7UsC+y40y3ttmkENdhX5be3IJn7spjbMv062w
T5GERbPgErL/07oIHqJ4C/QYq1qn/s+1/HrxlAdKPvz51y72OcF8eF/XMQUpspBe
+4NAEsuUHFdNRKh0tcX4Nps+oXJGB+DTxOGuvl5dDI5sDFNxQqg2SPWq2jS41qsl
paimeB3XF4S4pUzH/7AqJn7ry9XttaBxs0hAG5WbyGwW+vDC5wKCgZaRVjn5Sdvx
ns82SkKN+mUG3BQywXuLDm0/BDe+2ynYuBkMrGjbePdam5q97AtxGTNw3Y7e6dHi
9QHBcM7JRK5TjYFn8DUmi0IwMpIoR3PTO6KEHXgemedIJM+Sm8mJ+kVDbBPjb9ak
GDQmRCUalh6VShJtRztRrogDETAiF1UB7Gs2U6SxgMh7Pc2B0UezLUJmqNJAlWeG
MC4oe6bQMdqrtyM1O2kWcKFyuBLkcyv+ttPMLw/WgmhKdMncXLgckagvJPPO0do9
cHqTKFcCB6MsvCn7gx1caGdrbMSVY3PyYV2UmFnipIw6KTKkJGZQUeRRCD2EXo57
j/nQGN38z2chKq6Nf843d3mZmI4yujSxXVZp+U3lfzLeNmQEBVwojaq2FCSfkEAG
BkWZbyl+9EDsf/dFPBu506ny7yZAMrJhdVBHF5v2pQ3nxoX40lKjXVhYyLJxg+Mh
Ct6A1xuRp++AmFWeWe738pZOrdgu+PTwCvL7uzJcBZ4Mct9TcW2spNCBwAW8lyw9
YBsDbo/RUjVacjeMOx/umfGPfKfGIJElF+DUO1dgc18NR9h/g3OJVm4UDlT3z5A0
Dz0GDLW1TiC+Kjj00QvZJQillp8Gjd2MjBZQpEo1B2xVM809Qi/ILUlYUY5G5IR7
ky7n8fZAVfPo1gzihWs+hUByN+gLF0rJLXou+n7THh0625210lJvGUQqOFHlG3vp
T3HCL9XdTtnczf+eu460fV904JoGji2Ei6XQmghQeANgTihkH/AUHQ2SBVNjtWcp
T6qJ6QdHKkNwB1Vb06sxRcS/jc6e71r3irKQaRgylrUUHUhTQ7u0K9YEg8zj9X36
TiKCKXGmdEpZNp6bzmo67aNhFC8RS4pJv8ijSYc1yHpuT4EwVB1emA75Sr9aFnE4
GDXcHqP9PSEXCcLSJraj9feWLsvIgOv3WXEZ3QA6WryO0S8YTsooq2UexkiCMMEe
/Fm252bVYucuayRlabUOpt0GEIN+sOOFp+tQDsRjQl7W6L/4WG863M47wog4HT95
6vvLWLp3NlpJ3Fcn7wxfA83g2KJra77McMiNrsDCjLGWyix+NvK2277DAyyDhtlc
ef52ivMZGLVUy1fFD/mtgv7+tlzJ7izYbmURy0XcfqmE+4096E7WvG/1vPdi+gCG
Ff2Q3DPkGCT6F6hvZc5I79M9h1IwcBRL5+jgr72bpeFcYSb21s8sCtwr1YGe5YPm
8NI8Uw+0qqIVG0Wjjji3PwatbH+eUropdypj74sTPFiLkR8gfIvJjEQDSf2XyZYr
iU/g4NDg1esEJurW/g52+1fh1vNjpRPheDUjp3aoXq3S0L83rAc1Ev9A/L2ZK/N7
5gf8k5l0oi27Ii36T2gnjMxbZZfojuXomnfW3tf3TPWm9D9UcXaGKxlwrppmlfYJ
yBKVTb8XdRx9zOKnrMygvS/CYiWjdjJSm7C2tZgOjd3RCt79wwP4ngzg34SKvCYr
/IUrJ7TRcmCqHsvlfY8WK5Dl5voOSQjWlrH2g9vxNQTsdAXT9pH2flSJSugvfjK0
RS01N9j0w8flHSHYNNoP2hjmjspB66tNZWvWQftJX7FYBz2eCECI5Vn6vR91BD9m
4aArdZTC1742UfcdXLM98accA8RQAHTDjPYC5t5/95gbSzVvx5rrsRjFLmuw67CX
7g0hpdp/HhLKQPY/+scCphgoyykpabrS0FVYlUAr0JvG1Bzq7MctE75n+eo/eg/7
rmPsjjQ6ribLptXnqzT6uhlVOykqBgLlWvmiNqswUEMDamNgnZgEZgvZmr/SED2+
St7wLHxnJZiTQic5j0J1bxyn3w4kF4KiPIf67pZMIIcKmhWNz89JoOnnjWZhR8xy
k70LdZ+JzmERR6GawajgbkHCZaeRjLL9CbTXFq+mteKOLw++o2l+p+ho9/ZlksQx
18dKrBQuWXHptdp/2InhKbboanCnL8kOiVYnWrwJR6+5+I/9wwTASHS6lpa7eLFz
S672SEzZSbRXpJMmEymEAQB9mptnM/MnSLEIelklG3AbFdS5UDv+CqXrxGahGZa+
SuXshmaQxsPcbYubBXHh3mXKOHUFY4D3Y89U5l/matpe93lEvizpENLXDFmyMut/
s+ImO+OSONMFdD0KeBqRNUUDLtYNOgUzUIx1Cg/ULomwR3hpwIGPfvQ0wpBgCTq4
dyG4JmGzLWM01VVNUWna6GzUq4ysXTQL86aqUsckkfIEJx1vt42bT4l0F6OVRvHz
l3SsMAFapCnrNR+TMuqHwbcJm2wbJH2JgVyk2ryVcogJ2lE+cFVOpaaBJ6ZRHJzn
ECNqWEWKD1Fe0WX5IB/qRTH6cKHx5K5NV/rAkR9CPJ1WY/shUMderkmg5xnrYGJV
VX7JzLyDLdTSIin7SEd/u5JuWJJJ9CYiqvuByRD67vUcnNbLnsYtTGC/N6n6GJq7
x07UstM1PyIgpUMZKfe6il7A0p8rkk0NhhIdBPH0PJEBSjkte49DB0zu3ngg6glB
d8z7Pdm2wf7fV1FPie9AetV7a4opru3p8AmSGLSPY3/ZTkHOZsMTfy9Ny/uXHEzn
dOlUH/AwHThmjg/d4isChjD+SeOitI+rt5SVjURXv+NC+hrWnsh8frbiO9dnYzEv
7xELKAWf1aQOa2x0aZ1nxNQHwK8V6sGMQkHTKRWrWDa7Gy4yJP2HsUOOyJ2fR4/O
OShH8flDu2hijValDkMVN30TzEGf8dy2f/17fmu6wMKBPzvLyx9mA+++L8xU33kp
/Dw38VxE9UqX3c3T0DuvE12XL9zIRq7M9yT5dBo0iimeSnC+MBcmKBQIEg+VXgoT
tUA/WDIus8XZ/ijhV35kfb6g5XCPQoWoBwzbS/wLgv46rZm72J5F661BTbRtxfTM
6cFqB+/SglxLVO+AkAPG0DMEJ609em+cTLQ3f24fsE4EJARSRbANuXSKMtzSqbhZ
rEZp7XOQkcqC+eet98sXoObVpWGyLcJ3INuExZHF/P1gclYN4y2afueCxfwI0KzT
FQUHKvZjI2v5/7qSy/l/ZNsftUzYrUVEHwD6s4qapNnNWx1i015aUAPN89A70bQj
xB8lt3+219urnyuDngGWPjq5UdIGy8f+FtNeJ3pTcRRjYP/y4YsaBnxzMyi++rRr
uuQhlKwmiaJ1CYofRA8rXOHAz/XX1CSgqLBnieCX1HAXAH5ulmH+BbMFjyMnpZRr
3QQSNDeTz/YZE1yq8HxCwFpGBXz/tx0nJAg5rSby/Khz062qsuOhIurxziPc9EbA
qz0FMIQqxbvdiSLHHzw50tftzdFmob6PTj420aYJNeJG/sLP71Evqxr6ZPvuYal+
aqzQz7vjEPp8jzArE2CXkoep0PsSJOrD4YaO2JtVNC5UjeO6mxSMLW6aPKQxmAWb
14VLzXcQqO9ynDFPN1w4arAk3GBwUvB09x1siOZFm4Qj4e2xF6vLMVdxB9pkCxE4
XrVYYBp12QsQ0BhtZyjfNE+k0svsZFvarEkAraeFjcf8zWWHQQVwXRDx3ZNICSHV
5tZkWbJIY71sYJAdIYcfsVecddwEFwMrfVNj8hc831pf1Seqiw6GvjaMJ5kowTZl
I3Nd2s4vKGt9maLb5g+3U0cuzQ8MOwYPqU67zWLwQieIuu8n13jldIe1FRP0j6MX
duwMnkLB7AYuNqPjdQPZcByw+YwBWD8rP2jJgbpAjYenMcWW1P22MuYjY6+rJhaF
nfg1wsCXq98Lm+4dmgylhKdxJOA+r33HAEzNp+YYfOODdrJjJyG6D6JBBQ1DmQEa
f4mVS64eMS7+PunCiRLFwh/PcXmAg+UNP5YuFZnGn/SaJi5/0WZIBhlUdN3fg3rh
ybq0mJnLTQ/2PYs+I1bTmht/+VY5vXdoO68DQSFXuugmDxGY5D5YSUf3OcI0CY5c
fM059+dLJoH8dAhAMrITb6zNJKYwgvGCDGUJYC3fvjmKK0H0tC77fkuTinEkMxYE
oYKRaSThcSTN4Gg4my/QbEnQsgeQsWJ/beQTPi1S0oz9ZBrW5UVqcITCv5bBT1F4
X+PCvjqrj4dInj43SCmZs8SCOQrD2WP2Ag+4fNaSeFvbP7p198XC2d6A6WpzxaIn
+4h5nC95hC6yC8s1VptTdc5d/aqK89K+uk5ka+pO7X3NzL6kf6XJF+kyCqRzCWvE
z2mKgNrWwR+0DtMIBQ+bMnTac8RB8PfWyPz9tM9PA88ZXJY86G3y3RAVpsypIhcC
LxHOEogYmxlNFOQQUpH7QGGBFRiZ/qosQUgWW5J/3VOLgA6rneqfJ1tapLtUc9ui
Lf8g5Fqksc+5adqBLf4vX9ij/qa9tladYmBIyQKfSDd+pGhtCX2fi2MrT6j5k2aP
c0agtRwg9B/VIPulIzir2XH32dIP+Kia7zZOeuK5Cngx6mBEgbyzfLStevDZqs9y
i4TY1j6q7jegbZmwueVVl/bNvjXW3vrHmLLH/9rrJEPT7v67UOQHdvbvdv2DJvVA
z17xqolLBl0OFhFeH4SSd6gDl+9pBbhKLxkodBvsu2iTxNDWVeRimulSBulHk3az
tquG7W7vEKe9b2VSB6ceZIuCvvCdShnvjbAyNurrTHPL2fYeyA+/2+WAHnYsvDPD
RrGYpIPEONLRdYamOZyYmwBfdXHcYt5iC4nnIjNbhWYiJSRn6YIvPXZfxsnrmzc0
bNwH29M+z2kKrvz9LXaiR3TSy2XTAarA3ZnuaL49Q3aEp7H8MJ4ZeA+OjxSIpHT5
/1X8eSi0iAUzRXY3QoXvJM/ka6ZG6jP1xNmLPd0nnLxpqC5t4NkAHOXVxh2YZUgk
/SClwIRAgT9V0AtPlYwMWt3TJe17TjqmouTM139wUr9orE+npfBXgsImJOeM4614
v/Ptf5ucaK4GXKu2ofH5hD97WRcurig6jh/uBc+0B5HWqX1uNnxuI0ZcHgw9Ik19
BunOnGe7a0EmClN7EIgqgce9qgX67xEYLviWpz3INs9S2DwpgjiKzxCxvzTB2kGe
DN5i9GmqdSXmy86SYtQwNjPLUyFTNyrkOQX/f5Wt6c2UqaVR/ufWwz6I6oUnp2OX
qu6DAWDU4GdA1hN4FlXO1lq4pOqMXT7OOQQpYz64q8b5A4Xv6aWZD0/MMrTiY6nN
l607NC4lKw15+8Rg+xE7CowWGzuTqEuk/lkoJBtrNKu6C7qH4DC+Vq/yAXmsIB7r
p798TahKSGd65W5nj+0SSLPPebQbJzN0GfYlTidKtgM9p33DPd5yVNwIn/Ru3+M/
QjhLu5w0m9jA7p84cH+jySnRzW4QqGxKjc0h/xdWr4oaJziLfyq+kLQwsU1gOPkO
rn7vEMdxh7XkWGaoyNVhf+xusemK/dKtjzzTecP13RZQD95tPoKDJwazlJeJdHRq
vYEh2PwxRQXZsA7Lp4tHYiPZXPkVxMkJgAHqt4Ru+/zfBE6oaYAuuOfCQ0VQ6vkt
me1cEqpW79ohI5wzY/NQmS/Bq6x0RJ4muEMuhXrMRO1qupAIiVlDGaJzMhEsNrSJ
hfaAOXAzYhZpMeRDuitYwXue6YX2Hi77frfJb4gErP2Zs1692Y6ktoLPdg4BUISd
S0PYwkH0oUp2f6rmtWwpqnat4zDN8Wk8wfzaq4y+LLBmQNzSu047Zd8zJsamq7mb
cMfgJYU8Yv30yzKkmEHvuiwjZYzCD59O1RU4hadIMYTcQKUo0tOTVQbO7gK9nd12
a7BXe2Gh7BMx6p9/UwwPYAa4ElNV9AJZrk7m1AGLIcx650VPdghTb8a20ZR/5D60
gjHRf9LhA7HbupB25wX3Fh1HUZYFSpLD5VpefeK1EbjFAMQ/s42xQRd0qXHgJGy2
RZosIpQNp9Dyr18oZJ9oQPgb+gXWzcYyouUEJ6gKbTIYDT9o0D9spU2YcdpdxFNO
YY7yYWpfhW6swCJtH7qM5Ai32BNz9dIbjc3egS0p2kJJuWVLiuP9vgeXzKT/tZ+N
B3fmUpDblv2XPPQ0tHk74+KYodTEEVSXOTbNoJ7Lc7jSUMtN+ICwkBTd0jikIHZZ
7bW3KQjss/pYJp/b/E4JYvloz8vskoyTtMTDdMSlNmwBX5alKZnMsI6eVSrw+KvK
OvXK1Z1182fIffeQUM4lklGp1iQlZoCz2+t0M3vI63w9lYTfhafwW1IdcibHL1z2
mqMlNFMue9qRul/nrmafvvtnSwOv+EwVYBLMMBWkzLHhdHgkYiW7UUG1ooFVZkJM
5jvKa0k4kMDpm8WpMwUjCHmXUWmBau7voL2G3QyhO1QE0X9Qht9dhU7lMbJrjvHf
EaQorTGigOOwyEuq2phrFqzjuD23TBpMuxQ5E3o0ht38IPzYW/F3m5iQ6YMUYFbm
sodvbvVU3Tk2TsmzhSRIHa8QlHZJ91kM4Ig4pU9hZR7HPPkiJk/uTEFKO1jMN931
4FS9McbcdnoprNSz5otSzodWCFckudOcxDJy5Ej3rVvnARs7UmCxM5S+Asyu34LC
uX4C+/DdLmTrMFM8bHU42NCGLnrfdKsw8GLDJnF1UNryAsJCjb6pGgPBVyiXnMB5
SoqrJlu8hBB671gfHTy7pTYWZIBsA5lF0J+2R3Ntahmjt2JM6lSblmCeLyNGbEnF
ml3rgtgkPNsu4S69VlmGPa4aiP1/xFU8GNphcLBmM4/cBrtDxEgan2lB10cb4H2Y
57gMWAicqPZUvOmFeLKgDXUik4AD4COufLorpGmObjbrVfafkcaFGuKybaVSuFFU
NaJyUsj+bKp66t7OcHTJSkdedID/ktuwkFgWNe9JedrKSXZb6QRK/I6dJ91RWATu
/14HRWEGs+sL6e4ggWl4iJKSxfE9ZFjYbl38CFkkWyiSB5xZvmQEfGHgBT/Oj7rF
KHWfYq7l7wcxhrZF7VFme43taxR31FyU6MMRLsmMIj4k24PTRC3/fwVL3HEmKJdF
QlcB7BDdqdhv3u8EDSTn3ahv5Df8EFv7p8eNOpIEhsbJHyqXCQP9rXPeCtuQY1B3
8+UtoPTfw6i0WKU82MfoTtZDhk9hLNGnJigHqNwh2gCGB3xSNDwuI70DGjcjS/we
Zn+eBfJ1N6xOyY8DiH+jg6LsWVyYd7AkNsR6aPEDN/F7wuFcxhq9FRsa8vKMo0L7
9eGHNFmZOgbdmjbw+nlYbeXLx0855Y6YtB+Q3+2lRuE+aPi30kbRMokTH58SxGwN
okIds36f2ChKnqdMS4SYWCSyai2H0rocTGxzR41VVkLA8rk4zMitegARBeHSMitu
OkC1PP0MD7FKTM792uYpzO20uqCSdFQdM5hUrdiBBl0o5sXNsl0XT0ntrAfX9KOe
UlEMqF0egG6SJsYbtjCjW3ugPOqcOCwPjyJYP//kzBWxugG26PxBUzxRMir9VaR9
Jc2zQKOlQZxN5/JZuybuCdsT78ZmzTrYrLmUnqBxhdWmkKRHSvw65RAmlTik8qsB
4CfdKR8gl1W8GpYnAJAEzIZ5SORtGgMSJNr9tN+GOkUfdCb3fy4hEE7t9QlXDIQw
CRLxyADeKuKmzLD7arPgMDlua9zKsO5XKuxD1ug+DjJRM5AMVKDULp8cDxjCwCG5
y89TwhMAE4E8WH6vAdzJ5BMmAdEjQggIOHWOvhhf7N6WZYtOIsCm6IFZ9faFxb+1
SGIVsPlDcEVtsYJudQm3xzWf4/noslcOaYB8S6tc0Z2nQvwGAi+P+f4yFtnnlzeI
gUj9c9rQObEK4dDOJ40oYxN8WudRNKsIXuMDMGyFNqpLqkii1mD5WkzSzbbLY23P
4jMy0mOjMzwbuB4kzVsmlX/1DdxSLL+gn8GYxhBSQax6LCHGahSuSeDiTkL8EZjR
Ae0ggcoQmkOPXnhb3fRUOpHCIBi0Ts6hpD++jQedvoiZVuqT4DoXNiR+IPXPOvDe
2yDQ4X3+V62owr/mcSTWabYCwfZ4TSvHQkEoUin8z2qjNbxZxUTYyy/a0Yd29ULh
0KIGNZsvWFsPekxJhUBUPhEb1tTBE5Ihu/9c8sUvICBnpzgQA0lUmfyy5cY9+HAc
itPUTLZtATWLtXw2DXdNsMnZwKEjYj1cIa2ZrKVAB36LzyAwdUcMD925ooaH89wJ
jjbZKhGonTyX56PP3QFX31rWX9geO4aJv5/Ar2i45ePt8ZLW+1DkUMhu+wr3ymyV
i3L657eE9qfa8WAz76u+UShNQkZa0hItLKhtCJNNFLJtH0skNfNNg8JC8QVtpzpu
flnzMr7d9VvDmrcRquuhVEij05wVffKSNvKY2ufnFeVFQYEeFn6Nj/chK0ZbAJfy
NmbkJXUf6lcq9a+9D7nVQIbLwv2THTo6brGrAhSz1DZ3ymyfw0Z6KsFTLIA51aLV
kymP/SEWJCFGyiyVZqftZ1ghoVYJlUAUbaZtnEs1yCJemGYcQWL7pmvaaIWFk2lO
/yL0LcE1Eewu8LO1Q+9B+gz7Iwj3wY9sd88Bj3RswhogUYGlUeXiTVDbo0IRxoNZ
HI/Q01WuHdbaILKb3DbTpyJEL7/Q76Xb59D6qfVawEEBPqBRosEINwq+jve/VQFC
1f5W4i1UJK8u1TWANRhcfhGNsDMVbLcrzaWDXg+0/Ep/AwANoTX59+YNLlhwCO2v
7bS8IDBsGw/XMa/fgpYmIk9QDZn6jNkOrjg6R38KVd4GuwJC/4TD7mm4K4EO2+Yu
rV3ZqPtGD+nzHprkrhu82ibC1ixudRwO6uWUU0h0Z5w6cF2lFLMm7+GvyJzuD4Qe
J9Ph2JOxO7YLSRrTgS7FpEkZApdw1mSYfX37OPepSWi8zX1wEPug2moahLULvanL
DY98B6o/xkJhCTjZrmV0B6CgIntEFghieOD1NDSCpPYvRFvEKN8SogKe4P36j3Sw
lxF7cK7uFyahXGZ0hNch0UUHKltLinvezI7zP2YAu6vo2hxVHcie8+a3etBsZ0Tl
0yg8QcZikUmXCKe28OUvXtNVJAfpUTaB8Y+JV3ysS0M6N7lIwcWtteMtLuoqS2Mm
IVCKBkKvtRnialArxzF0H5mSuTp5eEgs/6fdl0sua4caeZ31Je54sMcVIXoZtumM
uOG7a4YZ9EEXlorrGp3yExIVfAPh+D+mdjg6Odx/amFRtOvg0jMSYeAmrmxjdeG3
I5EHTSn91xBeBVjGiK1G7BfDbFGdIIpt/LSqPHN7oup165tNBmkyV8AoY7hRaPsl
hUwndJyGcAxAOPG8c3mYCTZWUm8FbtIXg4QZKRzkKVrvzMshby79ZaeJWF1Kwy7+
GVuOm1mcn+Y/p4hqmrgZ/Z4lOSOE5f1P4VDnk0sRxEj2osfVpF+T4S+ARlLA+n+L
AWQZ9njevfwwqW5JB4jUINN95X9IP+Q5AOLXIxUtzTs1FAGeZ9Qnail+/vLOA6hz
uknhVHmVwa7UZFZKYK8rPDRYb98mgk86XveTr788YC/wOrzjKdGNiTrgFyP8Ea5v
j2mzIaukwK/gROjjhUj8uKOX+pPk53BY2Mn3kk6dVqf6dReGTEfom9t+AHcZi/zX
E4vpm+V0cX58viQ8a4Ydfy9xixVv8xnS9f25B+1Tg+0a72f411w29wB0x7xvqWgi
R0JyCzg+2i9wn/MaFyh7LRgrSQfgiV5s8sGlFo4ocR6jb4nUQldKXIR7+TLsWGkB
PRe3DDzt6CVbJqn9oxTSSOhAliOBsDgTQWd/TiPXTAJgS2gE8EO3vDrwEwS0R0Qo
PNIbJ/lNseBk+VN7U3TCQbjJI6eRIcH7E5CeKKZaxDtjmOLuzxh2+9R8dpqt5W7q
yxt3h7d+i5YSnTAy9Pm7Oe9ksqJ/plyu+/Jwy7xczgKWHS9brlx/N7ErTS7b24mJ
h4TWXfA6lMbC1PTzfglZV7shdQoQIdlAMdir7oK3EO1VvgvP0wzfwiydqaIkQImi
Jkig+mjxRK8UjvcnfNpG81A6gnOtHkGHc0dK3bQTQ8m2uycP+fYfBbG3JeC0/J6c
bfEINLfDhbnv9zsvyw+AxCiqmbn3PbA2p2GQb33P8ERNHOH8/koD9U1Pr//qinC+
mhiG9V4izK8Z+SK1+lyDjO0O6l149kWc56axCssQs4g1Le5+qcx77RYhK82UDGOZ
YBcwopCHQQ0tU5YxNLptWEvd1rVsmAEbmr8arlboEynIFImdZokFdMlQ1D0iiMm/
yOuVFFuc8gwEMQrfgxRgg5UZLiedcebLiKW5O5ANrpy1ODEfsFc37ZORTzPvwEie
PhmR0Rn3RAujR6vb5rWiHIKRcTwmI+rMDfIVNPlX/PLgh1vWq3r/HOLi/FSmZ408
jsIjtpo+gGHNwJ2+we3Xof1uU+bUHz2eQ7K7TZA94AjFEcP0vamDHwYr0IDzaT7t
WnaDwRhTF2aN1wcb6G0ZKs5h3k/maOHcnZCJKALtkr7IQR5xsk6nkuQ0XxkfGAqT
yaD1+6WVm+MlzUhNcIioMYF96iNwkoXMw8UO78WrZSEo/WygOe59r0Y/iBj54Z30
awasYuyPehkA2nK5/IFJo3Mqeg5GXTS4vE3+QCxvDjt+wG9Uhb/tzzTx5SwRtZ5T
sI4qQKZjp/eFFrH/Pta2GLqGSXaEpkzW4+mUdmbBKCE/WeDYtek4AtGCQdQ7YPFf
RsD/sjfu+OFDDfCEy+wbl1IPj2vGoTxasMqH3aJPqrkAURhcnaYik8azlmFQAiVC
Y7O4rIaBYK0IEECCBF15W0gLvjWhg4xodxDr5P+pC7KVfYzv+/VHsFL+Z+b7kIHK
V9BMt0Nu29sncOsCUovrzvlU86b+xOjdIEn8nsreAjH1qJHiBKlo4RPOzyNoEo8W
OCIMQAW69ffJHAz6Z1JCYv/ebFQ5hwRlK/KJIYkWcSSR2MWwju2NG4CzPUvbXVUM
+UIzRcZKhsLQFPLSQhBAxOghylToKC2LKMJRxEOHZGZUBL98IOf9MIbbNcVbQWv5
fZkCI4o+5MtubMgkVG0RCyljeQo/AsXUZpTir7bDNcBBBGON11If3RSomya8sben
niQeI6BL5GgtCJ2XtT3KOEa+gnz5LYH22bBL85wzUvArPIGvuXKjqlzKdRjOV7vX
S7eatY/ZYQOFLbj9ZT0OJNdchKBp+RvnISVvU45ld0cLnnCP7H3DaG+UBct5I2Ap
7D63wOTtLDorX0LmrSk4G+eV5Vc36f6vkkqAMskN9FVV8t+JQQDmePPwj1B/zLii
sZ+O6C6qNPRBciyovdGiN0MiYtnRuPYyLXMF/JtE223dZLiKmAsehm2eC+u0x+1p
3+2v4kbLWUxwpNF+Wem2+f+a4tmHZkX4IeLGXdjeap8fxis33kbWiay7OYyfxnIx
ZOs0UAVqMcVatdCdxziUJ5iyDlqhE3/dt40Njnm0zRyAF9BKrIx1YAKDP6H84SOj
daRLyM8qK4MESQeribp31k98jcerVO81owrNKQ2lDQ8Nh03rmBfFh+FjrNRcqxmU
wKKAirSOQe22bBjKrz/uNRciI0vZaKPy68f0zfspE/5cspHj/dBsAcn8pL8Ou2J0
A0rWK1V5CYpo95YVIesaBHhDFl0UjaTTKpMLUXnrmPS4vjGnuqJ/BdxqetPP+kEG
cLy7i2M1vNJppHRR2UpRtIIfLhO+/hMnfIK9xgFXLwL88rPz81O7LfTT8nhz8Fkm
HPFWst2ZqE6dMH/uUN6K/B7+148ogzCDStChf3XzBVnYb9wOkKT4JSNW3Dnb0riG
oF4bpy/bMRqJY8emChCRIwkovG2BODZ8UCPFMfpYLNxq7Tmdqf7VYAkTZKQvt6R3
okm45MeA3ropr/vV6ZNOBKIOVdKzPrPKhcPoO4GiyhSktVDjK5fYXJ82r6B5Ayz/
mG+DYK8Qa5bkD+QVYJW1rGrBlWxXpOanEVUJFlcHYW69+UDHbbgP7Qu39UgLeITK
Pggfob4Yc00uCKU9K1XLm55IUzn+3vM9aHInweGTzCNxwWbIPa4w56hSvt3HsEPx
CG4ZNjyrxNzRj1bqecNGaCTSvozuHuj0+/mIVRt2/EQsbles6b0dj97EkEzhqeex
xoXPK/2O51Ob3BHJ0tQECQwUWbcGIx1bQoG0hxgct/PDhWZKBc0T6ur3gfhvLOvF
sGJxPna0PtZikWexTlcO53hGSk/ORjYkGdnqPDabsuRPSZACIa18IUlXIAvznVPQ
oclkn9lVDZveFaJu5df4txUBArFV2d/a70EO+iTTPJkULISves/MN70M7GkE+uiK
epW1wsWA+G/LCUlaFUduhkFgDLoUBh4NaSbn67aeVm7GDsdgByu255L5VppSiU1L
3b8IykPDyKJ1yJkyINmZ0U/h5kR9QCB/0M1Y+3NfA8iyZqFOKgwMTft1Af/5pJAm
wzCSwBkOal86IpCAaKWWA6ppE3yxVmEXIc7C69BHee0zgUBo31XWC3P5CS7B5PAK
laTxiFDQxN7uhcgxlu1eJ8LGcYVPh3PBFlp4N8pSri8nz18dhPQTRmC59PiraNIc
XZhJT7AEXueZ8ZFfL9xrV1+I56Qtciszmc1liuLfuBdkCyIpyo8NXjU7K7M/NMjC
lX68tLQ25XYm1mJVSlOxtfYz+peQ5R00NpFDejNRviIIm5BUhG6/trnDrmOC6AEf
TTcZzLjQIrmKRGmLtT2tcwA8pyeUl/239gQNDZX/lh1bEB6XblNo/xRWlweYqOaW
3yZ3acKSqbRYijLWXGkR8b3ixKzF+limLA4clKFmIHpMLuOrdYZWavrtT6K5d3Yp
V5Bh18wXT6++09YOzNMSYFpAbn3l9cv4bgyKc3l8AnoYNvVuLEXNDjt4HmjcRY5+
AgIK6hpM/lBrugBOTwMWhIV3feZN/JNRgg7O43Af26kPfkuPAchIL5j4zxhKM8JI
u8ZfzDOsP+ZrxLR39DU5QTW84jpolQyq4OMMuYYJ87cAjx3iosisY+8e+NbGuKZa
4ZhFpyAMSDa4fN+ui8HjGjNLbs2g8CBg+w54EB5fU5qZgWkBreRf9zrzFzrNwRp0
WE2cZmuJu2HuenSryWH9bhaUpR4Bs5LayIbq18Mm4dFy7aIw0zkM5ohuam/15RLK
9V6dONXX+KjahI3EWvQFB6l42tIObdcPofluyfXpH/Hc0mDgnHhcMvr0uoJEcbQ7
XW4o4UlKkNUc+q1AOUXWpl6HZCcgyoWEJoAhomdJ3Nfn+l1jELLqqd6LhuWP3fV/
hPZrQnzjVYWstOYHdrQzm0CE+qHlf0ZzEZa5WMKpclniWt5cjFjh6sYdHrVcsWnf
dW5+RyKtBssux9gxHcax/OIXEPe6qEFPjxYrB49c0ceepOKxNSJn9eMv2NO31gHu
b+W0aPusW0qHNeKjxwTNKVScjL//AJczMJSWj/ZZ3jS81fr5nHimt6xheSnTSKZU
dAw8imCqGRyKkTRfLdCLcAre2Ltoogu8IqIyWkFnBYMUMJGRq9TPaNTeoT3B7M7a
h5mE8XtJHOG9EKKmieSekfDBA0Dqh5/V1IoyURySn0OVFAIoeo+awIEeXGc3pSrM
WP1eBvWRc+OPCKcrPx30lbQwzmcOIXZ4AkiYvN1uHUVgrcqo69J5nd2Q58CyBTjV
vCAb1M2pIstjX3oRUKIkTZWS8QE1SgJvYnHnx8NTFjQQlkIQ4Uj437uUGvl5uhgN
cj4niJta2hgAKPuCDt+oDsHvLqlGIDW96iwJ/b1ahM4l6JlopC3cwERKQ18+/biC
tgCvcTehWHzSUEA/vwvDJ9RGYpqAfPGqkeF0EtxbRxQ6YNUMhlysOZj/0xBDlBXe
9plfdixT+IXmb7F+Ox5fHVdRIDdm9dZJBE4C/K61qZ6x73J33sECtwU8RjwSW0XA
C8Zz7qeV78jLLs2kgKV66ffBE+YRNEIdO2+FsEaH6NOvkPPEiqofkygVk++bRe5X
fZBEB2XhT0l8u0FDcNDqulGFTBpZRhSOlxxO3OOdwsmEECc2ef2wgaxDWV0shKXa
9vp+8wuDdqVmGfuGqcbiwNMgnACzeBOKvY7h571Td8JGghxi5ImdzdK3rwLrDss0
iSHINc0ktkbyjOYzib2CXiNiN/JaOMZYKHjBrQ39hJZpMQmbdHQ2oROsHaNzb13P
kpaSmw8p4lX1klNAwWUtUgYpVNIhWDXOQarh7CaKQ9C2hkbh6m/V9ff8HlDUQuua
TBEP76LfUI9hqzph5GUb+2nV7KqjrDNmkIxwe+HmJ8qlFyxmxMbDLS3F00BLcG7T
KlQ8xorUFm3+zx3Y+KGL5qbHYmPcW7cpkhKTS8r1MEGE069VCr3vB9+zQq5ygwfV
aNT+dEA34DWch45pfGntkrRXk0G8vjYdFj6kkrvrDbi3qfJuj7psfpASfzPbRxPl
5p1qijdcUm8ocvcK4jxab2y2W+DeAKj9kFVR0/j/BNHuYpxBWTBFtqYeKHkz0tp/
5Jp5wiHVAGdg5V7r7D8ZKgRHOFZq1iIHeOlP8/KyOfOxwlzDAtQkyKL+F6AoIfnX
OxVb97AOy1o7A6zAidiz+HNrT5PKhBGloqLgW3fTgxUEqRKsh5EJyuKfqGTVmRbP
L4Zv+P4bR/eA4N0z9/5zuI0QkpvOVF8zOr/BDXu9gRUy0cXDMfIoiqm9laZO45e5
EQGu6gyNb+oKd32ufAmdTC5oXurREgB5ZIjTwnXgFWG1YoTCpKbezAZYVAJw5pcb
6zwMcXm2s1Fm5GFF0Y/603A/h7QHavC1aLsc+fEsE6k0ikh1iaoPU00V4TYcRWf2
5AR3avYk/CFmJtDfLRZ7gBkajbnpdw9ujZFU8SoVSo0y1arkafHbbXnem91h2mPU
I4tHDnL5QrIm2/QTxpY9khy/MKQFRVIGiHGa+3iAuEgeGleYcbAvWCxB9vKrOMnm
xWlfnaAN9mg2T2R2gTjNMp2ky+vzxzEnq6Pdsc9zclRlSKtsKcfBLw13QVU5QCF+
RkKwuaxZAS5ZRbCbn2TW5KhBBu0/GhjoVWrxPrrB5bVyFqv+ethqNTO8hxyhYS07
2QWCHy+HhhDeUhE3fKK+RirTIdvV/sJ79DV2EpoF5MY6Zn9G5aJ2i7K9nEOpFIm9
z7b8CQ0tI8WrRDGegj0Z2FL0X/YLcsfKNmpeFXa5D/c6HgR9EA9SqKIH+H4AhD87
e+Ws2FqfTOZ59cOXPFnXaZKYlNr+Jk8WlOzPmNtl/KsOcDMNHFcpV7Ybx3ekAevm
z/rRpszO1xVoTtEdVagpQAQqr8xmH9U17XkbOlVF1MlMkCJ29zMyABEpNCqZkvh4
0nYZ0ZtNePlHzl2ByD+7qh6t/ZbwqAOCEQF74AeN5uqxXMiLrIOrQP7CI/zq14dG
Ve6gBGzD1pgDZpYw2YfOVha31dBOXRP7hRPRJrx6WNxG02cduCUNtwrLazV5f5J5
+TW2CLluW7x14Paq22A+rHtAzXdu5bWluvaN3kW8nTNDCOU5X6GhDv4g6/9vWsRF
dkjwsmgQWqQs0Z47sP4+X6so11tpl78bn+L6lsV5tIWJgtpGz6ysK7bJGGHP2pvA
aMl19kx8BWmUrjO9BvUymEK9UJ4DkN0Bu/hgzu37VCNlZSWI9iLwQIe5boPWh7Lv
uxPKUWEE1uiWH57kWMKdQKvd5xrc6a5XJxxZNqSOk0AWiRKwySM8DAeS8GIWUE7+
TfIblIO7JAdtA/ymssRFeW1C+mCFg1/9M+Z2s5iqkbvreV9ipbfTzGD3yTpfjrVj
CWSwnc0TQIInCAisLd7X6RoNmukJGuZOeR6Guu9kJmRZ7UNMcqE7FbJieq151DG7
ccN4O1W1kM1STY4PcASFZyI9NRMdZQ+X1m+tbHNUx6khi+QRpTvo7Qhd7LT5lHQk
3hGJVBvXirCK7UNw8TTR4O6IefVV7WS8vYxysGOFuX18+PrOeYxECs1joYqtNc3j
pFtucB855qsQm6pyK/hxZAMePgReWDXu+wj1H+qq/W1M1gTbhVNm4p4DxbwTqhLX
0/yloepNh2Fl1ltnppEw24j2kLHn+ONwR4StEPICf0fQpkhw1aoYY4ZWLSwvXfui
HtsqYA6kM+0157pn/HidRr/kpmcFdotlgITknXuPu5p3terklqq6e3lcyiOr6xbh
fZ2Nqt8qZf3pRqap49tABN8khM4Yu0DQzP4IWMEeWAHbnXIYdBHxw8DCmHn68LYl
3MA2ULF3HZt+fsk7c6wvyg871Qw7lJATwei+4IAScDhgO4glGcMwaqWdHAPppzzQ
YDVHFu1cyd0RQ9Z07H/6ruVCRlbYspNuo2E3bngnkQndaWDCSgcsiM9S5UMnYXep
xQ3KpuDSkG1Lz4zc2T+Mo1djv7Mhhu/jX6p4Vyf+ck32fmIl9mQVxd5nhK7U2JMb
VrHFd+BgrpXAfe6lr4qFpT8pTSNMEgFuaaoIIs6ePfbTBL5KzsRBEiDTpuJu/qBS
WGR3h07lmcok0UtrjEk1IH+/3e7jGRS9vCqRcTfIgFaT1BxYL5hsbexrOtMsY3z8
KeD67XouvXhCGFDEmsglQTuOrsbLE8wUIDQC7zwN1AytFferGAe/PWXfvN+Zm0Rg
SeunLVOW2yMUsNsko4/hyD9hDRdOYkc7d+dRsFs42wzJIOewIxXfRisVptfawook
Mx/WuUxIG767cpYeOO6q+z+8gu+cmEGE/N7QTpzhHDoxK/hFEMpXLJUgOVk7RT7R
HpEDjygvECKFuVT3uQSRgFJZEgSOcet+a4F7+iQi4uNqAMClAwhvl2EGlVh8uBXq
r8MQ6WeeZ72wQS7iX0+PPbFTUtsKzE1zrnIk1Iwfs+U47m+k6HDzyev+5PFnj3oU
AIcubz5k9lCcGdBDnhV/FzU5LYqBMTX8KfNZRXSYDZx7vZ2ym4xABdvy1sy6LWja
Er5HO+MfGOiv/O2Q2DS4ut4IExh1F6XDyamTByszKnMAYlH7MwiJZDFQb5y9j/9K
mRL4Z08jjVGLD1e+jZTdIN8y2irdXEZ3fal0Qdec7M7ohAJ+sZbiavvZOFDk8sKI
XbYZ2Xn07Yok3NHiWZOEmQQzRrRflEj9aBPxbk5CS+HTELd/KnwMe8Aa2V3Uaqfe
9DsjOzAl1TvVCjJQH+vCdkEmRngygVT2PECA9Fmli661+ZG41oDFkA7UPdmZ16Sk
VG9Zgk7QAvZlVlmWCK1d3t9iiRCNfOb4yY3ecKggD8gsBUvkrRK9LwcsANmycloH
IVHIAdcahkHBSGyDHOiNWelQ4CrikLUZbNqe/+JN2zuwOjbPcZZGtQ6D7JdwOdEq
yiYrPveuPIHBY/Kda8cxkueH/QUm1WVoeEdl8SPaKIxZWBV1EWCfJpfKHgPbrXng
JTIuc19QLHXg2yOVG3xWJfLy/E3EQjY2VbRjYgCtUOVutKhaVh/17F8VrctgC/1R
9p5a8RIJB6fjtz6x78fsLSKJQ2WTBZjX3K8ifXb/rJ5ad3pF2Mlq+SbFGGaSOXTC
K32wRuEpd1Myzfwa3rYBxYs46AIOmuV9gtHMJT0JTYye/IWwUf++InQniX2C5kSh
UloxtpZygMFKDnaMPvr17FE7MmUc+5VeJkVhO1INF/Wdmj1IxUDQxtfwaTN/ZAL5
QCkGBsnB6E5xJYRceiki5M+v40dZ6z7ADL/XLLx5AW806Jfd1eowKA2/6cEYVNbe
F+pPoH2dfizFPbIkxN4z3kMlcQj40AnteoTA/fvURc366JUozpM9B1Az00sJ2gQS
WUzMN/iTreHMTA+Qfbn0SHY0ydMGuhiLP9UwM6fHNBjSopeuuYVmTNjOPErxdEM0
Cm9NgHzS7BCBXP4/moBwLN2+hAXp6+n5o50Ug5qzDjyP2vcD0Xpt2bZaAybJo1e+
ANsQ5qr3y+ZTbr7iEyzQ6rKr6I6IUhSD76tF7c2QEEqfRPAOLqR+BrAwsdFC5xwn
2ru5PrX3zuN97wCpf6t2j31Sim22OhBih2ZSnY4D8ob9LWi2TN5zxwtXqDrsj8dN
m6CcL7GGaGk+spXr6UO9Eq0xdZWZ94s49Ew+jrt75DxCtK2Ww1YdBRreF5MvWd65
Ow9Jxzlammw+yAZwAzD2VXsacCvLCE2yn9DA+F4pb4Ldq46b6kfa3rXn+YGBj8BB
zb/Q4Ns+4FEerqBpyTvFwKKVu4xDrI+TaeVqwQMXNmtYiwpd+CskFf+l4eH6cNbC
3Wd6jdQedgvdQKt802ZO4ylfKhvsYko0EXjWyxDWzmYaGqHKcUTkBeYQ5D/kNgZP
kXtrWSRiOM15IJYY32dLsKy2yFAwukhEGSxR+QEkB7NV+gUFuvdAG8+sJNnN7dSl
NDOBg4ua3nQATgkheFHIU063wZQfyWVfLFh8ijbRzRahGe8ucA1TwYdvUhpGsvB7
+0MsuLP7STJ1RKIKX0XMhmTYMm9EQ/Bb0rmqcJYBtyiWjHYBawPkGlwozi6rPJl/
hMqG+cNfa47YD96nbyWnGnDiq10+vrgqe9n5IOkzkixSYE9q2XW2PRhLmtl9RCvA
VGSmvdK+EvKOqGiLRQsHZ6SUECPmD4pAfzA2E6dYAyKU7RY9ngvENTMajLrNC0xy
GEAlhlfmqWwbhZSAKuuWersIKY9kLSmp22RP20zPbNk1lKGrT1G0dRK0BGa2pY+s
Jo89cTxKtSUMNG8kR8Bgft4bTUpa9z3no45WvmXovTpNWrMnU60ynGUWcgpC9Yz4
XwwZD4INXf19aK/emoD+LDdBr36pmbaT9DQC12bznKHVCpOPvwtlpfJwV1dE1nBr
H6JJWiJ/rAvbiXXiTalcE9Ooz5yyZtS9icg+jx/hN4hbufk8hb3MuSVcJtNHikey
+udH4AawOatb/fg8/WrLEhsMpuGNHf3/lvm9YRkNlvO2sfjpcMkYAk3IMBuntbkI
UiUR3EpcAxN+4Rt2woaIs9eKaFJeb45EsdMiukCfqexYi5mySIox+JUcRVgSGRtf
wKnG4rrp2CukXgV5eymfGj29pWAqaJMroXThP7Tag5UlT0g9X/FBarP9IYNAej6D
n2Nug7OShTfv7oue5va+IpoHHrRbs8ZwWpo2tQT2iQqb94evOQ5145RnfkpdscIa
wCCc7oHJ/du4zMJpLt0j7qqmQtmKIrNxBJ+AufAxotT2oyvip1f3SNJP8vge0CF7
yhQkUfyDRqmySMjj0Pdo4ZDk6uzp2S86MGY8LK3vbmT3/NLFmGn+1jgPaqAU//ub
6Bai92JFpi3zZFzHifYl6O0ZkwYvonqp9r/oE4u6NfOUvDJ5GKn+gcb0ql+zHQxv
I4IU3ivrdSG4sMwjpHZIviVIGQQ+BjODAMlf7Iu3pQQAeS3hnITsAZJlcmkRGloo
Lwg2PCZyfYERorO9l2x4sDUZ9VDbTtkGFgBgpJDYb90npDlVmsETfnhKBRkpuZ3O
YykLIyL7QbgSDfvL1+1gMVyCVMNRXqkgNrH/F9SvACHtJ0LyVWd11h8diquP3oyo
QcvZ2tLDhIg6fthbxp+O70hP3bG1OxopTtZ3DprZh7AnWJD5WYHsvmWlUoRtlXa8
+uSJ/yNQVdSdn9zsPkUG5LaOwfqRuyquyyRlVugiKrUc8rvW3nUWpyNEkMzf/AAv
Abt2OCuPZBH19yc1khSlGulDaWxjK4QGKDQlgPxAPtgm74EFTZjCWfCkqyw9EYF6
8s/9P/370xWjAZ3oCkUrfbK2zIsjLzyaiw//R2YMZFKcL4NlKPw2PFpVJiwlvA0j
QslrfSD2Qrq05XfJ8w4woSRCTp2wBbqF2RwaKPc2ia27tZVGBw2k0YTxbCcrZknb
SqNTaxnCrn9z4AZrbs+LcRIcqhu5jwGGPDtR6tjnG3LCsZDirhlG9t/PnDBGNnbr
7E8sQwmuFo+sZLUgXw24TgdIhCzhFs1Nuj3Ao2/N2kgqRZmhxXCf/sWnjGJoe5y0
JCN9k8ItFO2Uo3FCOLFZnS5Xt5WYxBjd3xMV6aeUczanW6QC4t4DXbooWlr8xO/9
ZiK60ctxJPJc67bkNC6Sc5v6OO1hz9uKznIEsfUdDwRCiVHttvVFCawJE5K12i4y
Bup0iknvFZSA/zLqSTfD1++42jXYSoJRmcQI7rwbvqhP0QvShXve/xUqRUPVHgPF
fBASzgcav38P0r29gGmHOuoBi3zhsMvfVoXmTGmuJjwGX1l3DCLBohX3NoCk5TaO
gJJuC8tEo92b02DnDbO++EobQE3fOXfezbBdXqcLGkGASHf+IBZXTBsr1tLRhEZ7
/FUXFrto5PTWZ2iZO4ka2ZuMz61cUiQ/ey7SJFf3i3VYfckXdKlcPz6LLdZHPaIJ
ltJmfnNSsXqLh+o3ar9csb6x6bLpgxv+Y2wZpFhQ712l7sYllNCj/lh500YdVdag
9BDGrXmDwvxnsIqDh4AxsKp3MbqrTzOxvbpBRDxbtW+QmFGgfz4FkgcYVZ69BMsh
6u0IJOt0LqQ82IX6HtdIS28zY26eMgSQPhYfhiyuVZ/Z5LFSYMiHoUvnweYENsZl
7Sb7aySwPvZmbpk2Tw6osFNJ9buvZsMKewcQTrMC39xn+O/NHQUGTNuEHz4b3VvJ
RWqm1gfX5WTxXSw71yxEVkF/DbYaNZ7xbWi7qbHEyJ9SDPXP/z1Ct4CRdnKLtRmL
XuVqaykSkw/df6N/14FC5BS8OGT6enorgD0eKjlmumU044ZfCiHy8zXvurmybZYJ
Ke25XZnMlkhUsuNjh4APk9c5yvO/AbcRU30hFd5b3YOc8C7xTuCqHMQHbSr7xS35
le1caVIeck2ODFtqz+etX/pLAQvkVtBWvRw3Vl3Pr8qu9/ILIxp6bibVZPeljeD4
FQEwsTEJ24y7D/YRgaOU5RsP618/trqXYBhBJpuOIF6RIDLDHBdgDGlDzX1Yd04U
GfMUWlrMGvh2c1N7DOKaXf5fGbiHTvWlck+3AiuspXMEaKVAJkbcHX6L/0pJJsO8
a50473OI0ErYPABchiPeUlxK17SDkbaP3MkauCjc0uKmyYPAkHEgLtOgIUCAJHdh
DtBysgdF37oLdPI6KVaHd/UdNIvf9Nh+PzFBQfwQhhN7A+n7h15A9rnY0wuKeCQm
3oiWSAVSeOpMnJHJUEDfCoKtCQtNCFpp88Nnes+aNPbL8CgKiVfm4D4yr+z2CZl3
2YJaRJ1/cf8N9yo+X4xEMJ9DONKwTp+5sv17H8BIYmhcfX0bfB9isYBrKzkBoMs2
hVjQQ/+MViJ1oh7z5d5lo6oHl+lDW5RPGgHcW2UxBraJaecyp0zhJmbPlIrzBOKy
VfVpRKcMhfXsgpYVMv24IB0VnmgtcoLMjcm1S3AsT6RxB9AN/EZJQMS6/2Gi7NUJ
cb6RoxpkhShvmwtKFemtRl1kyNy4jEroE04aEt1P2bQRRT15i8OXP7K1qvSvoqAY
TH/8aq8RpNsSPorTvLO96qsT4f1im8RsepGgTeAv3FUM3ZPMcO7oazZeokDw8MPD
Bqjm5QViG/fW8SEZXf/2ERBBvGGwTNsKNDSwkW6w78nbooA6WhjQvsz70zufWgyH
X7WV1FV44vLRW8cGQwNHpe8VhtEFTOFN8ZggYDtUDZimy/u9U53vQpq83qRByzRp
Uo3/HwKLR8FQtC8E+OEmzWkUnpRzYi2/NXMA783lt0NtClHM9qcD828CKzaULXIq
Dw3zIlrMA5zyZtwgJh7EE5L5TUaoTZwQzxWNsAkHx6Gjgb3uIJJGLVUh4D7wFCd+
VNbF2Kqdhs+7jNS1pxIXz0UD+YaghmtIVhJtlvWuQJ/mGoo0h5mMoVgPvnGBYZ9K
h8rSuoINkotR6asg50/rCwy72+OOipamYHA3gSn5CTGGPX9I/2v5Kr8VUcLStP3o
KQGL09/8oV9pvaLxpsfgIV2eUV3McJjZdeJrERGLM/0h+Ik3Ap8Ofz9g6sXgCJco
k+Iomq1MrS0Yc53fB3MbeGLGKojakYcoVWsy3VF9rDVpr5pvKNVrvXlqJ2xbv0+u
i8rv9Pb/bdN7Cap7qtfkTXvgh3gvBW8+WgCC0i5WlJ/TyQg+YZfMXS5a6df4/WB/
AJoe7tslOwJ2LHY0xP6F/AHxwWh5pSbiXoo/qnLyWmIVM3dT6iqMi/lVyFxDZ//J
lLpvUDCqnP/47hBy/ugmyV06utS104TpyABjHLUtvARWahq9DYelOTve4JRjCt0O
jycbF3PXj/Wb0bsKg8dcJIvTEgVL44X3Fb1DctWisEVXgMdJh/7jthrpI1Amu7Hq
9Qb1izZR2dPcPA07uKPEmI3fec55xXSZfsX1MNQ40M/DxdHAtsKeJIK8r4rYEOIf
lFNUq84EC4Z6ZtW6iIuHjdrE+VTjmgFlowUxFyNTc0NJMrZO5MK7E8gwQTNYasuP
49xIeqZLlin/MW262or5Fw4MJFRnXGeM0tcT10rprKZlhlGytZZ98hN1PD8jnqm3
L8Bw0loK9XD2+4iXvGawPWWMOAH6vx/wopBnW9PsHc4uEQByDc/JeY2EPOrqVN4m
DF5VF7Oyuxw3mfT0KKdexGxOeZ43yHrkeW7eGrRmLzaAZf6kjrPIjN8y3x5Pnzow
mA5JXXO5Jk2vvV6RbmtYopNjsywlSQ4/mKDlSEp5uCT4lCbOYPLcakiaT7FYoSe5
iUTMlolHJakiAfYZSqrfsEgLU0qqLWqOczXVwsRXvKj/crZ2fXZhZJZQaGSuArg/
VA4IUPzMS3IFq2bqpLaeUZK+PDnfI8gGS0l2fntUCZUXt2eUNv4LLrVhkic8rsjk
EZ+W6VLAh6q66wBVxTB2JTxawsQzeo74/ut+qaVs1I6eMSONIMo3djWLzt08nL8f
8G35al8nGc0HT5lFcIF8FLJJOYoFUbfhw/6pxwgKorerAV8ZD5iYTd9qiYehJ6U8
C9TiVhbobW8fG3Ny8psfMqRrPtjESfupv8bUpjJl1D8u5nVNuEmFUbaU9IVaC3Ix
0YjXrR4jW5JtK0j8mzri7KihL/s2mKZHVHB2lDRHZCpsMG9YDEflPUzdCwFVCeoZ
xIWxKFmkPyeqIY6ouZo4a822sUMhMS9KCI/YlcoriPkmScu52MYOncYO6BCgO825
eXVwSOT9fjnZM3TleSOa9xgZ7Bdys94OKqFfL0DoaqEovKrcwCSKmpECWfHMlSV6
Y+aSjqs3hbE1d5LmPmgrpFJi0OAhJZI4RLs6wkkmvnbaGTA4mLkrs8U8+eEzB6d5
iscgngMa8uq/gCfFC0p02yH/vCflvpRvigYTr1hvONZihPjdtObfmjQbDkfZdlKp
+JpAA9megZATCvWqXjok6FHR6LXXrmu7trQl4MXqUH4tPsnL0DgaAZmZSPJaI2Eg
cyLVXGUhZJt4Yh6pR+Ef+QlA2n6ctLdAGfSHCB7xqbXmqLIzEGBxZs7DivNVzW5B
ph3Dbe+6bN4dtWGEsDNCJKCnU+8sDRDWqby6pW8ZHb1ylFTzs1L8jw1K8udod9lo
4Yn9vaLDir2ZMKYn+Rl75D5ifJKpBSKJJYT56cxp8v8zy+tzHVDqxEirbwQQwGui
01nomoToqDBaXAHUtyXfxTgm9j1a0KT56ISa7RYMx5dXidOxS6UbC349/20WhEhl
ymkBryCH6PFeSX32RLHhwO51FDFo/dZC1RMST3qvWbhhXCndvCHq4Se+4rtFhbG8
ZN1vC0qGwoV0X15ppb8XVN4O2eoPrOtdW0cw3l3C/v4kcGg8LS6tMuzL8scN7RQz
bAYH15pwwMnQlQWQKhBUyiY50Dd2aub774+xDytWJjxX0KV1XOl4I61h6c5U1uVI
7fG9A29JH4v/4mwYbXIuyXYU797CN/w6OhXirI9ZcWobiMQS4bV3yNTZD1UT02b8
pV4iGacrIHNBy1jV171qrVBXcbAN1ocqR5qiSupyFfDfKaKTV00qP43Eqdx+95gc
1D6XkSQr/GyMNVPVRhFIcc27dpV2NWByFvKUqgR5vYMoQwriBVAhbWTdZj5Zd5Ix
+FHVlQiQZyAYu4R1Kb8ZrizxIcmuPh0Dnw72MpoCdRs/psWJWFFUbEVtg+Pek/a8
7AKbNWXJoeSDV+BH61I96W9bCiZDZA/HTw6k7a66gIwJC1Vw64kLY01y4ybIA6QF
aRBZGPnDSGLITfZDXR248Frxz/wCSadZl+gZaEu1DAzYiQJP7iKDc4SJl5onGXak
iQk8B2/Pid46bntJum//GPn5tenA61acbsfbGTsBu0/8bgbAZJ6g4RAR2kFYtG2z
ZfRRTsJsjaHTYwOee8DBmfmbthLIUO71toLxG+eRsvaMrOHMegdKzGvafk5kULPk
O4PQWrd4THexizsKnvFu8KU1Gt3ecm3p2+mJXYSjFjHIrDOSv3I1sP+kGxBMJ0lQ
SM/yY1HIn1tQEirJdgNyBUHEzyy1QWGVOtcYeRw7iANT/m02nrRgOE5CubVEFYXM
+WGeNIWBPn5wDW/fmI3MmvmXC8/6KcVWKgMHwQaEylm3nAp2449UW52/0X9cQiAH
Pe6cJBxclAaQ81DcKGXbJKMrZ9T4bD5EONjFtlHZDl1bmTjLEOUl1TiWhY+FccIL
OVzMbQpMR9ZCAqD/LVZ+PnMh2PeU2rXQm9s3CA6tIFYl2jEdo46HwUHAzQGL9UDG
ra6ZCT8R6dr32/22HdiMfek/GbwuyWHUfTUqJrm6RpQyxNGJ7tE35jAFFGjoOVPT
8mevIrNlKsZ/qhNS57MvtcHZnz2K1rW/u8o5lA3liUPgnRgFdKb2k1mS8h1ipMhP
sVl1WwX1owcB8m1f5aDBW+wxUWrw0dsyYjnYJEzYHlRqGxlKXn9Q71zoOHF3n7Jv
hFV9UwTrV9XtwrHc/CHEjzekjMoqL2/REHa6O6Tlr9FDaWN4jXkARqJgn//ggh5G
+P3iaIlP3yUsOU4M8xDKCCruQXCGjTKTgsUK8qc2eUUy+S0Nl8CNNYLQ4gsANp4y
IguyfNY27T85anJZDcSOu/wqoEKwpODt4N+eLIL7lkjmMObML9vIFALVeOV3CL4o
JZntd41BzsNsfwDds9Kr+E98SCprCAzOnuBKyC9nxnNdrarkgo+FcBgpFnx3aQ6I
gQxmEmOwLMVSWxh09cNFBNKW1GS47+4o39P82g3IjvQ9YY+WRiz0w3VEV3D6S9qH
/GNtcG8ye23hTWS9vYBddAt1yWiGa93BtVEuL5JWxs6N9fEJit3zd7NHWKo8LSoN
7RdcZae5egR+hp+/nkVvVxt81YCri7hOjbt5xCA5xLnWVkhU6UD2JJLtTT1avr0K
3JD6GET1kxASmwoOJ/DhkmZznXG7lIsriy721tg5thh6z2JR0QrQBjKoliRcvGT+
0Rk5ID4ZTYPbVzXOvn1E87myO9BqhbTDTRfJ1UPofHz7IRBN0Xo8F2c5+qTKBTzk
jiFzf9gIDHoWv/uZLc3QapDunBVfr9qefkgHxPeCQLv65mtc5wSDUf2BTo8F/JdW
DT01EjhzMV/wXKvNyXP+HLY5hC+0ZNzCR7I2WgZfw270aGj34SWNN+URyasqho9n
vhjh6tpWfda4iaj8WnfKLj44lH7jonBJABjDP5VKcvcL7z5rWEllOMhTl8SDm1d2
YPyyvr4ONdjoAkT0V8YnHE3Yx5gzfJ/q71LDCeHCyZHerW70i1xY76SuTdpcMDOK
1HHX2fXkg5Ajb+MrvgQ1cBRMkTR+7I2EVkxleJJYu9UPFlKgbicCVVkuUCf+jLF6
A5uQ+iEKJlW7bLRVQ+pqBbc1vBDlmEJMH3b7gQ5HI60w6BZcc8/A5KT0sIULqNne
uTB4E0OZU8Bb59c01RD+Xmw+mxm3TW/zIzVTFfHmmSNkvMAD30Uv1zDWejdkk+aA
e7EESGWLz08TJoB2f27qpEGie+F4U8tllriiyQSCUzN4KuOkQTovh1bHTLEgxtFX
QiI8zEnpSo9UwcgjLH6pkO0/hpcb47X+KAJXShKzAhs1lTk/fmQv8QyCeVFvXfLY
MRZ0kUiwpZM8Vng6JHbBmm1Gw9OLpt1xisPOki92nYqOj6Ok9krG3bJOpxsH9KrJ
3B9R5Fe+3/38fnNZAkF6rRjXgpaHY2NtamWWDzkgnsdWk/4Or0/MsfKj//3nLpCA
t9UlGVN4fi3h6+GcEJLRRke+jzbZCCTy9V7GKgp0BHuXYtIBSMczBEvA3geXfWMY
O4T4hM+trlE5eAeRCTHbheQFpn5Dkj2+MsMCq26sEctkfIMHkAkJvgwsJcehM3Tr
Zwrvm/E+G8tXvjd1PzDTLa688ZOc3sMHFC9xaxlcwHY3DVlqMEWtyxoJr4hpT3QS
snTyB4ZcS6HeFcVdrwGF2sTrvXYIrgKUozygKQSFJdyCryANmG/ab6Hoo3Uqku+t
5Eq0iLE+bgiI3UmwaoTkeMz6iCSIku/ns8qHlM/SzJBS/v+RbuIt6LpCsTpakr2b
b9SJyY1PgIdUUNYW5TzVmsqoZPDR36ucsiG+NOLvtetlayUIn/pJJ3rJFcQLZyF1
MatjiAhLvTdrX2zcMAIEhIfsMxLooRGUfQC2CcdzGxNvR1Hn1qiK3hqD2lDyZ7Du
XDuiRTkUayKE8EM1pDnkir7/1UXMJIcw4J4l4nHddvUhjg54Y6NdGEWb3T603CQh
FhinjGSvSi9v5+vC67i5AsKA1sYsioZL5PLnkLysigmUJgmkmGL11ZHbOKjjSA2h
w/HeFBFR+mtkRByMW94Bf04/xsLkMKI4JshoaEpfH80N4t59vKr8dBhV+/W2NNTq
zu7mRQGapxs3EK1BrFtgxxZ651kC/78KldoWftQRRFghgOZk8HDOmette4/fY6A/
xyX0xyO73pVPt3tUUlN1Gg2JcQy9BpHOpZjTa1IyTqUbAZ2aC4crF6FmJ37FdvYB
vsBlVTN3Qt0bVdR8HGFfhHnoT9B/l7uTL0+te6pE9mpwJJiXqL4kWqtvJe4D579v
7lIicDoVVadFq9m14SucItxk7v1VZsXQQrqVOezzQxrIWxttPLdSqNcqviBHegfj
9WSjeLGa/5Ol9wXSUUPrTqN1cOf4kiUcv3zz2YXaEwdSfvtkvcIAUSRIlrhXEz5R
/IpF9KaR7GJkwl556zDHwGmhHinrCzEwDn/8XAS/NsIjv0BLsqhT32TEYb3/d/0k
z57sWcBRAAjRt1rBds4/SVBz7EsCITmHvrfTRuelWkb+o5xSwrZNRF0igTODN9z6
nI552cqnqQMSJdqxE/v4YNjBR1JIqyY1PQr5am6KnM2X4pCFxSZ93kGhvP6gR5oE
y4qL674OIf5UeU7HbXackkmU3FphXPoBaor8HeztMb3aXJt1yJWUEAQHx3s7t5Ie
YfM3J7wMcquK5krKTdu4+CH7E9/9JKmDx/WWbpfIlWDmPJvhIm2fiJL/iFjDZ8bs
hHdiaL5c1T/qUy/ZcucqsJShwOsHGDGn0x04Gs8Ixp80ZXSjyRet5LCu22ha0nh2
rz47FPbW/CJDJhFPP+zVB92fHYoEf1WOtuN1+Gzu1T+rYhkVj/QObHaFamfch2rm
XlBo7LwGM5OLg2kknMHw60LMV70OUaAgOJfO5zPZHVLlguTWaCSMPPRinq9L8jj2
kj4FlYpW7sELBbyl9ScpHuesXZlpJqfHaogqBeB2l1OCI1Kd+SuZd6zHeUk3Lwdt
QpPnaX/ppaabc1SrkQKhhBIKPqvEXEzcV6Q5YyDQyXWtr16az2HXxjlkBVfSMZaA
ULDZWTPZCJoLyVWv57s34ru1SLonA/q1HtSZmsiAPU1fpg2SvJbCmCPwiUoZnqon
BKNYl4xSMAWhW0+9uRJ1i3SRhRzySOyIVraJ2crPpdzi0CBPygunFatPyKUvUdVv
DtzvOUDqSrDX2epaQR77cyYKejuFWDnM531LMUFMqesSJiv+L5t2CnRu21Jr7eUT
cocNRwV81Agb5YsEVK7UkWRSzk7gRm+HGnTsCg0Gthf2f9Equ6nDEL/FaXpVNqKq
dilCor1e+DRbccJ1UM2FlfbvkoM6q/I+w7ra5mstlXsW9t9I3WlgPra2aggxpfiU
ID9JQtrVJabiNw1GCgMQ7/B3RkZqiiKTbNPkphrlx1tuOgPsEV2U4msQd/E7JLDd
izOREwSnSDu52msvLm//tqpQ0VzOUhQCEtemBNgqT4V0IDfFyiLZ30F/L/RvtluM
0onlwvdygVX+8ywnpo2CBZUJ5pxSK3JnjPl6h91mT7SX+F3PaAvCf6rCU06mwJc5
u64bcfQCeaTAFT7jcC6iAHi6IbFFh5iW4bxHd1fr/uWosnEq3JI71wEWXQUW2v6Y
W5sP5FJ9W3hukXKUBSEHSAkjHJBfNogYaDg1xEIuDqYSba8Mf1DpXvheC382CY/A
YHS6VarzgGiMpV8mjbqx+QCppIln0tuS1nmpNRmEn9cdf680X0ZmsceHTghSW4Sv
JWVWFykQALRpFRAoZuN5olyKTGo9j+I8MPGQxIAXXndwve9gwMsDBc1x5+6X7ZCE
vo0EV6x+db744LeB7pfHwrqLzaEoaHdGsA6iKgaditHD3Xo4GsigFWXARRlp637q
JkaslrNHKUZLSVDv/1+xZI1QNgObGNEmTIuY4SyqNvkF4qo4E4FeRtc3qFLPKkJ7
7NVWjDUSs6UgsIoo/+UJHask1335puRSYfOcEYZlfffXpOSf+ZFylD4lRJ31kkTc
FyHdA4K1VrFN5DxgNbJ95QlXsFCYCJla/sAInS3fbCbBIBMSUZajuFhHtr8IZqOz
hGGprBP1vWDxAjoTii3s4t9+vvIJZmf2JLdz7BvgPLK4dLPMecJkQGjaXYn2hVAE
Z2DTEH4X9HVm6zSmd8SRsIQfsVW/VBFgyB2H84L4qxmjslqoTqaG9SqW69vcziUj
YbfzJGNSsm8wKuWbj1Qw1uHnqf5efPw5IItaOh7yvEjo6lWUNfrvbN9bfzxcksF7
ogQPv16+lu3oY4TowDfwI1zt5xzx2aloJGbCnDFGsx3IBoD/F69qHGnzAN2UpV60
yGgipxnGIpVnv3tjVRKvlybA3flpe8iRPzJwm46wZh0wAuc83JHxwXsxgQhfdPv/
rLA9w8WX48GAIOKsPWPbIU4ndYW0423NJxuCBrGl2ryoxPXp7LjP46kyQ1Cg/Rma
qhGtxEHeAVPyhRGhsM+H6+irthMmkl6R4jNtGJCWEH1Io/TB/RILcIEH9jcXDYS+
lwwdBzRZ5nn2rsljLAmU70KEYaXoaWJZy3dbdZdb1CSJWRfqxyNUH3aoBL1GOT56
asFFS+vek6SQQ8RpyvcGbOoq0nYnV6TExSRqWVzx1clflBVgy/BTEVVF0A9onIRx
13LssnNrlJ2FxawUMacYpiYvK3rP6WvFrtwlADvIvy3EvGZYbZstD4isaqoqzStk
uArQ+SAkcrLGf8KS8Rlg90tl/jLKw2pwWQq6sjP8AplfVmt32k3H5qZr18VhYg1H
SssM/d7xHlJlJ5ELuiu2mA8J1YOpWKfRTIGyG5u4eM3DPvgmK68SlLmafRNazZ35
kMZ5M6Px7ARAXd41jAVmvAvyWtXa004GcwUeJ6kVAV0t/3+qflKpuUThJIE1ytHF
2bDVDMmy/9GgmbGwutp4v79kux4wYOT76S746hhrQQlu4pxWNSO1w21bsvAnKQUZ
jyEMWrhMSKvsuAJN8R+gJe1MtHfLdHGdxPMxp7Owas7B1hY4srS2ceJ4AKkeEQge
ZwIf8fFUQaL6fFjpssNWFiyj+M4ym5VCfILbzc58qnQk+gIluf0GzJf40CC0y4ru
0H24Sg9FqPe1A4WGHcTzaspJSN3vAfeNQM0uKfbHmG9ab/lVEoNr5E0iMrZ/JMn3
p4mS4EA9PazXwxEVWPh6QzpzOfWETsy66G3YJ8+eZ/APyDkAVcA7m4ZviFEEPPQ9
kU33e2dKh0TCtJVGyll0ddzGJ1l0bNO4PoPif6PtqmtFSaEAwjmYrE8K2jrQ70Yp
W7a+q5HtYVnUCn1ndfM/ml5AIk+MhnF7FSz8ot0GGwF1uBmQSLee79LVUgw36uwk
KqgtPvq4JQZOTz07iPDEu0/3VWDmahiS8SPmxQ2WdftiWy26d3zKKdWdhh+tLIP1
AHJ0ad64Xkgg1OYWEq/fb6x+o9UprPRQwpa1fbRPxfvPIwq36oMTFLlDRTQB+lYh
pRWaBC2hBctxUZcWjzk+EuQBU485AEUBoHC0Exink5+cVpF5CuOHs4UfBWHVp025
1aM4qTVJFaMbGGrThZ0nxVKQI+ekdRzGptuzFwz1JXrIZZ/9TkERPyjhSJg9YJ/w
8zYEecXkk4LARNODQDWZ8N/490jUd4fNq8r+H6VZkyyi4umVlhDnnuwOIcJPqFDN
P+/rAAGvHrEbsXLNFbmR8t9XEirdu8g3IinmNEI9OEKPpL9bAcPz8fk5T4HqXWXq
yVWcoJ8433+a3Lcd/GkqK09HByqJ6+2sgVU5DMwcX3wV4YA7fBCQYFwA3Iqmskma
Whyf2tRAok/jv/UJ6F0WgkirApkL00WlfF+ILtGXTgtx/5dPhB9ZXOKIflkm0dL7
zdtx1w9fyox+KVXvZSql8o88UXwAEopAtjbIjc94h6e4quqjvqSzV54I2GoScc/+
9hoGJkt19jOLDZd5DqqknCSq3/tK5RccYjYe55iEE5j1UmONSEx0Kea9JuDKr74j
S0MAMizNoYERPzQjXGOEnOp066F7YT+s22kKJT/fGF/XXW294wRgVdn/e7S1WzTl
8+FrRhU+DNM6W6PupJ9IlV8o4waclIRNiMzcfLamqfw/+BPWatEoAELKLdupr5zX
SuXLqEo4RWsLpa2CWMYRIg35WHbHIrW4xBzNXMCY1Ccr+SleGTQMkTlwOGWGH3d7
ytvAZ+J3VU+CO7ak+lurLj2gkKiIivPuiA5f2ta9ibXkLHJSQSdea1sJvc+9+xP9
/yC19Fm27rmK/252vC3GGTA8iCYc4RA4tccWMBGk/5I6Wh8B+qc3CcAUDHjEfgYr
Uyi9g4TfN60H/SXjXbXLk8LmzQyINcA1L7O5CpJeRqg1rIEeEDdhUTvevvvQrrOg
Y+bDbCmrbR/PA0r182ucU2n7J7fwEuSPNcW88fMZqiF5TBYCdu+6DdinIWo1/EFF
zZAY1Eux3qjrLv1HtQD5SZNjfpHFyTlqgInMwfwaZILL9xVDdX3FbNf/f9CC3xIf
UyM/ZA0AE6k9N8RdAlcweEF/6Zeyy2bGa6tqpkHGeCw9yiazmNtfyXp92KM45EcI
PwmleZ7EBwr17ynS40rPzahQFYET4vSQEC0tH27rD+rD1zPpKg1IyYPnj3ae4K6Y
GUYLN0wvRY9yJiWhm4dpXW8nMMvXGFWzbBYGqkD2dH/FSfk9G/yE1mPcTzZ0kJAr
SHFaAIsJFDQ+VnPlIK+ITpnwKSrQlgPGyLVmtKgKLMOEKvNl2NOC4EneYrCMNUlI
k+1U/c72xVTV4H4BaF02cGNQSVczdbRe1UMDGIPChFlynA21RVSs3tYoiC/LTKRc
vl6T/v3PNtJ6hg20dEXoCBj+p8gp2VihaGf4xlkYnDRwEudGlgxKBYBZ4qFL3Gbt
yhjQdwqzBB8M/PESUzBIhNeyIwDf1eJbC5Kqz+9jJAAOvoVwRQcQsqnxND5f0xlm
KzRtXHAG17Q6dlR+nb+LFkBDnaZA8Ke39sZ44YMdazU5nO7gUbBNjPXsy8fR7zFw
HqzG6w8NPuAmrHgjDv+2zt+y6zdmUP62F/AkPlTruVh0G8Ey3XovsC+BJq3SrD+d
AprreKIIuMr7HeA6q25aX006TnnBxfRGrFNT9ye/Qjv4gYa4m4C9J+BBdbugSCfI
cMHUK8dzbjD67MwWexKnDBzg7uSuKNXKCBTutl80jSlsutFwhgfVHHyymFSZrzSi
4nY5e7ied7PAwft1P4Ig4TJUreyVe6ZgFd1xZGpfm95uCQgl0eGttyRZxlqxBpZn
yktCzWMr5Fuf8C+KLFrmwQOSv2z3HzeezwLEGR8dORy8ihTscxrztLDmkCun95lY
01pmsqXu6B/8SIv7PmEFLVwfUQN40nIozhRSxKpntYFVt+0fWSCrWPexpewHHTHk
WcuInyYW+GK0VQw1K45giI3LDxiYSCtD9FzVFr7JDuDHz6kA+ISQkNPArI9V+4iw
6Bodr0ySz1FQ7nwhKfjptBxtp4BPKgKJbJPLdljM1ZUOaM5aqPiuLydDg/bBjkkq
kMn1znotbbbbudDuv2nB/3Z5GPVabc7NSnAshAhZvmuvkxBC1Atg+ooygHtI/F8j
9RrF42IbRzpX6WL9G4t1CRERJkzldcJAL5we7LXuV4u29V6Yeb19r5Y9Zsx4q9sB
eXAb/1AvHk2ptUZXm8MEELbfrPUp/930UQzw6NVuNN8OL/31e+FwaI1hM8Wq3zve
dpDVHd+7tNX2eOBFWrRIaveBxuyt3g9MGm2CPWSkF7VD+P23KyeDETQc1WVq9RIA
VEVfJvKW8mj6suqgEBxKdjMdisPdAnMa6v4FfO47+ysDho1QOCnDCmGBS8UzfPY8
++lqtqpaIR6MrVrRJJXFp0NK3DmCG3Q/qzaYDxyiv6ICzkNyjVR+KSE/sfp0jiPG
ZWRp4QM80pmhIKvbhwtAzvoMlUOImQeLGXiYhDNqV2Dtxr9Lg1GPlfp40Si2HYDO
BsIATSsopjedl9w56PeC0Lfvazk+77meSqdTrImUTmYL4PnZLy2d3beGIa12V3TO
fp80jx/e3WCxCFB2eRo/dza9J2vWbmOJVN7cSjMcRN2vFTUug8qla9Fl/g5wG/7Z
+C4sLGuWYFB0R7DSO/1IVI+T9BRG5lSlfbEOCxnZ4omW/C1QP913LtLSrrc2C5a5
H1GNUAKDQJ1Menc63J0e+I+8whFrzin0Vpf8LZTuF/wsxlGVsiyvsLkQ2QfwLKag
ozxFvnHMnkAA/FKZCO1tauslfGsvJ3PP+uCGIJqh0pWnaSmQkgFW7TFNGx8tfQME
JfNpIDazXBfAecTgTLXzmiQomqDwZPfE92JVY0kDX6MzCSXlB0DCi5UEpada1QAj
KNpOS2IquKp1WjcwEKBV2eOVY2IQVheOzDwsZEnUjpUpl3yKxVBJJAUitweXMlgr
oWfBGNRvOteRnpJa732o/YeqOXEp2AOlCBrc5W/YgEhU1DN6A8BK73dDFL7KepWA
P/OoEuzx54A1pqBd5RQ5Oex8bny3HnUhRj+B14UG5zzJ+YArb1rJ+NelS/zq/ef8
XyhRpuI1S+bijB9g+0904RWRr5llE8cTHmw+x6lFNDF6zbQxpcnqNoBp6OAU1XNZ
kaxci2xQnsab+KXAKnSSKHQBmc424aOi5XYiHzik++z2ksIHrKzZkHVtiPezMVU/
J0pCy1DMv9lhGG51l0vQovKNSbKAZfagiAHPVj7cg82O2ckZSxtvbvGaRlzsCX78
z1M29QJvY1K9AHk1mg42qSRHamOHHGvkjiZ9ur6QGQB4184wiVf+RENCA6tJc2RY
usFL+2mC9HYKvH2CAF34gEJCkZ2CQRa5+XRn0rpxEIQruptWtOLSWo389gDciCMB
dC5DUcjc09i+S5snaeuPgMnZNYCoOBVqydsAFJVt8tAYuVp0Lyq/HrVT7qTJIGoc
2y/Y5EsZjTU5ArgE+LNBtHpqNohF/b4CBq8Mk+/p6rJVnzm4W0d/tb6jaXq15Jjh
SMc4eKGA/AjRn0kCHMwQXABkyCVD/bTacz1Jy/THwodQNv9vkMl5S1jHpduSCADC
Of5O9I/TqWaTAvqctFU/HL8VTpD78RwjIQJt8pKAJ1oVO9VmTrjtuOAH8txuV2jt
AqCML7VNsRtjr6CpZrclNxwU0zz/0+zas4/z41dPXY7NVYplPa83TevaVZuh1vaJ
6XFCWv1jajJ+QCpOYFQIAAUIXet/1LclqaFnnyzIYkB35cIw2De7u5AHbhaTaKek
bm+OMD0nZjVpjO+FN3OwMAeJVgmrHTXmAkiY4EsRdJKJIjY84JDJGnO+6XomQLdF
S+fHoGUg7bmsIb/YJHD2sV+KXzSJEetVUUrw1hxQkZfwKVvaPw5a9yTJSgx2gqMd
hGt2D+0mpJmXPbhRBZgfZg+fKUIlG+Yd6RlPVbTzuGnyI5MFj0gjZNXoIDL+UT5V
jfEWsll5cGVH1Fyh6aLvFELu8w2R+G+Nob43SXFky3RTfyybxUjrt41d0mrSHtiV
JkequEEgAHQ7Ojg/DGcC7oQTMe9VPdHfiEwunPKcAjndtIU+hAQ+Wl42lNG1/ZXR
uk3UHYUiykjFL1ITO+g9G7iWRI46ezNl34kVjRmO3NUey8bfM2wMiYlop2HO5iL9
5OHXTgNu4gj+l3ryJNDQIRGLshPnCOns8Cib+y13XYRbSW8AqXLE5tITzOxdA0FX
yPt4sy8/WVTwCJokqAJQNZSvwZ5yZal2ao/3kcKf9JCKSNKWbEutQzVlZ1zMbWou
dUbB4+Jy6EXcvEIj5C8O7sri1D4EwOuyjaUtMyfCpemGyOieR/I1NVpLdsagrch3
o3OSls04Qf8uDUb4A0spOC/JR8jAOJgaM/sN4PmszL2Sephfw/SqBfEjyFjTtE+B
u4XeMLNX7bLj5ya3qSprsZUDURtgqK+3xqinFHAlQudXWCmY0CfyvX0QJW34bw9o
V4GAfEcEmsPB+IGrKr6EcZR8gLcbAnVWZAmPCO1HQh4NpNSVALYdVJXLbkQxy3gM
MloWON5j1OGaWgCmqjxJ2VRj4FuPE41Fzd54wkSdywhVqwgCYIdaomw2l7UAgTHl
FDuJ0EEj0jypmqVsRsUepasLt86lcxWyxZPhUKA1kgNKupjSwW9yOa+tLcGiLCfE
56KriM8q30XMLSd7LxWPffs4Vsk2Iqr2BcQiSvhUjYv/SyBxHV2LRQNPHwd/za80
TAT9zAHTbCQGovwmRSLor+Xr5+W/qFy1upUU1PjPhOjYNqajBa4TRcHnP851SsOO
l8WIhTRf9HZOmJU7A1+rpb3WzHlLqdjPC1Q7soUv7gAPlxavCFUgNDbNvhssp5Fy
UkGpBIWR3rQONY1I+MVmBk9WABIy1ZUXKafD8BybzLORyb4FmvEmNkD9gmkJREKL
62EvDSugnUirNEwNogt3OPGUkFJPUVgnXhE/gkgTECOcTI7Cz5A3WMV6QcnCLJKa
dyCfQoV5So9Pd4u3+k/IF/iLGdW7oyTqI3Ewlan6VLWf8zzoECjTZmlnvKpaPIdk
bq4O6U0pPmWJx6THUOAXPLMrj2fls1Jsda/mSj2Oc/U4mvbRjYbzofKeLPKtxpVK
JDRhdc2LNSOyQaQd7qCnkq2xUtDZlFR7bcID8+Z9hd4ejwZpPh3smtxRCRaKT7G/
fCtsEDiRDdd0Od/YAnBsfi4bNvmDcSMmLMZcXh8PXnlGWTxIqv41iXNel8IL97KF
XixLf9uLHGIZCa9reX7nwWSZz9hM/T4rTPo+fH/mS24MzttGGvOUnK0TZ9Aqr147
GlyRC24yNKGZaQz8deflE3pQpocCM/5OHSqZcI8JdU2NL18JuZiFxxNsNIA6jPdB
9/sD3EIWZMIbxP2eCs3WjnK06Y96cMRCYYReT7xv+4cWVGt8IwdJ3ezxKKXfY7zq
cZ0jUnHUVK3nLSCGIqt/z2knzhFfrqB7tdx2X8Vv3Wn3ujeWlCSRG3jpE7OfUPKi
Zlbm/CSlT+eK6ZhjDKgPuz3bcgtNcyFYZh299IUxVCtjPs0TGVyCpsCKlET5yfS0
xkIN9zsEIaIBCh5ts4dNbOCizgWaaXmvaZ9F1f5gePP/JWH5igEuPKIDJ2jkZve4
CmVdzkMqvEnZnXgBHmxAQK6nTsUVXIE3ebRhYV6mB7WabH98ktUZ1E9ldOtEKpHw
bdVj5z8xCDSd093m0v6vqPM3nmK0s0Tm3dRjmp/RshWcjm+kegH4JUFgdDGQKH+4
voMIR9iDBbMZgeiMWLZvmir93bX+OYeDjJ98MW1pbrt73+b7AupbQnruT70t9Y+f
vU/m7FM7TcT67cOtIFE3ISM9OgRhWWLaRFhEmbXKiu8p6WjUYGZwCH4LCmU+KtgG
Lg0OoFj78AaZ52G2gqukiN2eTJdsLsRJsU4RDMVgbi4l9Yo2XtLD096COLn2zolE
AAgcI7P0Eiufw7MYYB7Ngl7O7SuR278iWA0l2za6LSu+0iHeK/OIUZdoQ1QuqUfH
GqgsssFbNNeZA45KTKReWvIzfrslgKOSJGmPGRwncgEFiyfCtCJSNegKb7HgIG1k
2yKfZ9oAT8LiLp7I3F9bfh2pm/OvL0BmXzpRsOSfhy7h2kTgCnby6q0f0u4dla+c
r+FJrBEpTHZgdM5iLu2+Dbt2fCFaGzvbrFiY27wu5bzRYuuq3NrsEtvOyiCc+toe
4aAj3oxRs6pfTHKHDnJqZQl02dSW+t1OeOy2eJQkS33T3q+B7CVkuvTTRrJ2goB3
WbxSa5HYpZZ/L7rU/OFs9A0o7i6Yucds6ysKnWUftT7zszf0EETisPZv8Zb5VBb0
A9pJmdVaJUR8AN63PDA8dU71/SOomKW1/bU6W6kwcdnH0NVOsTQm3UunVo462D3s
UZx2rmeW7c283sk/twTCr/k5JFKySk+zUsm2HvHMNqlKXmQvlZfK7tIoYdpffspG
67M1bFZscu4R/Jt//fI2JylEJlqYtcCfpJ6R29YeDSNui732ZadgTEy7v3qyp1xW
4BMRzWAEGHzkYi5UM8L8iOx/YWqN4byOJZFBcl89FVXbflq2sD2tqHNywBmGPXmV
kljUgXtJUfFE+ESGcyPvuES5gNj+ojTKj71bOyxiJiPsFBrKA7uHYmYmpFmcNVLm
TQJZeI8fRzqaNeb+LDLm1I9gJdt49+q+taC5OAzR9QvaaCNUN4ovD4aZ78lU5YoQ
9I2BYymqNBuRz4c9luZCGBMsDS1KCooq9A4HgLGGpuHHlaGSQR8gd0on/GIiex8B
IOAZti9GcWDafKv4kRy859Bns7UJva7jK4cjEGLm3Bodv+BRtgzUQa6QAmshxCJx
Lyc8CY/BsoFJ2eisNfrkTW/KRMI5WZTKKZwztqAKLU81chuZO3ZoBfZM21kyu3Ew
2aBRxOpxKl4p5TINy97QgN7QDLBHXODIWvy/EW9eSYEmxgeuRcLa2nRMZDYrOscC
mYh6IXrUbPxc56eOEvYXohJx4Iew5KzGwui6/+s2hOz5V8r1ro629urKiGyWBFDb
k8ejxAOjo7FbrmRCPE83Y/FTShlyRXcuyk/UpI6GC2HMw+5MAi7635UwPOPf6j8F
aRytgE2CvuPfNWiOb1pQ75vuzDGrcPO7vBNHt+YbNkyOtRzVkN7yZfZBBEsymFp4
Tc9M2p6YmYq+NkN6FvMJozEmGQPyoQcVXxffMP0eqqy6PfxU6eEcsvgQJDuYvD6I
MuPamsyZxblAl0aAZaRWVU7X8Hp+VEe8cQb2X69bKMfQ96P1tlHOpG5w6Td8FXIX
U/5is/djsyp4wQQoLDvOFw0OldaWTQNlr/dV9AySI5LDT8hq/TYL3P/qfzg4qW2r
N/m/X5unfUJi0Xyg8JQqLIpJ4/eszN5FBR5SnkIeat2yiEyJPGpdYtqDDkBW4686
D1AvC0r7HPVac+qxiYlu9N6A+JnMEx/SdfGFGrjlWu4bAdqOCv8mEttPQb7QFY/V
wgjHi90XnA20fdg1C77mpFuhYhpK8NxvnytYdJzJgzkBNwTGQI33Dd/Hr6OgAqkl
4ZUTrNKcjpfQF+c/B3iWEYMtz16YVu0anBdBjLDn9h6rlhP9ZrCz63O7dlN/Mb0B
aWEjtNCqn1DoH+r6QZhtBJ1v7r8WMUaqC6EvfN1W1JaLHWMVf+igufadASHAOSQt
3Yv9tGRINemNJXXKkWeWF+6o79OHNRi2giIuaEXKaoB4sshuY8uJX9P5/x2SPsoI
6W7v2NQ5XAh3GBmBFk8miOJ2O4daa5ct/NdcEHq80Oic8wcP1Y71+CxHB5kTggUe
i+vi5gxqzPaYdfsT/JDl6yfcNSEdAz2qmaSIUe8AKvV2kNSWmdwWbcLZNgVLhSJc
uUFLxmXNTAw56RH1O6v+29HNplO1zZAkbkVbR1McWfFhXy/C+NEsYyg8/GfXz71V
NkGqtnF8dzY11eixEuT0JUyzU+AM4mKvGWzfOUS9FTOzKuGP3DkuTeeSIrDRHnz/
5xRGAxymmAqoFVNIS1tsWZRfONL7c6qmajBaZzD/DInlWuaIDmOvV/V4NOZ04XDC
tb6Fz45qUoRUsIZ+Ouxz7H51Z32VgpWqmQdDtGERTrXGNp0IPLj2Q4oDWfytHqnY
o/Zrx7L09i9MXATY4+Fe7AsUDM/0S0LN1tj4aFfshwmHbBEtuniD3rGXCIXgIBlv
SNg298fIcL/0WQ04G5Oc3sZIZI67s2LvBVIosw9zx3xpqoO391/Suowe2+XaTOEM
YgTnWnt+2S/Hjs+3W//IIH34GUvVch//tdCnaktB8hqUkXSrY+2/q3W47ZF9AaAl
/aE8tYenhxxhgD2fMNySe4mCszSuwbp8mpfuy2kvd+9mP6N6i/wD8ThY3mklfJXG
oz1vhoGdoakBseAteiz8qU6Iw/CfqKuXCZP/j7xQNRfNUSGi8DxlnGJ1cZNE2GLY
t4Kz/S0HeAc1Jtl43Y2SIc4IHidGBjVLY0fxdqCZop04zKvQzIFbuuDeGfEKL3A6
nL58h4JAAaXB/Bx0p4h2L24KcM3O30bGkYaRFJuw2WoknsJM0+guolxhevxKj4c1
5pGyw1/UmSys4FZ3UrzW6/Mv0was3ABpFKJ0aQS8zD/xK90CSde5ZCPicDEKHWDD
vYK0dzirjZTqaCj+D6DMMJetvjxxkbM/0Dr4oWoLdPelUgsrM1DDQQyeYchhuOVP
L+kPsqmNPhWjCf+D1EKtg59MQFQS2tTKPRf2QoNE91OYyw/Ium4zMlgqHCk15gU7
hhPRuI34QW3JjiTjhJM+Ep91nNBOGxfE3JXrir6Rx2Wp3H1UUvTy8+kOjdpwLxKS
wAvQT9FZjJMZ6rrzNNodexy/ZxGcGzdEcCzvDSGoYc68xjMwRNAyEIxbA9HfrMcv
cks4A/2LcExqOKqaX/TRI5LL2v9ar2lpLbIdgiC9ujubuHiT/wVvzZbL3XbmGWGx
F5CC1NHj/YV4putXIntnB1G6/kB/9DJBfYRx8bnJ9JWULKTZ89dO155nYfSJmFuj
bcz3P+FoPAtCFDQy7W9scWQPKCwJCsQfBnDezvy0X4W2zsQ4fFzQ1gPscz3lRqhg
wLSjXh8wpEV+rNd+t2IRKCMxHxJ2xaaQuzmfj7UCc4Vfj2RJMTuYO+AJ3Nb6iG2L
qvD4oaGggFiXINMxpah2wX3ESFp2AkAkvRNWbta6QLVR6nn/HQIMns6KbQlzqJAL
9YP/9+to9c6s0bzv5qUuus8KTqHQYlEe3r6XxeOVhnIUznrb8F5QcKNTHbTABO/Y
fZHus1pGg/1iVgrQv/IYAE9Y6cymLeP0R1jFPSrTUaPcoAzow5cov1yUoZlucdvO
DimYGEFUbPA5AdYtEpyJZYtJUOAFz4EEKnIQWMVKUgukf/DMfm1rvUrsr14NWDHz
lSpg2BF7FVyd1ZWbsfVFemt5Syp9y6ScuA78upLFYpuqwUyiJGsVSdkoMNDzxLRm
KOPpMphmQpiLtuuymAO6Yys110OLFyrDHGJgme95n7+CheD0M4k+5Z9ScX6JNas1
d0cD4hXRkNCO6TBa0ivUgpc3Qkh6DEFItujbBkKAJMrsEx9/cQjmNEeBiYYaD+mS
KjsnkZL2oi3PkeOZG+/edznKCUSLmRHsYq+gNto0526B1k+tg4cdZQB8PIsQQwO9
cioMKYdaCg889Tk1mNIizsonPmRQPjrp3YH/HcPB5+uhNpVaPsxtRNRj5xbOyY3i
gNdAQC5dUbFtHm7nbliIOY6j2ReU5xlbxv3RT7CcEoYAmajq5ykx0zA+9dihTDGZ
4/ihtooTh7KInNt2Ue1BlZJJsIRangmaw/74k9cmskgESB2jVi2BpTml5aU+cFlB
wblAjJ34J0MjahR7M0CTjtnJYihTT/nUiEqiW+AfwwfgBKo7BcS0LbqTLD2RRxkw
LjDkgegQ6Kn3iP3HBn0Y2Oq6zYXLWjuarV/vNTkYbm2QDx6ChLA+XRWgBa2FFriC
GzMJ+A6+EsAuXi6POT+JsIlQNikLgNSWBQlT40a/67HbwYhLI9lSUguIzggSm15h
M0p1Rvy8eM05I8a5IG6N4hlRd7uCI0kUX7mbySh5YQulNU6Ab4zU5MUkyL0Z3MKC
7Ztdo5BXjeL5qoGBYTWAP0Ndz/aF9wIFUvfQsaLe5lYhNtOM/9w1VxWnDwQ4QLnq
zV/r93MTqhFHBi740ae50zuxDAsPpSnJXJDiGO7TdVzwweipKnIwQYu6PYwn2I1O
O+wIXktrwc8Jlo+1b4Wg0gI7Ig+n4xaTz35IT4HHmieqFU7aPwiu9DXufcA2luyN
EKdOWZsGazgqZzilmQCQzk6HGQkwlh2wM8fUFibrm6Ushy84BTxDMFmW6Texq4Tg
VEMdCaSvjsjtWUL5rOzCsqGXFvAnMUUBouPcUnn9+3cT2EASzfk4NeG/KhkQsUPf
FsMDMUvltEScKerohuUWNXodqDjCpyq8C30eInTjjwk8dierdDIhcTgFWb9ubpQ0
6RiJHCkAU4xAWDRdudFKAQbnHN8RCDlNJM9930xgEew2Tdm8fRBkE90GC4rAw3z7
NfnDt6RrL5Pfzr7O6zX805i0lJOThyKjU0fy3x+TOPuE8C/ZFO2A2femVakyUaiw
pMfhwQyEOP7BaKzoQ5v6dAGuc1xVzRrEA43lxYN/GCn2SK+EN1XYhhQUIUlbBT7l
jIU3Us1L6gUheOmmvbYlWldgTwupQUtmJczgnb/zdesTmBN/ET7Df6w2rxmQdJ8k
qIsB7rsxswbRmCmwyRLIBE/fRGnbFzRb1N1XJv9v5gq49x4SYsSBLsgzBH4f1eLW
UN/gkmvTgfnXQEjYdvAhs9U0CAEN0EJ9unk2LN7rtyJiBBV3KocNGGt9Gkkz9t4o
3aJvhlIZ7XqswK8ryZUvilQvjsjle0td53kBGxVzoqgENuQhxbo8t36WiwEI0ajp
vfH3D+GghRJRsKy9wNrNurNS0JlVMiNQ4/vbHPSJGm/ngcE1at4K8wu0Wn5u3bp8
idVTXqCcwIZAKfyE0Jy+Afl0BdqHVSAB2YPfo/7+6fqfrvOQfBF2T/ML4MqTh+Sq
ceCK5REC8afWWTJCfNDnw63WKIroGEsIpmSXdACW28CLGgtpbQUk/TQ3Sevq243F
dP0EccSxMeor5zCTedNg2Q1fbX4dzqqs0epBHY51U+knr84E0pui4Vhk3aTMMsAS
8kAjmRKSQAKjFj+UR0vEBsYaq99tDQnbEo9n1tITpGzGSUpvTGfl6qJ6AZuYRBzQ
ydfmo7UXSQ0wqLdMu6G0nWRPN2wIEYOQog8jh0vh8xB6u8VziPksD8Vfxz9IjS/q
j5AcmoKKpCxHySPMT7APvS6nVayf6Hjhz3Bi+NZX4rRGNU/D0ZrWehXj3xYqt4a1
UE+BW74YOx4qV3gzc2vnQb3udODnCUjiPlUChZV+1VZPNDG61dungBwm07Icq8Ab
p+zbpst2jM2skZJ9fx2JXv1QwTRK0iBbrRiKNrLzgPYVNpgh+12vG7JmHHFgD8bq
mcjx6GPQ3QEReKBbwWm6aKhvUv0jeMuGQBN0+3yEUMZVZ43Ak4FBdS8YMIAVUMHF
1TH45EDPy8rvtlDTTPvaQ+Cnac3ugIKvAkymx6dF3MwPomYSKcr7lwaCBTZnja2y
A8vjXVOcaBQCMkOcnk3PrRpi7XUTWgpskWS0+U5J5efpH9lVOCduenB4Sh6YP2bf
MwTwjJW2oAXO+d0AKimikZeM8Op6pDQOYYBtkW+FIBaUm5hNwwSqWOVTCmB5rsbp
UFipowakCUxAjkl/rJqSBGDJWPF8s0+9Mvymz0g/K0nWMU75qWyLvVR8U7zWZfE1
7dITOIeM+Mh5HeKfSfY7mX4gFG0Cfp3MQLR63ewN3KMkz2YtZL6S5j4jkppJBCQE
GhVNzkVd0MK9g7+bxZdGoZZvIp6b+MMmZDFu03ihYlOuzQeQ7BuZW4WoAMNZ23F4
hNpB0asFaxXSMd+uC/P3Y8JeEsoOizDt8lPfdr/izBUOQ3JU84/v3WABxzdh+/1w
6sF9Qh0k79MVKZ7zf/rNzIGd7RSVJU76PCmGxXIqxAW2k/awWMhFDFvQ3VkzhIZQ
u9rADDeQ0HM5eReY+fhYYGKlVMThUzYFUIu9fAEpVvLqfy/Xa2/nvn2yhosdY0RC
/qRPDYU3zbvzov5E7rillKBvLj1jjB/OvkogsYFSlNdMYPZcVeRcjW0oT9tSGm3W
ODCj6zU3fuv23r5DBTR+mrgio22C8BIfpdLXKgnBVkkiMmbpvgs1tsLBdzZx2ZcI
zPEePW1z7Yu0JOv1HL/ivIxIoKOsNu9KOU1wc7LfOLCqcnyD4Fg+pUyqMuMGFo4f
x+py5QPuaOSWUMkuNcM03T7ALYmsNdf9rzcZXClbo/BqPbmHpw41Juc7PoVDP+Rv
li4m1KYS0AD4yFlzuBT2KrRaDRXV61FUtC/Aa20klz8rbNuT36Ff5ygNVkcQ7k6O
ibZIdj/+55o6NDlHaGMbv4oaudlw8Nur/Y6o3a2PDsHmPYi+NplaS5tlZkVg7D5S
oQag7EyMkPbxY/h1oI4cNLrh0DWpoNn6GKxohnbLV9tryGgSxbfslheSu7qccg6U
we3rCDeQHICO03Oe5DxSAJ+rBBZTZQFHyCENfTj62M3YDj5joh/sGGJ4EHWIVDqG
i4kI0pKS2pZeFQAl45gwybvzhFttXJfcI67zOEqMB3EPuZSQNjYjzTHm25s9s8k2
GTkwvKyYMBMLdSUN87CIbHQImCRZcv7S9TOHqc4tSZpcc47jLCVArpCQ/ZiVSni5
dIPXmQaPdsbgi84TVb8bZb/A+LbIwxnE3cTdUc4huZH6t9cW9E3pWrEiOomdlPWB
qixMKok3WJNiVB3sQAUK8wJN8jQyAABRxy1nnENf2SAn5M/pFn1ohLvRv2JQ9v7R
ahuG5BpP3Mk0aR67QWRZNVpEj4nqAFtEeV1qlEUjnYcY3MCHgO7biVTi94gFLZ0d
wsr9KioD5OjEZSp06TOsgs2wsmHeWuZKIQ0m+LuNUnpS8ZZbX1i/WQr74sXFQugU
eT9yG0LzBR/Ir+bu3W5OV0x88+denYWhow6OKXUep5tNUUCf8ZuML9NLL6Be6zlL
kw85Ppiaxa0biPr1+yvstAeGwntXwwnPmmp0emeZ6v7FpcY1N6MdTBjmjBySa+Sg
jq6CKeDsyn3XjYy6swvTYdH9JWfgCnznm3kAW5L1BSj6uCNbvjqEveBIPICW9koC
H3e2Zs5OlkmkCqpOmJpw9kXfPROMM78ZRxXl4Ze9pZb1vqE/kUn5yQ/Lc6mf0tyb
CJBqgoJHBfBqvNwJlkSVjVITYi91cER5zqZRArgdavkYgb4wQP8+C+n5PjRXSUej
t8uUhzNNCLK8IIfLfsDCWELzR7d3QUDZzgACUCGdAYRs0f3HaEaFuRqbPRWllnYI
clheyG2mL77oefDovjYPQawc7t5/CTiLzSFm5rxvbvqQad6KTLRvxos3g4cgNjyd
x8kksDOOjCp6TatJSBcgHlSfR7zmgH+NEOKRZ5lP/v6fpK7hVJPe7UEHB08X/IVi
a7MBdgq+qFZRg2pLjebiFESVc1JlGuriAqjKobrhp0ZpIF/oU+1B/GR/xoobCtOI
kWI2ycoDMKzgpH6hzoYq99R6647bLsmtLAFmY2gEKCZznTmL8hymVFH06UHOtz1o
g57MsZZBfu49jZIhbCyF5auU3ri0eF3hqQCiL65Bn/82RfYTtlC3AQO7xKTC5/gE
IlkxRR0pHJ+kzVD1e70EgcvpMrsSCEsJ5mqHQ3BU+xtTHmk0rZM4Nolr8Jvarykt
kl5FcqQ5LykidjgJuU20i4BYrr7VSkjDYktHUDw6KxRA/uYElgAJvWeD0t4mMuJ4
1wXLLAiACSUoMVVbgudtxWgQ0oB/LFin2MwVjZNTBpQLPkJy5llqooZavsfJPWbT
1hHzzX92ItiQTSGbGxiVlT/emPKiAZ92xnIUvqEclXRvJ6zUfjzT7iqh6MzQaNsC
lkdOj7nHKbSHj1XD8yFRyFr2VJ8FnZqKVnmSG7dRSdNU3huLWwiFqH/KfNoXvw2h
5AwtFTjHeHmhDXtmw6pwrEBluE/xycvxCSAJBAZDbWuAREwqjO6+bbW6zzIEF3B6
KG43rXwafd6S9lsvXFnErVJQFIXWfz+lvt4PsGFmoT4+cgI2TgpAmgM2VSLWcs3I
Oq1la5XLixiM0jwDW6ccCZSADhKwyzFQ/Nm+MHtEfyR+Gak3+IVXCx1RkuhMDvnF
dSB0JyKHiOWY+iUIXXv4wYEYIn9frkbeWaCYmgR0QdMj2iLkv/LPhJV1muQixQR3
qb65CISb5mzFxGkrWIn2ZxDlLQ2yqtpg+Alv5bXvLBxqalIHFav1VMcfOEu/pHzH
J8E7KJ6cwOo/Yj/DZxjjGt38zzdhT6mu8z+C/EDJkAKuNOojpqHOx7Q0lKK9rYVI
XvNjvh98iushXmCVYyuckPsy50YeX/yfmyGo5eahYogHhqKirZOtbLEkiujICW4m
JSVT373ykptxQ/AGXd8uEj9YBJZf2JODPMv0ouRWKsXmYBIcyaM/xOMDjMLM0aWg
o+gwYL5wCDD32zL6+sfOU2AgjD/s3Okdgjj3nWSBC2ncvhnQ0jLWJgY+thYTBTBc
LpPjtI45Hp2YrNm4RAU1eMWTXMeEYIg6fb9YFSNvLwX6W8aKMDZ6JabEY9u6fgue
0Vs8zlnyXuC9FjnanJEC8JUW3uTVIYjncPCHZ7OdbwD4eEr1hgwcSsZtBK/2kEbr
UZ/Fw6UNctRLn39HUvUeHv0/uqomiJGBfOGvRw+3hFNvERWDCpn67ENRMyROrAQF
Us+XSrrIHKeAvVIn6V+AdfGSs/YCzDFnsT/9tnOAoImVNYPTDyDSgZcn20a0kQJt
BbeNczS9GN2jXmhPi2z8vOaTKlows4Eh0T7Di2HzWWUoGPdfC2TYvNKfcDslPjbx
hFEMIwkSBnSr2VEqA+NwTUIfRjwnliV2wECC3VfotJEubuHm7xM+WOM9GOO0Q2Lz
qIkP4lif1THwM9xvuCCC1sCZ+3aNQu1iHceU/6B5ALxjHHiZMW+2DmLwLO/3UGL6
EUJ/3DAH4BMoSmLLGtQR4p21Sd3o0r/nzP47KNOIc4y+N4Y1tSSt4rAu77i8eVSD
e3QSABIAFbxfQnIFaP9w+35JHUymHYWZIBPWxtWL/nR0GwXROg3dDHOjXZprCp3I
cPA/eFOsTH2alRm1RFqeyIMYS8f488xi2rqqdDMeCRxt0w0N754m2fu3abNlhbvM
anAr2TuVFyLTVH/E/kwmLkorPGshWcYLlhsR39/cnlGRHb63o4JvujaDxqbOFFXg
0NIFsXw7ohSqasDHgAWGHFGhM6yUPo4FtSjHzWrM9shAhKewWYHfYWMpRu+dEkH7
QBhIySiHMx0iTnzgEAyj84Nv00zKnZIZ9lO2x1+0eJdFnLEc8mcx/S3i40jy+gVN
o5fI5IqDvMjwSh4Be0ofh2C3xVM9HN2hggeh6iqvvtNlSdFKdrN4hCz8XOqfzZ4U
bWCUwD89JIvzl13QIYaqOKXlqQ0w49DHFy4d0zNDYmzxx4dfHwRnpea9IT3KZh6e
U6AjUPS3iBkaG7Rff8rxXxoiw/DW2vw87LMTDjOtqdWLAF/P+ixI+Ss0tMzgKQkG
kBPy3UDJnEFUAeNxQri6N5xqA23j7pVvDoYCgtktcZJ2Q0Vt1DjipyzS1b9kFeGk
XV7KObkFWevJUJgpqWHZhHsnMhYClVWlSc4M3WZaPgP3VyAj5xH1+e/qGkpNBbIZ
tUpNiaYRTF6xMC/9w7AYaGgTcyttGwvVf/5hVJFdyA8lah4kR1INGkVPght8Q1bX
TCSKYBnvTO05DvyjC9ZOWF4Dn/Mh+KSkbQPXX0a4vzhiAPoASixXZaRE71RBJpfI
TmlqSlUdkOchTmlpINmrfY30J1yNLh3mEEJ1L/+j0DwAb1EPa9kWYo/glpZ7kPKw
tVevf2acNk57oAqHJg357Lqs0Uem131MaTxq/839adrPNEo2BYNvMCQqzqmXGMBT
P7nb3rD8s+woEwmZ3GUaJbPpzdqOQMUkkI3R536ncUBwYPm1u32CmmLbHp1FiFIM
MUGD4vjRKOZ8BET2pkjcV/rTwVaBPapefENIBgTswFr/SGqbDLwLbZ+4z3mQXASX
SzJp4Xb96tZhluIPRc1LLUUzE1UoWmqNrmthKbVg08K02e0UnwwOoJiT7G5sPN97
7DMza4fqtUrdKj29exIh4LROasf4pPvxdC6cevRFNdtaUm3ytsBQgy0G9rjIWv4X
XvN8mZOgmEcBn9UT1p5rh4fJ9CnC2TJ84RZKOpsCzcoOjR4wS/TZs7A8C1IlMg+1
dKOpgkDusU5Mx0wou3QjdxHA3KRUZbshGWJuEUNd8wuRNZw8TVjhi5tqQZDc5yiB
rzw2e5WkAsy5pXcAnuT4diqfcilSz1Tmb/mWb/CByPtt7twEImEwTAQUh0Dz5/4C
3gOxQLf02WG8JXp6I/QG43xlKeWcEov3Fvb6ctNpmAVILnvZYWAeihwaIQke1kO3
XeiyuPRHGQeFPLzC96MKTpzj9kPCe9ryLWpAdu9p35oEYqhYY90zE8VOk3kbbwWn
HPaTO0y4FRrwbZrO0FHDQMlhJXX2t4ev3N+ORE0jvivmHPm72P3aA0ITulO5lcRo
SV/Bkc2PFJO83pECP18sV8vJbVCNfNHdjL0xnaDZOPVn5WHayoBejJ+nmzk9Dv36
WWyuEJwgrOl56FC6ZG8EiurOw6i7kbNLYtSJ+cisLNNqVw51IOLgBKhFG/lp0AHj
taGFikYdyCuKEvHqjGdOCNg/gqSgfAYQtwHy5YXgjfTZodM4jcUtzobPV8qM+IMB
Zp7IIk3hn+OyywRQUDKkEku/jnGuaaUS0FIHWxM9Z2dCVjOCJTuAbc8F3SJQlFrp
uW64jOy6Cn5ETIVX0SODDPAXqSfeU9mSByEb7E9j7r/eNNLxP/tZH5ZI3Z5jG1w0
zubroAWhAocbDCvdc1dt5uhcw3p6vS/YHa0XCE9NJ7cpNKYOcmgII84CVlbRBjWz
d0UF3avu3lMtHRtAloWdcMVfTP790g+LTZzUJEVmJpUaFJZXqIVaB763/fMc5FuO
oT5okgebqxqYF3/XmnL9AmWaFZDTZxiazvfis+ahTkPU+BsBoqkFoM9VhzUPHsMG
sjZyn2zNF3a7kfGKIfQDm7yRaENO2TtXorR/GO1VPaKSfE7jMaM2iPI1UFJqx7pC
dqQXp9591J8/WiQ/buwxrgnwcc/Xxr0n8V30a3PvHO7l7wI1vN7X9k6+ZfuwF9+R
2IJnV6IbFKOzTzn0irtV4FaLbDfdbb36nLrcOg2uxc3BXCn6jVVavxL8UDaToVnN
dEQ9uSu90Ac9ie1kHYAHZceOiMs+c6EhVUK0eoldJoix4bhf2EJmtzOc3Q7O3IiB
lnIBpZfR9cxkiXrz6w9ON1slCspJeXKlTOe/S8lQLythVY9k24+vpXhGLOQ/c5vc
3uumiAboMnE959aV47vg2D8O6hNlHRdLZfE1HNN3Ljl/ZXFbjHG0VlTpNYVSJB/y
aDOKpYm5oYVnSEpykqyWptNL5P816CKoYHbLANLlObkIRP1c1PmECBrKa8Hyg4SJ
EPhtgtGw0saedVmIU34Tdqrd1X5yJf3B0PHqatEoMn5D26asLQy25BkJdnhRvCp0
LQWzxqKG+3NC1JzGgLSRuSIK4vvexAXMAnSwPs+8zj65lKY4cdrGTmXclEeXO2EF
fTG4amm3Mp9Dingw6KNFRVp9cilXiTvUMRVCxKy6qplq41EZcFo/tLhO7dy6yEdy
Y5FEwhygdOigfklJivviuR3cVVyKs0UAIHWM5SOKpPGaApqpN4ZHRRm/mGaAuX4/
OIjS/2RQw1rrtFR9IkZJyp96XcvGPXJlyykKYupzC3Eio2BRiD4a2enmMdC1s1hS
KRho1sZrnq1giOrBWfagu/S9MsTRPt0Bfppd6JbDm0ctSEBJAMdPTxCjgnHwuzpy
27KA6EasFp6LHy+D8YrpyEAyF59Fri9ZyLDM3OojVbnUZU7qAuvjJ+C2sI1rmUTY
ixhDptEH2UJn2BZ9SsEJS76fsLVv/QYbXSyqZDf0PmbWKN20jx8JIpifGx5GQUva
0u+NcYyLiUA19HjkU1Bh2zvKlh7mv6GjLNp04PlswGIzoImixDTrv/UfRCsTzOh4
r2IJnd0ZUE9kwksiIoLSDHVL/m1oPdKn0w7M6LF3Otff0jptBijf/m5JcT9QiIu/
BkasRQjeDnbeygFWz4V7na6BqiqrJh2KQud9ru+13an6gJOQRoY4qgKj1RGT4+mh
Tp6NYNAuky8idqWr9DlpAKym58ffpUSVT8aFDwXmiP/OiWiIdK6+suW8rTOBN8Wd
sX1E6MRLQpFWkIXQpNpHN5z9l8CW5wCJ/rqTbKycCoeb2pi2pW1qNeTXRoumpXcG
RdD4+HAPza5vMogGFEW/XFulDe00dt6wTu249mry9ZcBmDW4O6aIdUl+rD4bLNOt
ReJCoIZwn8jtLTZmSMD8YELTiPzdqo4QnULu1Pf+FXDo6lat6V9y09lejG7qt2Sg
R4eVz4l8x1YhWplsK56clWuqzF8Om/8znvgGPmW25pAM7vne1U3m7LvaE9mlY82P
wB5EohpyQy8vQUmoi2UAE1kx0nL4qwhCfpvc34pzZekYxHAoFzaAcfDIQDqg+aBu
odg0x5VMvg3refKQGVmuAQVNg4lfrJ5RWxby5NfDYBPgDC/yFLV4fKd9IsiB2Tpo
G4kAtXJYz/XsCPBXu801I93IB4QWh+x0GMDBhJH6zoRJ5i2hUrytLvZCZH8hQAYd
RB1MK3xOEa4iroe7+q0rQDs+H2BDmZMx2Sy5OfrtHu9FYyn+olN6ywhcb1VOGZQV
fz3p+FJeMqjz2SKSsX+eveK0R0ctXpFnqeR5mG8bMD7M8PmLNm+E6Bd9M9uijepg
4FlFt3nCI+psBbxcMdCTmgRC54Rd0Dtr3fSufeTT5nlV/n5VCWKUac24KgwPm3V2
/NsJaXK7/VadAlHApCQEnSAxAbQ3pmceBUektiCgVNf5axKzsNmYmkefyMn52yb5
4j1D0DJoYU7MY2VZgHtLbGOXRZteuDqWgLYbqjF8C/VF89Yk7ddjaXyqYS9j8KOA
Q6zu6x/GvrVgjX7JnVN7801B/5PYVwIGvbYVcheEMTsgcX0qR54OMg4wkF2mJkXi
TN35IJfOI/wSJuCZXPyOJFCUJX4SwdbeOaJvCDUSeRhDRx4DuXQX00tVuD+YlglZ
+gRn0QX9LJht7+olaCM5iMgv+Vs5xv2erHPbbEkWoOSLsoyZVnRpamxLf6wc5h41
nRf8jt9a/igOke+UwRIh4SR+MhdsAAEn+I92joLEsESgny8ej+K2TCQFTww25mBy
7fPCRmpW5WEt7OQSC0O9H45lyyP4pmTIhW1Pn9n3BGkHRLodNWbKGFxPTaTeSsAo
AlhyDkJZ/6dnmJc98TPF8qI9UGbEUrtiKva6JbaPi6AfmRJxGhtD4oRXRr01r63b
4Sia9Icwm/KDf6J/PL8BGpiPRYv1hGH0Ty6re9HM93nfrzC9DUc1XXdt4SKwUj05
S7sWk2uujhc1osImt30K29Up8D7wZYDM27VrDvaY2SiTOjHY+J8msjvVRIaYk8Y/
X2xHjHsj89vQOnCGZ1bHfC6LO0r/T+nEXU4bwprEbTNmygPTZkrSPXWsYsMpDngW
jFreZutiStZpWTf2CZ8VX2oYEExXEmOxIiO+2lC7qWSQFowKhNidWwfDHx3w2xWm
lT036jbUfCobf+kItWGffa1Wbt2h1VYVbFYebdxhj2LL74OhHutG0DZLkobd78X4
UBSPLgGkQui0yilx1mf5fLg+4242FT2i5G/fSQpSncjNkrOgRF3Fj+f6N+6s9GjX
aKrKGUswXBql9CKSMdBYmjhxDviI2mpxDV+sddJPERXkTIdLNGy5hyAZGdav72FO
b7jJeOyNmnGKdUvyeSEda0D5lMHurFAwhZ6AZzTmUCPvobQ4PEo2QSKZpPDn7aPM
wds9BS0jEb5uiTjziwEatMi50YePWTaBbSDAl/sjggd81eXAP1I1GdJrIqWZtnWO
6oZ6z/FzC+p1gIwgpKhz+2rnMQ36MLHPkng15B6Nbvhgu/4VIe9LUGDvhk4EFXbC
FsFaGsCAfCCiSg39WUM/GFBlkJVCjMjmuR3/9RztkycKTdw6sXMLwiuoquHfEj5B
EoFZKkGT2oaOWlWJLmp1ZTGorcXhlO3GS2/pl/+4gG+hNk6lCB3jJvdZtFiY1dRb
FSErMQ4Q4TckkbUcsJfRzckEFXHPPV7w5oz7RcIgRPQIhp3IJUpDqVw2hzgbG+ql
7/SoEg+6J7a+J/4fHH/O51Bz/OVSIoy+87Wxjq4C6678iQo6d8MrZf8rPj5OGvIj
C18Ss31rBWAlfNJSaV6KS1hEjhxD0OVRN6CDPysfF6SLYlm0QPZ9s7QJlCbx/K0u
zGL68zrAqBoTKNVO6Y1j6B5rMAJq84DIrhF0w7ynSKulnjMOyhzZNogqYjsHQiRa
2jKuYgQHUt5q9rK/7FtYO3fSK9T2VBpwUqwleo7L9icn4xj/Lp5d7V+QbjeqQERQ
v+xekmKGRMagDfP0r7uqnKF4UtKwO6xAbRhrIiP1pNcUfH+QZyjAqmCd8n4+pNu6
kjVmwIM7wr5fgJaKWXuH8wt2HVxLjZNy4FZbRYlSKANxDKjGIViO6UGNomy1XQJr
Lw/5+F4FjSrkqml3qcnm2yPKVDT2TeFLYAlK2csjEv6ADVz33iisH8MkZvbY63vB
R2IOk3qZ/3gsJ+aeEW7XTgO0UZx2R4I0Hf3JSzYIHvaqAWJvMKiQTWwGcG4OegF3
PNPuXsQTk2q0J/LJZgVpmIgbXy7x76D3B/AUCGXEZNIncYpsJxxZbaCR8qLBuRuf
H7o5GRY+KnGgg78MXs/T84qXbLLdXXTNoncR1b3nWLupjhjkwVL/RrNznc10pZGj
TUz+rt60jSMDean/MyJC8lk6d3DKsZs5I3VMkpgyr9Bg5ni1Z8fCzmWOlNuo5WlJ
C2easYO1fDTlYr2ydGLirHeMPJkZrQUvuRwP4kp+u1loMbn/PJPCrI2WwbSelh0O
iMXgRF/cHYTMDLenyVWk+lRExRPp6dXlrF2wIqtB5q5azTIpNeWpEJHondfk0WNL
XGXjImzovBy6RPdJwefOHjlksm0mzh6KYf1iFI6R+3myfBDEG809hzgV6n/IilJx
iBukCs7VMwqxXzHArC1baJ3pvuBCMQaCqmIubwOEeFq0c5sUEtCENKR+ZrwNuf1Y
KFcbkI/7s8JGDfEEQsdTIAP7aT+dgqcrnlJk1GtGZASKr+IbrYW1C79en6X/wxlr
HQ43fc/Qj6Bz6j/QS9Ami188LFmj2fLCsfPnOK4PNhOk9vRytsVk6jJmsovF34zp
HT+nd5NWS7Uf9pIQQ8FAdrMsiX3NEgi/bkxldFSVdAPEbUiiuaCpQ5b30aD/EAQe
oEZpxv1OFbqn5BZTs4kpdBQ4wcqhK4FsRAu+eyqolh4X9UEYrcVP7NRLvk83iHHx
1JmEPSeNPd0tUZVTAZkLfel2zd8NVg+T+ohYhtpnOFP6ka2NItXOVFLCsDPNCjkb
qKxKnYLckxlHyYhX4xUxlk7zxBVFk79t6yAMZcbyLxktA6JN8IdE1tzjgLEh4zot
VVwogtjVoG68YvkICnU6puI+QH8WBRbM4GIBE4h8DLiUWC8l0xnOyGwJXGx/s/y0
7/snrjlMzai5SLDzdho4eRAwkRlqt3uIYhl1D2T3w+tghEV10rKL/RumfN8P79at
rw+pN+0gL1CdpfKPrVEpQllEYWRS606+lgSP+hohkK+fxF6nVwn4wn1ZcpffnDTL
L3bDhKzSVvI3DlimCKckS8YIB0aMDwJRWVG/QOh8BLt5OeTj3YQD7Yf7VuVjQetT
uG1oBjlArjHNsjpPuiGIwL+MQxBkKTs4xkOdFVf+40DX+ml4OhkYwa+em5XT9488
inefglTnl+5aF8RbWaW0hHdUaSMmd1tGncRwE5Rdlp9cnAIXryaI9HlTatg/F5ia
PZr3o65Zq8O123wLvzAevB5BL2Gur2kUAtgd9A6xiFWnHr33KqDiQ0lg/0a+L3Zh
PvzsA7eYI+1nvGfxfbG1pcGzoqWDLvjFCKCHXgC6gPCSr+4ZSJcjsid12cQYW9JW
PR86dSCYhe8L0a/5DCBw1e/WNQvVghV2cLea6FIEWT5HnTiMyV9RrzvC8gbcgKQM
4e0tsOP1y+qD7f1rdlYuvQHPXadaC0NiEuXRtwFbCX0zN6hqftXtm8ItGRESW13e
mgk7Y7hmrifXus5Be9IL+apnBEYtiHjXTYePZFeUIwh6z2DXQ+REoTq0HU62rUj7
ybJAIX5vpEyMzVpqcqPNLKKL2ZhTka6AsVCIU0jfoejMykPyCgYGsower0FTYgj4
AuCA9AmKPtYvCFghE1I206JTzjM1fzOvrR/odeRt+Wfr0npcJB2OQ2XTjrVaxYRO
UdG/cTgzGK0jNk0lcXuhEAphPonJIN8TfNRfObRWMDk/xi7LmCXnb/OT60CL9WaR
VlsXL/aGfsHf2UYQ3SiTQz60Kq8Jj3B4Z4YohrjsdUDrKDKCYYEHGBmY1JzbYpAp
SP+Kj7+/Fb36Q4EspXYfMn3jCSMvtAaGyXwoBKYUhKyPi77y8BMS8cxtwRHgu/r+
yrIZESW9gdeSj00DmIZbaazGbuNuEVblHZ/KUI9f81w0csCtxZy6dVpf9mukFCZw
Jk1EpVr5INzxrWtRuTMRzUjHb21s2VaSWFWAxyyLJvKG2K4Jd7kwIfW3AmykoRID
pN3IXaQJ88lpvF/d9MmbLIdSH62ANM2nJtpnX3xigQ/Cmxnt3rXa2y3impsdKX3h
TZilYgKx1n9sZxyZ3nFo8hBMOBKzoF/k4EcAeipiqG6ip9Pu/VnmrMUAp66IryLu
moTSV5s4KUOMTl4zeSwVHHMyZN/qu2XR7qTphacyqTGq5uc+d8nw4fe1HQVeoGD1
HQ9NV2BcJ91MaYN/8srfYX9DH6ozVPdwE9MB7VTYiFJSJAbyPacxq+IxRae9g3fj
p3l6UBFYCcLOQ9cVrK3U+vjGol/T97CYPSXOUjDxsqmnGap8GGuWI6usruR7vDN8
gBjN2HxuvaPP+A9x8k8BjfyIe8h+cO/+pH/QiLN2OOSAErLXe0fNX/2pw5XfCMVo
Y0JKrkpmTYxAtQzMkqXgIc1iU4FYdtN38oDRmiDM+ov3KSdyOgpEnMH4assSQ4nc
fM8UdU1Wy8P59Gj+lwEXoNznxlBqdgaFXiR1+dA6B90p/jnrLeYNE0dcTC31HOsV
9uBzKNPbhDmmyWf9Ai383ms0/QoMfq77xSmqZo1JUMOtd58tzCPHmzgdAKlxNnQt
OswvqFD+v5wm7/NQ39IaM1ewf99OaUCOwovdL5iTPz3HJPC82wdPMjMh9f60ZHqI
bMc5yTmuKkzqbeRPl5gC6PTU9Q8PpNLr4LVbaXkrtiRuRtCzi9oc9ONxk53qygs9
GYIztK+E+NLC0wuvigtrUXQbKo+/0dcvGlCY5B7YMdLwc4rjAlL7UVwBpjII34Am
aax1AdXgMAzMhtguylW4w01zb5NStBXjKdH/ezdq4wAbukHJlbkBd+9E56PG82es
/je0XSnWo2Eog0hrDu9/xgvOYTt5MM5gl6ny3AUl2iUwFVpMZzvZgBJJlRMEbZCs
c2I0CmokVQvS/JXwzrgIp0r1a/CUx2KXF6EIc/x8E/lrAUL/74bRPQcwQoYadVDk
wWyaEc4DgnZIjV3VDePMn9ItYzpCQw2+zMNKVxXRcdVDWfrrxFyJ5d93U2YpZtfd
lb+xad9VvkRHMsRPkoD6MmnLDyreKwuukJWUhHKfmTT/58bDIyh8EeRzbzj6uCDW
qit5A465S5L1lTutb4gb1LZGpL8J0l0AZra0RhNoLB8Itv39Z1tUXroZCmvU6ruP
lWhz05hvqZa48GowApjkBJhte/WEFNt6bWWSWFVGYa6WmA5zCVbLV7c5PbJxzm53
rG0PQwMHfvYjSYagVtBJsuSrAxeJtO0z+E3Rk2Ew2S6d7tvus/07LbcFOC+AEF4r
q7WFZx2fCnMRBv/L81JXbkbRwfeILqMN2DFjUjRGeudRKJCgrlEi93C70PESOYeT
3g2tSTZaSZtTbXByM4K/PzNXg8qe753LdhtE3NB0ccS3fg1cE2i4p5hw799os5ns
4p7pdFCxp1sBkkydpMyrI0NxOLJs6gG2djiOybQax3cFuyCyN0mV4fmB9DHhnboO
jT6TJSr52KXsEmbN1f12i0m0FRH6CrJJuWCwcmFA6oAdk0a8pWWJmVhG06dIWG+w
tHt7B2xURsBVCTbd4g7gj5Vc7ZbicFJcKzb1I8VL+qzjWsmPjuXpayB4TBxKG1FS
j2RuZWv+5cRl6e5HIy4yj9XUoHTFenaXJXli2jt8gYuUru2QEbLB5WZB5eKsn/f2
rerIJCn66LR6xQXED7/ecL6vzx1pPcCEVLu99klskUyhypHR4M1tIRfGd1v9Bceg
b3eCkDgcYP6U5QFaEZbTpsqp4UqYfzsZnm/q9/KsYXlZqE0jc+doJdBMtLdNNnt1
an8s1CEBpfR6oL8RBCL/d+ZIRGRocHnJ6laZlpR7LrbfwD83iM7AHXIohSsk9PYL
UF5D37qQG+3dBnMj28h7sRvfR+Ij9+wWfBSC4Ba/ud/xFfICxTXWkd8DvcC/dZH4
G8YrfHKcUssVatDpgphlapKtKHAlBjNpho3+ZNDyTv9vhkew3yJQiGZT0IEbg5+C
TWqoBuOsAQxva92BLi74waM6zUtQ+9gjCRISMphleECUpZIcsT0zikoJBopfeu4V
/XqSXcFnvzV3sP6KoptGfXKYh2kgFIXrCs1ZTQc2JDHGR66xLg8oZf3NxZJW8jXl
bO719X/wDhhW6ctAbWogJVLTkjYS83xTQ2NpV7xrU+7LMOhEYCUyoqTOabjj6g3Z
wRpbBhSm3/JzQL784oz27eoVi689yHRoDkiqfvwPdUK+XhWG9jRcYZYwoEv7XpQf
L6Nx9yzI6lE5MYBH3rTsOh1L9obygIYqi2JuZ4PbAt8hQqEn2q3ay7ouH31W5+vp
siN6WfPPUDUdw3/u+ALiNNvFaPj53h4yeTRoviAQgTeaqm8oD3D8NnSz43F1MEs2
daM0ULVvoZ9wz7BRaXqeSMNw6m7k8qGtX2oTBQzKSTuvgUQaIh3HzilIhM3lyjCy
jH0YWbsyQwPygpXZDL6wY0pGbluKZisrtz8dlycXA5YbSUTO6h9VrMkjIHD5mSy9
4zEbUXGUGQYLmFAqvRSwE/9h2uHZ/CAk/gfat09invhZ7X/CGO8TFcUH7mE9DDLF
UxsmNyEqLNh1hfIgeuATmR4z+Q10RvELBSDXOVxL/pA5ilo73p9PCaAn+2Og7LYT
Nn/Me7HD8kUf/XXlQ7WNrooOHA9jLtstbljZl4uPrdallndPMYtK3C1cAC0yyGEN
xWn0/nOduVu1hc5a50Pfkohyi4Wu5TYOX5O2zm9kZ4Fuq+NdptVaheVLrGoeYVeo
cjDNJniQYG1sQsJNEefFEXMko3zpnn4Yr22xPLazwWnOVcRnIM/om8t2CwaLqYJT
jejQbaVY3qG0VHVdkrwAe6LYYzBPeLnl/QyzfZ4+YvgWGzVLQ+st6D5Gyr1ohxHm
9tk5hw1chxqgj4L9LiFAUyBaxw5eqzFBZ2z10mF7POZ9BzzQlmk/hv2dKQM1+V7C
R3ZlSZ2Yba5gmKesqRnvtVw0BdH4wex5e0dEbqy0faUWQppsYP1w+dDm6uZMqMEf
LQtS2k/xRiaUKyqL9mQzWOngkQ7Ve3Q9yPcKgnQhCVK0dJlFEGPxEfFePX68q1mn
8DM0Jwtke/leIC9z4UwWXTkttH1CxxssLQSxYEVZ75AMsvPI2+ZCZMbkOE17hAL3
3MyXJzfVk7nbAyJ+zhLut9CvDSjMzv4gYriNTSACg7Ty1mwfGOFtOoLqO506rBZB
ynzQuXLBuv4lP3FCkKBQ2nU6WvDIARgbtly86etd457yD9QBg1nz5iIHZ/Dy2GeV
zybrB8TowflU/twb7iZHD6IVTkCH8OBC2y/D9Qq1AnFN74oF7JZUd3zyfRasxDnm
npJHznrUj9eLy2EYPQhyWmYkiMqtq6vDlxMU/EQVzco5rUyWKNMM0v4L5GDAO+G7
+lp9VjrxeDeFsxvhkXPEq+5EL3KOMrYoPrZLRwnZ91R6WO0u2obyn2tmQLYBaWEE
Mn4sp10XMH8TS8S+iybKI3r7FFKnXz7ruSvJzrrDosWtVlNAlOEdxqLgq6BBCVNy
SJYI7EElUUXcBz7sL9uukX4Io9dCWNrirJY5HOjkxvksaiBf2PoMMnJO3bBbfnSU
j4KyNE5l//s8xZ+GmZ9GDa95ARkVaMhUUKiHe3rRTpzUAJrjfwPjA8ulSM+nv2Tx
NTTYvmXKq5yfoio4IPkDZif5DcLxgpkUuWPAotJbiqtp7ojOAZNH2QNTyV0sI3R0
dWq60aT0peMzzmSYaO1vzrw/jQ14wGTig9ikDSVNm/omQ/T2VOtUGqwng+wLUzA3
5Ka9F/v5PZC8/JouLH2bhqAl/bQRjnQiYTChjq/M9fRE+2AJ5ROsXCOHdubDWwyo
UAP6+rvmNq1XM1E6z3fRl/y7XGW3hqaaw5iWbnS29aI4QCkCK20hyRJAdcF7tSem
2sMvN7reD44FfdqhJbHAAUROfpr5huoB5obaH/f5w6Zj5g8x1TWaiLzfELbsOrxx
XwzPMxo0hrRsbLPABdHnDTRQrZDnVd0rmfcd2yT0z9W0Rk02G+Yzuts54SLQynGh
J0mVpDp8Cb3rpPtiTctTi/luBPeoB0aoNGOn94qzqua/dSWxOA8kMS07RT6Pg5Ku
V0LZ6+6BjCGY5j6pHmmJFrOiSjjgZNOodWDbKnUh6EpgOxEbrOIQl5l0KXu4M/Po
NQULXf5azo86rEYVlvEV1KwSsycCxEzx/Nea1jtO+l2arQAcupZDguCqlhQ6U/QG
/8iZT9YmEUzwh8nJxZ1Yoh1OVBqyaRJdyuFm6w0m3dCdIpr4Y5kQ9hNSRhF9rqLA
KKDKCcBJGNIep7k8TvScjzYMUK3yHBtKxbidIvPAxsuL5A2/R0QUuhHCir4RBSk3
ZluCSyyLJHUqcSUZ8sR2ZKb+sm2mEZKGvLFGg430wWcUDLZtFZdO4V62SEdSh3X8
HhXdRblTjq5dsVbCwbeZnLJ5s/KohChU5t9qQvhF4XZefuOtxfWQU1tSODHjERQw
vI/5m/RVUiHgzjj09NYjhsp9iNxeB79lhmEg3MGPs0O8E1W1kGUHZf9MstSxR2bO
HVztuvde9Ykx6U2txZHfuG4bciE48beyDV0FdaHtnOYV6sidY29Qq7PGjBm/dbAG
vo8fj8TjqtnZZwL6YgX8fwDBiollK/uvbnpCG4CcB9L0gRMT3vIeiedyM2rlINK6
hpF1nsaVI6xr6n7AtWwVkM4IdFXnul7cFOmXj6XvgrxBeMhbzHNPB5t2011dLX7P
9XadQa6s0F3JE8d4ZgduC1A+4b/3b0cn1o+BOQBIBJrRTOi0AHGK5gkrE4rI73JD
jROtk+HhIiGQ2Pfnt+lyfoDV6UbmdJ5Y/y+bxUrUHyDrOYx8SCPUWTfASTZ/IwFt
6w6pux/nqg/dE9WlNFg2zQZ+N7CeVimW2QNLZZdXOMlHyEYu5KNALRq/Tflyx7iZ
w5Wl7MFDKc6nKgAcolCKeVNkUoTlBzQEAktubuD49rfERyD/1YVOUk7JOqlxaBAE
8satfH+Oj/uhnMXc/NK0nMMt90POUXlaX5j6iJx8WEObNHhk1NQKcr+jL5y1QFxA
GpGlfIIVoP+/oHwEaZKMEtCNjP65GiNAjH58KeMN8Dz8u+ZZSzAEXSjBxUSHhyVw
xn/dmuQ2YdOMojXRNJAIHO6y2soh5V+9NSypjQBTIbVUQHBGlY8dlYQ1/1iBuPpH
EkOQ6d+aBEF432GZSgIBBGiJU3yGGpasLy0sVU1Yt7yB0GzTxItK0BGGZVTsZLjs
c+5eytEf3CQ7cRfqffh3rlx14WYoK/0hLSD3N9GGAN1w1Fg/8J6cwF4ZfcHnJRXI
58tiNsbUCnzMuzm/eWVlK8jbsnCUvPzHv6u40ayvlRPKnXBG8qDHzxqty7mCHhwL
bXt0MGKRpA5dLMDL0RMH7AZriw3mLl2kUBF4trMdVGU8eeALBPAb3MNlFpuwaDbq
lkFa1hCwPf2CmIyK8oTe9AzNrBGUyKmCgU43FtgFZo6WE376AKfNTVnzHrblWOya
x8bidr4HqsAHsw3BTZYw+hVG5ciZ9Tmzr5nLC3uJl4xPIjCf4zsvd3vwI99F2z8c
ZfwgQfnYtlc9OZiuBC+QjauIEJrk3kPHUrPvfCF82hQPnHogYt8K6xTTWmV27yuR
GKOHWVJn/w5InBXwtuRyiC595rKeZVMgeTYYnhwJ6W3hJc1lEGyLrGpRL+xl4g9X
JgbM0GYvvrOLbKbpRLdLnGO5WFi8Pm9mWPssVmngbPgvsiNOTT64C+4Hl20cs89C
xkPupNNBcl+yvcWnpkEKB00yiH1kD6VcFUrmz9YIiPUOz7OJftxskTu6P7GKIJbm
cpYSMnuZKAuTJIsU8ujteghKewudxmVY3q6EJ12cs2rWHwQKAc8Q6Q7MeBhs2YeG
al5hHzCsJvqtGenFhXUFX2FcSxX7sbAszOL7NgAyOEYx5G32Wz3vJcNYipeZPoyz
0ntSkjJKkMKhyMbWZyky3oXCOcT7WptulUAuAQet9kYMCV0WDHnsErX0uC7azZyV
Kvf8d24Kfit7zUz9bc9CVAVCUgBDqFqGELJRDCh6dppukGXR7f/lWRn12nUe7Z3+
7WybjQc5ZJ/czMqXcbJIn3l+EWKgqsAP6Y0MxGPZVutv56v73WFGloZTN12zZTzS
JtUiZozPHf6v/5MvuQVdbFRUnjDoIhuaMmDx1+lrgcIlUmzCQxrbm4gy8MB0hd4y
VmyMW06gI1NGlk/96rwjlK/o+4DOPh4lX2Xr9Yzve1P76kQTrlZcwQ/yjG4BAguZ
8xYbAjvjwjav/FkSJ1Ovh4LTy5XGYu1rFm/eUYjsvAtTw2sj0xpGRk7qf1AmdOeu
GiuSfPim2dX+BVSXKnL8StcN2TwSML1JCZXpDI0GJ1CvyQ7m8bEDu8z2vA/s3RLw
+B9TlrG5zbIIAdPhoUkXRPxex60ljr/KpRbMyX6D5augS8AF9u9oMXlTpUA6/p2+
+PeEIfBYGXdtzvVAHQy8SLOoNIVF0I2E5qsJ7fruH5/RlqdW/0DkAm95v7VuMpDn
QU+eVw2Es4BMWKiYQmOBZeV9WxskGjKugLFhbqx4l59a0vshkCVSn0eIo2nF27Iz
MyjZaCW4juoXPmSknn68sZKYgsHOlk+yERJpsepej5jtpUZZlRxuQjJHtiAPpPd9
iKrf4Tw6pWsX2i33phM4hsyeBDMIl1rc2wAwHRwjJGtMgL61C5FxXDWKUxpvu8QF
vFDAKkLfXoMi3xz0JWKDu9mUw8lSp7AD9eeEkKJOLXFQNNCVioudqM0F/q2aM1wH
jFYqxI+6u8eSj9JbHybD+fg8w5p7iMtHPpz343quuT8NJTjaE8Dhmy4Y6l2NtB57
uQz26oa8XjIiS6CRlkf/edlzfQK502fjy7PTUWif7qGcE0tBX/5DN5z59oTpGn4u
/xxDepkYfMpQpEBclNRHVA3Ou63va46CtwML6s/M6ShsEHHbNzVJ7zIUTwaxDyQZ
p7PUS2khMSWu7Ovq2+UXiN7HR1cwDFzgWH3KY6/hw2qUoLFBp1orl7N1+HOKA2zq
v43FXHtCeBVW1uQ3XCR0w3ifJW+c2MLqek1QeSfBf0APxR4rTr43kqvukgGc6APP
wVBnR90wengOkS1Ws7QNHZOIi2P7McyVv1RGHULgNXHJKTUVfVbaFkbb4J9GFHuz
sNd/WWJeUkRQI1ci1WfdjpN+bHzM63VG2Aoa8tK0mlVoJWjZRgcOoenxby9wAM23
qfN9Yu9jnnxTOgETgba08cKS5JnEIVz6WzVfHwnC0nA7uZXcDtda0y/BQf1rPIDn
sSS0yXOcWLuRxrpQBSKJ2UY7FN+4X8Mj5b3mJ7F8vYPjhuyzNu+L9ltanngDMM6t
+tfhxYYCkCbxL9lEDxpCpnktlOTKZL0L3uQ318hCcLL5rwrjMrwH4QkLkMgJP53r
1O6HhXX2e176KjRveftsvcVh4qa/iuaJeUkddKWYIFyffKvw7YbEuBeXMfV+9TIO
Aj89zElIkzm0r7Ol15h6Jvg16QKzcFqPBIHye3AhRBZd3ByQWeQwyWkFYlBvBS5j
kt7hn4if0fZt0eECfRwkhMtZ2bDmzDpn8SDiI1BInOxr3jVdOCci/TiJSovm7bdN
N4BijyktT4K6oTCM7PezP1FgyU/VvtNQrgHstg3GS1Gp1CLm0aeCRd0EmKNcQKjb
9z8Mr3Ik0f0IqVIfjgyHFi+r+h14XiU9fHWXQpC+p0h1K8BIwxktdA8vXyL4VDq+
bDjhRCN3MVIFi5vTejdtHUwYTRDO76wUX6/q6L8X+z4EWH4cJTSsolWBaYLpi+9q
sJLpYq0DcbBYNaYYVsfjMXR6/TjkQVCxjeJCHwVPaSnMc/e83t65xIrK4IwCl11A
H6g2WzX9GbRBY45vjFsIsDY8t4zkABA59DTO+aWMFsoNIROVGNDL8eQtlLHlw7lE
1fPn2G5gbvGh2A19Vl0fm9d9cPxwS0/fI2+wYGR6rJAPH4uYpPN0BtFEKFTRuj5g
KbC7yel6vYFDwxwfgQUob5eBqohVvOVgSdh5I+I80tWGGjVocLJhl9xvcliXiOWv
JjPyps6LdZ6OG3BJD3H75jzIVYlX1xELKmGGSIn+LSH0MLNl94Cqc7fpDdojGMky
xzM6UaCCAopHHqVILeU6RKD3U4DdBqGzCrWFoTu2QAftCt9W7mGRthWs+m8wmNw1
y/MR2tTropm688Dbssgyv5epFVUI5589PzJJZbGchTrcJ814czWXnyj2quoLgy7N
KDdrW+3dJu4saieC6pX5Nnggwt9UrF0DL6WdggK37gf/HPvmEsgvUcUjgy4bsQ7I
JkBHgJFq9L+OqxcebdV5v79XBL8TrtYTpIkatZ0Y2zq32t1I8oyr5RWdCcjXxikS
OaDCe0h12JczorNvqv3aKb+A5hMV1d8xxpfk/Z2Ds7Naj1ApgGT2hjcK/wTW6a7R
72eD7wItDX15A6eIApnlw/B1ZMDn+bMcPFhAD+DPqQRQ/F/MGuCSE4cE2QAj0bTq
qtRubVjIDytMRqBt3YANp1CN9n5ELaOmKtNOjtV59aa86aRkwHjegusttDc7JbOW
7WLxjfpZxs/W2FLQKUzKbuL2SZBfdC3rhI35+scI38FbT/0gOXa1M5v9+myKpMYW
mNMbko+9/VOYVcQnKikPmmlqANfAcwxXLgrGn4+r98iLEmaluocMXepcFFXvfzgq
Q8/c4SQBlY42jXtJWLmzCUspWg6oUmM9X425UiYiWpxNSPgT7qs4ofeFZYyQikn7
t58o3li/kP6uhfHtGgYppZemSkqRvPvEW5M6lJlGmGnB7L28i55gV4fWtYeUQa9e
TZsZWTeqleBLSKGOSP2TKdRGQ9VhJQe5toc4q9bsR87a/5wtJaRPTvav8wODW8SU
91mSv8SJqLifY7f1EXBsMFiuQt2HeAgFqe1cfcp/CR+jhqUnDx6FZnNkcjG9HwfT
Y3T7wSZp973Tw0nF2B9GemAvQpq3TVI47GbbTa7ogyUW4Tls81U5PhNtOQntWVzb
/TNCNCA7gzldhcKUj7PCEE3dwzPrllft672R90zZDo/8c2ZzFbblkLxm6dOahTxO
eaqoT9Itz2nlaO9tGViT9sfm4bcfQJmk7rxxgX5KuvoiZwKL6YJRkU+jZXjaJvmb
Ya0usX45zAsuDTXB+lRaAiWNV0LVjgkMK8FBZIJ+Sutfg2pYa7x2pl+kotDuKVZK
dp9Fw8EnwqusRcliFLjW2fi25OagaIHaHpPn/XSs9H+vN/d2gtPvWJZ8MCaKyFAC
BhOnlLZqqBgEQrwMtiGDLso71hwNl+BS7mLVtj67cXstessWerniZXxs6v9IG+LE
IQi6BX29Ui3KQvTSHYMHD7M+oKB4cKiWiI/ryRtSzJtTBsAS/z8G4nwAIepX5Wq0
+n7bLHPQW8YTNUbPC5+oQuzhQuTCo8/673Jh4V/NAQ2qrt6/iLkeC12XQQCMLdsu
OjdivVb29qc0gNYU198q4Xq6vUuSS2yUJa72RUnKbKCf7Cna0bO7gP/gSOpqu5hN
N7ghGqjshX11w58V1KXnebD8/89bsbEvcyFtbAlgKf+32AwliJ9j/wwDdNKi/axh
LEa/JUdELLXo/2lIcFw1udtgL4UCypsHz1Ps4yBxfSPEmgYt2iM5NQYAM82TBeuW
mIlrpN6uDvY2CCVxHqjuJ7GWYEgUuOu5Y7LGjSg107kR4e2+CWuX03A98HyLfGK8
1qD5HnWs+NZlznnwpJdWfGj/xOAoynZFd/7Irdv+GBcjb+JP4S7psCXlRLS/nYsw
YdxmnbXuJi6sZ7WTWXnncNR7/dCh+oeGBF15YPM0t+9o3FEJ5ER/dZy3mmklFElZ
7M5CvU8oVX7LMKSuFrPadsrqiEWk8knAvBWCj1QqXsLdio5rG8VzN/Jdrc5xvAGG
nD1S4fBvR/10AtAZ4akT2O4syVCMJiQ6tDgsZMuOEhIS3qzNYM/XxIdzMO4E61E6
ckOLmvmCM8XgfvzaCvRZC4qkD7A0opkHkiTW9EVvFft2hWipsspu8edwDc8Q2dCA
CMn1qsKygQzgl9VrVpNTpGlertPlLoPNt7HtLKQnqaZQEe5amWm3pFgnEicJ3Msc
ypjQOGtMeufK5UopWtg/559fXA9p28QpdTOh/5Enh+TF6keN42whyFdVGrkSqgy0
DH5cAG/1564H9sLhLxvVNRxztVTFmbbviwloRhuZgwaL4kncZwENCjfJd8XbR0RD
ZRxkImHcE8vxvmT7R+E8wOzo93ILKdurmJQOn4pril38O0ej/88+5tIQjWyYso7u
vjpujfTjRZxzSwDV2yrspdAwfP+zomzGY2QNR6PbBr+dbRLIdJDCvPKTkwBiTaOx
LRMzQ6nAtAld0CGCQewEZIffH8QU0qXmJDGKxhZ+c2P1VH6moI9ix7OBeToKlBDT
j5symgugoOqrNc2F4yqXsufO4EDWUpT2gBzWo0c/q5mqol/yUcs9aPSC1YFtc0/b
AKuMwLXPtydBt0hbGaYAY44lFd0yp3ircJ1vR4arLQ6RKUwRf2GnJ2OYetevlYAL
CwcbilhgnwM3gPj8hhKiBALnBvXXIOwz2jghvEzZp1S0UhcpOuukuCKbTQEj6nQd
vaT26GuiquS7PwEr1vBs2UUIJTby48a+CLgfaYBd/kNZF9bizTNJZfsXJCIGzHHG
BY8YIFbj0GM35NsvPhpqA9th6pZno1DqmjheP6SeyfpOFifsH/URZhlVfD+w2Vy2
w4JftaJjul6aTx1TbduwhYzg1ppPwfGZBiE+xWbjac0+wQJtfxQaqM64GYMmk/7P
La5hCURyeHqvQfuwq4Z1E4qjhSTr7nOAg5NfyF+eNvgUIcZ9+bdpTotIgL925vjT
Au14k6c+XN/fp9UNnTxa9KLskYNG2bXLRsI1zYitlPscuJpnmfvOEZxIPLlKm7bg
gzR2xSdHlpVhDOdrJiYeNOKmM5p2s+wCyFWx/X8t266mKeyXG8Gt70b2+21p7x05
rNwqnpPbG5LKI/vaLTNX01fMgAeMPqpCVzHeIG4c+Kw5BlyKLI4UaLGnMZ2HufhQ
4aHOJIRnG/hyE50NnK7NN4AwLUsyfenR9dUJbMDMjZJRh1WQ1tcFAvMKuWySwbIN
hoEBritC0yshcE47IKdYsMB8FwUScgIdd5QIFX/15yNzvIWpN3Hyn6JfH2p7dUoP
AdqTxNp+jEQHCNlfcpG2dV1+I4SZk6C1JlTZ6A6CndZ5HMI3wkyWB/XQyM3vpBrj
RWNp5NFHulxkv6qvpL9MTcDBMe9VS+AoSXAcQ/BJwO75qbb8DBB8NXNhXg7sFuJZ
EPWmdCrnHQOrGctQ5lnN/O9+riusmhmZCB3uYidY4u/1rdZIODwSCB0kBKry5APR
9/vDar/AqSrP++8eZQfeMppZ64C6M7OIkyyHt43Z36+7DRLJBVshXPkWtRNJqWAi
qyryRaeEpVwMOFKo9OVYIXzl+MlOARY9qItWMapwFQkPBLArhsLL6tWUuwusCq29
ztipC59e0ExezlOXC9GIG3D5bKog9EvgTNS1V4WTloJymWkZpk4qC3g8Ux7t1tOH
bVCoLNpltHFXmNx7y/tq6v32JLlI88J+eIckNNUE1WtG6hUGSbpXgsp8I1HWGnkd
bne4nXAwqC5bfnMe1D2Ecm1mNPJ7ShJE16sFVkoplkslVMORDAYE98ohpEUIKZyJ
0o/eh3tRi3a7nh9caGFnaO+60unMAwmYv+jC3WoLYySiPHE0egYRjpFfi8nLWZNp
cjrSleZMdQbTGfgVYiWTXbMsB/zbhc+0FkgRhhYLfOyvbUat3xxJ+X6K6jl02J1Q
1L7wC5tPJwVULQv6f7O9m3KTWJLQEvuE3NRQxyaYDuEjaT+xxxi1n2WMDAOdVcD7
JtaaLgtTEFhoA1+vt06mKwwJni5HYFZW/UmrKYqzDKuY0w5qg9t2pyQKSVwz43bY
+v6wCWkFp8axFnNOvBrbcAlt/FmS99CA6ke1wwEQuX1xT0wHsmkc95bxeXotS2iU
EAgFiP30w+a568IbTzG19EvJtwYeIISCHCKOL9r3ce9E6Jdz+tr/Ud19ynmXdq+e
1rjQrE6lP/wotTL6LIYffjVnLQKQG5Jud/U+hkxZnu2/eIJSLJ8InNXWtqMXydsU
YJ5PSeriY/C65geNVxRvxskOwyOqHptFDe/iEZJrUD1O0MUPZVy4dYf0w4nht1kv
QeMVuCr/heYAjnNwmnPMuNLiB+NMXsX7WnEONc3NQcov7jP99q/Us6IjwDoNlmsO
2ohZW5DoK4tavZJgxwOX1UBHm/eUMYQLYPFKhaaIWph2dmVa2l8Cd6eIxDChjrpS
hulZo78sbK/p7G0o1MQfbTVUGMF5hSC+wmVvjVWvUcgZcxmjqy5J6QN/n9rqVfeB
ealscROo740oHeWRviDGXYOS7oOR0+2m0JyqsX/xPgtysfN5QJPq41pJi4Yovwnf
pQXMJ3/JCAO0PwIpsx6FA8koxtcFp+Y3/NCvDi30graM5jOLBFsa+a0AiIBpkBsf
wBmrC7s9Ksh1l0IqGfkH2IBZJzyUNKSUA3vcjQGBgzmKbwIy2kId33dDNTZrRFQa
bsn4KfVKKnlRaom12GAz1yBupzEOSehsBPM9juawb+phTRXbSrOijxqhN/yiGeG5
PD144kLZMpUPoTIbUIb42dFJrdzagtzRn/WhG9GK7rU91/otyaAfc974H6Nmf121
FfiGlh4JP3WWu8wnY32ZL/KY3YaLsMjXFtapLJUCdkjhdYvWgRbrjpGpVzQ1J6te
ODnAZt0JUTyZbqOtTVh25EYtrLeRSA7It/FN6WeKSIlX9auZ7pCT883mKAlllWsG
J59tOeNxWLkJr9N9LYcMiRvJGupiHKpmuxDiBxGMxeR7V9NvMKKJnNYrwYeU9XV4
mUDAFGK827Ad/XywaKPoOyZIWj5s6c/phRBUFglx4vC/TFSxWAKhbxdgt1/mFqfo
PIMTQZbSd7QJJ8706XkF8TpLMSEiUAI5opNdELB0snscMWg81d9O9hf6Imz2vaE+
XF+bMIqXOpsTqMQLFEod7GnajuIlTDIKea3hKvEZZuNLwq3DvGsTKh/vY9SF38Wb
b6b0haN6pxBMT7exDwJqx3unjqESqgBbkmBBNX9McYU7kuvkwnhf05IvANphWHvP
dtPVIU/9W/CAATlyQ2zGrXT+USZ/JyJKy4xMU0exyFPkrq/x04nzF1bPAfBbSYwh
hrGPtTwRClCEFcx7wfFf12jfiCpznGTjW+csTrrlK/CgycZfX+ZRNustoPHHHlbY
ugLfR+ilpHOpgm2he00chEpNJlSW+shVTtS6OlwnV3r65iUL4HR/FcuX+AuBvlce
qqts4rR9FZDyRqeZYKSIkSjcHou6WGDgrkv8d8HOVyqS2QNzPaSCGoXNZEVpbm89
CxbaHQfxT+u9IVBGivQ8ljs/RZyURFUxWln4F3Vd+Ngy/apQTzgq72xz7omSXS3p
7OhRJdE1sd03SG6oVi6fsEwVc2QgydBe5GTcRi2eWmkhuNgISyKyB28+fjEWYRQs
psjB7vza5tuJzpHtDqTk73ZrMUJuH7lLC0t/wpEZjKLnveqNtAEz/ghpZPHC2W4G
XEZ12ZE5alyUG8qiobop4imJh8hqwv4pEbcOjIns3A1MP3MQhvtvv7VJ8lxSMxH6
zQzoOID/KEh2UYCKJytTU9ofr6lPuqVxgcUhyHN79XrdDV4f3f25F0+ufE2eLzVf
tg5X14NzghQ2mOiRUtEOmfJmHTr8m4ggrjVoK5Ja19D0aYItJGcCodtnSj2/zL/j
UeVBzx2ElBp5TtFq+UOvMM1n9GkHewUgzawrjFbu702CkrhWfmLJC8EiHuJ8rUsE
QbDX10kKy+Cygxba5egpSn9KMFUZiw8qCE6wrihLP7v4Kgh0+Bv4lTzsOgWFf+jU
OfLus5u57caQA70G/WeUYMdCPE1XcZH6AMCqaiDPBz8pTVzbOqLE/waSQN9VeUmo
ROJOQQOf3JY3sGVcnWsaS7D3JOU3nTO59LZ126Gg1Zk66wRD2hiJQZ3xI/stUS28
WUsAcoboUV2H0PQ+XAQYhqdRQ3ecHiAiaWUavfqlfYtwhfukgU0awapfybkzKdId
n8qiD1rsYXZYijAgTB+M8OtnR9X6KHOWPnIpsEES5QXAXDX9Ufu3CDc8Rirawdsg
Xw3A+BgYeVizEkBFh+KJb8+UiI2IjwzuGr6LVFkw6CWsTAowvTzWRtnVJQlhsqDt
9L1rEKEHjNBaNu/gyZJ+CTcfngMU0FmSqrGZcPTLokxQYWYpbhtGuY09IIA74r7N
pP1wxePuiztkWocXhcd9Y2VQ3aJacMBL0S545TJ2WM5Y26oBgDg0PdYgG8TDE/JT
ZklH3y7CnKJy80ubiZITVP86B8UdLWyIMZ7ZjMeuCBrGtg0YNPpxj3ykK6OGzkx/
r43kW4SLFIlnrLYyZ2jt/Vl8Gogv+szglf57RkIzx1SobTJhLW5vDSqDEL3gcmK5
C+7KcLzHzSoITsotWg0WP2vPy6/Xla1UfkBxC0RxfUYLPbZpyDiUKx6AKlwGoPoR
5D7e+k6LsoGN7BBu9rSCb0y9PtcgCFOe0ip0kVJtFf9OpBiHgLveyzxVcn5eQrCa
mAOzYpIRBVw8DMBFV1HncdLprTfoA0crppr5W1rO+TanMobxwrwIfmIETKCVDMFY
gQq8iIQOcCw7Jdrl86D1xLeXmGPefNxdKD6Z1nObl7ccF8C5enn5CxXg3x2bwnTl
iUobb++Z/BHA2WbvQhG9E/2wJtgXHNSN+jTWsRDomRY+X8uLk2KOphjh2LwkVr1N
T/Bbx5sHsM0S3ih8AxY3V3ET0bg5hiStNTRw5OkqzktWSP6ceKt0yAu6I9E9NH0Q
wYl00T1oaFwCqpJmukSVEijnFZt5CQtILsFWxlFM4irA/yCs3R2sexcFFsOOQOnn
hdYcmN7hmm2zhEpK1xE5XHNSzuNKQN4w0wqo895m8mJL2oXmOD/sMVSjvPBBN/7W
cA493ewx9zKbo/0Ws+0TYlHj4BGhcpeYslczvxTLQ1wVvr8Z1oYdOHc0+/dSyjjU
ahI2zCm4LD0uOvWZkM7VoXGw4pynxaaVOfd2wXX3xlXYIUOh+OjBU+WiYdH/UFut
9XjPl4nUQniofnsvr8gbbwTKpv81YKx5+XwdPcwAq+e9CVlZ37hUtoPOcmp7YEcV
hJ0ubYRSP90Ts7wStIIF3iqdJYBUYF5aHkFmFmcxFbz+Eb3Ol/l+Ov3AZtI3XnGu
zECz30HP1DC3ckSEWp4gm0I8HssEzPl4oZlYdF/clIul6UbpdAgAQ12JeTJFW0Qt
1xFIJ0ziRWmERhq1ViXqTDQ4b7IX3eN+fE+1nYfynB5n2bs/HOCZds7+VnBoWqps
FOAKG+ar4SW3FWYZrrn9ar6cjkTd7zeR4gNuYzzKcLf1Vu8y5tSjRrYGoCEcaQ8Z
GO4HYpz5+XnXn+XiIKWSiWfbIEe9S3J/nWWOGcNJRkUlng0nVj9rWlfcR5c5vigj
b90yWxUmoNXmlG+1FUBMJHRPvZH1MYMAUGyLHXLADN1Eklik8SAyR4+/nyqeIlNf
ZBpkOTnmOhVwBE2HqDuz1Uh2U9ruIuEwUGQg9flInd+fHJhPky1am5fm/Pi9RoyN
ROkLBtIeucZ7H/51D2XYY/ISUz8KlQ1j3tYj3B3f/unaaZkClSW6uPI14cWUSSa+
FgJfbx3N74YAhpdoXJ7wscl50/6v54LQn3cOMQNsefzuMfL5nzk1jQOcKn5K55XQ
ANuct02zaWx+2f4YDcWgMw3HLN3vX+yWLN+RnBi5DLWUaK3z/cd2ApZYYypOYEUn
lg3zew0SXer5MxEX6vWoUz5Q0ICSBkD1+7ctNkYtC5D8fugSrULSw7yr0tKRU5xL
T2oSI0731OovMeseZJ32ANZL3Bsk69pCqWtTnCdWvrCLwe17gt1TyEikIxVPNDpY
R1yPFv7rw6KN3dAbg5JagH3Inld50wzmzMw+o4BfTKrU5hDYXYK6oKBuT5jm9gdz
zwktrTntDl4d1+cdUPD60v3XtdJs2j7VRtd9TOUUtvZ4oOJXSzYX7EGh8JMhvyao
3Na4mw8bgXtX8cNGRySLr8wBjwIRpo0z2D4usHXnQ+yqaYkduaLnqHwK43zowe7/
cv+vH+5J2DlSVmneCfP9f8tUAcBtGqt2pL0OagZ18TNzn3firgH94bbROoWMPYn2
4hRnRuT4qP30P7WMEjIvZlVTjzGo/199wpWoRFvIZ+wynyiWD0ltFpcNta7oObMM
BzKyjgkzmb/dlp2c/WdsIhMdyeYxBj5TsYVng+mG2trhbKErzBWX4inv+8bjaK34
F7wSnx82dTevOSP7lzMBDYGeiwnOa7YOQ+fqvCzWjVS7+h1lC8zWiGLDFesnGc4c
Tm9TREDbY8T/Shvu7w9XJjqPnmkXczMOTYqZLZCwuOSMasr5f6NAt5DyJR88KZad
TtWcGCLgoLfhusr+ysEyHEB40GM7fqQZtnW8cEjVkR+QdtGXWvu/ZtxcAM3Xpkfd
x8b42FqvpC1DtwKirFMZZNCLZogspdydhaIdbFleppV/PuW8K1YK6izrhln+xzDi
/jjMu0zi0YIkCS6DdMFoeugxWDB4lvVvjt1AH4WWbuW7JlIEpsDpSlyPeGza4hNc
zqYroNYnXsO8zKqqY9wKFOiGAUl1cWDZylRZ7YTvHNcA0EVfrc/0ErPGqGznBypS
69SNneB+BSYCd0pquZt0Ke1iAvQ+4sFAU6g0R8Ycn+ztOUkxndlhsgHW3cRFBWLO
DJv6PTRmqGQopJpqkJVQ2tCgHBBsrxcjogQBoxB6FsFKdYXDFN1ZCJBaH4WME4of
wd+ypq5LS7sTXyo4SuJOTSE+ld++zqunt4XefxPeEVQlNhAcWTuMv17F1CQv6oV2
fX8SeOJgea4SzDLhgxEK7AZJoW+pQxdcUrOq9guDIjMh/1xp8juRDBdZN21lqIDx
Q1Yc8hXiCqIGxUVShE6U2pjJV4dCkXvv6Bj/PZqBXqQumj9vZ9fwARl3zEZwFu7j
Hg82v5SgCiDUYT0CnVdL9Wr2yN1zZ9T1rwzdjQ7jPjJgKKX4GO9GRmPnozH2+d2o
TtUT2c4kByONR8R7/GR9euMaaGhz7Qvi5NlpCkp0LyIYhoGX2fJECvMGr+aI2JaH
oWPKOtK+dwByXPn+7uMNcj/hcO+PVkLqsQMe3MelS3zTGKCP4fzJGRNYj/jvEv8Y
MXWiEZugPRpEWKN8xOx1U6uexWP4YK+wNIjoWpKsC8YN66X2e6iZscjHjMt/aJOH
UpH5uQTxbFf5Qun2eXjR8bUq+FRvQr3ROys8mzeqrtTjPK8GuXvD8tFF8HhswBrW
Z29GaGXUqs3UZwRP3QDjTUHmZs8lgC2PDrLeVlneI+hrgDZBeBpwWR/Upe9BR/8q
vtIyZIgmEVe1501vlpWpCtzHMfOCBKcanEZB6HI5a4PpS8/UIjeMVqlhXlmtajFD
fBUp1jVQCUTQjIaJo36B8qybnWw/psKFRKJtCN/4r9nMsKXAke5MkQSB3rq2D3Iz
IThvsO2jEU7YTj4rE9CFbk1lHOUBKhKy3L3bcQC2Mm9nEf48RnS0DSuDz+xdRf31
QtqbIbeb3Nb8ifwTvKtGeiQZk+bTMOt4md68qSTBY+HbunP2bkuoD25bxIC35q/5
fl0UJTjgpIW1p3hcaa7FerNwQPvweLdN+blKBYiDhy2xDNc5EZidLMJqMJ8aPSOW
JRVbNkJqcrxcJajsmYjMF5kSqf8iekzn3faxB76pdnckEuT/YpUzY3cqsNJvURIi
QT0AdBSjOFABwIdeUVsvacUncuFjicSS6lhUo5B5K7/UJ4fQhL1sU000AgEdHup+
8Q3LTb7i0y5yw0uKvpZl6vll1rp7BCVgbkfHqun/tLyerZaCH7lKdO9bqFEbEt7N
4WvpTgy2y8wdN88crmQL5Jwf/QaYuM99YrnQWJdmVZ+bxmEVePLayb86UPe2I1WZ
qFA8CpS4KvVL5hFAZ0Mtev3OoBzmWL4fh+StrVr7Xu8NRfUX5xVBtdpSE59uw+2A
inHfM1MMxjP9W/1slzWbcYbg65gEYDXHZyg9YYNiYvSs4zIPz1mTXbwZnoBpMmbm
8vO5A+dnrEKFqiiD46esQlXQ8hAFnzzae+WCdhTNtfoenJ/u5tFn+vEV9yBTMOS6
GbMS693WH/iBIpJRogjR0SRFQ/ViLLaxhJPQgqiBhfEc7d1D1UIsONOkKIYrdPAF
TLOvOG67lkzN9/Ifhmdyf/JiCHmsMIjy7qBo/a4yr1Pues5oY6B66ioW2IXkGdN1
Tulr+vXda6lfIK6XMnBpT9lKFIxwU8fmUeG57/nr1Uoen8kYIMR3z6wgA4oe1c6Q
7XiknxtyC5DqWNHHCbJ2Zy6e/y2/wfDr3kBsvxw3R7Lew+wLR6r8OgzLmNFDlgfi
BYF3Tp/KpE2XKXIV3bwwbABxaOzAikPMpXiab8ASAH4mP4W7n/7U2jAaaKZ5jmeF
tocgBbEo8LezWCvdGDXBkgARi/qWaz9WNP0m4FetXUEZCVN+nDaxipfohqSF1DDr
/I2bF3nTfZcrpZJA/41191wtU89XONpBvXt4604rh/yqKwZzgA4QdGiwdkGacgv2
w9JtcUq1cmx4NzrDKAPVCM+f3rDnEjUloENS3ZoBgV5vKfu9HUKa8porwDLz6aDc
CetMJDH0tbxxj2MHTv5DB6/rAJJUt8mh133aeqdhwoQGjks/MRVQ3PlEIHnMxMTk
tGScS1HZwFDrrHhhhd1rUDrI8KAqb02hWvCNEhLBUTTVZkV6zNWz5U7Scc7C0yGh
neXYPJIy+/KQMLsGQaq3htqTGx5l6hEvFLIgzcZcDfQ/G+r9LVf8hZhpzp2S87q1
zpNrXQ2+1TNRCymUFk2P95tCXupVKX8zlMknVfnve9svHWoUFIECzWNnhm1dUM28
5p3Mpe42JGfzyq3RX2yAdHDif03+GTY90+5HEpr7HDKjM048xJZPam7l98Fcz/GT
oJCm0+lUsJJC9sWCqeq2mkgPp8TF0n+PcFDgbXOwi0w0BF4GLxl61yQJFtz0wtx+
m/H+/d3syQa1C5TyxZIot1wqlLJKyGpb8g/GKA8wcsFAR0HsSwWzOBRlK6uOs0jw
3+CLbYublCcmLFn2lmJTIeo9ts1mFUKoxB7cPjPft0n3xepr3eBY0adgFTVZCcUq
1rAPrmgahia3RHCdcpPVVSrb/EfcrXJ4wsT385HAQHr9hm3NYrg0OSSJkC06pmjc
SvLd9SQUyMTfsleEgHydvMdif01lLQjP65MztGItH5HXkmq4pjECUQsg8NUp4CFG
pZax/68iwD7T+YTnodFSnWkjySFVVvl6l0uJOEZIkAUkBs4GZfAXjHoCXYp0ITRj
J61MIy/Vz8AuT/iGjqSjkKoJlD+onp4fhk5Qiz77mJq5W32LIWXgoGYn+o+lUTqf
+hduV/XaXJF/AjIZpznzKPUQbYXQ5xGFm9npXcykLT2LimyximSUaMYpJnVdVCEG
1lDuA+0qd4FpSFmZ7+qSG8V/ka0WRJ0SQty10sjv7lkJZ4X8qQszLgDSEizjOR0n
BKozyrRH6FX12wetMJei+rR0oJ4N7/ukIXqikBtAnxuNJpqlIAPN7ZPET7ECg4fi
X2p34/U1noL92TNd0fpuaGRzN5llvqFc5kzS/iYP55kAlZBTD3Wjz1e9e7Efd6iK
95yv4Ey8Wb+DPmd7huKHHj0gMfuZGFgzq2OB3CAKKkTeKaJC3nRzSOdndSmnyJy1
uhYYBIkNn6fDzpWRN0uNwugxvDNGwyMHH8fUOrSPokJkeuVRiknsJXW9q6HS9t8e
ZK7XGHyWk7xagQ4UucDxBcy52oKPd6aObFfeZ+GJTcL/v23+qyYUfyTIKaCMKBXT
VS3Mrtj3aiZnzHM2KajIKyjkwf/B8LGl6ieWFEgpjKBXHuQZ/uL2ymUmQV0CtLB8
nUg4CbHT29fBfNEYzLe3xWxgsysqNkWAlkCFpqrTRPVHtzS4/hmfNpmaYDKOxY92
xlSX+5Ep2aVjwm1RamKqtPnD+HRJssXFW5enVgtd36Mb1OXa55uN+GzsnONA1dVT
kHuKxr8+NuQy+p5Mw4rY0frlOcuKunQZR0n0jds/v3csqKQJcUHY6yn39zqS/DUF
hj8vWLv9gMgMZqsGamCgLq0k8TX2wj1/EWngXa8MyTRW/0npO1ommMvHb5eqXHh4
hrgy1I1E07mDONEwdhq6kMZBnwIIjvjyXs4dnl2vK4OkZHDmQ3NjEnbfJYz3Huth
jn94bfTWrjWpvsqejH0VmSVuxM2r3qN7X3RvdbHX9KQ5wZbKW17/9S5UNRWWHnF9
Pq/FbRKO/NhGMZwGrGh2/Iar+Cx7JDoddxJTh3lmDIgQZETuZYF+l5GuqYtRHxzF
nJlo2cbqDqGn/qyJbpallOqTQC9ZmrDSU2JM8f4oYhxvHEfpimSxZzS7xGqq3F+t
qB9fbJQZ4wD31v86Iu7SV5dEf0eolLXC0VBrmsiOgrRkVSsV+BjpMjIgsl5prxxV
xWdHXu8pa8G5+tNbNaLJUuxsVh0i2bCIQROFlfYIoDHKKd/AMiZF2tQm6UJNNAxA
a+MHXyr2esbnbbmZ3ytmHvDhTLU9/FbdhBbItX2yMzRd7ojrK9d5y/lwdUmgV8iO
xlgQakU/OCwCr/F6jpKxko7C8NN3RbB1CFNxoxt9J2FQzFBtmjuQuxBhvasm4ejx
XRfMedqQ1fQGQ056zRYe0OphybTTB7cV4tCf7XXJWheD/4ruZwOfDHAP9Wwjrd3H
iet1Cx5PApijtA3Ao7qzvE0LgM9PMDNyJarrE54pJWIB/iXkwddP3gexwaW+RNjq
T6BTR08zJgMv894jYqyn0w9DmQZOgrjjRPcQUnqGhwy9/Pp6MdwZ6Vz1B2q5fVqx
t6I1+kHgFqoycHt8cL6CDjAESjEcej5s4aK3dpf3VF2MhlDtJvkePw3hu8JAWdkj
sK/160ZizfIckHGVhMp2BAGhJeTDQDEjA3W/Hmbbv8cTcDT6Zu0y7+WQ6WaiTOei
hmApCbGY+5L0A7Jhd+oeac4qO0x0AlDQfGaiTvx8Z5kyTz2qGg9Gljct9Ru66h1J
Bqtz3QOSsPcptWhngwB9hZt4ZisF7GWH0C7ASmqtm7fIgb+VOGvOJRN9DCGPXVNi
FwtSuTN+8ARWG03Thnxh6HqzSLrmC5y4xLoKEfPLzu8OavhliFPjfSmPZGtuPxfM
H8zdYnxXDNIo8rjlWm0tmjk0T9sHKvDJqfKBhI9RyH3pB6JTdtDfoImiJSQZGzrQ
WYxyXYDJbntdz+SsFk37E93VqG1Ypo7CxkLixclr9u9hnAKI7MPEI8H9P7fbA8nK
Q0uhieh5alFk6NGAGCpSMHOuuJpLWJHEEoNtqSASx4eu/tVFiAjuRHtZrWI7ROiN
FREvj44V+AkKkfVuQCFzroAMqCMdtML7msMomaKAVAYwy1y+byo+7KOwyIB4aKeD
1ugyehYdI1esc+wDrlJbuls2XE7xHUxeibR55x+4LUuPrDLcHUv+QTGY+h4K+bSx
9rrREocmFSA2d06zki1u+i6lldinrUtawKiONwB1ohbRPt1DdVgz/9VNLj3Q2Pos
osySEsriPa9sokiK9aNve4dHcfk95d/JnqxOSHeINu+8fUhvF6ijrV0NRbXoGZTk
os2EgLcnUWiQugXCvVw4sU0YPq16Mmed/OltF0fDNqp9Sml5FK9jZpl2k+P2m3x6
CXnTZMT/sW8RmdTkesLhGTM3A+VPUxXFC9HdVO3JKBOj3mdRrWubS2Gv24UGe8Xw
Etr5y4QCWjrYBMvdLyRVmhbfongM8lqlbHrJAp72V+mAggG2WfV9E/pNRyG8Qf3b
43gpldO79gozREdl7uIiFu2fR8hmd71hH66y0ANBt62dELz2ktPKsBBDsyN2h8JU
ZOtiRCbl4aXP+NoGkmOEGolKUiU+6QFF4+HTxDYatCFPxhInxuKa791Woq7LrbQw
+Ex3w6P66eflVo67L7feZr0o1SI9iJTV3vA55n06kQhSvVjcKVr+FjV235wKGJ08
A0dlmY7s87q2V6V4o6lNAUzNfBcEujGKXx1ClxlEyn42orJuA0Jj1niH33DpfIOH
faAZQlOi6j04YvsnHPXlI23VEIEe5pvPRFoJaCd0WlEatjXG4eVgK7/cEmRfX2YU
kaWKkpMJX/ETJclBa9UoD+kvB+S3A/A8wF38FV4PL4TLPXyULSWb3HCey9+yG67J
l+XkgZel6F4WMpj+wG3TyzM3n/IYuGsiPdbAqQcQD/5rdcAMqfgupqZ37AdUw+Vi
z90elJ1otvhKKMf1H9fDNlEEKzQEMKkUxkNC7cgwJixtQgxOXPixHJLYB0WAdELA
ciQa9OTPjflWoU6Ou5bBG0CLF+4nNHJho/aVcN8xbhsmqMhNYkMsvMwaa54DUoXo
xXLH88cPAJD98slfEEs9JAxwtRFFTPAET7NzQeVF6XQn/GJxnTpNlOZRb1X/ykIt
0SjTkWcmf41LfNVo+v0X+lq6sF9jeV3DEr1Otw8clxJXjP89Fy6/hzv+85TL89UK
Ug1Yh2uDXffu0n4ZIlODiA0pIYQEsjJlM9pIWqJz2rhAvFRsJJjxrwa3XGzce3Bc
HuYfWDz6kbUt92XQ9kaBzLMSxEsttNoYgnUDRLnoTxZQkSLgZL0BCu79tXDlnGBT
`pragma protect end_protected
