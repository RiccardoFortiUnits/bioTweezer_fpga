// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
mSDqHVqUcnnM1vKroHr5LWtEZSvI5OpRcb0w7LZw/1xa3Fto+sCpQSMTRpAg0MRRHQBKkgEMPoUk
r/duaaBSnRIUY/9+vq/NTLG24xUJUdYiIzS7SGrtraxfbpFB+qF+aqpNpp8x4FWnJU2LfwwU8KnV
IVzh2ZxOJ2BhtP4r7A0bJpR1aPt+93cg5YjfXZjtC1mRbFbcfEiB7THJ+DnyqL107EmCSD9bRIDR
SD+Qdyk89uampxSr7Qby/adqoFmB5jI8NHdpJug0nb1ahxD6f1aaD4017TE5/KYvO3cpUflRd3mA
la46Kqb5rXzGePeeHUu4D96JL3vmDgb5E6LB5g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5264)
pZyUcr80Nm+v+Alk/g2BvyKntJjVkas0UEVeGO7hSdiRVpQN9e3kHwlJXGjwriZvj3kNexfK2i2L
4l7mxdqr6w/qapexnolLQiuBUqxgEKwt7vQ+Qq2VKC2iITYlm/MjCYla4IAUGyO21Py5YCJch8F5
LSO/A/2xu3N4iI/+BAv8yUTTeFqn6Vi2aISIPmevFkVTtAZTsNZe00B1lnQcsrlMgoOy/BYfmE0L
hppcGLFF24EBfeDcVWSM96QX2K9cXhnWxj6kSlMHfOZmV61bmbFux1HBGzUt4s3MhlteHlG/w/KR
4HklpcitUWCKCsuaU+ARP5gogk0T0k84j86SW9nZvfuy2IMVTNMZBQy5NivAraLY6TCjgEj4NCHa
MwfaT1HciqKGKrLl50aUDRJ6IvNOWyI6ri+Z18Xr8yuY/rIN991E6s4CCBqswLIaayarSCnfuGej
Y6+MmZWQtsxQBex84BxXfyGR9pkjBy1TRXwOY4k5geDm5VefFiMIp+Vq+5bbe1tHlNxDo/u/9VFR
t2eAklk+9eZ2qn53IacrEvfzqY8sXYqCdONhd6y+hba2inQdyfWUR5B7vH/0wTidVXHL3DTw13m8
vGP+yTMQatKyPRcryIhBS7DyIIMwEznjlVn/5hkbi9wmxP9Yg6IXZBS5MpBKpiLME3B2eb8V8Bbt
EO7EsSx+SvWMvPPDJGgXNchMXs5x9ZN3ECSZcrsWnOtKZBZsf7NmM1RqSLZJhRzCiwQ5ynT5dvl+
c0GrU0QXn21nN9dq8r9PpUdgYWgqhwAclWEIrVg6FMG99zSA3oywNC32Yt8M3UDibVvutopCZg/S
0d7vy5vIfYp04HxiQZc/4AdomDNtttK4q1nU2Q8Ibt0ToOzPgHW0tzCfx4lpDtAwYLHzKk/PNIQC
Ae65pPOZwXYOE6dZqNyzjd1aE4JJ3prba9BYvGMmCb+kQSPN5G9lD2dc1gDkWAsWlehG4dvu7Ii3
9CyBGxLrwBB93g1C8CukXpaB3om6HQ1q6zALqVxaIYJTKiuf+Imabxzl3clkQ9Djx++a47J6w3MZ
MsjZAp8lSLrAYV9h5d1/tpGN4H8aGFxIUTZiRk3a/S4EZ4WzKeIZkzMjNEbMcMJzqVar+wbDtpJE
xtRKwfNGZBSCrfrZ5MqDm0V3+2DsUj2Ajf/Lj+Qhf7fS43+fviJV+fT8PQW+QgTG2TkP+91mEbkV
JvW5KREGbBA7YaC06+w9KNxaezMDcjKBG0qg877P5tPF2vrnwFCkz2XfBpM2SrmsDUgPNYf0ei+W
nI7G7vPik7gg7EKiv46cBiARMUpY5YCPG/dw2jrdtWdC1nY4gW9gXvwzIKFNVVu3pEF1Nb5hWKFU
TlSqVNKXvNZmwT27dxSTb/NJraAVKKbgxiF4DaJQPhm6dLeCnzcTr77ssNTpfdzMDx2pMb2fkpNU
eCq7Hir1X0KgsQ42lBhX/tr22QZrwrOa8/Kno6ngUaS1jLiuh53hXAWJxq9j17RnBx3upE02ifEw
xW+S1Z380iOkb/Vmx0OFKZExQAqHKOT3dpQUlx/fZ07t3U2Jw3s+ZKvhFjddQMUdTUT/5cFsztGp
PJdfjLqcDUGW/DcnWo4fXCyIg5qr+a7DxxwwXXnCAkaT+tP9F0jdFerIbLuX2ezcVwOezLZUPAR+
xy+h7+s26DnmrvPSOPqfvZwueiZJ3Mdu45OF3bcKjspHyh1VgNKZ5qc6XY4pttXVV32MKY6MMSt4
45ZQlTps+cndqJi+Um7bnhNMmpXPLcAVk6BJ3ZPwXAAq/01mu0R/eb6wNOUrvREDbdQaG9A1XBUS
agGjidwTcsMf15WtK9OrCRGg04nOkzjKeVZo92BxvGzTJo/UvEuYt35gDlUZGpiPvHTHRLJXrTqn
Y7SSssWqUbkIGBTS+2aKaxwwetwAFzy8su4wNVHb2KtbEKKsM6LYr0z+KOnzvy9sIMSZKbFBReCO
oFjlgOcmhwQJITO9W8ifYN5GI1EFX4WwNwA3jMdTZu9NmaMFmd5Oo1xL0oBctRgyoksLNZQrv4W8
wwVjhn65KwJZMRY6zNOhNazkTO06y4YwF8LJ2+LPryzTvdqQu3+TnaX8Uz7b4G87VUTlmsmEDUoR
b0ANSfgsS/pUpe3OvcwQNVngIf7tBA/fRSE6M5XzeAFcWLM5C6ssF0DvbxXEAUZQZbje6cxdUJnD
zX7E/MRy/hoWtEpkVcBldiJF4HKso2pdmhETtggikq6Jg+svjil4SSx82/hn8CKDBCuREZz3BJMo
7dp5ZAn5tiYVZkVtnQ3hJFS537EwQBR/rmxpRjQib1Ba+I54ID8XU5tCEi6Z1l35JHQRurpjC+UL
qoczEgfHCJ9UP85+SDJ0wJdONQdzJETmkVU5ETd2GVr9qviaAC3Ua+Legrud2L+rsvhjQ5cuKo+b
0jyVontfwkheJ8E1O3GuvlqXxc+xd8CxZYHrcwz42AFJna0/9k4fyk3AGnu7ftIvdez25sJgHxfV
jLnETDfyjMIROSRSbBs8Y6PJgUN61Nlf8i6Zub3zpTSAngyqQJGhxifYYChoq4h4tavUCZf5peww
HQcUKBJN76YLxAOxPDXIkTpyelHVzBLGNvYO8oVRMRO2eViH3Gx2BWomi34d1g2CzbsPC5AfbSec
BsnyTqJwPOR1cVo99jVxPup5C29fOt/BENIqk1CZByojKIsVPHzbyqDnYyBoW7DuvH1N02Ud8BsO
1sKNk3ISD/5nq75VgHt2YTShHR517U3Kb6e1T5xJfSec5THom5pdrws46QEv53Zqjq4y26aD9IFs
6g2gUksaE2fQDNhSvENUniUnxNB+2H8e10zpRMDsQZ388NGcTSdVKf8GjDmX58yzIvTFqaOLOiap
NZFYEgj9DRsbMVVtSupdEvHQZaM5NxO0CD0Fry/OtV5JoMtUGb/RwFfYAgKf34ar/bCP4rwnYaxW
iETRvVeGvxDTbWcI4eLhzCAe6NP+n/LKPOlc/Q88arvA5wKYlbF757SStkcsgRFL+6dknZVnAlMr
e0H9nkJgLUHlH3zqZU8HJd0OrJaZg6rl0EK03WGr758ke/bfhXx8prniFXoEoZn376WG1g+8rAtc
Pl6Qq7hwdlDE2YWXXW13z/4I5NJo3+EfHyGLHYoXGMmpAtISNBgQD6g4Fo9y5NcGAywMctr3QOYb
jI6LUFqwCTYaHzo8pqZT9phXvWPf3NXme/mIeKZr8wGkZ025ncw+zTpYNNhHeir7Qg0T0kF5HTIy
8+UaNdISNsc3ati8C2OXjdFhsEQwNVX2jyxELcr8sRXS2QGNyVMhaQTVfH6o5m1fRM4+3cZ+IcGz
3oHRFRc6IAle4YwsoHXnF/S+IpI/+uE7/E4EVArV+u4ehy8fBT5uI/V6nG6ZZKCrNL32eI5wpFYl
+khmJEyBQbTkOrk8pAG3dPhoLvSNdJT4KNhC75/G1EQWofxo+FxQQYKiRiudH07w9kZ/NZ2C4uXJ
e/6g+CaKoKspii7k7ClWcZzW/bycmDLs4T82LIuvvdEZnVpNo/CQQVYpIOEBLRfqFVId+3OTNvHX
WZnK3w5OW22z7wrnSDm+jDuEnJHthd+xeiisC+rp+VsxLTsaoMC2mL6fJdFCu+ivjSEDJ+bemMB0
hnsO2NRjcjIzFgasi7aNNW5u/uKV//NvvCYtsdOHBgKxtbblP2I4cMjrVEPofRq898xsuD5UVax3
qFRMUgEyKBVBkKhdbj1RMHDEJilPbykvcEnviAJ28UMGKL1rKmyipJQYxgqNz9qok9f2RDuhDGP7
H+54VQkzK/Os+xh/+8SsmawBSDh+lQzY6BKPVpEvtF8undp3mMHEFfvWQgyL5r3+yX1hdFRhH5g/
1Zn3mJ13/Jvrfeii932fy4JzWqOw7QNzK58u/p2W7mvYA5caJDBsMyy11pnMNTaCYhErAxgcdjCI
/A8tGhOw6e0LWmIyk+3/vuSL+33Sm20xQLw5h+cAh3CJruk1PI+uwFNbLYEUca8k0XyPGWKskWy6
aRGKDxCNYYO2kN5f/0+9ugYOCvLLk0hTGhIprh7MA+4GVkVfcjP24FeC31UnQ0j0iBU6T+iz/RoO
R23wSAkgMSEYfKQ0SKLouUrdsJCR7c/w4O+My2Q9N36QT1gcTaN4pMK3q0WLckqFW1c3tnyMGve6
4m3x84OMdmr5h5aP/bVBRLtqCniRU3wVlYcs/tVQyL2A4KHz5GklQ57ceDRQvya4XPIIGR6SBZKP
pHK1UdylvangkrbTHRlx9Nr0XvRcqAqh9GlpyrPp8DxtiwZH4lPLVfMdaDHlhNw3SjvNPGL7eiUg
aN/iVjpD6cXx1oFBBiwI6IdKfnhXndOq+eP3PKTZV+ljG14GrCKjktyh9JnwbSoVE0LGBtvJaZ1J
8h7C2kO/osee5TKxP2ChbuDWYgUSKY7i6GOh4sJpLSfZ0lW1QT/noO8HCYM5xOr+VP9t9lzpH43x
4SQxd4VYef4nxpOAM2av6FTK3QrcGuZEKlKfW8UCTo/AEf1Rth7+e3YLbMHWDu43H8xDmjfzA3hF
BlCUtHBlrgfcHzZf7zGDYffNxPs1oEkVGDQ1FoiF74SYEXrq3PK4y3ve2t2CGv77kFCz+aljRoMa
MgZe4rHyBr+QMjBx6rHZvCFnkUk9m1pv4808V/sFyOfH1mdQRtslOPTargeZK8uzFJrPB441OjKO
TwGAicq76oeSyV1vwfHUjImT+ZLnpGZDi3a3hwConvAJWcqrr8LF1TlKtxCY/jsD0cwZadOdR4RZ
AvVY+6VTVWFVPN6DiYSzuXIPujFjQyr1plix13zztm+qGp+91SNIRWxJp7t1hnHrTfW2USZJyqL9
haHZtCagE3sg6KrSn1+NBeN/skc1d4UswrlSMeiRYDzt31UEYdDx6edZGVq2p6e8A4XdY4/y67nc
rv/4bigYaTZaxYzeNfaIHb5dXKa7vHKeEWlNV24mVTPTJUoPFOty5m1m7t2mCWXjXY6EM6WfuR1Q
dxI/8pYi+A2XLJOh8u5Fibvw6UGv1s5etucOgdKLX8O6oD0K3ljQRVpq8ET2JDEHYo1RphH/PSt1
n5ubB+tK6ykJXPYNEgTFZ00kqtuOZZt5bTTKK8/eYyYaQ88GYAkBEVBeKY7yUkrJOMEY9hMQMePD
Ik95pVDidT3MYnY1SjwuO1SEk5TR4ucMbj4sVXeQKqjZ9ZgNUh5k5f5OUiHegsy3y2CDFV2hed/s
koupUtRwC/X66QsCIH7XjP2BXce6AtAmF0Lo1LIZEZ3vL6h5vGXJctEyTfxIdS5MjZw3L4c+VjQM
yId1LCyyiAjlGiBunYU80SUawMj3rAN9vZf30nez8fk481bydpcLeFLTM6xHOYDcfyrl/B9xVl7y
TZT4KCAeuCSVPo9Y77upvScX2N5ga5AveAfCSA1lZjHQKIeL72adESREapS4PpBrUWTf3Z7QY3Ln
XaO0gqE68pH1aUvNsm0e95vfW4IhQelcTos2RL+xtyG5Gm1NhccPFPVj3Xxre4KZoESpc1ZnmP7m
1RAwkUG/VOsY/66kps6kqNLL2aFSqqaMWo2LrC5Y+iu2VquFPfRTEXLb9+Ty0X/TyvkLh3g3ov6h
ebpQsosipxLPNDJPXZudVMYlVOswV39i4kZ5FbjpJfGl7kCxvIk16IY47Y6UUzl6sCokOpmy8Mzb
sOGKEnOrXcpYWjVEB68TlJJyEuFc0hSV6dv1+HgloJDGKqdzm/qhGvErX19uaMPMcX8EGulQX1W4
2WVKkUbydwLwvqQXQWUzN0rKqK4ToB74bPinFsmW1SmuAstWIW8/huR17q7mQHTOKKdKVEnMryPd
qhxOY9ig9kpfYpuHsKcjweseMa5C2da3EPWbS/eFQVHP+EYf16JuAVdAXaxYaXSfH2SA6DU7mkod
zKbTTmYogFrVPaSdXWuiqkmjTp+phhbQHzFYNV+/taH6Jtjbc2hYgeniyyjTjeVNUwkveqc33vtk
9aKttaiLRhRRlZehIF83LIk70UkUxe5ccrRcly+cpYFif3vsqALxn+J1KWNDufNHjfqf+4zKDCn0
gNEtgds19d9j72GmRzqJhlMnlXqrkRZ5qlsj7GqDkEPDjp/Rhz5YChafbXwbOqO3z3HbBugvy39G
rm64DR/gliN791qpPKPmqQ9mpRMgfhupKXEqiKh9QY/9IJLyq3+YdNUtN+FW79BJHqHmFJsygShL
Hp+fcq7KDMwmSeniXqZnAiVW5IjN8KdMhklK56yauNYfKwRJlZpKRWUi1hUwMyNK1PCMpTPmkw5j
BhGfYqTnqafoydjYHs411MLGeLZQfqXnGy0oXzNu2KqZogNWdSI0nUlWlauN/+wbRRDXry++7x8s
Q+Selmuf9ni5sFodZs6opmZt6t+lRz9yh4erEwNpFyBqV8BGZHLA8uUph70/YiJqanpRjlzIsVF9
9Qi7OWIfzRC/SRdWXxzMMytrcHSH5r87Iu1FramOIsHHJXCLmVzeiUd9nrmpf5RY83yMFTROLMas
A56uz2xwgEIFZEbDIUAIYoSchbeWBdP/0m/iifd9bjUeYWa5tSouKbzLeS8rwZymQ/sUEYQelBEz
VvwWZirbDULESQLzfJJ4k4kkNBoCU2bQ0m94LFLkXhoKqsasZIjIPY6QpAe/omzNp2p2KZhAlPhv
wxoI57TbEtSIPkCeRbCkRN0/vBDFwrl3jT45wE/+90/qFRD83BIIyVoBRG+fFgwn/z++PqDZHMWx
QD7o56Jg6/XXPfpFVac/dFcqzKiIlQyNoLqAF1EuLXeVYxyA5zD3tU0HyJDC2IWRy/2vRhm4Eit8
ib+nc3kZIODgFLO1BpM6AQnEF+mXKU8bUeXyUHcUdwzZiSZokrHmKTT51HtUunzKXt2tjDjHRO2B
Wj61sPpm0KjnNAkWmyiWqKhAl36T8ZlZYDJ8DMfQEZBipHqnSRtPtIOakqP3emW/oiQZjlCwcUNx
8agrBrNBNnwvr95i+LUH+oqFeM8=
`pragma protect end_protected
