`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rI5jlYuBUz8DXW6L/Qro4tHg9u76SzUnQ/XjqAgfP5WphaSzwvZUQBOVp/7NxXx7
Y6i5OIrTf8JeYmSdjJA+4sghY1by2r61ndBo2u+9RwX5dC0Y5swuqnJ2ftP8+dNZ
1n2rhp22ljgDrV8QbGENF5t2wnXB0aDzH5MmZ349vd0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4192)
nQ9Uzahc9HTyWH+DN5Ibvwx4MonMQqIj67oRIfqsGvuqJgvXSzh5spXNaILaAPPy
5Xj41o5T71KkY9le3McBJAu72rsS0oVgD+ZQ1Mku+rO3ryRz26VXFQpK3ftQoMKH
cPwLut7WM4cu2A4kGPZdacWtfEikb65ubwA7WEoyRLJam/UwXGBzfsmiolK5JLwb
D/ZaLJAv8vaqwoXACGULyO8SsG40GF03zqmU7KEVswVTkKDq0F5T77bbhl50JEo8
nFaxxi2Au0D3OU0jFe8x7PFpXEtri3l4wNjpmDKMj6/aT+HXspLkTBkSWH05bk1G
EnUFDdF/5GCrhkCw507+Sx6uA5elFXvJdlKhwbPwPuPzKzOW0FlXi4qqE6FBUxb8
E3QFOnf/p5OBAZit6LnPqdK8Gvrvl6K7b2LGzpsBLfWQEq/531TAzAQTB7QTgLZ9
qGrXTOcScdCJaaTp+RtCs1Udd/YiIXQjaWiWE1/dbVEw/pkHVFqOGQ4ic2QAusgP
pDU1LfrS4FW0wBCAINJmskR2CUAGWi4rVYxjJAzLBInHLJ7qymAMOx3H5+bAqZ+w
i2QF4DfOfgAydkRsrOu6wYdHMfuvZi9kExh2BO6F/qBB+4GE+LrqDNuqta77dVxG
2FXtD0GYHE26ngwjIpdFpE5HDBmJhYydtj0VmS2D1br+aVrLoJmiZSfMvYAzVzcR
bHgh1V0vA3PCPJxNYfubOnWkxd0opK6eHFfGKLjO3cWD4BxXNJAmt+0jb/81F6N+
yKYe8hof6Z7GcThtpDDm5WgEpnyu8r6laShagAWwwFOI+nUubQbJZEg88pAZ6euZ
brBMkz+0aMmr47f1xG89t5ArjaDaD+5bLLL7t9ZosnD5Ha14YoEce36EADBJVeef
tvsdnfJGrG9+q7Gp9K5jCzHXdD+3iT+KjGKjDBalUqx+YZEJWK+uRsPDa5YGbi97
9IPhtm05NhYkBZMa9nb8PUV4tk2Phs1QFlg3eJWvujbp4MCnM5Zr8xnWdLdpU7rB
BZ7NCET4bARJZR+rMX5bqRMLDKfd6SHBSx9rFmlVCOGXRdyiNRsQN/TIN8SNeRdk
VHGRaggbHwFCu5tGh6wwNceWk522wtmw44M2XVNcjvrKHnb5FjSjD2X6iyzOhMCV
n3waVS5BGLRaL0V7JZpe7m0l1+VLxNdB9ds8Blg5axqOSFVgXaUEJHSqBN/+Asrb
RWbRyZBYzVojk40Z+pJcG6+KhiC6USUu2MDJUPSND8WDDCfZ12+1+7XMce+Qa33s
OuOAVKjsyiXxQFuKYdqOG89GiFFMg3/S77/OUC824FDshffXw+lgIN5pWb39WBjI
/eyQV+5rBIADYmCMLPUwsYz1WV05IH4kMoORoYY1cWbGJlMCyUg9UgOQiqj1sizL
0ffIfoJYTwqp65VgLhEICuItg0e5oylmOhuEZ4GuH1cKztrxbH91HkM0A8ov4n/I
SEgRc2ozn4f/2rOYiSvwdxkEAgVdBIAiRzLGGmSjj+ExRserZwvPUB9AyHXMJfSU
n57KD+I6U/TBa6dgtRojx5xWqOdef5wwx4U0AB/ydU1MZtTGQOsesdY3A5lghOYk
1rPn4fiuBdL5kheLajwCqvjy4tvu/SZ4EbXOKkmwFj/WDoaZ0aDYnL8ZaoD5fN2O
mtcZXoAbisEclF+zftYk8BZzHu3L3UeaMcAKQWH4xjiJ4uVrwoZyGURtuGs2RqKI
NVz2Ou4z+KN4LCtL9DgvpaStQmaSxCiYUvD0UNhPTgvG//M5YePX8HhA8DDr9Xbm
P62k9UkpqnVixkUqfEv0yCDEzc0CnIEV2rJ6XLeISLTXFnqBHoV7JMd/dwBFODMw
GprbKk0pqONvvw4oNvz2eADT+lS4TOJtiqlVmarU2aM46umXcxGpglsx1XKx6Upe
pdxBHCzM2eBrZnhomM/Hy1aYNpbJb1+9FxIjL3Hqq4kxiqYRApHJbEJKtAxnnorU
HakuFWhsj+0Zou/XtGm+PcCdFymyywmZWgAxyWqRxWZk5cySTCteGwBgrkvAe1Hu
hREnqKF3IEsHyiydom71isCF3D9pq5zPwWGqi9Dw3M3SW5ujEL708CTrJ923EHFK
v41z3wuyUF8Um/YVXKpxsa0JiAl/j9sLRwXtGSJ8Hambb28SiQZU9PVKoAf4+NFE
LBQw3rGYGb7pGLi0rZH3p3bzYALgzEmlF2KnrkpJ9o7Jmp4YnzfeV7UvEpHxWqvP
V5jAtIMlR4yoJ/2A8bf775Vi80ZoTfslDM/PiX8f8yRZRZ+walGLaCGLuhvPa75a
/T83HCPeaamUvjhHlS4dAAqWNfT1rrch2BaUBlKJ2E7kvHsrN7SzxL6p2ypcRZc4
mD7Ydrp+Ob9q/XAG0vKCqAk05ucHvSpS645idxjtVkGDrykjPuxVk2MbczFVnHOU
domFuZrvi2KNGNPK0Kririfx3MAGohmoJgO8dyQZafoEfEe+oSyFz8pzDo7LeLCb
XB/BxuABqbM1SwZU8aB739hD6Jo6ObgQFZCrZp65XU250687BY6SsI9VTcVTkRDm
C8RE4tKg91Ioh9K0gwNHVCM3OHqiba9qaXe3oF7AR9YJeT4o60FCGgcqnxbwAJpc
LSnLOiEjfPeCWjs++Y7FpCG51WghP1NWrAKx+T1xmUk33BJ6gn+EK1C7D1arhMmp
pb3baupz5JkOICDLdvyQFp/aljIXSep5xezRrh4qXRnaLOZLnsQu1dbWrjGkTSaB
EwZsZpulDoNyEvppGTQmK0onpHdGyAKjOv+ZaPA7ytq+pup3dpqm0HGin9daB4Zj
AmL8utNj5vu+dJ79yqJDIKljh6/laPnplcEX/sSzxogusHkZd8Vkk1hliJsyjfGh
OR+61BEHJPm1+WleILWnJmU3Bntfv3XgzvKKFCgOBHLoP+uIK6B6fWw9nijo0QJP
HWRlf5vGzPoVbnDSRI7em7uuodHD3/GDlL/Nclpyk4eJqn/uTGmBtdZtddP0iIDM
NdXgm1nvitk63xgv+xb4bxvv29X2PxcLO1JnsJ1ZcJBmHFcLWBzgNUtAYu4lv2BD
LDAKkzIeQ7nBiX9e3J/kKOOLBBKIRggYV1/EJq7QcP1/RhgvxgOSbnIvxluTSXFx
zNXZLcfkFMc+VKjAOd5ym6IC52lpFXaQT+KnHUK9PgNDLuCv/S+7c48OEJ4zUy4H
/hKpjNCwRjBpfut0K+I21tHsI1KviRtk9Ih3lkpygpTI1rhOhJYCZqmW3F/KxOX/
Em/Bu4TVbswgod32gYUkRVQYyzL0m2+oe0zI2ifww3kLpaEnSNCINZGwTRlfF5cz
V48T66psSJ8v+/ep5mkC62JdrccfyybuG2hYhbqgrnoRncDQ07k6EkII+V6Gn71m
FZ7OjuWPA+lwODm8koz7cZBZq4HeUwOoACd4VKd5oId/TgJmx1cW9ZLpD6N9OTao
3UTvfm6ec/jMyuImQ4kw2QK4uiUXeasirdlD1jHo6s3XbLU33jMt3VtjoOZHIqPB
D0prJoqf3MHF/B5ooHUVUYcTWqSKfQOl+hgzfGucgG76XFgEFC4I8NVZXaCJchI9
9IFfCSIfwPeBQaTiKu0wElUvFoSMxTeOB6MNay14YwaMg462ivi63aM1JRF24eKf
RxlAsKzf6DfipeTO2PIEtMRUhYx5ATmak/gMEdgXQFeieGt2AgF7ymnMqHjg/AvB
oygF3sSwcJSv0gIzSRCzMb/1t1kAAfkX/CEeOeMUVAxCxZcwIJglavdlix+mbE5L
5EMyJZg9dEcnNyQkUwzn4Sv6ZU1qBP1GukUUt88qHVyeSX2tDMed9pAIPKp0VVG/
P0q9hy+H0WxEI8zrYjnboozReaON9PqqTfELtgyu/76mMgUHQzI0zGL91q3ZdnHi
c7HCnC8dukvxiX0hGGV1K3ajDldRGdIXflD4AngGGt0+hwhdBL+0sV5MwS2L2zov
i4wPk/mK1ZFLCpiRRGD6NRnlk0sXER/GEjAVAt8s7OM7x4DiwN0mYlmURw+pI2iR
VjcyR9YX1O+ioLkP5wehOhJQd3Yk9wmBqg5IJQhnJy8Yz3HeB8J/qAWz6ToeFhET
q4o4sFacoqufO1gKewi/XgwFkzog1AiAuhbooI6tUVNwAtbG1/2uDTphGHQV7uyZ
ndIVn11bF0PQZkzVZ3MJCVuoHRAIMbWrEIzncq/onAJ6Rwa/Xp8xO8ACoL4P6wAR
tT9w9XsSOcn8HltP8dSeZsgsTyImPuPY5LFdvU/ulsPAaOInSY0xzsQXvjsZ0sS9
+V3hBkV4N+CzSPIcmept4m3UqVXNrHdwW3RnXPKN4NODsTA/9lTXuT/f2pdyDa80
j/Z4y0Ticec0h9NckSgalRoxghlBK+oPn4OnE0MMviXbnWeOJd1FNo2suevDjYo8
rmUXwRmjMp0EWgVG/XJlytP6JcBRSHezZsQKSQPwlve8n4dxigcLw8c2rIcaz0Z1
Gd8CyBj3MbqrqITcvKWm+ruIqpEKaa+Ga+/kj/Bk1zI02LWkAfhaeDjae4CcVPo/
mPzeSOW1WHXFlNHwntVl5KpGt7RdV4xof8xTWz/bPfdO0No03ZCLHIsJZq0RwsEe
DUe1Lr1HpPg7Howik90/gWJ+jxEsZE9YIr2NJvjflTHCkpUqK+bGQMuj2+dI0r1U
D+lUdxtpd2iprUDkQJ5Tsd2QpwtvpLiHrkVBkeFg9NHb9oScmclu1e/pbUZ/sl5Q
LiyM56YD4oS4w5oToqa1yyyDqyL+2sJpW9XBAEwLpeH7fc/7EKCsA73GaHE92h3n
lgAoAkzCTbZ7gVE2TrbTmnno96RrLo6Dp/Yumg7vxDqmcIH8dPv2yy9BfyxgPiGF
Xg4olbTDXBj3S855bHNIiq691MQzYkZVFl1ouyXpvfidn0zTFhINtf1mSQPHTR6k
lnfnPf3gPMLXFz+aezqzqVWbVhVfG5+OHZPNdhth+a8VTcRQy1MhJumh5uQ6ed3R
3XBT6fwieFppDgPXa+g3uqPzQq6K1MYm4L0xgCypkZjD6qyzRBoTvNBg0lZ35I91
E1hUlZ5HuCUupAUAOMsJ3VjzkGoGrEdKIowTTlSQIXMNgnETPipcT3j1oIanrC3e
tzn/ihq2ezyzw6+A6FgJwgK26pC7a9cBTpWvHMZE9XYleE6n5lKMOzJPbUoCbbK2
15kT43niwyluGoMz7V5tLiRUbjwiXN/lt9Kz/S0b+9/qIDu+DNSbNfPkp46bu2kA
3lh5YduCgro69PVs4KNicodrpS81/44w6M75Giwc+evKY8+VYM6Vpli1hVIdhvaK
y2dMHhzTvFBPION2XiFzqTFWxbozT0Z4BMjWO2W/Syf/fXcqTPNY5Vv/TBKJ5QgY
ocAhzTCYtYw8FgXn/GCYQTHaz8HN3UmBNhaxjIXGRwBdWnAJNsByxllkNUWPosKd
1KDaD76csJGZHSsz+rCftoXy7v6311e97zjSbHmhqGyPMdFdDzcPqbPcPeUCG+cZ
Z/aSG0+dG/EKgiqTBjIQyo52rbltEtw3KvEqrI1YP6olwS4c+kMZQpHG8+kropbt
CMQbuXa9fF6YlIvcHCXxRQ==
`pragma protect end_protected
