`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OdeWiWHaHJX10oqCW18EEBZujuWHBxi16aB4Eoqd19kRzwR5JMGk2MWHKwtcIJ8i
3HeFFWPS87tAthejG43zsQAlWyldwGQgorVPYJW8RH1TYMR44IPSHty61ic0uI3R
bDEnha77IcjP/5OgsN5gnikKaU7S3u8DZh+CABoFV5U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48656)
7Bww39kP61NZE4LDwWREDr7uQKnE412bfUjhD4d4H2/OJ5DdayoPk9EfivEIU3b6
B2Kom0d730c0ThurJL+E6AfcJ2alZFQKeTHkIzADjRFmyuXDyjJN3DLywhYcHbj/
yktpkaW9mG1t3LuBN0Tq1soE0SO2vPbJJ4gXtn6qqN01gvY9dzFBg2463hU3j8gi
b/pnnf6zmHi8TbwvYb+A6Oea/HVRPT/rohZweY6ezwajVv7UXSivKKEzBoxEHVo4
QhO+oAULuMa7Gfm8sHQ6tWO9n8FYzIFnp4/mVLl4mR45Vyec1hq+HMe9NVOLZu4Q
4YWHtUK2NSCqAe2C9YSOipuzzrKkE8Od7sRGgfpFw/Wy199Q3MjmGgBka+BQguYc
ckofjvTwWLK9T94n5geawwmvohuxBPHmz86hQLBc+3D77ofTj9XKa79QIvhAZgk2
gtYK9jHOZNyvEFjEbcHkVsJnvFMB3ZZrTFJnJM4PNMmmN5y8GkVLH2BLMudZxbmJ
VFRlG3VYUQtLvaXQALh6A7VFYSRhpeciZ8JsjKcnxmNE544EEMdNbd4h7dw9upQL
7swj+RcB+SN0NZ2UVyZvkymUBRF+ZAhMam1P97rG/7zOVYKMEfFv2qJ+Joe64xZB
vJlBsGcPd/YIicbtYC2nxE4VCkfLLgAisOLBCsb0xluy4E6OJLT1WAG33gw2CGe1
SM9iS68i/4CA4gC+a6gEraT0ip2AVtSb3JuPxfYoHQRkt4K3p0a//PSeApHoDXSR
OsVRlku9ZNzGo/fIWwHvWhnwNji3Na6WPz29nyBD21hF8ccbdosIa3VNyoyVzqNA
OtR5TV5T4tCEdlOHyolgUvcWASZRvqrDrgyUiinEPzIkhBzSJ2DdOLiSTfyGgmXN
f1MyKGjHSx6MvQQ4ukGKgZuWvFe7Uqe//yFn2JDsHtZA2vkXYqERCQg7xMse3o96
QRpA5Cx36CUe+NTTqDj8ONbjSyLxQohak6i501sTuPcJfdv0XnMAfxYsz422wmlM
hD6dHSKX6wBNnw75bpeC2dSGqgNMb/KQ5BO3d5UPiarcTtxflipcccz7RiCFPTma
4H1PxsR2rZ9Rma954Nk7ysyZMZwnYtLInzWRKjIKtiePsDohhP6gNLiDxXexcNuL
IQKwnv1WiEL4DqUI4hAliFK8xY4Ke/KVZobm3cwBxIlZlejQkMDo5KvWxdzC8WAG
cy8GRhCKTHpXmR7JBNrewNfWGTONg1aTf37dq/BTgtrVNCJru3WFQ5A7fIV8Aaqj
a8cFY9ESL378Digickfz1pQDaHtPiFBuqpRezZXtOEEeGIbgJ1gO6QceLIh1TOyi
TL7/DSOKRDmdvFTfZrG51hxeT1l4PmIOHzFrLPAkPKDnhWkPcsIaqMEM0ypIr6yf
a8GT1jAUUvt+VbE9e4xo5VL/lHj8x646srV5xprOkX32X0FL8G96ou3aN/Kt4fMO
2VdBXlj8+dPwbjcHrUTfM5AVSXCA3U1/2U/MIxhASi6m1ycA8SjOzyrLumTn6vrh
PBD/wpDfuUdexiaChXUpxqPRUm2XxDfvMt3qAKMabbgPIMi7qRSCJYP+ETDSu1J8
OHOa93e5Muv2WnkAMyP8xDh9OKWbwdyL/EZgNLV5wK2GNyhDetoyQajIA1Cr4gQz
lr66w25sRp23E7GYX7mOxDvBAwjL/VLHoCCdleXKw5Uf1N/3uS7mV516Isgtc2iA
o6gqYfxKT4Hcd7q0BGsm2tYKnoz/4uv2doiu2Iq9TrBpNyp0z99BgysBOkzLnTFR
eusr0zhu+7bsGr4jruPjaBHLYo0QkBSO2WBrfdDEQESDI7JH1fUZacqJRl5Fjo+x
h7YeJma6KiThxu2LCqlBbCbJDPECGRzE26wp3RmP2Q6XWRuFb0zb9IbYoAesAIer
d+AiSOLspKzupws0NgIMQV+zjijUX+u2A2UiTeAliUE9EgBVziPTg7mRrBaxgnC5
IwIu3/5zVDY4TCy6P8oc7mkPeh5DNmIUhqEJ94RcjPdilWGVSeKQ0+Ow25wiU+40
Y6RzfTvz5nsXT9e8t1+tHh12afU9L/fdjDzeGQjjgMxlI64/04qgdWunkqpHZlZc
3mDGydtQr5H/fjdcscYCqDaZxzfIOfXIvofVpFSkQzXp5lSWb55w/fxPi6wueR0J
G+SfDek7FSS+OsBCQP9R21ICrftQygX7VwyGvhDWZ1qbuJz7ysZM+7RVbrLyT8m8
W/jutQWKNxJ0ZMM6vKW9bNLPbftN81eDhRYnN+AHPm588wPQ+x0rhVxNzHtmmuPt
o3aFXQ/z9XqllH6KZ0ZQItzzcr2pvwy/Ak23XlGvIrX38zONepMVjh1zN25n7Ds+
Gihg+hmx75pFc94FBiBPv3vW6+wRxtJjrfTDT9wMFZfKSUAATnoaRfjCu/cpYoqO
iURTerAimGua6QsfC5Ypj5nUUXId5OOcobQkSfBm7JoLiBsUjZrNho/lKMEeQfdP
gXGLJ4uPnSdXF0LH9zr7bKjHnIdOvX6pmkckk+BiDquLQLhRVa2pBLW3Hkl/qd+3
iwjFH1LlCeVbg6nutFsp70QH/kJtRTWYe9OWhfXdiMxUVBeRG/QNQdb02MOgu5Nx
e8WojU/OrlWgIdtqN5PVRe81Xy0e4VG3IQlBfH8zx9C49yIf3QNP+xkMdd/Vq402
XML+d/VECfjIH8bt4d1a9PB0ZmJhR7yS+eeZAWJfbJdB8Mvxy49boLpYNidXCpJQ
gPK8hoMyYO3gksN7MZmFV/mLvUMVh9t72MW9sI2EeptbCkJ8TTXs/E5/Gw/G08pE
uxXtzeO47GZFu6O4BS/MnoFN7DSCTb/dsWBP/OkAexKJ0y4neoprv0Ggr/AjqS+v
Jjt085hRXQyZi6IbGmoTJaXgdtgLOtvFzosqpw+QCKL3VpV93FOwFOLl/zhYe8/h
GJju4kq51PRi/9WbcmwiAE55tkihzNW6Yels4KkD3AnVvfDJQ303pDwURNO9x/Dy
H5CP1LllBOANW+v3hjYQTurwD/tHsMLp6pu7lAML0xCK0U7OlPn9BOscgInKB7C9
1cMEMlbO4zZnon0h6nR/CBu9ihnhPjoxhkivgvBvNFT82cQlJJUtruczoxlGjz3g
B40uLS6JiRjsV/vwpYDHcIqhAqRX4nonnhAw1rdPUsODWCnT7jqjxj0Uw3+dg8gw
5W0TtlVbJHym9dUYAaegSXhdz0aKw6ZvWm4s4HJIXkOUOP+8uDbYe7sZLNNqrtKT
rfPSQR8cVc7L+Ts3MYglNKGlTnaxMMo6dVm7HKXfxIVCY0WGZKFFqQXLDxaiWmKV
dbt0xvJ2K+l3vs2IJm4TpbGCGzrPB0GqGvjBS23ygjQK+YtVuE9kl3WU7RIPGbqc
myIe2PJ0Fo72PlU5d+td3JPxrkQwWCm4wuVesHaMvMOKxOEnb/CbIgWb1WX6HL+u
hjoKNdEAhqVOkhDrVTEyMer6Zo2915Df3JXFv4KdpGld6Nb+uDFKISVELk9TbOFQ
E7A5rn1YN9RcmHdSf/i/yRYAq7LfOdjnGpaXVJnRYA/HUyP0tff2G+G0cLWFRxfF
7uobyBqvgHOm1TTAk3ObB5qXLDPm1y8I23+2Ga0z/4QIcnhSWwFcFyUCKvOP/Pr7
pWxBIFx5ZY7fa6a5jzItiGZERv7iVqYc0NNVcHs8TvqS+A6sD5Sifdf4Gzl+iv41
2ovdgBm+wAdEGWhovq3gOO/v0etllFdzJ4mTzEfR4VPBE/PiuChOX49hqZcufb4s
Hb9B9xgdYz0UN9EnHF2NMrWo/yMVsgw2bN5AzY912i2nBBIqHuDzfTmy+QoF3VO8
GVpclgc/2qE6I2DLc1sYcyGhogasHoRx+Nv32M6/DDrli7LSEewcZVlWz+pK2tQj
OFnN7vGSlHIK3i9+yop8oeXp/uGHe4Xw9mXpd0JuIAVDb0+EZExwJNnZwH7herKg
KYt3eVSb38I6VTwS/eouQTK2XmBEBAQj6c3tKABaE/lmHg1OSPrC8RblDw97T98a
jVyIKvECsH27EJq7GuIyddto6a1UAgtG/1nFVpGsgsFwReNcSbhPPFlU3n4Vxxbi
ATTJN+kaouGli6N1aBscUwHl7zeAr7TCUtgrxTzimqP4FbwRSmurTPFbVgWbqXEL
AVioOmoohQ9cXWAHYDt9fIoPw3JpWenrrGwcZd/1QVx2zMWJhYGlIpRfQOQbtKYY
6NeppogtSyxz7k7UzRrHstnFgq+yzDv99BiLS+RJtGH1wtHFhsu7FXuozidvDgyN
IoxIkjssbenDUN60tS0JgFn60Wg3baMpikkb//FdqsILdLUwFzJM+59/EmpSGLxE
P/uk3zvMaFqXENzjpUD3H3befcK1ys4rTY2NJbd+kBzwhc5kziEceQIxHsIxQ1f0
tMz0pkQDUX+eJTGFMfPsmMmHQoadWlNMBbTJE4WgDG2GFxJTpBDZywBXx2UxF4Oe
t5jpLjCFxvKzmkjrVC96FyDZmQome1sdlxKI8VyMasmL/VjHXXKBoZX6bIz0wX2+
+T8i9Tya0jvvPLoBKGvbHmopImI/pvjDHi6q89Disd+asgqZLspZ8KU9XkG3F+ew
QxmoG2oW5zAua2Dq9EtmU7cXTUijjIBu/ImjsvFpUeMEd0GCXomvTRSd6RaLS3FD
O+m/DAxiLMByiOXaZIxXBoWtxwa5Nuui1SkLtKlOc3J4uy5zEBIMgpSZyDgC016O
EnGa18xCsiud1JFf9SkIyEYLe16G+xoYNvHfuRvzu41cgZhpqbWrPl5QwlZmD2vu
TUM5eTG6CDiVV9TEg7p7BwAQjR5n3+OrbyGX8nV1MI1dWlrB1FT0nwqWyYL1Z2Rz
i+BzGZz1hN2pMpQIDxscrpU22gCdWW7wZYM9ObThMICoVug42YOcJ/dEH6wBcBE/
O6rK4SJ3PqYtSkja7aEzGZ8lL+ZYMNVjvIYOYvstyYvOb6H6inUYIH8OV2lhrbi+
H7tDh31UfASheMNNSd9aurs9vDltKXXU7LfgLCvM++zivzAz9kPpqiXFQlFMz1qo
H226KFF/qGth5yKJDR45ZZfI5neSXE3hEngGr1K135BFYjLpJyzQTKdLLh1nVp1x
pjkqoUjy+sFFAnki5e0mjpdaqmO/ma8oD2OKq2EZsYC3m5TAevWg9qHvkFPZGoTZ
YJhVuvymg4gXNhWfcQwftQnw46j1WfmqcoPZZmzQMGnjRI8SgV6/DRfmFpCzWZjd
JUQXybwzL2hny4CAzNfZqTrMfaC9pnCdOcoX0RXzW1v0+PsSolV6La9MOS2zzcwr
9tLaVTlGMal372sxf2XJUhPIDmxK7YoksJVtsJzPpAM0WQZ+WyhbC+u0Vj+lccla
NbxVKBxUdtMZco7XAs7B9HWNszorI7uImXkJ5oJv1dZNAPrIXrsBxWk1xsgk9Cys
fcoZppQ6xMBp71vaHRXvxbs7jvIcgCt+rP7wQlnGLhU26eyHC+yo1+921FtNgVhb
M8MJjKlNYzihAHG0lA6lKt6gvNTQq27/Ph/oh6B0JbzDcXFopfIoYupl1hq3JeH0
Ken8dwQk1YUWUt/ehfM0HadjVqDNzIrMCf5nTrrmf6+WJVkbS2TdtOMglbTI0Y1d
C7sV38hK4NLuJwA4Gl9yoI8v4JKMrJseAxY5JdmxQ+JSJcQGQRaRkPUIGE0Gcqn1
CAvEOAs1/+fp5q0e/aOpQsU7QpZGmE0ppVkLTtdgMOMU9U4YfYMbFiLZkCWnt9N8
pSgmRp6va4ZBGtYXBrKzRuAo9NO2Hci5QU6bZfCAo/secK6NOcZD9lKAwPEsoPO3
0jMe+21D+c6sl1qgy3/fC5AnNWyph/CPPZm//Iv23BeqfYLWc6sp66o+NNPOiGvo
Sav3wF1estsVmGWYr1yePOFFO4+SozxQSDJ54x9t+7GqrjZlSDQgKXXBf54mPHYF
tOF7AhzhgI/Wewj93gafR1vwPxlgiqitkhKN5adCkV9eoaGK3bg2MZtFj4nbfGE4
oelfbVmRWnFOmZHV41HZuCCsP9xkNq2bg5/vxY6oehqZKvzt7AJc1t6P48+kIeyA
aOyL1LT3PD1Oi9Qg3/azl9aG9zQj90EfyQmFfJJf982gLA4VHFJhpnLmJycEvXn/
fRSxU7joGtfBdmRxuXZwKFU1vxjnWeZhHveUbJ2sq5koVCb+LgL7oTSP4/W2xVGb
NZhwgYcNch/60FHCQ9Zza8mQIkpKA0u/VRc6WsrBlFu+OcFGfKF8TnQcEWSzMOz6
G26w9lhlIJfqtlMkxshUdhMyuoUMeBaX9xjaukG0gDQ5tvGdSC/6xUwq7li6INvF
J2FD+55h2CJ8WkYCwOsuX/mMaatSkaFGY8lTu1MJWd2sdNpT4EWEQ1ciNQOzZH4G
8Qkyxsb/RJbbJzs6na2p4+XYLNPnfWFzpbFifNgM92+ehPaTw5TcxqV7eCwLsmSE
Gthpy3f6lbpFB8OYmb8/RRYBlPU5SbpOvKdVVLQGMYmjsBAZy5a5g0KCIKYsj8KU
QJpK20VJpNn6z0BprSZ6nQoxqgiZyiqB0UjgXPwwN90thwGviel9IvtZkTHxL+gN
bKp5ZXaf9NBrJY6g5ZCEkLGT2y7oFt9RktY5uZzUtnz7pl7G+GWLX0IOy3L+H+HO
+ceh6uC4xttW1RxYbuuJv/akAN5mkkXup+0iONBm6vNXaML/9Vix9h+qXyXCXPi7
Z/8D35gHyqlcZBi9VNBDfcqC+YDum/grba1JnhFj0wrtjB53ySlk0vbEooOd62v/
Hdw8k14acHqru1tUqW6shZPQKXiUcOp3/LBYu1/q95j7bFfV8QuJG77Cd3/9hedh
JUUtQKphjn9+1VK8Hnw1bN3D3ynwL/I5jvowAQO1yBxPmG5FCX/xqfcgjyryhAJv
RF3c9nCQlspohufdVKjeQFQw6ytAMDQtQ33uOiQ14v4BYTMtQDDuj+UIwqZJUnQU
Y9/94LBfmJbHtSMRqFGtGNq/7EMBRFhkhHvStYEjGcji5BD03B2SyL87VVwyYiVr
QG41FhgqeBF4w9l136WeEklIVugrOPDBVevtycJlVOKs+VXMxsIgaW/TfuGphImm
FKVgI2HnY93GrOPM/5e2/EFJaPt53beUZRnk7uEbdw7fuQmR5mLs7kcgIb9JjIGa
8rD+pcW7Uwqi45XcvOEZyEraGYTpoYOqBbPlaLDmlBGFtVXh0hKX/Djn0IhzZXLb
xopnpfPhcB5fFV8DuQ5uMagWMMz2Cptgi4HKLFWjKrW8m5PcFyaFuQQ/GU9UgIK1
BB32Fj8gFdd8iZ/vMubgztx4ZbpZJie2rs1uk6gVbEh72i3MZl5/NtbXldifQdcV
ksMWelc3I0bEEdEluQtr3na0cldaOxm5gcj0AefJlHXXifC/MNq976ZTl5IAZ4+5
61XKqUyKYeHt1GpnBy4DO5cixRg3LFO+AKJfwpWx/eMrAxkld9fbD0/JRpB0tKOM
pW+wcLmcwuTn7VLCZCN2/v5NLmtXIrUhnmoeHlqvyTyZCp4ICEzMM8wZFvCNSEmf
AqC+tfZPOVYWGMm3xIDfoHOkoflMfIp13uP/L9NTopYdZdyuOI1piEnXTgZwzsVn
0Ja2Jz0GM4A9rVnevJkp4srf0orqPpzYDYezoMbk+9RsIW9XaJcGNMxel7dHyVqO
Smdm0E3R0EvVRSGIioQMGajLwGB1PFIwymIdZ0CbaXB/MUkhmQQvD/BlsGXy2HbV
urQcrEDEWfIZR5bPhqF9IofXbIzHRu3gizE0mAyR5/IHqK0e68XFpVMeOB/3pV21
s2inwPEFB/3FMpKzTSrSa7SHYDyBH7L0U70Ep9QS50IIt1cHtQ+NbiEkAnbZz88N
5YF6UvjheBClU49bHmjEkBlrGf/MiEzh+eT6FSJc2E7Vi8qFrs72AubU0QsAwKG4
VmWGNAgQaE3VW2NGH+HFwth+2xYJ4cDoqmd0Iy0TSi9gKSQuGUQIV66uzO/ZzsSK
rJCVe+tl03C8XqmqXFvgq9+CWOjs2rCtKtkmo/OuyLvVcBsUXGztAphL3UGQKGPK
1oPwDjpDup2GzQCBH7XrCNZhXINfEi+AgMcoK/9qQNO1tGMMjnJXe+NbYBKxuIta
5GTJ+mXNbR5cX0jCdj7nHHwtUCv2LcfyKvyf4F8XpFUoPR7N9Et5Peht/HU+W1lz
5rjb85TWPy1eSlTeO0/9Azn2art0eoG947NE0z04NYugf/5eHyH5V5Dhwmx0yGD/
+3liU0lM1TdoMfbwzOIuV2i2fcx++qF9anYiCqv/uC/NAkyHOuDeF+l5FFX7i+br
WG8FqTIEGpqnhvAay2Wcz3a4trH9VnZXwU+5xvfU33as8iQItN/KlM/dGOPJnfP0
PtTB0mtqSauFabfGHsiVGYuMXkmpmKPEJz0cH+nu+amS7A1mMDB0w1LAN7rFQ/uL
8R88Cgqz/MawBJX9xVp9VEovR5XDbGKvU8N+aL8kbdPei86Q6uZzAbZ+899jI5bf
2ZfQGrJUEi0/T5OAnmFfO2rz5gj58vbAnQlQGWP8ZiurrPFbP0DWZCULj6AXog1Z
k5KcuQ4spAZcHjMFmmWWIfkBS7GodfmTFC+9kpvtIimgC91rL1zPCcy0r0/Ou0ly
a3hn5bofRekAOOiiWdZcnTfbGWwYsDR/n31S0GgKJ5FBLHxwNTET2LNkBGI/8Xum
ZSyLp8qE8TfSUmRzusfjbuC8YYdw9BQxtxjRwZlPT4mZ4K3HDBq8Yt40IrM6EEjs
1b4MBnM2JewfDnGgzBgmdQDKKn40Qu4ZRqyUglx6jAIamvxVya8mO5TcVmMe+qVI
B720n4MFyx8zuidaMZ0lW04Xx9cqN85PxhJ668nvH/jGBvUkONJQJYrcSomB3wYz
5bCkbSaMMSXJoxZLlJYN4XtB/vmzB9WA9IlCBkBFiTNdARqzztyn/NsCu3ytwf3g
IPTKZimO5J6aNVC5Es3eYVoGbYk8/P7YGjwqHblR7MREoq81Zkt3U/+Jg5ZH3grk
fhCs49l/Ka1/+5CrkPpfvWV5gSvFg+Dez9V3Hay6wEw4B0iug7yueWWsexEyH5j9
P73Ar4Hh3B/ZruWLUgkaP5f5ItpiFeQPPI2yyCPDccCxv3y4skVjeS40cp1+RPsw
OO56l0tVeQLzri5ox9zLacg+5RmKHdE28On6p70EJ0/ogfOm9IHtblixdRWvnQmf
UQPV111+2qW/REPTa5q3g7IKcPNeC6ve9IQs3E8bd5SkiOl9lB5VCIKreSVAqu5J
JSCu994j4ODi7isq/V3q3pmX47oY7PqLVkO8z+tLzyBMjb5rN0YaQpjxNZ18yK7y
KimmMhYKkQBdEOwQJyRO+7RRk3PEBCW73160EJBoperbkhSCKEnhZL8uwXjJAPfm
yegPKh2vVf7P77IvdIUa+ONI6LFfXcUeb79BoBa/HoeJO/T78Uqe1aMYmWfVVCL/
iMjGWZCRC/Lld0qBBMqxkDp9cWoq939dpr1moUjDoeeOFGGWryRAoI0Nnv6bF/Tp
4Hqa9sPkrSaBfPHOCYssNsKN7yM3y5bxhKi0jCrf0Y1m2AYSDBG82IXPtneSHxzU
F4u8ASxlZVdsBUzaWFXcnoKTcFwyZmdIPd/Y8tknaf9rWaqBX9UwCJzGP0LtrK9X
TIK+2G9emrN3Lw3tMafG4JlmUOK3l5KXIL2faLMQv2FvCMNjkhopX9Nohqqkw3Yo
k/eUFgpIGwXeIqxA34DnJBf4S9zBvUeNG6SB45MGgEvnCpqDpvOVTVqilfGczGRf
3xypWHH+xVL8nOm9JI2L7zvBtKYpWwpXdk6aerIrIUVB8iWRP3f2gfD5GLlzt3cS
IL1UlfhekPMF5ewr7ztStaicUXrpFP4IMSlLn6LJGfwf+YlgcuS7mWALQSMgYt+A
lZG4A5z33DS7DnYW1VES9jM90xfpeC/As5usvEfXHic94eQ2Q1JVwyydYs42g+HA
1d9po6ofBJNlvWyQ5FRcX0sUScHin36JGeGWSVnUjXAf2MVUkdW6kBrhkIr5SOYQ
mFNP3U9nfNhyS3+9icYLewQGrZRT1tAtPc+msH7hgksiDaCrpaShq/ieCCbXg36x
41B5yYYhi7nZU34Q4LcMb+pcfqvRFBE6beiMUG5DqW1IJ0LeXk3Muvw1jxsMAbJh
nVnks+V/WrpaB6g9h1l5XzFPJHM4AuCfCOyxuZlWADs3m3VldI0SQ44oqb1Mwjv2
83eJko+8hBSvBB3HhvDvyVJ5++uAf6fEgf84CjK4aFAiwGmHSNpFPvBfYvpgWjng
lfUaKxNf5GCPX5hccFtkp6EQQ51T5UqE4cBBUeyxCuufDjbVm8tOWGp+8mAp0lgS
6uAs9lKekDhEK2/++SBwCm2qu0u9ODJGvsuwrtYAlQihM41lYC5uZPE+rEp+PiUc
lWRJRL0VMezaLfr05s2ZiQdBarkm/8YpBZl97lhpLuQMq9NHtj8KrjoxsmaFMsLA
b9hIbhEEf8+c3Q/ltNflLgM1VqN0ZPDqu0lnmCnMsqrMRSNwjBWRKnBOZUKiRbCn
uaO84iyq4qifWS9wZeYVz9gw8svUnSYZvGBnTBDw7JTF+CFwc0HgmkcaHoj/X5m3
0RNmrBw6mIRWLVCCoNvQM+q8KUYZXnNRhg1cRQuAyWKcVOzw5n0il+UF/4zB5tHP
veuK6lTC00hFKIbUqT4KhcskxPKzNJT6KZfXJd0hA5SO+mF8GZBXNWH73FkGLmYY
OMXkqU5lTXC7BWhVEZRBN0m48dg1/VWvKJXh4VmdLDSZN9+KfNWL4QMeSUB2YTjM
dDIP8lsfOBLqnsjnSL9fdduu1L8XLzxDmCyLSrjuLMnFeFlYOg1xMJdCM6GArH7r
6Z87no2BDWcQcI4cxpeIxx2emvTqccFKhahp22XiRjWrE3VHgG2wg5rGH5S33Uk+
HBMALustZ0arO9T/UU2SNIppTWRazwADa26Z5y/TBPOrBMP72/R5YpUog8Ck+s64
ivpLlop0qGSY92b3XcPzvXr1inpUBWOcG7PnwjeCKUCfo6m9nRLQkmOYkr6ZKFMa
bOhl3BaXWeWTkLKn66+pcHG4Moi7/PwsqKGugkigH8zV8DJHGBOSAakcWzM95DV3
H2yDBGXhcqdNroMG5yYYUedY5FgCpqsG4PurtCubxvyQew4MBOrjD7bm9tIJ4dKF
rz640vjuWRmatSJUpNW4ZT4DKCbK0XCWdPAmDFAkoEubS7xxhlFGM2zEFK5/i06j
EhJg3UN7WhbWlV0y8Dupp0oLXq/HkWAV5ZYe48o0X+717BWnYgQTrbvJ/FAuUGG0
1/jF4x5qiAH1Uvd1sNepDX65nisVE8fk4lZj9yw+4nOvRQaYiNKadFbgy5oYKiYx
CD1Mw7spe6H70eYjrcfNoQegu9AJnYE9tyELGD8rI87/IHIm10R4Axrrhb1uKjVa
uyK/cwTcZ4N879dLfL33FC8Tx6Wn997W55s4NpNArOIPScx6YUSfcZbmcaiSu+ln
Za9s8VP3Q/arrAhXftAlZrSwkCFBQGzHXOxdYymb53lixHgfKteuH4JJdXihIsHq
UcCxlVGlRwtTWonzLc1IJygkUYTo3+M3ts1JFaMNQMCo3vVY5Td6tSu2sEIOi3YN
YlJgt2mlYJj9NRPosUZ9mJoGPShhu0RS/T7GmkVBILHU1zqXH6qCeQRBXeKKKWHd
VwYKxhH1eWGNd9X1XwTmBfGv/XMMBjoPe2i86j7GV0wgy0C4Khsv3ufsp4eY3Vqf
NAShZ8WxDKZiB2bD5q9ELFliAo8BPghcFeiXa1fURjVNwtngDSAaugWzZBeCPsHG
Ys/qN8zDSLRWQ4Zk7Zvv8uxwJ/nNnsFrqIDSxFy3Ycn4krc4CVwvQjIcTZWLjii9
tTgl9foBVqIfmqe22c0pFcFyE0jJsWP49WksJuDC7nfw+s4A4+EjK2wjb0Y9C/Io
drQcvIMcfpcqoHX1+lGH78RtqzHhJTTI7WyG5ZbyoTAyamIeoNANAoNlflWu1sBf
Jfp4j715QQjLyD3CUgLCNNv54VQMYiAK2a8R6o5OmPSpoEhr5JR9Ex4FKTHIMzpK
vkrtNFi72oSSly4PzJ12C1G8H+shlxWUWOW6kxr0Zn/d+36wh3QNKYfoGoyC9x3f
IEUw1g7BWox83b8zqtZkfcJvNrgfa8bllwXxk+tPpZZwhHMLKjbu3Uep4gCXnKvk
qVRXssdGAYpObzmp+oXUNV5oSg1ynqsiLiHK9YvP0SuBjjNgnvT75S0rXtUnw61i
5k6d8u0nN+1OpCnMJCqExEUK5ECqn9dXeFi8ObRKrvqhInxcTYzkczqeuJuGoQWN
4cXyly2UrChZAYCwjtGWycdtrjdn26mFEg+V9hP0dDlXd5tOVyxNE6KCM/jMa6cT
aB8ibDJ9bIxGhXu4X0Y6Y8frbkbWWu0HsILghKicQAZ95+WCCcm0gET3JFqxtjc4
A1910G3eS0StZKsJyOujRHHZ4quwbp3KiN+MOT9TAcDsFftOHz6BNsht4cS3ScWE
6xH8J/7yPPsRbY/Ktub8XfzdCOoBKt9bXf/P+YLaD5WYXj9Ge2k0/P+J0WWlz5SM
b7fsat5cUqkrah2WaxmTiyyGLq9k9+5AXrvGtJYm+Lh5Y27HHZmW3JanV10dxq3g
FH2DJztw9LZwrUX/SBwuG8CsmsVaSlu4Y4GqmOwYklr3+75+dnYO9jm4dlc5uTgC
XAttAULCdV5rKN++x/0huG/92deZ8/JHwRvNQK3Vb1FWA/0nsrLjT0YSaRats7MY
9ObVYPt0ipFOZ36q9Pv4NBgxXNdxh7+vEmZmGpzQXml+DzWqs/rXD0NfWPCiJEkH
0fHjkAW4gvsPMvSipRelUDnDkCnlu+hGnbg8skEvIdsyFWb/zxqhm/9kmiJYtj/5
8hM5j+2tPrE/x03YhsVx///0YVm88qlyLDmlnmAYt6fe8b/yHLNsxDzVHbnteSKY
BThxMV385hpzzyck9okNAbfWz379fgGo+YfhP55Ryh9M9raIWYElkvo/+Uzdm3UO
fT3bHJxE5pBYvDrTQ855NAh2srpsl34w8dJMrPBMl4wd3wfE6SwiProJ4uQiY06Q
ffpaxTKSQOrKQjahekko+W6yE4FWyHwJV7m1rCbQQCV0k/644nzfjLG/jeePBAl7
+IcWOnEUAanPLLE9vblKMYxUYSFUdXM6tPPJvXrzD0nKqMZeHKH10exii2p+GqQg
kjKRE8N+IrBCJ8E13w9uIkQbzFky9JH8DgRzsQFbS8H5E/BlWR0prPz+pnceM7Mi
EjoPoEK9oBxtjTm7Cm6oo/GY8O1wPn1TxT5AYCv73BAVq8qqbd2lCYKh7XcR52vi
qrsF4THSVlkW23ycjb/WtNDAjJhNKqn98CTgPdITAOYFyQHl20Z6SE7fhnWrj4yJ
U5FxC+cHeZ8+R1d1w8APvwAjm4AgPLw7UkVjvBzPHKXFddX6XeRWb0PsQc1ownBS
UsU44RvXLeeuSPybh5GcRj6uaOAfjA0cvaWcQvYnXSIT6WXk6623nljVLrPnCe38
vEtD0f46YIVl9WpF/ktcAL7q6MC+vRChJEuCEtcKsijy2rNwFILePCPr6dinjZfq
wAHRxFyGOWD4VUUkhVEUbSIyvWk044xcjF5wTGmO22xYd3zZh24DVh9cG3Y1gy5N
Wp64Sn18PF7eOc9IvqXxwoIoVS4j4Wgwm2qoLFb65gmK6t9D+dnGb1/a7b4rJ5Lu
wsy1aG2fjMJ1UGw5yYDRyCA8LS/66yEHtx7vElDo/7Cy+kqR0CIxu/SLwF5dBAgR
NoCy7H81x+b4Ut3rUw66P7vlwXcbSV7oHe9sMZogdeXSUFdvhpy4UoEXFY1vmQ2W
bKfr82O8xWIJaMnw+GAhQrB7/4Uc2MFkWXGn5lxKJg+97bCJZmT9kVgTdNQ4q6PP
TZ3v4eGWVbRPN1UZEy8R4feZnlr+6WHgc9h5n+FqUpDzq6E/CiPz9IKNsJvNys4A
dwxLtnhVrw9XtjIK/m9Zk80FBqSgptGZwR0ZJ85Dkr2T9ROljkjOdLmj/Z0v6Yxm
LYp5Ab5vIhoFddMPOY1FldQ4L1/cLrPl9+w8rmLnxLShTGlgEcyObGb4Z222bhRx
VvqpwqzY8ojvdRTAeL/awaY7rqNIysxUKns1fjePgopVur5CdS3yH0pTSBKMWS+Y
E+54+jmWLHwMR+gfj+YbFymj7d9aZgjOpQd1Ks96vnh95ai3c2QFkJlPWTYoLXQu
bQJYOlzj2+IGrdZgaofuh2DO0tG9I5s60WLlwDWjsGiZ3a0x9chHyF0H50Ysz9vr
2b0Dwc6dErIoMxl2fNGCjFwaYR6PdQ0e/5s7TkpGNZLTEZ9ixIZpIZj5gcCpU2Wu
Rtcbji20wnXJ8t+bfDG+y8EppkGTGCklg//APuRwR4xZYq8RaXGFGN/mTvRmBg5r
WldpSsIDluwNCZT7bfdtCJyIWedp6HxHbDcRLpvByuvbplLutJtzZQmaqD3WLOY/
Nc2xx36OuG6m7cmUSbnvxc2FO9UZJi34AhIlcyfZ8XUvwmx6eiDJFFNhiXGIhGwl
tnhNpaO6pZ/uGXrGKFZMMX6szGswY0qtKTDwM7mE3qHjjUl7GHjR8BczpUwxhkCS
s+g+AsXgPZoigkkO8btUUxE0jXlWZR1oxpTr0lT6pMcA7bWM19TIq2HpLugakwgE
PZJuXaiJ9b27uPt5wSBb7k+FBIVSk9rR9kVPGSHlEjfOcetdDXSAr9kVfpH/i27W
+/TyGQoBLPxUmpjDqCLQjL4FJbtbbQLdZdl4RIVQmXIcHsIuw5YrxXM1uUxnXSoq
ybxI7az4O+tBmgJ2BX/XAG6YYP8Kfba34190BF/tkgesKwOc1fRhNQjca/8YQaW0
Li4pt0+YOieSKt1Pdcrj0wSdc98BiikUE/9iBtehRImEoC09qHzBSwJQeFyAC78M
2ah1SG/T0d0iolG/OKe20nJbPs7wPcyFIdwR9jvrr+3ymlqShE9LP61bMoqQK3Yg
YeLS/eVMytj2zrew4ZvNLuPCFD+8iZugeR3JbFU9SttcFpMHNs8hAHxupIWGRpxc
D2GlE3vuTT0E2HrJfUPoAUfrnirI3gzU9cMjnP496lR80RhClyDTjjp7ejvZLYvN
iy+KNUWekUdRNfWcD95hQaSb5lsPumunAQ1SbfRZf8wCYRgVvJwY308ok1wRatUq
EJHQP+j1cxq8Ls8iH8KCyoGKLakx9tIApijpMUuHrWYjoe1BmzXLZMM3yqvVq6Bv
sow5st0o969DhqDvNcBQFwX1mfpjAxBMdJDO9XfQh+r6DjYvH81Lnz0gave9ZG9s
UtU5gAeWfXDg4Gfw3qdsIYmXjP9MoZMbBSCLP6mD2y7posLOzAhOa4ALBuT0s1SF
QcNQY6VGQ6ZqJjQm7Xfj6LNYdU700pftHuHk1z/QzT7OJc5TVgTYbJWOlFt1RbzF
IXfo0ED10HG6qhXWPMbvyF8WQMSAWG/Zyf/Jj4OMXNVk4kz2TSyuPo1bEmTUB94+
7TZJjTg1c7Vaw/mH9evPK0aRFdlBiQRsUzmHHEeSm+u72HVuBsuPcRmM/bNklyIm
Bpy67WhMdzeYXiOFOLOMuvHx1ZdBueW8ZZtORaYKLjXCqLHZ9Q7hGlknsl0XoDxj
3q2FwD6ScAxljxnkTza/svBJXr+YjqH70dvKXMJ1T0lVY8E7tMVgz0fVdaHQqNGt
WjzNkHW4No5ZSIhTojeghaGIKQKkgjMwqgomtTqQCgeVCYJrAo673dnPqLzn11n2
qU6nCYQbXJR8ZN3dJ8/SOOgcplP/5z+TmvxI2dzusxB3oYNEJDJ66dzEkbyLz2wo
UY1xI47Q7TErFFzWDYOPfZ3SaBcM7O7NgXHqpmjjAFJ2A1CDwO3cxjHdXxFQNelq
HpL4qmwqbW1GtD+TTMfbOkTEzmHf5fx6BpVdw2k1JgA4Jxni4HcqEAer9XiUPxW7
xWzMpqK/XKluj2VVB8TmmmcsZ19lP++Sv3XwsKkGTw46zLpFKhyJ6RDQ5CxW9Zm1
2jBkEjRXCZ33aFPsallVazHSCeq+YNXYDKr6hHUv/rAuHs9+tSciRCTWTJ4sQOw7
Xpcz+l0qp+VJjKk+t30ohfzGZjLLYRnH487Ee9rPxwe42moYly8rJDrrPSx1jl+3
6wPuKufWVhCj31IVFyzj9MlnPVrNe+3k5cCclsFNAaYNqQDVa3vyuDM+mqoPzgQa
NqpSnSkHJtsDjBHG+9mjN2q2grJaAJ+5Fyjj4MVUkdK7O6dde51PzSuU0g0mCu27
D7JDtMt+EJTQUkkjWqjPlHEzb56JgwDRcxg3iU7AHI5BT3iaK8ufXuGXQoYk4Ze8
MRM0FwJQzHUSVokKV2A2Rh5wOqk3yXhAMZWZBpwtQDj574qP7rDs/hQTccMhdoHS
KetZ/JEBhEBTE74gdP4O7jIXo4qFc1Uv/dEw+sfbCRvo44KNHj6H8f+dx+E6j9rX
vetTA9Kv21ngTsOiJiS/x34f6ZR9g2vDWu8F3MbrLfC1ewBYUJOmTxFN6i0Mx8Gy
IdfM38uCgVop5rpCo/IAzOhCL0+wrCsnOXHjsQINPqpHCFTwOU3+Ah16p/nAwqvH
E2fxWBeoOaPo4KsKPUI/Bnx4WmsV17VOnESv06XcJZ9HTV0XHFtuaJVJq/U0q8fd
HUlc3bC7ggwSc0Y5B3s/Av476BKMQx1tYDiiqJEZqYbvW/i+xrTLZVjXzYmeLLrM
IYTxPZ5fHT9XxtMk+JsFGa4seOkkA1/PT0cxFHC/TK2/oBcuhS7ZX3ViKBWf/eoU
I4jGvsGgzAP6fZQYOZmCEpmdWzgMTs/ynQJ1sWNfLhF7X37HtI7jDVBN95oymV8w
uyOQkWxBrLsyrFKkNij9VWHVVvbHBdee4BWBBGykQsXYoOU350mb6PG4gtq7k3We
pm79XmaDSqc59tNWKQSkNL+AfZcwEmMQMvDBi0v8K9kK3qFzxP1n2n07lBXGvvpn
8iLy6pcuji1wfeAWn3ReSENabT3tw8Epv/vxi2j1fhE9UpgRkSwf5NQOoKyiS6Ml
7c1n5DxcrGdwBTw61axNUHmLTCLeAhooXE7wBScxXZGCkWM3Ju2wggS/LQeWbdum
JnSy4mGFEj3Wrv3kcifP5cF+WP/4tjK+DwnrEyZrUBTPIsGlwZ3lv+IXJmIUi7/9
0mTfeJXmicQeGHW98qZpgHdKQjOJvKHFJwiPfUOPTJsvuDnAh9w+88iSXSDEMfUX
CQy2ci7HXUEIbbOkEOoangc0USZe1j1VeKzFR1pCCiurvodVORplzJANE3YNUvU2
GyQeca5OYsNZ6zwVoXjaSrUdsfCIFMA4Sy7wPZPiwd70XFVgeQ3UPA1JTgeVmsgJ
NZv51yQtbMR91+wu4FVSd/eZpDGL3E47L2DLpnzSkDOn0xxC8ktSwcorReiVI7tP
yAjt1qG1BnlR2bN07EI7vyYrqKeeCndBRCw8IuCZ8N8QDMBvaRsvx2jN0J54kjtz
W3jN6Ynnc9uKSVdMKInaZ2EJX4bKpBCOvT291ynDPBitVPt7mrf96wKISAneEhHe
d32kd4r+vibfnH7Uhqc9MmTi8syhq7mMluWlyzoZ64JgHj9PI/X53yiFiAHzmOXH
bKhb8Z0g7SJghvjfnFf7XOl807Z8vnFmDh48LZCeKWCQ7jHxDB5G0FsiTbcyBl/H
oS8IAEaCMztgCxRWO9yWnHvUAUzXPg4ILPR0kXigaLvYexS6XPhf3I6V6//risjd
fqGNr5pvKd1GV5J1kunByi/dfIHCBYiaD30mTJV9/0D2OnAFIOtvzwKKiUDwN4tQ
lOirDb2AuZAsK6jIQk97TUrFuduFZSTVBSHAkr6fMc9bNUCbKaMzIdlUSIn2cdxn
gsGfKBff9THb/6bVIfieZhq2K7uvTYwLBj2qIg586F7e7jIJqiK48KE6gOQb+vzD
MAqjeCXpV7fAY0dlCp+INV8jEHjBw00uZQqTZ/fjwXHQIRx6wn7kGTHdCBiCjsoa
Y7bXSyNhnbhKM2VOp523Wz6A9sXLqjw2aUjWITY4xgfH+eD2zWyZ6RYlAypOe5nh
Of6ZBr8ebEVH9f1Kdcs0vSSlC14yFUQIeTH/V9+7/4LYC+ShvWxqYuNAjnMDxvM7
rSx3KUUxS6Eju9Ps9IrshciR5YI1I3JMFHyUc+o4Y9s5KkFIAqCm+JXAUaBIOEpS
jS9xb18rwkOlo2MupjxlHg8nuO0+jCz7SY8FuxcUjV3LX/ZeItlT5DCjBGk9uv/6
emlzbq+uAYCpyzX/GCG3oAU+MM9bKWM4D7SOunjOLUlOoZAfygAazabsXnvhgfBZ
Ag37aC5JwQCg4tNJYWvY6Djx4OKAzotBIdlv5NFnjZOjEXs2MGJPizIaQTqVPw0k
qze24OPoYqtQBKv8Jc9Yt9tZxK/hURiokDcbDY+FKN0VKtgpi4tjX2WVoPBSjUil
pChYE/qwqsAq//gWviNtwUCWYbkMAFZJ9U2wXHi2vkQdg+UA/Rc7EOEMwTBZNOV0
jQ78uNAIlloAN1i4UUJgSAtNKjGwd6iddD6OTzzN1nCCgPuGstTibJ7RbYKwkAEt
eregSBLSEYbBO5Hf3TwVapNmlKt8hmzIswMqvyTlzHdru0OtP18ZWc6V4pKBRORv
1F63aUJCmReEEH4QaCorM2diqnOtbqoT5KJppVQcTbRKvem5+Q1858Ztv9kVgwic
T4SrQVtmQi/u22P+IJorqS4JpfTFbbkyN/FD4Hg/ItU7Prmr4m+v1nI85z9VyPJC
lmQRyW7O7owarDjA3N+zIKyxbf6qJNSXFP2DJNsMV3djdffzeNSeky/jwUxNL7uS
m8e/SSfGcolOZzIz4K3b6sLKwD+xT/pNAwZsNd/ZpJEm9ARbyaRuQHWizgNib2k7
kZ1Lmq78OmpG+N9I7zKqaMXl55N27NDOBd97JK8niCvLaZ1131GtVrVoFsIkqIDf
vHUn4ExUs32RvJbkst/8F2J7K92ffV7MI7JMKgoewki+YV42+jhdeRjEjjsFaMlG
ipTAXFFjo9N7CBoMYKEOK7cI4tNCMdYwkXzsAb1ahl3TUG0WVuvxWyH7eKwVn6kO
8ohiKyfEInTgBEbaTfiiPA9ezkjzv8kkxRkAYHtMfVqi0JR5OH5AwkQIMA6u+JWG
4ir7OwHu1wn8YXE/bpHVyIrrf2AgF/JYzSszCzqZS8cQA1TS2EE5JV0rPtRY3FtU
QYx/rHtJBviTsBxT2AB9H0qDBvP/NPM2Od/aX0wHvytJTtzmfTldI3Dl0UMQ8Wvb
uMrAgu0gvn60dBcgBK93DrIYBpUk8k7a4poUWYM9wJAC54fJISfIUzntB2uxz8NZ
VFyhCAcHXZql/KVN8Q2bTg3bnjDJRJXyOEJfnQbq7W0yRNwzWu1so101s/ohd0gA
3bEAhM9nL5HfW1OXWvR6w6BfntkYeKLi+dc/jUa2O2X0fe0+RHV83+K5cTUMo/KA
ZUnmv/Bg6kexJFrZt08nsnyuUXB+2VCQbYwPypXiqeLdSj9/LgyPKRtv4qpqjPPI
9WrZd2x/Wy2a+yy1nOyFAV2aLvhzf1440rHh+0+2R1eHd0eug8lXK+LTmxnOzyYm
ykx1sGlv2qRCOjbwrGoLzSyvygt1qBrPAGprGubbRbfiMggsfg/DfymWqhbOW+8l
i/1bHxbK2YrI+Q2Z4FWooG77Ur+CBizr8jSs+3Q64AVgdrOjTyF/LfuMRMh9dT1D
yhtrEtaAStvPDV8R3jy+BrdG/WlTzYy6FgXvzZAjp3U88TmF6m2eCZpf1xNySnmd
ex7aHawtpRLbMaNB7iko1dX5emJMl/hnUVhoQDk6CFChT+PWfvftmetQeRvjfUxE
n5XFDdcXJUwa21d0nZqeyBnQl0MeWAM/hV1pwZnIjysCPTHkK1yFf3wgemKjcSC6
6h/LU33NpMgIerrUsHmq86QgkhSw58DybpdSAPZim5/xEzVPTPdAbipmepSZAwfc
x1CthKef/EwjrlnYOfAMW/BUqos41eVi1TtzukSHtrz39MuPoTX+Ry9jFNJ+dvHb
SoEqlcBeqwq3zfiMzpiS6WhUdQreQD1qF6uiVJVChfsrht6gQVL/IsjxW4NTbER8
qRQEnSAr+rwTapVrcT01BE6hMe81cA8effJdPdPwCV9FtnqoW2iUSC1gEWSN1z/f
GggVKy4baITvA+wGGnznA/2IB5GuLq9uQCbqmGEF+8hMny7i3cuxivAOIdKcLSBa
xwz2qbuxWB/BEYbiVNEEXJAEIsFvk1hmJf2l6I2PYihlNzs7pHa79M8D/VOc7+bb
BjJyutU4doEgSZvAnEirFj7gLm3XKCvi82B41fjd/Z7sHTov2Q5HueORF8HXPC30
D0XQLuYc9L0jwCpAByB9VWMAhzflPXnZxAKku/imojv+1HrHaW7oZFrGUWtjbcir
9Nekzuj17lnnYJ23QRZ+1k33OILbaQe+VSi2hQYH+M8NeyjVUgXD2QfC+t9WTWP8
TnyGIEhD56yOyqoSzMU78k5W2H22avLTqr0CZOYSg1tXRvRN2T5LFX3Hfjf5yKPs
ZWX16ALLQBImuVUmkiOsXsqzwE/IwYGiQEKl+fcwo74Gdof1vg/K7T/kiHL6pQgg
qPuG8SkWxVMFHQ1uK+wvecnYDe/3lFeiu3XpdQizAJDSt8tmGDvsxlwfZLQ8gKs8
/2dGJ///SCOHyxj/9wM+CxRF6gsTqzGgPQfeX0ZFBbc8ImaNVD4uIHbWwIibEslx
TjBdgi/yQqvna0wK1c4f3lGiP//pGZEJwXdSNiigFMpjN1+yidGea0LjdJfc3TCk
9ekBH5+M0vl9Wub4KT3I8WVxXjXC47C9bHrIBS/FqWAI5H6EOfFG8T+fzzG4Hv4N
MCi5BZSFWJy4zcTuSSxQ/k47SrAKpBwN7GE5MXCnZ7Q+dj5qncU7jw7tYIuA4T7F
ECByWTUGdrtjzObO4Ud1DjGmorrlTa8RNG5W99tynQ0XB0L5zuq5OLEL/lB8P5tQ
TBe844tPpPT1k0+xyRKdUahx6+XEJWw5UPd3L7vz/6aQGksl3IZGRogbzYlsmCgo
+Shhx9SzTG7oiJiKNyPQyOIIETDD0X8UYB69YCcdWcjFGrPlIf6OEyj9mjBhQ22x
HAVH1BHQ2+bG9vAcVVj1vtPT5B4gsGW4Yk53gj2/h7992hCmafaJy2+gDVL4krF7
usWJFgr35XpzZ1yO7jI/4v2BC9qF/Iiw63QGpdh6PENHrD5eYAjurB5QKqO8e8Ug
nPelx2Ok03gIanb5a/weydB6sP54K9adusek7JMentIxNnZXBGqiC90d/lx+iLlO
T+eDnNU+4Qd6uUovVy/i+FbGDCUQzufD8Be4L8hPgeXqEPGK2NrGK2IhvYvpr/zx
iEUkIcrO5ynEr25CELNhFrW28DVpjUgqi4wZ7dxNu5iVlHAHN8+WBncd/QUTJL4D
lC0o/IveqrI4WugQ+VIwvMr+Kq7bDsIvRSK4jnHMK1dIMd8APLdkWCBmQ158fWDU
AAA37aUv3r4DVMQYiSp/gBu9fKros62cyNCxxXC74yH9DnZVoJcM/T7fe0aY3vR4
rgM9Hzfeo5ej5Nd6Lb9vyFk+tQqeXrlbRXBn0r00UBfj44zF8fIvlmoJ+Yo1ILrB
I2E+hY2KAa7Sb/Ad1oUZKK+O24EC1cwdhXayKPlnE9QyKcvuypkhnbd86gaic9on
dv7r6U/4I8da8CDqiG1TA6anM7ukMRRZEZW2G5rlzhTGxKlTg0VUVla4I5mqRgAu
y/qJyJ/orbkOAGYy6hhEB+tZTcVe495VfqLwRn4Q9aWfG6zOGv7nfNaBdQh4f5I+
7z915bYQXelw6wzoKtcf6WUol+f9bO6IGy60/9Y055XLNnY/dA7XlwOzG9rps9jB
M11DPJRoomgY+kiTVKIm0lO7/ap4tDbmLTikDLvnwbj5yLfxCcmbux4pQ11k0O9x
C0NVQolVyC9PuCPES6hngxKkM41nVoXbV9ccsnm3M2m+NYKuazV+Xb4LBd2k5GyO
tDX/nxFgk5P4Wej3mDa5gME4EAUa0CSCVymAl9yI1G3tQoyjmqAJTkCmtcclOTf5
2/Er4WgzgghnMqzNcirQSkjrDgo+75m/O2ObfPE1q+z+IN4y3JTdsBwlnMtaxJsF
8haE2C0ScKC3HHFwxOsm9hHFbjkbp8TcQtwhbHISKZ2wvAEB2eqQKmnn711PTAbg
UULFwKo4p3jzDWuYSo0IF9usS1+lCVRqxnuuAFkiGBPygnMUDGzKXs7Wp3lyHxlO
oFaV71a4u+AcBka3bX3clDp4nEh7CiUUuP92OCgvrX1xp9Gs4OGDglVUZolSNsex
WkEWAp6PaabnKDldv5nfz56c2opdySoWJEXfZEgtGyHOw8PaW6H4b3uKMzMr0rUl
vY0iSrQ0b8zBJPQ1XqzDHUHORb9BsIv9QrzUWQOoB2R4a4wCIQZ11E0URbkMGhE9
O40JbgTGToX4is/1i1hTg2gp1nJ2oaeU51Jsc0BzOlbzIJSbe16ahMO4LBK6TotC
8gSKiWMKXhjLiSTwCPBSZW3HCVDs1KrbrgrMbdxFSsbhK5REHqAbF8FPjP3v5+IL
pAhpp4j12LEdhWHLeDGFjkAYDZadDucFrn+KiTW/+2JVxZctN3QyPVh5NQSqkEEZ
fdyAmGhnJWCkaZnWqDPUdSrCuomwHyUhCOt0Fy9MQyudDwYSJ5Mf6AAbCOp3ALDk
45A/IxE/01+YFRnB1TbpCx6owjjswjOOb/euF6D28c9aAj+PAC+L5UPKQG5gPf+n
ssGGFxyxqhDwXkHDTcuRX5LMcoGwSmYVQpsriIJ4bjK3n5GWhg5sW68n2T03zaKb
4YvgBiZ4xVqi3zYYrgYwZiFYVUh7vjE/pXtlzDfa2QEZtl2NuMXNk4TITiOEAx8S
UZg6ARVyrMUbZNXBlAActgGC2Fni5MMruvqZtD8xQwOR6pqXvnnI07Eu0RgWV/hy
tWg79W+5pivfD+UqrI9T9T3r5tWKhqlJ3cp1wq2R9TgLtuXiOd7eNSVLKavsHfrH
KYyJNe0XeN7hZK2SpP9zZCUwfwkx91zUdFJJ5+7K3AmtAFCsiqIyVxq6wR/GCEeK
uv42GPjEGlzhFYLa4SD+xXW52iOyDoKN5FbK2uarq5TNDBsLzqj0v+x903IE0fNI
oVC3PbO7DRm408hxrWPfZLpQzq/UOBxvR7lgMBrXXcdtCSZ1wTEFC8b8I/Ow6WX4
jM/qCnjiidFYX6tU4pd4maQT3//2v9HIVP4uHt9xJvLSw8VUsSr5IhIcHO8FLsn8
x+6ubwmBfCKZtBUy2y5q3Y/6nMPWJ6iTQi6b8sq69J5pgjN5v5Fee5yXg2dIasmJ
skE9tLRfc70duZ1kmg7p22cG6b4Wf21tRAkqrI5QYNaKSqMKofkw8z77mr+Zbwtu
24JBLGtJTHvSSaACxDtPduBFUatmnDD+xFyapRSBpbNz2/K47L5HBaFZ8fDQK2RF
u5CDjHrWqx+lQwqdU4YphP8Ratiz1s4aPvs8z83aQcS8xhfRGugpedJrrnLTFvma
5TAS18lOgM/c/E352bZWiqMbjbXkDMZjENvpAzegtoHcvvSdE+ZDtvagCQTwI1c7
OfUvu16FA7H4AYmdGPoUEnnlGYe5MnGa08n3t5CItouvkLIsU4k+PyvpLH3hv37W
ut+KeZEXyCoL9MpverHqu3lZGa4zrJRChKHpu8y5BqEgs+NIKMNvYp8pGf3b41u4
rq5rdaV1FZpOJ5FkTJ6S/ROM6w4EyqpeqhntIxJaJchmZIGO3pVcmSXO5Qnr2EMN
sBSjQ7XZnP5FKa6Z2T67KBZEmQp4ycNsdJ3qKJhJ482ZXAgRIwA+GF/KBow2mSA5
lBgUGeD8OhzPKoZwF4NLDyXaLfx4pp6kT1CcOXDqxGvlQYD8dBbPlVreF1vNL+AZ
Xnvmba+Yrsrlw6LnbShSe+6AntjTY2y7ps8ktvUcU9BacjsUdYnNT47uSMAVdqqY
K77hYPaZCucnbY5Dt+b1pJyc5MLCyNel1TWwctUGSEZmdgoDLvh3xU0lRwdH7K2a
kITXwBNN3gL7DOsb7rk0kedKRwuCXuxfYrBoSi/AurYC5vCbUcHKTJFagHPAZCIm
4eaT9ueZsQHpTZ8qjD+LH4s4/aW+j9kli5QuKU63wrVDW4YgIdw62Hqh/V6nA/X9
yqGK+28ONx03Pjg5EiNBpkY4PnTLVuWOSgGZCLLU/pZkhYW7XYHSomdJu6yvxhtU
XsToGFQcdH271geinj44/+u3JjCp4c9rhWCpmcFvbWhlwmA/1QhLUr9I3Jnt6oSS
SyMaI/YN0uHnZh6EYG4QjrRKrqDny3cqOlToLqZVC+Ra/FQwOoK9C+cqi1a5xjeW
nFYAsdiztt6CYcForIqwPaqSRAwRsoxVkCA5gmDOIsyHfpftvv/tUq+cRDvIrnfI
5UaoxAu/sLjEwrzHxWl7WOAdUXYr/vSla/zkF8gppzXHQyx8hhC2FSgkgGF0Qn8X
wlUxpilDlw6tLUL4qvpQLlxwxvPvflQMQZTSnE+ALUxsygKU8dOU6SFOU6Op5AFw
Ew1lLaFCTQFyRL347no7Fx2L2IdTRRtOoaIl47bMdmrSJpQmikehSZqUPbuYjV4N
bmywfJPyY6Xv7ToOZF9iuF+OFdmivxIyeg7FM73Hlhs7heRSVZcdCk6pDh5MqiQ8
VnkK+PFFZcoa575xHvpfVTsdse3C29VlOXenix2ONTsF/UNFGTu68hfw6hHkOzaI
2RKOXI6a2bwWQ0pOkEOgkE7JaG6N/bQKwNyZ4ul+y4yJWDJiomK3zLv8dkViEE9a
Bl/+hA54hinekUV3jGFSageuLrmhuCoXqBogM5a4GOFsaVxlFereuFOakF3icdbd
Bku2WeDHmVzFN0qr7s7f7JocW2SZWMBoBhbpsXhQwwvAQX3eh1uQrsCDfnIfbyOn
nUknZgVyBB9vf8wStuWaWx2OKSJapVXU+NCd3bHiE4i5ksbHPxHYLzQ8rsNr+Rfw
lyueg+ZrZZUUUjXJcRGQcW4BrntvUqm3O/BWgotqNL41Vq/f9qnlBXHf0tqaTXtI
fZWKf8m3iIzIfsHdl2PlOp1ZVbznzCVm06gQDhebXMN7T1oBAUJHADberNkdLSn+
lFptze5ZKRaEgQrEWP0Fx08thH8cIr6RgP7sG5Ioml2lEUD/xCo6RoLrU9URVYTJ
krepXimylb38j6bwgR2QXbVZvJIbWiyYGhMvPY+BdZyuk7K87ogG8A5r3ZTAI/Nb
n7BDLPk24UG0VoVGLxxpihFku0QT4YHDJ6CuWLB1Fa4YHaJnVOc7PveDIWpJjeV5
S5CEhMllUu95jF3oosXgW1UycB/K12z5ThC4Z8JDUKbC3TCJJTPFgh4m54QMuABk
8SrO7g0SHGb1oawZ/W4RE62vVVSgrXyxSeZ1rOfSYfRJmN/S7TRNaW7hgIVSQWRv
fz7ilghI0h8zL7R66SGBsnNwIcylfkW+ddfCReeAXe6xrUTVkxW1VJc7FYvzWEQ9
rx4g1xLSNZNcT4psIxtqNUx3Xx9zjv1ALy9+/uHwFYSWitkrKgOlWRGlZbtygtyb
L5J0Ylv70Exhsk7hAfr1yEvuaeeV18GX666tGjyt/GyadmJldVFx+9TmaDuJbagf
RU6Lw6mhVGtFIcE8q5smdT1m8WQniXfA+2reICPR6E7nT0UWjfW5KRXaQnKP/bz9
MoRnXGYqSLRq+0jcu7VdjMSibjXs+I+eo4xelrSAtq2CH1BQ44g9Af3p+pa8t2j4
Q1gKFkylmgqgx0+ehW1jKilJb9JO83cRf57YnAUMYDog96Eu9rT1DwwT2D2wUf+z
RSkH8cifM0g7CoYBkWfCl4miupHqeZvPgwQy5DKidBb+M9+7qZ0Ch7VMY9tlMVc+
yBO1SkS0anhW/+YLN8G+xlOSRz5yIy4eG4qu83r9Pxhzn/pw8XSwSFLsNDOXYqAF
M8ydmJ6exlLyBHlM+FSsoxj9b/Q8ey7NBgwECO0N1vUtsx0RHk3UJ9k89T5QajEe
6Ftw4XMn9ynBg7Ruwlj+WZWPNi9obkrUH3YObE8i4ladcGwZxFwjslNooCUZO4Yw
shinpViSc73YrKSLYSe3QJ0P2cD/5x61jTAW5Fo76ul4eqmQJ6utbVVuHavuc9rj
XP6lzSBg6Qe0GFOmh3t44yUVDRf6/P1JuUr3LR7iHChunCFAfe9WEH51BxE9yWGe
mOBMXFhcZMBKQESSxMQEr3w1WO6KRIA3larytTaLCpr2/qzHU9P7oPC3rlrPOAT7
8CvSir56vm14FOyypWbrvd49me08pVQ/chU6vQ/I3zrWFeiGWyEpznpU7W8dTFDN
JJq7FxBLZCiD1jr/pk6CKyBKzHrqYYwsmd/Vi7KyssvwUG6y5dHd+0NqqgOMx6gR
ZkQqB4aB3PcbFQczzln96XyeTPOyZpYEltgbaqHnSLzzS8G39F1q/+Grun2EZ+GC
RO+pLlOQq+Ku+gDrteFhpjmv7o9QuzFTPkTP2fuEOveucaC/8asp+nPilSvpiI5X
UZuM7BWEz60IpAwOJuYTX5pCon0Hj63eX8RKhZiF5UTOCVr12WNGb0K7PDz3aJFf
R57UbnX3E9tOVVQEn20I/5ob5UDTXtuuB5iFhnXbyk48lwi2FDW3xOukM1xstAs6
5EWHEM7IS1rinHRYHPp4wUVHFRRkGKcYqGz35IGjsPVIf5Gjvn1aQU1LPBbGViDU
CjMWlTEGKx768aH9Seeh/W1OYO9keRuJk/LcE9lkMO9d5+E3W7bA4zu6z7mILIwN
eu+8FZjOKqL+lgX/N5jgq8Z32zCDHxHL5ygBH5OzA1LvZLiQ7foprGK2cZhycA2i
2AtmAiDDn7/LsOtMRneLOuwxTII0mJr9pXsAOVw3VYd1+Fih3tQeOweDi+mJXSDL
u1FX58AsdPcRjkPgdhtEZs1rYTKPw5KSilfq/XGSm95oukjO++PJsvRrjr/hmwwB
tc2QI5MZy3/qs1U9JU92PzYV7M5SvlZxvlFj11DwQGe2POPmGa8asiFRqDcnzbOq
UUP04ICmnrg+UJEtEnnU/NbDThLF0Qt35ii1gYdGhd7UEfReN6UbWtNsgyHnijO6
u54CoF/FwLo0QBpmHRu6l+w+uUcY1nSzv0JhnhIZJnjYWELICDda4L97m+pmtmpf
7y6agt9oRRR3R3jinK6ctIehwDLHeS5l/cPYrCnIxi8bc3LPoiIAWOW/r71HV93k
3lDhpi0Ic8ViVS7nqO21NOdHCTTfgQpnTLZYNAz0RPEl3YkT5l8rNpDYO32GBzBu
Z1Hs9qxQT/Q5+VCvi1/NiEG5b4JJwGTivLfC6OQR+zFllrBrcwHrOITCoINDyPL7
5M4K4Fhf6ts813z7Zj7KcDAFA9r8F59e9YT3wcZzr5+Bx1IIKh6JUmBoR/h6qsIy
3KEIKdXQqkuvJFgCIA9PQeenXwTXjamCXA4oWLPoJO8P3/uwGVKO1slOiFfgtPs5
VFdjmciHFiPGZrTduJQLUmrl/dPYLvSJWwsJLlXWkJMSkBGBh02LodCVu/NpJe9Z
is3j3RyONu86uQnnu1DMUv2g5NLeRV0IZ2UwIcHQFrXVGRtCBRFxKK4jUgnIls41
uxM5BFP4350U71X4JSoDQbBvFRIZtp3TKiBGgzPKw/sRsUIVkshRySKq86kBjUAB
l98UnTj73U+EM+uPuQHMO3JnsOSNFdxE+tDALIAd/EUiAdI78WcCj+CUNCRQ32Tv
b+H9aZNEPxmGF/SuEMimzMZe7SbH1vF2SrcerIe3K0I9QafaOudvdkxNnUjCMR6i
GuqMHPsp/eSOs9qE+Q9dJomE4qmfsqr6Q5ZFvKtLJIWNHMMBi6/0h0xpYFQRXxmL
IEV2A/ckgxdQGLRMSch3U5gkZAOD8NBhibeNztfV6M8DwER4c+4f56UYVSPLNikZ
WPsLG7qnFH7YA2t6R2TAhAKphM/WRXnNotcxnPU8KUzGX5Qetf3rr1ykEN3VGXs+
K2Bj9p6XWk6qwn6Mv9G14CYNrUQ5TMzn2Hg/pN9zz1sA3rRybHnxNNEQ+khPcQA6
HOceUZpFKGHT1nZbp8z6NblvKw7K4cbCyEREiSVG2uqeuezP1S02Am1j2HntyRFQ
Ri7Qp2WV+oEfxTnGrkmwPyoxIQo9Ggm5wUoopznusTFh+UELDXpIi6y9P15k7/Mo
Fpwb+3nJgbd5P0HeCkWDZaijHOKFfiyexjR1cqiCoi8Ospn+U/UClDXlwt2W4h5n
Krtql29NV0i0pXu5eM6cZK4bUDEvzzsyGQxSCxH1n8X1qQwwOoLGoDLr+vGjB0w7
pt7/FZ9r4PkLGxfjbqckamttXol4Ck4rpkHIUahre63/Pmomtpic/YR4TiJTAEZk
OxLALU0WAx6gk5hETnU3Aq5nGVnXje+P0DYhVYXiPoyh8IpZzHXX1l82Z6odC3Rh
I8tDd1EqOdtM4mEGDS42bweajrifTRg/uhziELAu6/djW/Q5bZA3BQCdvqe7coht
0OQ5cpiqgzRSX1xKWgXokdrGTbGP28r/YloBq/HCTUyz/OAwT80S3an0WnJoC9HS
LcqCpFhZjiqVrVYrUgpzLv5uuaJzyWGP7ViK30dMoEUplynNXqFflxy6P3NLSC/k
K3hjj+tDaPLYYKRSMjN5sB0VszPrD0IT3juMJLzZ23LG5IuLXF24i1qEX/JGJsEg
lN7R7AjVkceKXRIyMSWsyuGXGuu/y+zPSR2Ha+NFN6Bwa5AGpLEEMy1cz2T2iZFK
Gwj+eIU2xVA82zMPBCZBvUfS7TBjBaL3fYfP/w0NlsEVsYkT9mRm4Sj27rx7kHPu
1+Jlp0xn4GeId/byIzGzm2Ti/9oACs/l39cGP9Sgs0olCY2E+12fKwSDrrm+IWEU
xjeAHlYyIfC+Jveaj0pjd/GkOpHpUXDrUMBaiiLtn5nDf8fruhG7RCAu0HRSVA0I
9WGEMX51y3WrFXsFRpGy2QdXOZCRn1SP7NzVNhVV8vMH8xbfQ58XTsh285dKxFbg
2HROtIvPX3tbpTIJg7lFbWYjrRYXv2EqSmNp6SSzUsYM5BddAeNmSg9Qm5/6gq5n
ls+80ecqUG2VpFL0BTYP4NHrWhNxBDGyfrOnTw0mmUrOVdpRzkzMY/DBluia6UQP
lOPzyuGxx9VPEeRUcOEaydRMRj6vHJkQptC0M8PNxqWSgRqN3YyuEPPrpXZHS2Ir
AcJMVPc9MNQAkRk+qzX/feSBrQjkNg2QNf0csWj1gFXRVlQ6Zs4wc+h1dXPJWUxi
IRHu3/Mm9N7YXwiYt//nqns7pqYcBY2Waj8+tTkW4C2INm5BGSYg4dJO9Zn+XKlZ
rtkZae/RSzEJMpgtH0qqTozc1SN8uQgwrygpD95cf86bWZ+AcPeOFkg2R8O06oHN
4NKASm8hokUp59nlbSX2cP3y/+POQDWV9JfsYjnWPS2MG2EGVZrQsTuFHAs/7gtX
6mulcr0WquwRv/WyFxF5dqzqjR8yKJ8hG1ohVqSdgW/1midlcAwOHWPaCQC3vRvd
dfF+E4EGkPZp4ozG5HyHcMp0HfMQHbLFqLwNCVBgcV+ceXKujXGR5XQsbDxL7coO
Pbn5t/ekynYsdQ9zho6tucM/bE5b+Sakn5kX8n+nz7a59eoLCdSReMbrKxgnIqz0
wpdMqRSuoHsXyDZtCjcXXW+2vuMl5+r3h7797qy3Fhjy+GcsNNhh1ezim98I/+VS
j4mFjrdWM7XGCG27Cro3chTdWvNHtc3OPdMXN3q9t1HPR32R8t49VgUuIFHQzrND
7PzM0nxMvX3B46VGEmXXjA3ticvGx2IjcXb7AW+WhbwU+Ct60N0tBOEHo3f2r+Jd
YbO4CGm/+bnnDHt0f1YmleNy3xEjfPgLXnoR9uA/mVDYTQ5ZPSK5/LA+JpR1E4hX
drG8tyBmhAR5QaPc5XYcFBbGbENM3bjjy+ZuFOOfEGf67HxOogn8Mf+P9VJmZl5F
wFUx/UDAeNI2ETeFCKTdzHFBU+jHTyZB8t39hsrXBlSbrr/EGySUpKl6mAiewQAZ
i/kpL5YrKJC6YhZEqpSokLKU/M95J0MSLeby81pAekVxwHx44uHeP3kq5iIi4umh
HT6p9RNuujacO1TGW5wn7IHCdPaXBEdb3ghmpBXWNhh6i3XV3r5miLQGUr5a53i7
h2Ib8Ygq2cd6xIWe82MnXdN2gadFynydHtffv0UIO8pu59m4GEj8IEcNYu0035v4
Tj/cxKeFwLzrbxssiLYE/RkOhtYPw0oTnXavvrJfMu30kemPRuDAU052necQA96i
dig4+c0nbcpcYhc3d4dpYy+oNYiR/ugC0dlV0PYkun6g+ArrpVdx+yZ7H6y9vcXI
+DSQy9cC5Sn0NyfEi/ZRNpVl/cZWE6trXvzbu8I80cEweQE+qREK1uw88jpgyR2W
wy91y5/QIxijOwz+olfiaat61H5A8KPqbMTrsHtaueHkPNW1YdaKvK8gK5lhEUEn
gCc4ws8UQe5EXbUKgEt/Jb2bZPEFq4NMHsjestW9w7eHfbLOvfJCDR2Z19CPMDmw
vQCFPhThf0iWJgN+Cjh0nrnnclQYDUPs+Mn/aSr8UjUAEGl902kyO/rwtQPEX0c1
a62TDLsmU+WQOX43xBvLF0iZIewOVU9AhmcK3cg0ScNRmrllUVp9VLjWaV/0Bnbg
+Y0dUTDONSdMks06bnYkFDcoplGW/LspsgE2PmRLQTe9zcAsfq3tHHOcIjmIR6Ci
s5Hrms/yfeVfpskADORhCQmVzh2ptlPZD/05qi+v0NmjiYlY5rFhpNO4NkVJivVU
LRbGmqMKi+1K7kbeI+fDvhtBsj2vvXN/40VhsPMSDXk7EoSP9W2RcJt9n+hTPWsM
Nd6vg/tNSdCBtZbpFbE6gMf4gmRYLn6OfHOttopOhmKdNckuXt5y5h5fzIX8WIvp
Xspf+J/bKEZbcEDWWlLPUuv3vRuCRfiEJtKz723cabqjBvNp5F2ZHOFOLKDr7thT
UBlREbzF/tveNqTfnPKTmS7RTlqUuZ5PH+7tbFSkNMbmKTZpRIHfPW1K1qkl+XRv
QbC91bRarJ2xO/NOhq1aOb7w2Kq+o386B4QgxTQbJi7fixMmDjc9UiW6Dz145caH
fC6sZf9/5UZh7MimzWuq+xIM0CMTizdfmSWPzBawfrCvZ+gUcSbpbLP9V20TqYiM
E3Dywkh2gr3RhG6GknRJ3tn1pAsuPclOC3m65W+5+cCelmtDOhRd96fDk6qBsyRS
tqyf2OobtI8NCbujZWYqpytsl3BINYsP2gBVbBUwlctBVzdX4P9idatGgHzcVi5y
rj+WSCTfQDIaxhadVj7whdJFFCGv273Oe9sBNaH7gxFjLkj3uqUs9eDASrgWcs7F
Ifj0Yy6+GnIMAhy7ABhEIe6saiKfHa10MvwHIIbknbUPylCIBQxG4zlaHgV4hnfy
bIrTE2eBH70dQFDlxDvZqvSTMXAumin9icMkAEdOBSC1uYc1cca2/og6eA6fTO6W
QtZeJ6S7TRAitlq3LX0do1qlAt2YqnrX7Sy1aL+j14BveGKpIkgqrtrKNof1TrgI
1xSH6+hOicRDoQUfEqU/Wxruimd1EN5hxMbgGjJ3lbYPvXhF8mWkVD2Y0R82aJ+u
gGGGYbhkCeIUEPfp7pTuz50dBgudowdCCnXXH9z3wp8nLcIGyjl5NSazG9Z+TE6d
UERiCjCcfVaK8v7SV93k+nGuABueA0/Xsk+kYITTV5PHTBpQc4vt1pulwSz7Jz0C
g2UrCWVPBOfONmjBAnZyW0MhX91EMeZcP3yzzhvaZ6xJ0eE8kB05xucMR+/yES+C
Ce22efp2iKMytmM5xN3u6uAlHt/BYTngBsZpcz8YqN7Ecouk7GynWbYpeOA+DEC2
a1CSHHqL1mhbi4fInRVoICyo70E0moJusVKFB7rAd7uofBXc73Zr0RaKZperq13t
QGFMCnGK6VkkPnjsTrfAkMI2XnojlnaJcPUjAdjnhEL2maSEAMrWs8ffV0LfG+ny
irP2XsMIV5L3s30sPdZvQVFqs9lxC+GeUA6QsD8pPxHEDhHrtoJpF2c5iIPGXtMT
P0KRdBTcbyCDd7wZwNCbI6OgD/NByk2eTUcitzk5/JU0Y3HeMOjjoxoLSbnR8wvx
lR5hrokOMVnuX0Dy+kevNh0PAHLdMN9iuRbX2/6OlYCXXhSTGf2YukEgj5RHYzEg
WA93pvViKqq7CJZZphyLqGQhwvBIZtNLmek1jXowqRUsNfbDEhLzm66BhOxRTJdq
2WJAeiyb9C+6BQ4z7BZWTKRH3bkgErkTXkXd3Do+MykmKeSC54HrdB9Gxi5czwhs
K1F/QcXfQWPG0fMsaCQNDckDMlBbalU5ZucmAbCbTwI0S4o5uESDhOt8uBg+6XFG
aLvtnuX+Rorsa3cX8CpwaZXc+upR+ZZsUbnlTL0SUtGfdiZ4tAKiaAVx7X/CsemW
2cWECbGBq8MmGMt4CT+UPMqv+l3qfftSSIavu1nILunh63XILyhh7s5VRccTpsCz
EPM8jphI5kA3BqdiD1BzX1f2Af5H0enuhpzqW3pBWuQs57ypxrKAgWfdf7x2cG34
xa/B/BGQplOOXHMhJUOTy0dxOf0+STIuTyY7SJ+aus2hGuZkr9ZfzFIpyQoMykD5
oaSsnrQe+ongG+JOwUoRYETfefXf2vyGGSKXIVnBScMVF8yGpV9S2V79japZ5HDZ
jA0E6y6byoJtZgKe/Vt7qLxRE22vCOUHIidGOAa/k/X3rl2I3IhbNZIy5HYDnrxP
L3hC+/b+UVAe64O5dITZA+kFZZNdoxv5eS0PQ7d2EcoXymXu55XEwldtw7koV9cD
XcQoe657DKAifLErUDHaWwFpgvQPp0JbsewiqtzeSTne6kN63cPI1tMfClaayCak
NMCmJi0XXvb7eAgwRbnyyM29NPQv2SZTYqd//34NINWII0S9IEdTzVZTWL1kdvmV
XSQ6bmaRuJ16i3Hy4IYSYmqy8+IaaWNvzF8EY2BVnBOCDGWEMdbrCYvWUeqqKtE6
XS8ieWFf/M2jYpnd1OwfXGdTYs5mJTRka2GlyHS9uLthNah/YrPH9aJUc4bD/urZ
9CsRenj4tZcu99pZ7CX0TjPzwHvYPUPpdl8Tv6Uxyq6dgA3Qeoc0CnA4cT0dc/7T
18JOy8vejn5uiYawTavUq23UfGfvY/Y8z7puXV5qrmx4SjMh2L51TYkKwTWFkSUz
QCugmWjeqfM54kqPstjucpnmcmzeIy5XhkqRywz4c1qpMDxzLmodjqsmBf2i1ixk
3WQqgjna6HZM1acoDulWxMqbKw/qj6IbRV7bFV/qyc/JdCL7K9ggbocRQpBryeVz
TI9lPawRlsE4w11ozyC1tQcSIiYXkIXPX9VSoRZ2R1DnzjmzwIrh9GT+zuWlO2me
V5XEE52AUJyrbBIAP6uRuESoRAYKuQx8vkQ2jy6oYi56PNAtEeRM73+NKuygF9+t
XDjhsMSa72wyS2JZYndDppGAqGK80ZWeBr3vDmsMQw5/8UGbY6r+Ig2h1liSVauX
U8NJEGu27vePpT0VAGZy41tB+MsSCUEAYJ6afRtOk/78h6y011yHi7yNZeJ63hGo
Scs+sGSZlvvBYf13GXG+GriHchNybEHhOZ3Av8uZ7bqbeYLZuSHsU/DFNw2RgPN6
8ouO9jbhKJLntMuK4AFA7sANLV3FHNsuTALtt0tSD/u2hZwKZKuQtz5jl/9qoO0H
C2Hn/HDNHcrkJImstr7373ZnNUtzHHnnH3KC2jiW19ryexwvhyp6oTZfTw4P6tYC
k0Vtm9Ht1TQ6LUOlmV7HJsnvTwxGuuUAFXKlzgNdKmfUvmNzsqbx7f9bLcv/g4zs
puPcFMDBGBmfZDUdEbGLMxAeBJLAWs6FtOJDu6ZEd5bFbV2V+yDgYqFrAFk0zHMT
U6VTJB+2d5d93h/XdJ4GGXDSfD7dB6gPbbqgkIjyFe8vYO2dxwI+gZNm1wSCVgVs
EFiIVSqMzrG1xorIghrmWUJtVjvChH4hOHhek1B1LIUFrzCQ3iVKq3Qu2MWzfgsG
7ayIUkQ1rwnCMcqAjpW1WqSCjoMO10cLB9/jGr9UzgqusFsHmNzCT8TAb3qYWhG4
sXGQLgFVJLdswFwMhBwjgR6rKT9VeDIi2N7jnYGdpxP9P9+Zlkamxm1GoiB9vqcg
t8WN6OgD3UQsfdPA+nSOGvgdHZgYE6/bkVmevPlLM0z9s6TtXmLfk3YgD+kmk2Wz
leBMF/oxKJX0vjL+D57MisOhSo0ti5SuMFyVH2bq05XtCOiQeV+6S5dU5iM5Q9QA
lltySK05JEQzKs1tR2SBLKfYLDGmv+ZKuiQwbKiLxACbQYokP0Q7+cunIf5I3v/x
jmlq0GJNMs60XHZPvvvXho2VG/pYGodyeIrZld9F1b3IPi66+/Gpva6a2LSIHPwa
mZ5fPXw+J6vsF3wgY0qPjrUNOCzEAtJEtDH72RFKueE8cRF0FmHkpV2+4hIU+iz0
25+K71zgEKc/PJV9FQaFbg6XMXJcAm1yf5zhyNjQMbkUWjXqQ8Y3KHeSxG+sYqb2
07jzKHQ/hAXJpMAhRMPogmVf5QAxu5GMf9zQoForUaHo2Ceevj2ym0jYPNvjSiph
Lmy1XF0Bb5uqiy8aepufLfAuXRTDM/QrTViTYPWKRDG/qowd5pclOn9fhe/d1QbQ
w0RkOlbZfgfvLUp5I1T4rQC5KcK0pQePR326ho0/7ogFHtGTaAOtTTYIHYuUBxdI
Duyhz1drDrp7nuRaLLxclqwvEkyAWjssyH7+wmcI42s39+BZCRw4tvF+tUjJ50J5
QiJrH+wXtfxa9ehLnbbtf5iFYIkpDQiQ8LCpd0Ft4+MLWBiKqHGiL+Fi6DCq6gND
Lqfkm/II/9MPq0FyvFl5I5izy+v4xuP47k5jrrpJQuMm2LGpIxujV4VLCwyVLxkJ
5RNiZ2p5uG2A8tuDwSpbB3VG68mWHpfOwj21xhGg9SY/QFLEKdZW+kHlIhSg/XkW
tOFxHh1wQAg61drF9o8PuAwmfg+hVQBk1j20cL5LwfjhzevrFIGyZXtyD7IxQamw
qyGmczpXN2epv8KO1KEZRkhaDFUwMLNjkFF5y1HvY5+XCgIEm7aqGeSTuvNV8HPo
MAw0r3NU5LB6Q2jq61jLffxXzG6zMafakNIjlpu0kB2GM/8HPi0LgECnSd1XDKGJ
7/tU9J/wQQLYoJoQJMehN30SWuQ27bFKHGGvhQm0T80D7aksrU07VD3qz9bvjeG9
vfF255S79Ed6epG6PYhMFtjKQQN5kLduDs4s5nNeIZTCIUgxXOEjz591OrgulHX6
VKo9JFz1Qivw5ET6waAw3Y0dUL9DCAwKyLUdD7pTLVtMj8Ht2XCbkZZXKbKwq8Zm
ZREw1P1x5QFSEFRpe2daNa3UhHwvnMshT3QePMM6xpNkOLpAllbetBRlPvbBmSTQ
g8cEHf9gNieTHVUy3oGZIiyUTAq+LT+MeOQSENxejGO1SUOuRNVW7FrT+A9tin1s
4WhZuiKhkWx5+5zmkOoHGcTdZBfTLkjTumViOT0frizYStZhtNjT7QcGt++CUjOC
wyKlhpbGaYdf7HVCBLJoijG6lMNhcikj69TkxtqBn8l5fXfJpSLYV3f69bwZVJbW
dEE9LLEyVeNrq2Mdx1WqQQYnSS5DPFPCxbCllQRssEOG4qRzAWF79axGPPud4LFQ
dgIEV40ex4jaEAkvbKZXgyFbcVpNHrDKXYJno16Vee17FuczTq7AYuDTQciODJYG
ApSJ/m80KDvLtyTnAyvewOeePR2C1O2j+d9yVgz27mB6umguxiHMteHkEDTcV42Z
6IK3Hdyr/Uv+SzMUgHzkTQ75neECvPTeDfJuxc49Kud0F4Ua7XxdqFpVkfe9SFtw
Bc3Z6XAOcZHwDflO8cjh8lwLLjUNgbUJim7eQo3eRFLDmd2KbJgAGXnPF5PsAtdZ
7Aegx1rPSC9AynfuWzlHpKGosQcMFqAK0vWPNVRpDFWlKrfWDTufBByKhYFKei98
jM9QWnAQp6YgZLFCp1APHEl2upCLQrSleemcNwyUICoE+JzSsXTStU/WbeMbWByW
JyxwxuJm/9wB6LX8Bs6quLci2gRHR2MBu665ywBk8lH0iatrbSxmW6t7y37KIy6l
JbKKSUBRoCloHtrAsKSGmhokF22s8w7Qf0XhJq3dXtauREG21TvSx/+hLcW22NyP
PAXaxGFhZxQ8vzOyfojAigqHlAp8swP8t2gvsjVqpn6VUjzfE6KSPHa4z2imgdku
oWNpe6Wl7cD70o7F5y76gf+ef9AMcr1+50wkQ8ooZbI1edyjuIn74eZtIXtIZFiv
k99ZEArKuyw/PRa2jlvg5Dc1vpowkvleGV324pt9RuWsrmaU6RiU4gymkz9wq0l5
X9oNhGMNNiY52/bI1JdseF/nBf69A6LEtdPbqcVQBwUAgUBsytNakGCMJ/a7dNpf
eUxtdKmTlZx5BYZs6jnEZbm1o5jC7iTa8xkrpmCLV2ioghV3n962WXZYFbjq0oFS
hc8PvLtnC9NlfhVDrjSVyLlHP8oiUG57a7kXW0lQjrCDqbVu55TSO5cIWyQ8THg0
OxPNyUpTlbPNwUb7zV2rUkJQfOiHSJ/Wdeh+qi+RjUEDq17oiSzxBdB85eEixRFb
w7bPPXtOraiUbFw4pFzno27diBzI388vFix2rodZTUsRUL2Ul4AHoKSh8iFqEv8R
XYtcOVm0GHqqAJ0UpzCHv+hsiVTUkt6V0HZZuCBjM9kx4H7oGZPd8hewBzxmCt84
tMPImlnO8ERtSpIF9WyEQgHH0fcoEUlAYadgCVx5rCYGGVUfGB2eeUqs5DjiIr2M
z4t++JhddcJSeO3oAb377Mbo1riVK1W/pDiQ5aB1L+5M/nc8LlwuH135l5sPEGZu
8ub1hZ0YqSvo7TzffPlPDva0xYlKH2+De8iHMXRjPOZOIksEggXtcVqnBzqMsq9u
3nHZTc13ipMkbjL9YZIrfoJMtB6WZ6xzosqZLRh3ZPp87v3P72ngiyvmXlIhuosB
9j1JO4uNbS66HU025EvFaH6LrG5z3aNZTUFThbQbFdwg0yz3y9k+gv2P55MM0Lpq
tYjqIfKVIziZHP1qihUuJAe8gn8Cwjp+2D7oIC3A0/ryltR0f+Szo4ZjbqcRkhOg
Z2Wv9PKakoWYqEAoaEcBsWZ2EMo1FEy3w04dkeeLXcFFaPzRbzSDAyfxChh5hHAX
rMCD9CuUKnXQelZHfl6Jle+2gHqaWcLMnD9sqtVXmwMUc3dQHQLw1rC6qx2jw2mJ
KxW+0qJJcGraL7kuoe6QjvkAN48oPrJcC9YvJUcKcxc/ngyIt1BgU49ZBQfaDC8y
3Da09Q4k5dovTX1Mj+41y21jZFhwYLueeqQOpuiJQjQxi1Uw8hHqOMEYvIM+Jozo
2wORbz9e9Rb5nCe2i7foHe042rE+vgavaoh0ZzO9cSX4hyMScWbKKm0OkUT8FNRX
6+VWPB7s7jfzM6kACK7shPSAiVb9v1yDcOUMnHttaXu1zjvEaQ2GoNGkP+5k9Vcp
OLGhr7UP94l+M96cLkcyiZhTOOQi1rQyMdSxKo4UsFuC5gOXkbVPfCvmSifNkyzA
l2FZLB70iBgyG1oeDWlRmskMK4TumY0rGNloYP1Off4P9QULLput4uDrdDNsZAiE
yxHr3XDAGyEFIkXv78xGIKOQGeUNbzwLvq64qF7DBMEpvXwUnsqx9NNeFaXoig8S
N8JS7XoNCCkRbMhGV8Z6xZlLPhF9uZyrhFFKTZv92qmIJJ9lxx3WsuiMFz3KnJLk
ZVYJlFqhuc50OI+UQZYoMAI0deeISXpoycGJSO0sjuBrjCBVF/bD+2XJ0wbK55Yz
Mz0pJn/zLhvdk+thbYrQ6n7nM2C7xmbCfT1fP/5ET703w5dv0Li3JVjpHfZO9lLw
Zq09PHgdrIA3nnXadwsZGO6LyoCU5BJgrFWrjYHe0yaHKBpSIQ0s9spjNDdhxmOw
GTHDGLhk5K+fCSLYUNo9GiNxKXCnpLPXyapYpNpI/ZSMG9FshhPZPOZBzbC+Rnfk
yeplKlDd6uAzHKh8mI3tMoXjjssmMiBoF+OSD/BKU4OZ7Nwz8fBwVUmGd7CkPNbD
RuLfBZFpfi7qwwmBffyQbgQ4r9WxgC3EtNBr+//gE0H8JXlVboWAbqJJwJ3cL73v
QQjFP1eyfpzfA3XLVfUz9Gx83BLo1ShFgRLTydGGB1zlfMdAF1E+wHB0+in12ff6
YdGqFOLbb2vCzp/JSemYeqhxGmy9Q00NeTy6aycLAWowB08CRmbTiQg+Ch+lYEHM
xFpom3EXQHmyj5Cwcz8dXfFRaJav4o73+Qr2rh80bvgpcOo6UPm+XCo631CnSLDx
mQEia/ywqg34FzEfvznZF3yYnLz2o3u8XQs9RpBdcW8vAkPmYptkflqOAKow0LpF
4WxBnZfJTVxj/F4TtkMrGSixgfitl95XHjclCw1xQ8TJS7iFU4pmdq5qzHKTWhbO
Z330hiPt/+ly23IdFEENkmi+P4VEEkIh7CdxA8SnM7IcK6sdJfi7ADGvq/aZPE+6
5IUiKpV8p+VSxLWoy7SFoWgXlJZAu8r296P+JR1hi5MHmsmMcszAbJU8bB8VsKK7
v5R3uV1Zn/R3vGIJUapKlfYUvEQWjsMO+rfj9/dlofGIDYrOPMCUszD/3Jidj29Z
rUymlpOsjoAnKpEJ1XqdaDLCuR0Gg2YSRzZxFXsKxTvezu1uBsQGAWEDPgylNGH7
h0xM4s0sClJxcmWPU/qLkJUVA2ry3xW9tkUAfzw7uTwUf0j3SSJlTfTgk+Rooshs
iA4iODH7wg6njbdooMSlzIBqaMLXav5hyLy8v8ivAe3yKK5t0L3oAVKUU8O8G/KL
Hm1AmqYWEtGZtAkUxjJg0WTRYhCznmJ6T9yVhmhM63WTTg2y+smEXBY9V3cuCAGD
d2JWrp5UB/Di8rtZ8yzKc2eRF5Kq5E/zWGc6uRlC1q4ndQurkEaRNyubogZJWqNu
vSEFgbv2tySgvEORJz59/Yxgaktq0xum3K6ZuEefixKnp8fRAy/qEvZsqtpjkYcI
nbvkh/qBT/pL1fJ1psCPAD9qwH6mVdtMjywAfTI6kGKn9xzqXQKE5FkH4ECpUGqR
tc8k7pW2czGDN/NqjJ41Us2t8c1EdI77iKP6+h2+phtM5HerBKoud6AoMLFlK1AU
e3emizvbO9rTNPcFyCFnIaQdx5tobS7z71VOCd90zeb41fCh442wpjIuzS8BFZXo
3PJfLQhX8yNdNt08UuL6SCkwmaIZhK1X9rlJ57o+qJ3L6JhliDNGetDE5EufNlhx
411ELdr2Y49WQ2Gh0kiAcUH0v1HIm7eExkzcf4B6dv9+GJ/wkctC7JaD7ooWMB/A
o1ecEZFoT8cHeLNbhwIy28iUWVQ8hrlENL2+wWZV8/C52ncsDGXqC4W7QuWLPKe7
5kf7nVR6EMjk2COJ299DiyfZ5jU+E4jB7VdtKc8uESVspQnM59KtGnrKZRPQ205d
PXuPi26OOwIckSmUwAz8l9tn+u2t+X+UaC1Rdkcc6fP0mDueFX7irRIFMBliltRb
MyA7Gxu98nAZKTPHBphKTHNNQb2LgS4vV0hjO4CPISxRupDDfBJpdeYDKnMmSxgx
CCp4Qs/FudxkAlHgPtB3S7OkNlyYvbfB+Q0vBK5/Il164kznxW7Pkxjk4/FDSA7W
11gTnatsxMl9qaJVr/IiZW5pbHXG6R6+6Ebq0VYKha9SGqqY8Y0wRfAag7kFSaew
JwZgo9XLyQYysnZPtowGP24pBdml20QxRM1UcfWxhSU3gzWptAS1YWKQTo5M4r4x
PpX4tVPzzquF9TI/6E56S+bO1dxNRImpU1hkIjT5VC7T1GL14aLLWp/AqF8balap
dUTKxX6F0BgSmo4xe3/nshbrNa2JwWkw2xuXVBpVi7i92bX8akS2nZ3xcMQzRwCL
bLzHcozxpxnEYHXSZQI93DQSeTQBdozj3B+EAiKUPwilwjgQfPTaMM1HxLCjWphK
Hnb+1IIjfWgNnzRByAY1z1vEOYh8dSjvbErSjUFiV/ap9pjZDfuInimob6IFukUd
gjELj8C1F2Eu53E0LHkJjpYYsIce1UL3b351DpuLrCDx65YnyYmL60DaRVYnX13H
b9rysYq1AST9ifGH0DlS9quXkrWS4jKJHrezylSXp3WCmYQ2UjMyopkDkkB6rtT4
YrtC5Zsy5jGGNfSkZQe7CM00cAIMd6NW+CeqL57p4/pSAlbY7jSefNZ0n1hgw+I5
LRn6mrmgWbcnxEvDKxSzBJcvGqpjHq2fjhllDkYlc9YPKOVgJanLIfIOJXpNIkTP
tJuN8gO9Sk8GBJ3dlKOp+h2jfmIHTm2t5XdVeQzEr8eoAT6l8RQ0sqJ53hgmfc3T
hLqhZOSAD4VrkU0XB8xfLxYpmq19HAI+qySyqJsz0S9GmP6p9/UzqzGAh/7nyN+U
URh0wpU6X5pttw/FIAbIOr62K6rr8AH3brFtqQCpH4KO8elPQu7wN66CvqVn5JQ5
w7iQIo1eM54uE62qMoFqklCCkTY6w95tzkgTbVc5DE5ECtNA0DmYl68K1LnwC9Wi
cDBW6f9gYG4tfS7GlqsuE3HZOlp8TxqAwDeUSnbL4zxuYana7ytizVmCObvlk8Wk
5H61UyYMPBRusFx02QBJptMWlc0C1mNt8nfkrOAulFKGXl9T5lmISfyZ4k6phmyE
G1235a42XIS5j77EbQ57VwSIgpfk7RxsC7WpzvzPtdCxgbrauo4Ohi9UC1PKsp5i
ZZGZC6AE0tdjmQ6JF4mQT0HTzDzW1qmCHYZ3o2/xy2wrzbXL2awhqCm85ZFvUdhm
hQkZWAeiYUzfbaOBfv3fx8SN3OGpyl1JjcockLOrVXv8cV8HkxF/4vo5U6der7iN
sO7dm9tjirWexMOxDxxeiusaoJNeqouSumnbzvhpescSpPIZjZSi6S2+Mx+zmVX8
joLSXUEUL6T9kYqu6V1Ez4464oG2Mpbe7WSPF75trJg+lV/9oqnyT5USfD+vpkmN
Cs7WsPlK2AUv42qR3By6N4FxC03Z9qW5OY9QNAdW/zYKaghynq+4zTqgXqIHvb4v
R1ZBC78Q2p9KaqYla6jU1RK+ku4FuyHl+45E69+pM9DH23N3kvdcOwhyaDsf9jqY
Wehs4YCVXKlBeGf+DUHYyracLLRnuKGqBN29cNYkbzmbFBwx76oFjRBx1ppPEsJ4
LTBbQBcVkeyO8ol4MPs+MdxDyBt5pLVqL08bg5mIXQ+0xhX7kRMIueyKJYmhoAUR
eIUPyl267/5xB+w/EHSlIGuaRCjTKVNqhy+ZuWsKb3/4RC8iNqPyJATz4F5qOaHj
lrZKprI7DPryGT4PCC48lz+Bf0JClTF3B7SEJb05h7H03OLJckXYDK75YXcF+Qln
cVx9WO3EWlpXsju+WvFB1vjeH5+yrkBjxfUXjVWttR6CqQy42JucMxBfgxnF3aZE
3WBkB2COmFvE45rdNnfZHYGfn8DeolyqnbZHLTjkASKuiTaiZ9FMHMlA3NUrHlYM
UYK/mKos/+4wQQTiA9EgQWkfxC29IPW8RW5X6DgF1a8iSJumRL5uvTh4REQpbttT
1vIY2tTHBPG/E0Sp6Uqw6O5+iYeHGjXNjMHEOkLz2juVLWk4MEUjnk3rXwtwdHeC
vHij6UgOm5IwBcHXch6D6PIxvnQg7Jp8ucnL9KvvcpnVmsmgs/k3iaFrAIjIe/gg
qidJ76Ktk8QwiE/gpDvVYoWoIO+PZyWfVrjjPk2zzGRzbbONRvtJKdH7zwiLQinK
cneL6N7HlbdhCE2laSoMT2i9Twgg7c9tsTKgJVcdPUHesOSkPe2WZA2095iOM5Mv
+S8TRqGDf2WZk+SLRRuy/Pm6EqZJws+UBQlOjOxngM8YZ6foAwQWFoWeVur12q//
Cb1GgO68R/TRR3+NM1ezm+RBxSPHlpa+bwy2C41OIVg8TrZTFSxHEsos/wK0ATx3
2HxamhQU4KieepWoLX6cBQ8kyMKWaY+GDjWc3rkGHdDKfUDBLqcvkW/NPF44Ee9H
lJJE2ReaeU1ztjmHXgAfv4tkAgai09Mql/1DPgEGbNQ6USv0cPu5QN61l90LWpXi
+z3hrTh1ig546w9aVfNh28VE0jQiSZWHxQ6LOSBMDD+TaLLMXN6Txk8F9tvD9YMD
JaJlTIRnF3R6yZ+zVzXvD7Nk5KeT0pyhynYYWokNMQE3OVVxIqNWthauE60sxWnx
5XDiVSR1XtiZoJOX5Kthia5oF2AR6DVCoy4ufX58sv0B4VAkW32oKLEFEf9bJdJA
3+aZkEuEed6ECENNB1LCFGjmG6i721lrAdIW1nC5qpbEcBz2dqjEwdr/NjSHMp3v
n2y/PqxlFGRU3x99BNtA0EsKuawGJvVRT2lPqgymk1X+tvP2Oi08kRN7uCqXBhMS
Ykz+R2SzQuQyT++U8WBNFB5t+/fn7bPWnydr2vUKZ9fOIZkZSQBowkqpQ2pJ0APC
340k1EYDf5tUT8ApG+s71ytmKpmra9EJZXb1pLShHVVw8EkfxqxLXUt8ZcRX5yDd
w7DT2OenEJESV/nsPoqjryLZjg1csJ4nZpxrw64IXHzmi3Lxl+Jt8zd/6D7qtuSm
JJGY56juDSgzr0y6hrfn4PSf19mEi3bLdz7jNsBYXzrfsHnDyzZwTB4F4aRLCdqY
RYUPdd7Grmfk/LsVfJJ0cBU8GmhclpcyGCEmro+38HHJov0uG69ZQG2WZzG/uNTr
9/M8V6C1aGjbn2Ew056Hqqf/WTuveIf22RzrlI8+fuLjyNHu0hSt5VGomI/oaeIz
z1zP8XTo26seXcd98meB8gtyI0g9lNTe7OlqphYxYEly1kymWYEFOO9X30yyVJSL
KCVnv8ca7wqZ4A7/8P1AgK/fZBfakvCTZIP2PIU3TbcONp86IL0yvfzqCGq+jUQH
5TRZb8LLZa7YjFrtF6K5G9JX+XtTDe4T2/N0qSLhybe3SdZIqNdouPHHp01noekV
urgzG4zu3uYEPXha+yGy+gHRCY5rqiCnU0m5154segTygCVpdnuldCXcP28U4XqI
vt2nxU8GSqJ8hZf1A11MGtSpbSHK3en7rAtuRv9TLaThWK+G5A5+J9FA7NMEeJe4
qQshiPaJdYjgeUbcRkmJNfWX7PSGPzWBXQIdsO+0a2IyGZ0xPOYBI+g/ZIEBgTff
L5i9C2ekyZAqfVGUF+3a2OxKwV2b8wgdiRfgEYObQdmxWiOQRG2ddx0DV16Aro0L
yN+RtD6Ra7yODH9T+Ay6hGt3mDL5m3uzHdB1b23YUC0I8+6GDZUmkkqhiWHqaFOE
jHEXgGHv2Pr5qIb6FbyRLL+TI0FUDwMCL+ZwuOfT3YCyc4h4tRTf/2jNm2NnHngP
j6CEy47jU3rPR2TcMrZB4s1wvEoq4XUUM+RKD7jpjkS82iKQQjBLhvIbTAgi8ZlW
llfOgNqSMgOn1Xx7LAIO1gyvT0axy1vHQTku83ejNOJ0cIcnD0w3GP+DUsLCzr5y
aOxoLrYRh8TyTII3MbQVcPfxdHiljpy1VbJF5UUbmmdoSaztv/Sokzj4mx80rG+A
d3dgYywuRRtsX4cYaaJtQDwfMH5vTyGPVvZbgXkXt5CA2hAjQmbjSUMDVysPa8tD
3xP2aBEHxiR3NVT+oothohLFvIVAI4nYKrTwZzcKNZgTJV5xE1H5l/iiO2D1Yi5S
mwDdL3urX1U95nnmyNy2UhME/q+Lj93voywUeMNzHD/7SwKp1sBLIOftCsSqNTZC
5J6autA8P4/Pb3Pwcn/T3+pMIMx5NG3P5VPNogewLI4bw/NSQd/yvssekHJsyfzg
HbM3rf2Y5YBuep391fd5yXlmYw4yRThgQCjOwwkBoBZYYzrGPpoL/RFfoDuFJcN/
SaQctJqFhHUw2dtClny1Hl52eER3O9lHOw20EMELZLhVMKxpd+P5yGe6i21/Njp/
r8PUZu+pVr8UdABkz7O//EhBLkorgECIcheeo5zlXlzy8P7KWV9uRnglWZG3ydjA
dZYSPq26EtBS1jwhK3xpSswHTY4oKfENIUPC5y7caFC1VCQPF0b9bCrH3ejfQ4ZV
Fs+NzD6ZZpWQbAFxgEgsEU/jJo6Q7dynI7iRKhon4qTJiOAtvhqpUYF5c6azpjVR
izGxAbuWRYZZK4hkPnUumXtreuMuEPg7BfNs7QEBVPYPjO+Wvyk8nGsbqXHp3uaf
hFaqCcFE39EaPvcNy1MKt3R3ELylCZtantFBfgCnqqRlDa9A9AhCBT9PvO4gr1lh
1S2Im8y0HiLqp2T/WbjT0fVJBPvNoYANdIn7D4zxepDoG+KCblwO01JSbZe8g3KQ
9WYQA6a7TtcEVotjzPuX/SuLXLnd+7ZxHAr/9kv+Zdb71n8ux+xyOmgeIAwi5Kcr
bng48o2intOQ1bQ8o/NsaUXizNzlFXsLBkwxCvOwjAXMUeNcNrwR7zCRtm/5KNo6
1Ws5EgvGlQmToLmOKY1J9Ubshd4Ex/HdAmhInkSDYV+oef3PNmTpHocuadkNsZ7I
9gyOpxrx5YBeKRIEJ0xdkN/kxenORJKYT9spOlCCugiFsd22quz18tYMd5wNyMJt
gbwC/vZl4JGnjSecAVg/hsW/4TxmcG5DYB3daaeZwj0rtg81qA857xYeOV0hmEgV
dABqFmQmxtDyk9DEPvAWOLemn3WPJQR8Kie9nBjqL93SLg2YGvtPoBxid5jukXoL
JxFBaKwxJfiNWIlnig8J9BiAmuF2yAyVRfstQHMPlQHFmCRsVvHts14cwRnLrZnz
ic8irsKj5X7/P6K2v+dIfmfZW4f956WkNsdKeVhuthlObSjAP7VWpk1TDlQQGhyh
yh/u7osLa0nKonryjiV+cg3LsWdFVo5B1OO9+pzDLiKoozHLA27JNmVFZV7IT3iB
kdsAEwSzOjNJpPt9oRQDHXDn5UW+ZbfDbMe9y5jyf2VOjSmPlP24D0BkxJLiugd6
EfPxw8B4OTCAr3CjuIbXU+GIaSg6FXQPGA4PijP84Z9EyXiTeslIClt07+Pdkfg8
y/gV2t7q1hs2ukHPcY0SFDmx2bGDrwwMoOaPxV4J88VbRyfwMWP/zchOTOfH1tqd
Ef2/tku4XzLYioVNG41eVSUE6mVjc3KEBZNULHDxEXqvbGRN3ePSO+EpAnXzrazD
vftt5FHYvbhFvKSHFUfoefdwLqMETipwbRV8InsWYzLV46ZdK9dR4JYAJVSpUwFS
2vQnNJ8iAxQ6oFyBnJ/oqsDvIHt5XJ58lO2fpGirP9Dar3H8rxj2Kh7WvgoKT6k/
ZASY93R9NI1ZhRtM07TzRCoPL4qgXkrotCW8KPdP4/IlwAbR4pVuYNilzjdfkAE4
QxjeFOmLgI0GB9zCmDmF8I0C1mZlvNAJYKj8jMbNRRZ88sKdAadowEnXhtqm5KXq
sOiWKezCSO7ygE86N1hU7v3Bgnifj9jgvbw3u4H95FCpjuV11NjyCkJbxesnmHiO
tefhLtkU+lsulL3uLEQzA60FvEyFlxzMQjofej2YW93xJMwkHBuYg8s4Kj3EJZ/D
DkSN7n7HXB9XpWjhcFxivATn29HPSyH1w0qxG5JvX+5GFFs/fohUN0wEn5cc0gCH
AukDsFLpYoRP/MCTYo5qQSWA/Fmy9qdGBUfpZeCnazoWOCNh5Ss6KfITrnqSFo57
VO8smklNZA5AaHi/QNxbknmz611H59p6wEFsZeuw7RhsvRUgAE4if2Es23M2aBsv
xKZpp/cNRHVsmTvFlm7SHECwhPbCpe9vbJuYAYILsVTSdeaCpszcnqfNnnStj39B
E4N/ivDgLBQz1wlPH2mh7Ca5Y5YiccApBU539DWrTPxwrzX3ri4GNqXqP7ntkZBF
wTlcJ7XZbzquB5+ldai7SUpvK14nkNkaegjAjHeBtuDgbjkX5EMhel10H4kjc9SX
Jkx5y3zg2d7aZ2ubYHxE1itfVgzvvEilssmKYGdbD3YoTOjZA7e0ToNfH7WSmHxY
XaRJQWhaZNavL8TMXT/SXeUCtf7KpBZE6qaw20qxaUHWAu/YXwl6aqFpY3QBgqBQ
tnlBsclznwedtHX7xp42SAFyHjDxRVnx2vCa5KauLmhUWQ6TYEUurmtxdU+YzSem
BAA7ozk5zCnCPmOsRrw9m5C6SWGA+aC9OmgMSy382fChS4PSc/hQnYtipn9FUD4W
/M7T+i1pisMQi+JRVEi9k+43X8LxyJJw0MyFvo0+aFdJ5c+VCR0X9eDgqSFbduqm
1Eeom+Lnry7NkZPDYbIIZCY4aPLn8SSi9+ZHKnMs0/Qxr3wNRXbryg0D519D/EHq
E585DyETIse/STbhnO0mS3x5TMSM9Af5dryfzUZIDmsUNv4dsGQ0pv7NsDHxVBb+
4B8D0mlpCXC3EnCB1q21olIue2zDMvQ3+cTsMvWuRiwu1oknJHBmAkLdVSDfDHAH
MViAZbOP34zAVd1JC6saQXM6pQPR03/nFQL4QSG+m4gKTGM1UyD32L4uNO6ckkaQ
ZCjFaLvtt/ldA2/E0bbR2+Tqy3gzI2tfaxfr0TuAT7J92DpIYIU8H5okdQDADAJU
KRX1uzFNNjHcQCP3P9EmIFbU6uzWkdPs5irlqLARKBcN0C8O6NDESBHUNNN/WN0y
w0Jwt3xU1IvNPMFOq2uJ0miqydkZ48WyrGmjKhJMZCRdWgUrXrDANDJrDI9gKgui
A6khbEwdF48YHeQscFpuLaPhUqthwApcGjg6PXIO6QUBLsNwuVMDK7WEV0vkqyjA
wRAMcN8C2gyawLclKYm/yZyQnjmoVEMlFYivSaXuVd7WX0NphUCocKMaGEqHDcbw
OgVGYJyN2ZpzQwy1k3kpptCWHurjHe7LYbEPryvdDcsGnQHQfeE0RizzIrRUN7oM
19bVfZlnv5YB/CrOwiRIoJz9TVJH5/JnUY0Bt7dAwD1M52fNMm7bu7Jwwlov3e8n
4P5mo0khT0PoIFBu18p9X4+DJTZnGkJBdjfoyluITXj54ZrpUoXYCVfii2Xf/jrq
gkTUG3aOs+rQciDX0MmKk8FJb6uitQkojmsdAdQ8UYpPFiAVIv/0fHI5Jssb2Qzr
Uza9Czx5opeCi/J1eaKWSHIxtx5Cw3SF/dy+/HpfqLX5lwxZ8YuTpAgWbGTCoKaT
gl1suXMLbSoYZL1pyJouk6zGAWHm5ehFShR4EvV6984b4CdVJycTUaMp06zQbBSd
fsR3QxPf3bXGIlbJNPM2GqbOD4Or7flx6R8YH5RuPgwVjNxhknf+1zn3yXQd5u7v
ijF2RlhDmJcDRvA9UHuUoAWZISesNoUhV/4g7e9j4cYazqUIoHJ9H+IU/tjKM/K5
4xL48wLISGGmQ2V0sYrIcNw45dbbuj81QOT3OmPvnWroTFtl3RWt3+pw0II0qQ6V
2emIlO5I8fiOsPYiv7nxuFYxyibs+y4iLOhZ1QHv87pbKEV4Sk45Qxr3VdhqUp7H
BOaiNNtASQi8UHkA7P+OOL6bhM+ScMZmT+2K6uFYmvnB9fHvAyC2DLZOYOytoo1J
IQRLsxfR2pMhgCSAZYEFCyZC8v7bmR5UoIP1YAPlBafoezFbNt0Cwim4CxIMFsPm
mTzTDZ4MIUZ17pTwp3/W+ixUmhojpYcYwVgOZ/yYuhcAAprlcU9Vr/9zrX+Lg0zh
g6lfwaTLP3SDsIOEpiq6IqnWBPrpaudkE5HIVn+pGMeitrN72AHZh8rh0qlREGLJ
rt71aHXGeQnGYM1PABaPz/VIlpRfgcPCn7pomlyfjwJu9DJnHFFyX3jwvsXbMFzQ
XrkjTjOao8hL5SWH1P3PYoa6vtyQYk9jzbKJmlvOB898zqZbq8AWmKwjif+sPZEL
odg+kUM0ULppKZOCfKUBkoK+WfHZGMbLk7DVnPuQWMpIj9OD8vIhje7rViQmoU4T
7M7wyYAI6n5hAgojb6Q104IusUDSLELV0RENfwXL2c+X0jhMhZX4dlXKUpLMLnb4
hp7LtRNoYrK9kj9PnZJm+aNb4jY3kJ9v4II60dtki2MUoQ9ngfoIriByQleNn8cD
SVcRIhFGjYYAPPC5nJ7cDAcCjwG/hJiRhT6ZOo7ARNXJoDxjfn1/R7EqcA33CYDe
15K1F2cVpJlVCCIumQjBZEn0LS0jfk7xGND4SNmLBMJGPwyzd+gW4BNUbWYlE6ST
FYIs5jwjUJSdJghp3B53C8s07xyaiKR/qSNQkOCTm45Cla9/ISRFLqd5S1d4rUqh
BUSyltUHVKIyYFgHajWESnxwGHEDkwwdGppN7diJp/juQNrJrqh2bXHMwe4UoYU1
kA6nKoeN1A4v5PoKXheae/BZj/jsp9KThDw64ywcjWt7oNCltdqDJDMCg/RfCQAP
zXSJNGKim8ZQehyb5h2pFtbcnTNl9Kj/yIIAJ0WBhIMcVizpxbCI/RXWPQEtM9Tb
lUEcRgNw74e5Xfn5Hn0fTf+hpOayzxR2qXx1Za22L1bky7CM0N4XGMC4SwigfeuU
Of1IZkcGVfs4sCJLZX+fUbAqwSmUBR7WqixAZFsgCXgdrsRxKrlBY1nR4j3gH+lS
OXp3rWAS5w8McEsH95KOkrmk+AOZPq4los2OBA89UKeKPRBRHW048QdE8nHYfCvd
sxZjp9MkAWUgU1Czv5TISriN47Li7DLxTs5SmVtMcvGbmknFvB/I4m7dJwuMtJST
5B3mqan80maAJoCV8jb5biyTuMWJz5f25Y9+P5ZrHhxviJVciJ4dKhuT3NEFRus4
7mnVXL/zGupgztGhmgEafVG8bNYiyHQEK5w8ns28/afQNgiQ3Vd8FVQw4qD8EaCu
ytaVWlDZNLbe2HhQYWG6FtvoRQQSp+aObHJpr0VwSu85UL1Gk+kxeqNC093tSszB
ZvMoEsCso8FbY9rE/+AwoWhpL6gGZW8cXvNgCRiGeR83Xw7TeEDMeRpPavb4DBT8
pj9PLnfuXh6+QEk9psNBTYdIAvkEXPIF30lpTp7chSuCYDOFSMyKGMGnw7mxcKUr
/F0ujKnzRINDDIPVTrlFpgTXr5lCyWE5+5Z1dJEsSBk4W3P0SDkvwFZtQL95TtN1
34ejwsHWwXbkIskFRVgO3tGpjqEDHPMSOAdSsY0HpraOYZBOG35djy3KXF5DaCmq
DLPrWUbpwwkgZlcHW7WQ2V6BR4b46gr2unCXO7r/iDt4W3xA7RFAMmOMMagLxt3s
MInPCLo4woJky51hUw9cBVirq5mRqcaMj97wwOWY/pMW6Z3hMYssc6lXyTcCBAY3
HUa6UvwllAg+ag/iAxOMazurmgHfP/0dBSk2GRJOL2iUgMYu3Kx87sN2caBZwB2P
QNDX1eRDuFSr+mDDIigxo1q7RN2rzd1+iiwf2Q5EmD66vNNkopY/TIJuDtWzJpIp
qN2WIb1GdC0XgslODB/IyUr3YBU0E/MWEeWtpeavfZknCB/bhsGByJaiXTHd2S3f
l9Lx4MzLi8tSB14j/JBFGXtY8PoU0Q2vNldB/Kls56m2+TCqUl5axopXy361Lgr6
waSeTfDLVniF8uj8sjyueVWhzB0P89+8Nhk4M/ZRxgRK80ZQ3rjs3p5ZnUuXuWHl
Fyr7y3y4GDTb1iilc26Hl9l8Z3E4AgbaPu0oXPeYP6wfiZrUqQsCkR5TmZg4hCnw
skHDKdD2VM+B9s/SRf8ATi6mSSdJtBBKRx+xnbb02K4UBBH88NQ49tarI1yuAMad
0NaOhTMBC6maC7hdKzsDxU946K36XLSe8lwb+x7wvSHb7fDPC3fj8txKC7rieGCa
CDiR0VbRhz7NAVjCj6+Hp/DbgdbyzJoDBRCwuE5y0vjQbVI97KlU/Zcehx1SITlP
C4O+ABWwUSYbqmVNmHLyj+ZPuc8XWgtkX+tFCSTgbQjDaP8RAcpT22Aul6isQZHo
fafwNBm7xuJJgLCvmM4phtz1ojv5u9M0EDgItlJC+QKe0PkktvBrwvzi6R4OlFKa
tSUZBVoMI0XYVVfZiareBUyadHtkSwtPN4h8DdEH8/c5lag8+Vibawj/Tp8SK1EM
tByI4YFvpAIbxnFYqA4q+SPxa8MObhk4JXt969j3eFfSPKZocYhnib1/girjjdb9
zBRosDuwfWpIlAqkXEMjFfSlPGTBPQ534E7NnMD4YGgxiDH5yUIY61RMbS/dxRHT
iMkPjzMl/z3/bBsVabsgAj0pPHnmWfIsA1QJ4K63sPx92yqkhAKS5BUEOYzikKVS
Dlx0/kTDIgGfBEoIiI05x9kclVRX0T7n59yhl6BC2up0VBMRDqMz3+qI1iQgAAhj
Biud/EUm+5jrheyeg8Juyul6gcNDE67WEG5Q4WEmW8ODnU+lHlf7l+v8m6rOOtKk
lyXaIO3psHPzEVygtWzD3PZ4Ks8fwZ8fZ1ncZ3/HgVM4otOGAMrNJ2LDdsiy/t15
G7yQlGdrLJYdPF4F1m9mnkapHbQa2/F7IXsKHYC5dQFc5c3R1zPPQFipwzG6sSF2
IJRJ2dYIZtYd48YAwkIlr6ZVIGvGYHYkY3SCk9YBlldndzrXXhCvN47CBuUeuYrv
0gmdq16Q23tkgTiPPdHF4MPST6LhzlcHh650CqS7vr3T0gVqfq5glTvqz8ar6ld+
4TtX1rTdiml1wiy/bZVgrRtLtL1MWXhmPw8wAZgrCXrGD1r4ZwPUlfExXO3zihpx
VVXHUQS28Ep6GeRrgtD0t2zeyK+2AW2IVkLrcETAdLAKsPA+nfV8f+q+hO+qotRB
Bi9tTS2EMLN0GBkTba58WYNzwodUJz3clRRXtoHdadw6J6GznJAhVRg6zfr28zVE
pjLsjxe5Q3NsKb3g9QBX1Mxl7EtMXzgUSv+m/uCznNaOClSFa45lxyPze7STSfAp
PkXtGVv8a5h2FfzMXNwQXQcr7MK76CrxOGdZYnFUvR6QusWTZ1I0x36glLOpWCUu
qtFbMMqw+N889ktjbXCyuUpQpSTlx4vuNR3r5q6lm+uNteoDVbySwzvsab/QSUk6
C2wykQH4dwVaht/x7ZwFlAKgGA/7Ac2So0xfxuMUHhMqpCLbApQXOTOfvSQ695nW
D3bJNaaFCh+qx2McftUX4zkgrXXXjeSsaxn5cJhTPf7hTM01d6sccmMHHEvu+mjt
SxWPE8m5MqmTgSZ5XgzEdDwwHGHXQHAyOE8d4oDFeEnFoJ/ZB0Lb4dvYDNPZ3wIq
dH4Fx9uF909yX0/LHkOtHKvPAKCBRt0j6K8Dw3HSLKyATnxrXrt7k0GJgZJUTuyA
efq8rBnWJswoPeTPEwApj6NvUmY+w09a+cOLjsda8zPqTTI9aYxY4nVz0C5S4QVo
igvhDhE+Sn0gRYeibPdeF1owrg1sWTroYyV+5cl87aXWz6DFS6K/F4PLv6Mj+Pjw
W6K1WaYcLii/8f2gyHqS+ZQ+2+pQ/oVbEdktO+8BeGlHEAtJKOP5IpD1ER0VGxSb
7HoAbcIU1l3xViZHYIG6T7ecs7IGG7btF0Bnix4Hh8P0pEu5tIEximnwPnR/AHJm
pDsisbyQtyhxxM4XwuDEy8fldwsvZ2pmTstjJ6jWdzklAUyYk2VFILh6Zk4CCL8G
613LlVJZSSr95Uz4ax9RqZu6Ukos3FsdQPguqw3kGJPSE1+ZnfCcBeiVcWU2Ha2v
/PH8QM5J9XV5avdWm5u9DgphZV8zYM9WPj4IY36TVNDln4mplW8uj6mRPZ1UivpY
yklDj/yOk2rxXoDrR4FHNCIpFh69XObMb4k/j1uO0XZkcuYIuWThSbW0FnzpVSKl
JoIMfUkumdX7dBy8XkEDBQlnuxb6VOVAq92WfXHM3uGy75Yw/xL7KVbBjUnumzfd
F08OWxTveCkTRVwP9Ml943txB+V1fRVB2595w9+iEfSKUVrjewnREmETUt+HnwqV
Nb9xOAKj5VQPuFEC3WNiSKub3rf09PDRMCtPv3+CEuM9iTeOfOuqdxO8dFqytlE3
vRS6L//dKLzK0w8K2bw19vhqQYyODahDaFgB6IqaBpv3oNv5ZP3XmNP9OtWd6o13
i5FD3CDGgliwk0OweWfcXVbMbVlngBn4PM9USBT8/MuIS6xmwevATht2hUwURFnc
TJp4nsk2biGpvZ3CziKGmYMHqOkbt1VE1+pbrKlV5+so/n53vgKu8FRgF/96gosq
lObMp84qyEFoJSWbQLVQD/67xmfF9vRFGhTnS5OZa6cbV0jbpGtFkXHHiN6F07Ue
skl1qcFSxjpRiu/Gmp/mmZDTSCDzW/NDHpI0XUy1l38kgmF08L3+h7rgoKXoS7Nv
YZ9NIdXxMOzISstxK7uo45kC4LJECsC9lFwIwKUQ448xSruWDPprLzkJn/kdcGNW
0xLTmMIgXj7fN0zH5IFknV9FgaitJNnSoj+102x2s1xSs3b++xV9AAdZu9cgbq+i
/HFkxI8f6fNjz2hyCbsr30exHjZW5NVbIxtXV9nVpB8QkOHJ8SXSAW6n0iBk1ld7
J2TcwcLFWpwSC/Wb84vkSnLo5JmDolEOAh6eKl0XNpazh9GrlJszYSLQ+SDmcdMw
2vJbfFIqV91py+eXKeU9O4DziVytU+g8QLzW3vJsmGZ7XlMx0cKme2nGY1QCFPhb
A7mrb2DPqion4LPtUOwBk7hI4w5EGgeVi+GRbfh1GRztZGuhQfgmeO+PnsYpU+9N
hx8M147+7cC63TrW7P5l4TVgPhTtc07wwmduDAbFkduBpaHANlMh8iLRRcvyk4S5
8POZlLVbkicZCd6F3qAZMSY4JeQvSFM8B2ipOOCqt1Sij7/eSbZYtJ9hcHG+9gGk
bwqGlxwYj3Qug+EYUs8fbwGEZxs6SG0xXlNzriU6K/CR0bOg9hehO1d8GjM8lNae
Iw8hixr+PiDWwWCC8RbIIkL9ds6mULujrAW7IwVuQ0gRYZNBMHN+/hHLCSeQhes1
6qxcJ41XbDAhLoQACLMTy3kLYW9p+ToXNPX27TAU6ckmbRYMBj7IBdStUvLYzu+/
r6yCmkYLSsXSaM1qVQ7tg8/j3qTXmaQyABiVFbfF3/DDDVfT0lkqySmRPUfwErm0
BeNDG/5LJnidW2ls+u7Ct1Dxbi4NaKrTqbbwx9o/BBHthnOimgtIDs1b/XVnGOy5
zJlzzfwCtxY7iCPef1oEyt/gU0+cU7vQHeMmWs+gMZOlYDuEIlOvVl8AVt+m/qLw
nOhx/ZqDYoTqupLassuI3X4bVkpvfXucyIQFaW+oXnGXMyGcR32TMQ3VtbmhVJGA
2iOD4Eoni3MTlGZ/o5sH/Tjthg2g+bRePnDojf9BxUVgpq3SBs7Y8DX8eFon3eJR
YU+GIryprg95v0h/E1aWOy6bH2u2RdFBsQkYtQifU2ViRqeKxnQsh1TPBnMG4kfW
0Paimn67lxzaKEdVAoTKCyFe/w26FRCY2dS7+OVGEgAmnByPrYjf/aYVrg01jmtl
SgbKYOuEZgtZB2McfcD27J4PV3ki2zkVPFIt9cjSpJZ/JlmxjOm0Ye8LbHlMfeyR
qgSXPDqBgOyXYzBsJUcHt+wwj4jADgl1K6ceJjkYGI88qmfeZBgdbezGXMLLtSMK
YjIl7fG0aNOfKDRmHcPH9F+pUb+W6nEMyqguXZqosPf9qsMLq5aHVzGQ9n7ELCeJ
laviieSYGmRmOgmtnozgmBZwQCpVAnLRPtLZoej9yJXBqTEy+nzRpZbI1+M5stcS
9ovAlRGS2NixTFy120peBt1FiGQ8q+L8MMYoQC4HuvtDfQFNHx+TrUZJg2Ni5AWu
zRDKBr1xky4fP/e5BqBw4BdQHsnT+ja/InPSCWufhbJ75MKPvF+9URD1l/VQPgih
9cTaM8EJ+7dwCosEr+UW09Km8eZ9ld7J5Q0/lW8eWVCuUBoMMDvCITqnAkvz+tqd
qVlMdkShwZLOdWcG2Zig9Iw7QzDNrcS9mtqFRgdQPt+tAmD75M4wk8++fylVjy2o
YsQAxKESkCvM9AFWHA54SUoFW2YARIAwDovWSJELD27zTxM9lqgwZ5qSAutd+vNr
61KvegDmEG3jv2DfzaI14ZNnu50A84kt8G7k+PLe6DwLC8KPBspGxClbHd9ZGURt
SazSMb6lP3NS0vIt0wzqct7iTEzSk6qmvpVuRB6rcw+ZYyQgvZ4sXX0I5En3Zn7+
2WNUvaJTjsNCY3dFNRj1nhQxQQcfymigprP/G9rd1RfFKGpUSOD6dyW4+WvDtayt
DPN1jDIH/B2l12HnR2cOlWTpQB+wAGSoG44dDQmNmwySlA72Il6G19x1n4qwof5s
+GxXZAmm2ZbnbpSiOWrMXCZqkxsnTTHDPmY9wzl7cWrCY8Yovd+eT3f8WKGI/Mqd
WU0RdToVrJ5/ZVlJPIuVuC/AXraMHjssc8Qf1IqMCcZzknXaI//cAfg02/2YoaHY
A5sCAVC92qFU9nPEARksz0iiVXvlvRxz1jcXRIkDxELu9efnxF8vKI9wAbqB/Wee
o/rAjGi0C4R0JHwROIj1iOoY61X1xnE6I7gil/UM9aKfz6bpdLDWrkIpqPeaakm5
Cumc7U8Ddy3gfKL6cLTsRz1M/9fiolmPvs4bkTo9ZKfjClwD7bvNkUT4Nq8QUHJs
DtWOlha/aMLCTye6sk0hF8SD2aQG7ETHaoQ65fe8KGO+aWiobDiP3ZzsUPCyXyyb
jYibR9BTjNfnUSOgqTfiGA7srkV++yuBbsg6LVQh81OiFCz8Be1SU8gON7WnOQva
wQy4O23s+lIAoF3wgve9ecH7jgaUfpgXjGwUcgNLv0kSXl3Ap3n/ZuVCn4a5JsSR
cTZyyOzFFnUJ881USXRtHaBjAg6bod2ytH+OOhN0xxR084ORACWT28kayyB7qrLZ
V++EnHfhtMQ3+lQqKXXlkbBGz5+XNPeMtctgctkPJwXYYGjxstC8Kt+qt6WFKR2U
UMmLmS7QprSeLxS7Dt8T+rHMQ5cVXzoR/L0EnwEZUGUirn8T/M9+cOBHe6OdmvZ6
YF3I6ZrBHnmprj31ZSHvs6Tansm3pJ7VEDqTTFMSGObEQOMyXNGzSt0C2Qpvwyzf
mRG/uLjOJLrYTIVdVandJghodSS2RBk72mgGcoMoqwS5wuaRSay55hUoFHBgxz9H
3y1lV/hJjy9WzL37oNeeQvFovuu/hpBOhGOxaDJye36OMnP1A3jIV6f0agJEsqR2
mQrbdvRKA2AySC47ynEnmCeMxISOA84kjPxV6FcY+w9/g+rcrRWYZ2O+qaOpKVYV
p3dcbR/VJgDUMaYuroiNZ3dVt3CzDqm86IBAfuzpDQTSF8e8RPSmlTOmMcwGhEUB
wfeVdmMM5Ed6k3x9ySss5+yboaT6TuocbDASvKJ6Z8+CqSj0eJjUgEHjbD6gCsqa
IC3XyKVlVfsPqLqc/MNXyq+Yt8wYtQHzwDwfa3nmsZHNrkO3fG5+tdaFAgqeIjfN
Vge1r9uNhSb2IvNba9bVryDoal65twZXTE+kmW658AenLhCiJwjVa0mFAN3BSGOt
WxZl79FnXMljRNyicENXBP67CJejWOejWbiNEuhy7KHr47+JTdHQljnsqEMDT5wx
ntTNyljMzzSmF/Z3YFFFOrXM1yuU8d64Vru5aqlQGKeRx8Wnpq6Juj6GSp/1esAZ
BUoXv9McnN5PXu2Um8OcK1SJwFKwQnbA6yjmljYhmy/GL7gWWJXp//Ti5b2yXqk4
PVhHH3Kjo7eE3Jppdi5mNyVkGo8ZdSuIWkmuxO67sgITnsyeziWCK8/89OduAYAq
JEJ6J6JRzOGVBzVTBFgGbu4rKajbhfYexxxNDMeLNjZmoS4rvjt3ieSGUIsgA+8l
301x1gyz12DRHV/NqpBX8iCmTsh1SwwbeIgncNPL9qHtVri3QtBgprt+gqSmXFSq
lx5rx6BSu0wjZ+WV/4H9qR4lno5wHlKkIsnNnG1jLByvv2XQ/FdzdxAd937zFPRG
jW9UDZ7Nz6s+ymq+2HNNzK1h4koHYPCnv9+DMwEFHIcunHPsEFXc5URLYwAbINN8
4FbWKeWfywVj6+2o7N4VcimGmWMcmarPH3cNRpjtSBGh2aW+G/1JFU0xJ5n6bNfn
w8K1InGWsXqB5MJS5JV5gyIi8uJVU1NDyLxmgEsvko0FHMai0HIxXKyKU0KH2tAA
IqZRhWft3PiMQCwJAiMHDE9M+B8wa+emsuiUd5rsSAU4IpWsTNO+VQ2rtDHfg/Hv
I8dgDicdEpsFy9n7Mq8BBvfumXramvGTRY3cSPDjJpXqamvwzJwUjBq2LzStmUVg
NEey2B9aVc1/7NE4eUwAzGqFvMrZXjbI3P05w8tMNLBHQTkgmLy8hc96tbFVPUU9
JQIZo1GEoI2mxjPfY2/RCGuJA7PRLrGQWe6q+Udb0C3vF6kzbYSUxJ8EybLAT1kF
NzmjGhHeuhRUUMULUKxMHqZc8VnuRhr7TdGUqoQ4P7vfbUOo5JNNIJ7124NpYTVa
cNKtb2I5709TTlzuYFYS0/K9AxjebQpEAsiSO8LQcpi0S1YU2xJ6tWCQBjE9KU4E
xRpKihg8Y2gLTbaePg/nQ3w6+OYriXcJZXRRpHgIX4aVuzwkADWdyP0sgB5rcKuE
NMdq9KFwiHIHIKv0h4fMppSKTRCyQq7V0IPuujd84ILH/S5xqD7pyX+k/cWz5+Oz
KRfXd6F63gZ8+ON3x/PhhhOi1SQRTFOHs6FOqneLvRsG+Bm2Nf0Li89blJVPT57C
59dvsvOyse10MpxFTCC3DlmZ5DSkfN3XBTPMOWiZSJuiI67pXYRUOEf7jmM/wkLk
JmZdLd8ae9Bw645ByabYb+eC50ecmM8mHwXrxvZkEKvbuR6KDUd8+50y9T9qhwyz
ZZ5QTaoEOGKlWrweF0p6nLDEdrDq8BULbxkZVJxPlq5YFzxCA+oOxhdnDcDA7xjw
Z5bpHBp0t+H/0LbmghlzBeTLu3cAccD4MDN3oSBVfspLF1yxALwzNppTmSjk17rK
QYa4vzxBVH8GMnCutZfLuFA8ipjydYkgd77hkoJTi4jXJGKQ4EYejbd7xgrxzBrY
3X/ArWfLJ2gGY5Y3kcwsqiHHZFHvJU1BuShX8ayw0Lm/T0Y0zl9uk6NQ79vfE3Bk
/WBnnTkP99mgAy5HitHRDLM5u1Ld5DwfcpsfJI/b55M6zhPVFdp2VPuYtPyxYwqV
RcjJo0wJMclVsi7w1Ct9DRpYkiP6IpO4E0vklNjDLLuHGRa3JMJAPqGUMQ86LHE1
aQHCX5iPZQq/Iyg79SsyUUnB6kjHXH+Hq2MdiVWR8RScNuZ76C56xJcPUBmEnC9T
/P+soxzhEbZrOdKozmc1mduDdL0PmEtjWoQr8koOc1NWh4hB5A1YmA4A6t5bxXrt
QDfqVTAigwTygrSJxynZmHzn22mA7UuLCaHXdWZf4uGUjrOi5Eq+E6McWyV4uUFm
GW6eNU6/caaDMLSG59WO8NPDT9Yjm44fxPzrQwSoK2h5wfXs3QuKS/QLjvo7omWR
TE/ZeHhIfpMQIZd4F87NKQW5fn06P6E3But3owR4vIlJoa6Uri2Mg2fZXElQSLMv
aFY0YfrwyFb/pzaK21rCJxWrS3wjFj7tcr0W/6YRRIyeBnxOStUPlvsILJsNBz6e
/GZZox08jYpRwyHAKbg4FpKaMJGj7g4IGtxrX+UGLW6EBu/Rs5dhu12Iew7t61IA
K34IKu8ZYYWWMyyZG5EVulEBNJPocIrt+bdElTUjVcEmoWLep3pWl5Hafqq25QX1
LjqVjiGHLZ5L0M93IZh16CjsjwGQgehK4YTwNj6RFLrua9nZQuJ5A74u/tqNxTPa
ZOcrEK6hA7HNtg7TIEaIsblO8/h8e1eSpm6o8hW45ZXZxANLLKu9B3aGhzP/kolO
ghYbtTDkYZvwYytoqfcm8Y/aNlMr0pDEauINnqdccaXSQ+CC5mDJ3R4sI5M2i+tp
Kj8mKw6cdp8L+woa/LRGbF+Wf8A7ND3ojioKx0uIBUKVU5OtW+P3Q5q1dxQYFI2T
VhGmHBnU2T0rntUAh0iaHTrk8mAdtDpgvCZj0nW2Z9NtrbQgvspLA+70u1VqFu4V
ydeEkQSLijS2Aw3WfGVZkaT9wD7Xn8YSuYUJVePNw9mz4Q15YvGJla9fPkP1otRM
/vR/3pOWwsZamgXupc3rQ48iG5MG8B++94GWTpm7P0iSKpsn9cexZnbW+e3HifLR
/ilVKYGUWrmr+keKGIqzf7JVCpFxmg1JGBGN+TRdAh9cf9F7CGxiAaZ6FBMv9jep
4eVkTTjf2sWEpXerpHNfbT3e03DCkgjSmC4UH+8pSi84+XyKru8R8iL3413RYaQw
S0Rc5pdO0aZFgnAnG92v86BmQmpVz2IMrnan8//y3OkK+D0wh5F/Lj4TZuSyMMvn
Q9+CC2B7ZrnB1XBLwtQ3VwolwKAoXviA1XipIFitz2GYZvBUBidU6RK4HsdrgAmF
okqIivR1paBcAR3GsFpv41GZ8a5b7mk04FSgzEfV0728JY+t+of6VO1IclKOOvMI
5jtrzDySIcWpjij0K7m4d6Vc9SliEl4aQjubpHrZePBFVax5Oyqc9ZcLLoPmixHw
PfG3AmlJrPGmvag3rqHQDOQGg+abu4YhcZOwvG1m+pVQPLyQ5WP55jI6EzymoWg3
/sQ9yjI3HDmOvvcLZps8x9EG9dlYzk6tULEE03P4Ov0jS4ebo1EMvKLSaSWxcvM3
UajAmyFOHX4uwsD8tode/kZS5vfCKbkXpSC2THwcQF7gImIFm3LS4fDK07CSTQOg
NbH8DRNjRmDzFPZ/PM6WvwrQXoDJac1AJyiEypO5VQzVTmBfmGhpuI//GVVdum2R
B6yTZaTtG7n1+seXRG0Xs3fA8NZC73cdUr06Gbo9ivAGTng6vgpLPCgST7eD8ArC
qwSjtGx8+AsNC6WVDew5FSGW73wlsbqvnKtLCnco/vJxr6HR3DEqhSi/WOK5xHUK
bS9bBvNp6eZQtRa3RoTPzzqgu8lsUKgEDbr7Uql4d1KH3CFD2lN7R9fHf08LRoKp
aBxsQReoVA53998L02PCXW+wFmQ3o7zvK1BGEME7of2oUAw7787mPJ1roI+9JjlZ
pnXv+BRXa/NNWi+4o/Q/jyqbqjj/AvhX1tz3oj5E+TS0lkHDp2pRWsY/m/gIHeV9
k+P2knD0Xd+Drq4I08ynfORv/O6vHfWcowbqKbq+63/OZ6gZB3XGlzGAmDnI788a
35fq1B71/MpbDw5jByqzML6sCU0UUozE4N/aWEgghOzulnNvfhPoy8zqEIDIYTeS
/rUgk4glyM9wRa/pJvtGMRq+BotsjTkyiYG9AxiGSOfbIs3PM4lnl5NsiO/fwb+S
lcNOdblUjhrqohrqlgnh4+QLUoxoM8JWQkiUDNFHI34Bw7C9bkCJ5KGGPeolsuIM
tq3mNLeAAFfQnj+TunAhefBSUFSxrlBcageCCPPkJH2BJ8b8tg+GEWD4SyHAKCMR
jzAFPmBVTQgsI8rbvOtT7CLFBZ6uCA7X06hU9r2MdoeTNC3MAQuaoZw+a4SESpMp
PiGaZNKOmQR8zOBsQLTgtF0lYas83cnEqK991OA+8qKuSxilZDx7TnEMRTmeCUX2
K4JQ8maM9gUN9c1wJZV/TxPDdfunQKVOffXPPkq04t7o9kMgwIwN2fuy49itOXQb
3Zagiew5b//ZHY9h4DUgvc9A3HcD6ezWJC2QoE7o6sGWchaHTz39nXMUES1+RwcZ
4kh2/+z3mnLw+NOb1cAT3tt17F/PXrHD1gCQKtUtFTawfQaGiESa38NHXgoBx2Jm
JxkVVOzwwrLLt0P6lFjWIWHPCn2VPtG+FPhp6YRCW2H8Fu0+/aAWzKFOFm+qlVzE
/+LAg0lvg9w1GUl/EmdxeRHLyEXcnWnaLjgXPrsz7Y77fS8c9C83aI10zeU1tXFp
0W4P4hD52szBk5OHc9jl8dHy0KuGc892sD9zZs5oWkO1gh2NBjdxnikHJ/eJmGul
QiXpvlQ7wymcYrcC8jMq23sIPAriLN4S+QAlCTP99CBkH0n0e5YmjFtBazCAZXIp
7u/usd20Q29Mu0cda5fJ6id+twGy7vbzz8KNzhGtPclH1HsES1DKt2RrlaZLvrN6
lyWO2RHsX7Z9TxRhha090irGURlPgWrzeJtJK9G/5BZtyUziw5VFsZhPLe4HRHwn
1KBN//aEcv1R1MQMxeH+umT8+Mdui6M02PiNBqQmscAtmk5bsPpeI50JFIjT/IDi
6QE1rnL8QW/aOk0VM+8qww3olPYNyj9G7tY44lB53jM8kFOGyi6d1TKA1QEwUyyG
wvp362N6CjBWGV61MWaLKo71pFa+tIbSVI0obKIvA/zPCd+A8oaBmT4Fjh+R6dfo
matqjmRJB4XfMJiAdebESOcn14ejqQVfnHlSO/pewoZldfDR66NL99EErPtt8V/p
gZLNjpEswyto7gOiPbbeZSy5wOeXSPp4j4aOR8w58JWRBOJn8eS/b0skj7ha+UjY
uMzV7rd8PUrgAqTPGKNVxSz0JOBBk0f1rbAxzj/C9WGrgN0byv00jFOsG31g2yD+
0ia1Ah0eOSf35QurKGVhN9aM/CtkHjmHA9bRWozrVAK7a7iR6rbiwXPY6o89E1zb
SnPlPQkx0orszALrAImiwulI7YGwktLfbecK+dbxhFLgA5Qqjm3gMVecsdjzgT46
t6vjRN5MuNv/DXyqSCRYmU4d9dBon93xpWmGLYfcxD6m719dYrAqPskNTmRGNrwq
sJxaWoja3SF+QxQ6T3O3UPSXbB25yz+OC2bMYMIzBdKAe0CmLMLOCwpyOfwiZF39
Un5Yn20sfLBSPDIcBAM1Np61Kkq4O8Rtu98gf/9ItE21J0T8wAGDvSHEzCmZlkOV
D9HACao0hI4RX5tdc4bzZYodGyHRWH2ud07xP2S0Ysv9phyPXgPJI/L5KM7dWjOf
LB2F9DIjd2WXgFwq3yaFci5RfMou/keq+HuyLrBDBoTox7TAaz58RMBnZWR2I2Af
Vb3FB8SErg11wbb5tAV1bS/T1+QoC2jR5n33pN3OzBEMjHtoK4K8QFWiyGcCTJtF
330Yc6bOhpiT0WSCTwXzmZYUPuFjzewOdueE8IoDLaagmhEKfnsofIzSIzVRDKiQ
PEyYPsqZKQmogeTRZGzEU2fqPrj073W7jExv2Yq88KLCxG9x42nagkMxHZpubxsy
1udMoFdn1AMc3MSxrJlfKykwkEfFGuNzk5HD6NZG85Ig/7X83m5M4k6jeXE/s4R9
mUqg4uyse9QLsArApz+qsEbLQCSuS2/gPx3EoD9isR2Vz6jE8ZeD7e3PhiRJY37S
G/+Fqu9/LkpdtEKBJNrGslXmh9ry7zrq1pMnrFvpBzOZqdPcZuZNH5YHZlebA9Av
P9XMrqqH1BMmzlX1/P+OvAOyH/c8dSPHToknlJoQCPMmlT64jUfGUwpDRMyZHoyl
yqFSAD+THWCbSCn9xxVYekeZie12pKWerH5lEFdwC7vA6Ni1ItFgFdYsWZY2hNjC
qz2AqrWRYWLQqr1bpPlmoL1xoZNnhnZLje7WDIi8HARPEtkVZW61K033rsJRaZBh
mBD8C4r7cewjctLl33GhV9loi6w9WgwthygTH8pEQ4xIDUaX1NY2JfLIffadugu1
Dyx0G4FzfKLXX5MKyITM7xN8/SoJ6qpJfaUQ2+Tak7R1EXlWok9Ar0rBQb8Dfm/C
RiTEftku8EUdvrf30TiVlQol4zSumbIHi77vaYnoqhqnGxERtHnU9uamUEXh085Z
/qnY7yz5H+r7xsHoYhajWA7XZCaksdpmDDnkGST70TCjt32YC0eHZomKpX9TISEL
Dq7F4WDNmH0vJPJZILH65SfPwbqzR45INvgdz1FR4quycg3bHgeuIrsz3AfZ8T+G
AhEATCqIe/ABL77HoMae/khrNwdn74VuI9nswTc3LPwaPRwbDL5u7hGr2Jhrnydx
Kx32cuJVrM8NZasTYL5xRZGWJXCe//we3HCCTmev40bQEk18vMHjx94wCleL5Y1r
XNqS1FQ+5w4maTQ9iObkGuEWfvY6GRO4q9LcgL9c+R9MZZVmOvSihAlyEPQe4/uC
m4zPICFuNFAdYrBdE2u6+LO4ofsx0Xu5qsc1Zz+hbN88ZRJF4DTUz4n6TXjiiCRC
UQQPYNI2gq1xfB9haruhR7MCbe8AZRvCdQl5gDdfC2sy5FrPJ3RLIOUSL/X0ENM3
co+Gw62oyLnzG1a8Al0bbxEViQ15MQh/8LVYU6VfcUBwgY3izMtrhXxkqdV2Mm/Q
h3UNOGIMiY5PoyE4MB50w8TvI+v6QyaKT0V0KIAK0dyLLJcpCR+X2FQp1r14ZrMC
Csa+O8JurL7Dez1eoHzMYx6NtRSriFY0UNpPFAPZe8c+444XQNYjvewEHFbEHg9j
+aWp9Ws/9XpxTEEBnRz+e2e8SVlGSWj3qB2zMg3PbdD7UVk/lbNSDu+CL7lG3NVT
vgH8DYCBrNeo3fKo4ow3peWM5FB0Z105QL1qxKGPdgnQqv3NT5C2G8YJNHppadga
AuGSK4rEm8lmMph8KN7GKfVDArYyzezGc1ANWMvbSCSy5RjKW7ZPdLeR9c72ZIUv
DP+awp8FD6bAIxtr0ichrAtl/U1q5+Dqr5SZEgiDbOYhDdtSFCD1bL5sg3qsPuSX
sQMRq1jQIMeH6WenFD9hO3ahkcRg78n7DJEBIDx059wlE5/33ygxK4Q14Tg5IWxh
UICANA8HJsasgxjVYwE6J8d6zQhLrlbFg8+7zcpjYl+m+8kmWyrDW5G644rm6npp
b3idGKsFPARMIo2Wj/P9RO0fzL5RWB3JlrjsjUHgha+woUSsqcHVXZSkk+KahO2/
Mls3gO/APm1B7kWopnB5n/Y0Ppv+5uJo21jP87pJlFDkj3XVub2FwMEkM46wTuQi
NsQrFpHeOOk7EWrWTB+rlCaQxSczlzpXwJN8B+fw7vQBiq/J0ZEv2K9z+6UO7yew
HAsMTTicCKmQ1wrl0irkN4SGyxUjlne5Hkq3AwnslKg/7F75dxPJnWoLQUk0NB45
VbeioXVsCcjX3bmZa1ZfUoJCaZeFtfnWvh3/2MLtkZAEKPGBeH02J1uGqwncnvkv
R7BtkNQ0A3EdBuQjITdTIltvmO0rZ6plfqiiz39w05gi6GseNKj3SmTsTyfd3HEb
cdUeg8ADo67eQ4yLEsNYcCGCYfJVadXxsx7hZ+p5rASl3pMKqakIqhMk4zUqwtvF
2560ASZViwpiKwy/dChf6d9S41kRk9U6yI2Lrj8Y6GAkIATQqBCyB+xR/s4tqrtk
K+4Y+qT52BMz2LiZ2OkLyk7ob6x58luHgxHObIo1msa8rjDF3PIXZjRchlYQ3/hq
UDEMJKwh8KT2cXwfIv9rAv6/xoy5K/RhceDTOXGYJzcl2MV4TpYiOKw7uDFYIZSM
Shv2k75g2WeatCIRGhTeTlCNL2v515zgfzCZy+iWuOOOlgO7U41KHWT/rYhQIsZJ
Mh76/w4t6eWAEEaAJD85BksirH1qvkIfimp+xQnPFmuk72bDFXmOHoSuzSchTbnz
cKHj6W4bjaTG7BBrXqdLpg+Z0iWdK2xWgn/lAHwYxXN4jJH8QBBzndnY6S+jNCrV
sHtWdRcFqXSr6AO/97YXsGb4l1fB+W+UpE78UX/fuKNPWdjg6qVi8xP2XW9EPlKE
KXUDlY/ljpR3Vyr5qG4mjfNKCYHFZi+nxir6PYmHQTsPIc+SB6htnLELlimWR/4w
TYMrhwRHdAj8brRXtYzF8UDVziFK4UBVGAASCB84G5agtNLjrv5mNwID+P0Q1byT
WUNsNgy74UUZUSGzFE8wV0C1IkRC1+PYVz7LKbkATTSiAgV/hMG/Hy5iq5aSXJBo
mrpezX/Wk9AuHYgYjI+N3S6iGSSky9LJHS7npGlHJA6qIu7+RkWviqqniq6KySeU
S2Ny6/QRn8tGj7OpYRvDouZVwlPT3l+pF5f9QWv/McB1vZo+n7h6o+ClS14fx4KC
sr0SxsW3Ovw7vLBGlIdCe7V36uatS/aX3IbE066xD6VQTbIvD2XdlihXWIVuOzPT
8RK4Hu+noa1SDcIaonOn3IoEbWyO/XKOX/Mvg1NKOl2XEHP7G0yIMSp3ni3Fsl6h
ukdZ5ARCUWbwH5lKu5HrbYQ4Hgl0etVfYuIzBlHXVkZNeZzaoxVE8pw2ULVEW3JX
3yp2rdCkaX/eZ6WLUFyEN3woUW3/TXZOHJ7u8WxqZK7V6I+43b7CFgYM/oskF150
wbg9n6tYe9ZWswoQPKAZ76Rsyog1LJKduEINt7wXAFV6Vf00I37ubcBzjZfGGHtw
WMr+odtzNHfgVNuhgCBfAqcuc+ZFQ9HCQ+ZrGXZeSQcRnAcJ/SfRHxLcG21BHu1l
Wj3fFCYVBHK3Bplw0uexb4cyyv524wnc7OfyHfD231y9MWLzjb75a3E50ol3ruBf
Nv88wKdEXurzrg1enRKAvIkYu0MfJmdJd61qnne8ZBEKQWbj3bEu8x2Dd+gCkqYw
xuWjQbmvHRtZS0pRjL+wOR7rVqLhq/7AZyfo7oI59tVswF3VILUaWUTI2qL3l/i9
l06W7ycltvMTFIngTVyjKdEgv1CgkvXG6/OU1nVc0Q7bWYRNyiPxYb166S7sNxbc
X63xVcnqFFAu8eLJiIC78Kfquk94B7eLKzgbmkya8mU=
`pragma protect end_protected
