`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QV9cbzIQYZbTtMTcQdXe/eqoGp8+O5oi6sRg9Y7ckly6skaVLdR32P0bVYdPyNSh
XtlWJTR2058VPGad2fEjMIdA/NhnGwU8m3948Kom8D+CaaixSKl5dSfotVQFrUwD
kE49uIMmN9dVbLy/We/q24mXC1IPfDoZI+IIouXu9m0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3584)
GRx4A9U845MI3ztOV2iJ7/7snNW+24lUBtju/Epk9uGhbfcVBk1J5zjmAC649pgC
W2HX34BEPrypbME+ceC5yVA2266cQUQapt7fotAM+34EuQlwrfWA4jQB6A01ejGs
UMuDDRddATAfKYC2sKh5jfWAwU1moossKyoMWmNXMHYTfk60qt6UqWbdI9/qYlwt
DlRAu4Tw/VPHG/BnIPKZA5q2ZZhz1plwws2XarRj42OKJ7lMSQpuqqh4P4PyrNuZ
0YZ9/JjggfyoweuYcEPsMxPvP3aIkbp2fdp5vy/dQ/laeJjbrZHUX5L7z3zD/GxK
9gpoF2zJtd4KMy9aAtJsZtCDCVpKoNTcPAgqg8fWm3IukGF9MaUSI5D0m9qnlL6X
vRJOYUTu5XCTYO0J0M0Y4f+ji9GUdc5I2Wnfl2GX3VRnemceZe0w7fZrvCx4FfnC
qR5AF2AK3YRLPX1R6IxDYzutoD4tNvbTs8Whc507XViPtPeztZ0pkGRv/ujH59Pv
1TdPILRmWiw2XlI+HIua8l4xYDK3/H/nSgeyTu2wLczuW0PjacTcFRBMujXEzzZy
XA1CqotGprYAOS3iT4ZUvieKMAZQLCyl1DZRS3o0kKiVYj5+5N2+zowV+cvITA/l
vKC95OnGzru3SddiUmW64F5lNE8lODH0GvoSYMH/fXohZ1FBrw7yWbpZ2vrYpwf8
ZXK3onL+B/9JpsFtGTJNBDVTdulAoXZJ6NOcwjnA7lCNhE+R+NZGjAzWXBaECtQb
8M3MyiRJbhqYNPIysYc7rfEe5mNrz2rwLr8lC7ir4Y8wbS6sYG4aW5HRYlqst8LK
2lMubYcgyel15tQ2AVB38Vo5ek8tjL8rynxeUidMcAN3oeaI1dC5ls4k0LmuGST+
QtPrjsqoHlZUQvST+3hQpJ1GWoZcVLYjbTDwhMGs0zfBNSWW0gTbkHsmTYQ9BqqO
ITs2EseSRKszrwxe5/yV/MXzTvhfvu2B4Guw4bb6pliqTHMVyoj3XOM3K6nKvOy9
GncyoRXw2LhGC1CtWosAcauLcFpLuHzCaJ3IyeEx7iJ8EucDOVSi6hjMw7Kg18E6
X4CF0Az6U1FXztscFz2aR3NK4y5xQEoupxPKoprysg3fhre9UzXi8xqpsO+0wy1e
pjOrxOwoEU5eWvFza6kDAMCtbL6xDSk4SpX2lmK+YLhVUHV8oZy9TiNff2AUOQwM
4fDcQERDQHU9DkqbNKe0TU+Os8RM2b+f2FjUQM3vX7hije3g6IZtjIKw+7efMxZr
6FGeIzAo4Kr1BcjIta1uvTxUokjdrWLSPY3AurVuTvAgi97uvqYgLVK3AU7dqC8I
hrRZ4Fnh7VgGhoO2t4nHR6VxpEkjVu19BbTgKagsw+oQdm5OYWAMOhgkdU3oEVTp
wVCRFYPQ1pmRisjK4RpQl1p7EGO8tVwKeAsZHSvXVvyqeIK+hq5++R9BX1jqrTJz
n+rJXj0e6n4NQtHIZOMxk6ejL4SiNyDzJdcs4MX0aA/S2zwFLng03IKOmkv/wTYr
Oy+pF6d2Dq7VqAJt9aJNdo8WgQvFGOU09X0UlOnD6Nj9V9/K8VXcIt73fOGrOho8
Lza1hr6SWz2paQmRFFxYaGNPoBaF1W0/uwdZtAWpuKWF3OubeEaKJ5m0cql4hGg3
52AnYFc48V3hQFfCxVXlo/KNAgmJ2jDetutMRsGrWUYQZjh87+PGEto+ga5FjFEx
y6pfcG+YxaRzsGFSDNmBlApEz7ZfWXht0stFBBZ5TV3hQ3t/89LObuRHmjbYlO/T
q8P3JJvI7hqkumbDjUXwMGEgtKblJM3dZp/QmIFJuzN0KOvzeh9B/hr4ftNNmkp9
OL+gaq3gQfhiHpgu5nV/FGh3TV0U/RGqO9A44trDaLsXWQ5BknsGZqQj6u5ekiRL
eXtGfAdv78Ao5MHnsGKhEjQXqyoiizudLqNl9u7R3CzxKoG3Qk5FYrrqymWJvTTR
qlueHpCQpJtL1hJR6NydOgKH/+Qq3lDIYSojdQ20kH3eOBWwE7RZ9MwlwMhxIt0W
/4soSfqWAdz/898feqjlHV9ObuBLuWa2TARh7J2NlU9izTqB5mHogUWBgaKeTsTH
8tqwkwrUxgAxtGgXPkGjYagQgET07IBnRXveGn+nubwHhZb9aDUCPBYIKEcqLPDk
HGMfZzMfo/mYfS4EPMxhX1ZwCKTN3Mt22G54CqLtlSDUP9x61BEv4tj7dYnWDXVi
dQzj+b2CvVo6gt2+BDeGjCtciDvH+I9oS1QviNFxC7mrPivGYtwxkAwbn+hhwcqm
hxpsBJ9fk8gtI+kZcWJIGMRd1EwBjE/L/7apTZcfWQGEqNf9h9/PlLCZ7+2GCmH2
wbh6PoSYuRA3ROQH44pKkk1X3X2cbEypHQYTsBVCzsr0CvAk8Snw4fRXUy3gakJz
GqCuk+T+9gn8wf5BgWunc6ukLg4msLy3lhWzYLlhf9uTBKTZM2RgLgCrUWEwdXWf
nKetIPll9boEhAMNokDtknvRWg046dSdpdVk285zZ19bSBynlgaf6oerVRWdOI1Z
9a64ZCWuWT6CiBRy9MFl9WkTV29kU3aRoslVQYBJkMZ5QZ9ap1zX7xMqUslzoHQi
Y3IAAM4mKdtfiyHMFBLshlRhcvCoda8WoSLuaD9M2T9TBmy5nfyuO4M8RPYlHmai
h7JR0fFBq+eVmUuh+1cBKZyW22J5rtmo/lmANnwCRnRw+z33p7k31AyR2d/I9mCh
jDP8q9z7f64Ab48wOIJrjxS5BZgjuyBdQ+LZJzvskkV4l4+j4ghtWYI3Kqs/PW5Y
ms3AGy6JPV/XgiHKvtK7vfqUyUO/MjABF2484d22RcXPlQ8eh6/NtFBKIO69o8+d
sFYrW6gn4gmT2RPAKYqzGfBekCw8uGrkZQy+p3h+dcOEklFl/1z06l6RbS2XdTWe
bfYC8cRRMyErl1OL7Q1CP8NVzFyHHx8+BP0pfZ590H11in8OP3zoaVhbly9q6ilf
qMkfCBlgAcVpghXGxkiFh6OG7FUuqB4GhWHAwFZkvjEbh9Vn7k1slwBLUNMKJW7Z
sC2Of6YqPOPTT+9tWeAkVePevetn9UtXaKZ2ij/mMMCuCmJ/VKq4V8n6yuUSJIVg
CGXGgk+t6MQAbBwRL9br77ogPyr5thalQnn/9Vc5XO9gaUzjv3DLldNbIZ0IjZPY
9Cn4gN7+MlTcI/6YwzDfAQHZ7NVm8VJe8OV+HQv6H0mTOJfvhxiljlj56dTQMUgT
cLOVHm1r4u5rfKboSDjGJ0W9dcGBPTXnf6RrDEe5rDtjHFZmLaxSBOh6JGk9FDI0
+sNgeHF4q59yp+HoIXINq+l8K+Af2mNe0WlR16d7Urf5zdFpSJ0NClaZDeNQDZ3H
QlaQrGBVyUm7SAnn1iwa7uRcQdzVPftwBP6Jt7bwXKTJGvfZvmE67qFmcN9EGX6z
JmvHshL1kKk9dSjzpJLEAg4Vw6+0jc6gcBRYZJWX3Mi1LUgq6b/xvNmZslHbfdx/
r55iWDtQKkSMNs5l3yEPjFGtL/HLBIEO3oS2ihM04kpB2OKVRYpWTvw52SiI70m2
oJ8dt13GM0yXIHDi3OBKFOvsuQZgqlHTnFE/++OtqQT8DIqP931t12UngRX8bQ4w
7P//w7bVV+H3Vgl5yMz1yVO+Tgyf2+c9z4A20F8v7IQEA60xUkrYQ+kByeabVX+8
0ODpTBKoIbfHLUFAsoZ8/qRsUGdD9qx1xUQoYdw8cDEPGGDqEYzVPcDtbmf5PAAb
D+vO9HyPiUOyR+pUFkUlBar1wkN9sdZLrZVtTc5aeXHGF2z1yOSIAWUv0CdpENDW
jOev7AhHQSJGeI9AU1A9F7X1G6N4qL0lBIw8LXuRbcC2kPI/NQZQpb5r3/jDDvpn
RSPMAqz6C8NfNRveEAfU3uD1mkfJtLcluWag3+TP7izQVaubnKYj2kGuFHjRl20b
PkAhqrfe3gTNlKHM9PtqvRsrme4a3PcTAFgs+PSLgm9xraqBRCb0tps+YB0rtREu
uAnyE5MepVxqqWWQmBrkk5G5KcGKsOhL2zaiD3H4If3ruld3Id56oYO0/LpHWs9e
IRJT1klpmdFXx8hMVQCIjZgu5RjvleXxuemj48kMIFE/KoK0PajLrMucaS4uwI6d
/thvXxdQ1dMUcwpXJ5kTWMd3Gyv8iWZ2mS+IZIsspl5BUuVatel/DxDzpliJj+Fq
aX0GtA8FgNinwHRsYitvBQ+pgvgaCX/l7j00emj2KYO1yiJVFx4m/uDjuiSwGrEt
oIX+I4Ihuhso14fABsWQhA30xvRTtoskub7XUhCUFz48oKwsL8l2v3/bi60RSF7r
A4BvvM3Wy3YigAME1fId4N+twr63u2gh0Y/sa9RTqqqPfbmS+HEDp9tcxikoPmPv
6jcuwcj8Y5m5mtVng6bsKiE/U58NfSfzBzVYLlna1ivJltEXDpsP3S05BYGP5DxY
ZpKHrxI4CMC2zgScxboS/y13dTOdBnUzRTj4oOsyFtd8lj2+bB4pYkzpX31SF3tx
j/Q+Bw2lT4d02gGrr729kcod5r+gN7zwyF+sACm/kEltegP6ibzUD3e7AcLeG8LX
AaKLuOMnzDuVlw/tzgo/xPzIpZthdGfcHVfy/z6GADhkSe4VBIA5CMiRKIPgQ1A0
TU3FnZt5qknYQtQPufO46wuetTEzZpqvyDiTNj7C71ol+DDO5U3e3J9NnkPnU9s1
w10irrgZ51qUjUBaSRSvfEoGII95RQ0kRiBO4cPpl8w=
`pragma protect end_protected
