// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
lrmsx0ZXMMc83w0fsXcXNu7ntk/CrWo1SVdnqztBsV6/MhZoU8W7dcUBt22SG3I2FWzAhyhy1HbR
Cz6G8wPxjB9R/uD00n23FSOsQkkBikz/r3qlftz4lCZ7+hrztEqs+e7w2ekxZbdXJQa3pU5Ps2YE
xNCYvIXw5HOZ3Uj8jqpceEK/r1RzB6Ffels1SaK0owxw9wMtvIqDZdKeegp6kFMZ8aeaptLpPLhq
l5O6Q+nwrMwqTgw3wjWD7+hTz0dEiFk+V4Tnwm2czlZe1Iukc5wkBUFGL/ohTO6N194OAhV6Kymx
m59oTNumoM+IKR7xOUbOARJ/eefuv1oRdSChIw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5264)
ztTZ+s2S7waDGcKoDojM/JMV33IiG5sWV1E5tgSyXofuJENNv67IGj6TK/R1Qz2yH+O2leU+3OIp
pzPwlSe0/HQrSrnkA7p7THxLy4KB8zgIXZd/UI9LxUPDiMe2xG75wIR1Tsxp2A6qFC/bF8GQc4oy
vAVYXY7BJfgaohLeLl7Mu8ldPXlgkm9CCX/69yasNmYPnCgX0FKy0EU9qLkhSFbZ7XWYyXlELNYy
HClGGi1WONl9hhyGZUx4EXjVvFDowgIa0cYsOXD4lMQ/pRZyBolQFK455yy7X+CiHNAc0Ql5qfx7
oSustiKbBT8rokbKKrKRzLn1ckBF88UtAHIEkf1mX7q/hKSqkN28c9OSYdhwaLjfTp34piYd9RrA
zjtu0vCN5mG5qsXe5wH0LGw/9Y6guwmapGOV7OISxLei3dpYfZdGFKXinrMUxCBVhk2A/8VcXcrn
ANe5DQ4fGQ5t/slUdwrJ2/PP16J7CwPPk0TAgcxpy19HEo8KizQofxvomXRC2iSWcL4djYpi+7CV
9sj+plmL8IanNOsaNv2XtdT9KoFin4rIDLitsENY7cpqWMZLaS/Qz4P+12E1Jz++DxJnft8L2kYI
5D/14qZe4czvtYBfu5FuJIHCltzuDUdnUzC+WJ8eU6YaUOpXTTJlJUOGPDFylRVVbyAHRS+b8964
/JYVWgIAmpqI0FO+0LUuIuyl1wV6UrGC5noag18M2bwHAaC+yjhPxtr9UKP4y2r8VVjbUz7Utnme
pVjdJeYxp5oYh/5ebmTJU4GAFZljbWT7qpTG/zPDQyH+mgSm+jhtskhskpNdur3UtBN3VH/sA7fX
xMkhcQaGZWmjGJ7bZIKi0r4mFjfwcMNLP5FPFInqQC+NT62vJ3Xd91zJKnx8EbUuSeUNUG6Dz75D
URrj7mh+ZwiWW22BNgGYBTU6HbYso8pCeK5dktmGUaAm323vdktBuxZ4RJ4u1UH0a5o0EriaZwft
W16TmLbhrugsT/sKv9b0UpTrJqXVKAvC6/HDwnHuWSEr8zJjXQtzsAS7fzCspLLk4M2rNsCFblCF
XhCG2Ckv2j+dHn3GLRCR6fdp2Ck/1Vx2VTkEAbQpL4VpDlnP7OIX6pqBQ7l9XSJMwa2mU9SiBd/D
nru5ZYvQhUzc19xye6sW2k5CmUEebiA+E8CxIAR7hiDT2CvNrNRWjlt7kmCSjGilvS/054RZnuM3
OgCS459NlIHPIa61a1NWoEZ5xjlDGqJQTE9s5/KdkrChMgXpDjWyum9YUhHqyOOA4N9z6ZiwmT1V
rKdXUlL+vLGWpUL0A+RnrXGPN+gjmcl5vmpZDh6vmnVg6faD4JZSBQmTAK1j41Ced0SrX4+2NtG5
RAPS+KbOP1SawMPp/+yonmIwJht1BTQQRaJ2LfIi8Do+Z20MGI5XRWtBspgIZTqnXzNjpIRn354q
TBVSPzJreGN7G8Kvr9PHji2xM0VIcn+l9KuHMkwQ5By4Jfsg0s6YYOCHUfjsnyaS/AoFBkEC6KGU
u6Ce6zdxJO8L9sBfEjz/92pzUV7Rq50ZEnm1T4wgROpYoDdLX56cy63VznEcSnhzj9Deq0nw1vBP
fOJbb1wOYVOpq6088Zii2TMP1l22Ioo+1Lw9dYriBGh0g2fIAkEKT58WX/MqcUpmM+tqg58aE38l
ULzxPM3IMs3p/qA+eA14WNPy61zkQmUQlXu7SLdou7nrfjydrr9GwR2nZcwIUtKatOzRNV4nviif
CTKG1BnjWkdVm8URM1kmyWhLVfLwL3roC0wkB3nwc3ybssPtraQW6FhdKhymbD0G6+Yb+zgRNjQl
LtplZ2dJH8eZtLwzOFx0vnD8Md+RF57Plc1wzuiBF4R5hl7srT7bP5UwwtC+7ZvlShQs8jFwLCim
CjK0jW4sEqMx69Qzn+gwzE43HuQCke68Fo16bYTSjE/54ERvwnjwVA+Hd/SLRtRUb0gfmeKtgdDt
rLyYE1qKko8jWJCpqQVwHbbDeDGPbMmWmOLfdEBOVXbWjHmuDEUVx+SoYZfIr+Coo5EnAq9r1Qwm
qSEYmzINsoUk1wgI3md1/wchEOhi4e8WoiMiVagP6oKJGUBu7AViX/lgIBDBrnx0/zYAM6IszxSC
z3WVGDExMlJShbJmKJ/GcoB++fxsW6wgCVY7lz5paJGuXfe3VZ2oWSsKFZ9vpX6RD3hEJQIDWb/n
xXp4BxHadwysaivMRNhXzmbjTBqrdzx/lRuu8DfF7PjhpZLhzUTDZ0kglfrDUFi7YkYy5mZOL4bp
+w1yAxw72SmTqea04ViNyWbLmxh6CIB/vM93OrLdkhRsq1HCxjuOf4cDQuee3qWAWOTbiwIlTe7f
AN/437UUlryoEjpLLprLrXziHNI7EpTE1CVyt9DwahUdSW7nBsmTysDW4HrolTI0Y/nhVicEmMHf
RrBOVj7ph+o7DIJxpzMk5aoef4UCcKNnbCjB5203eZrPOlZ/9PRF+5M1e9qeurlH6SnBPbbe5l7+
KbwLOSpeebfBEc7+nyPMjicQ0GvKVRyCfwgn5RZ9cscDbrLxQIcVuTu5VUBgsyYEmEIXNScP5yQQ
ZvsPBJM+tmik0smHqGqr6MHWzeVYWTEd0XUlNl8y2/93DhiNdNy8n6HBiE/kQnS3ALXqqENI5Z2i
KQNArPzB0N0m049QvATqGcRGUyTTp/2MQ8OSAdYiqnUTCKWHx+xjOpWqu33xdvuQpDLEZxPXoPzE
Wo1EiNFxz2HI8UA8tauepEeVWbSpyzhjEfoNquInk5uQMOSjoJVszLHHZ4qTE6L7rS9uuIL+YbQU
IMgYtGn5ykluC73K4yEOg/4EPlINJiZ/CUWYrFtXC1DcxAn8kxK5IRuCno4XEVxx3CV3q1O/boZo
pNEO86KZy/L1C85k1uyRa8Mw9kMq3MOANA5OtvjUrz4VXMcWnfv/rRHqKbMxx6VuV1GEcE45Mv8G
GstQQ1GU2CxQ1KRrfOJ04odSJl0qHA25Ki8h9lFbyy4LPiDx76VZo3ceRtmUHbEC2JqY5qlDgDnr
vf1AILkK8NJTOhFx7egjV71UvCBL5G0f5TDrH+fAithdf+OgNNgbLMCMYlh7sWthRPHZHFuObNXE
L/TuHLY+Rw8+j1WMcpzOk8yoWWZbaETJOj/wEsHLFW54m8FWvM+Jo1PCG+0Ntrk50F3XOw2CoxSd
qNIS2Za3jBrHGNXbKNd0nO5cKXeayonZwJ+ceioOE1Xhf2hKmTztqxIq1N91qMzb7u1EbRijEaEY
CepjXZt4uDK8ZLqr8BJML4DJYU81QmPlDOqGwSVbTLXIeuUXOa+O2D1+/OUvcFMFX7RPNNr6Q3yR
AcNP0e6wG7tC7CxBustfdx55qA1DgpSKvk/hOYTYlT4QstE+HsrkcYUdH9aiz/DP/OlmhVIedJFA
OAxzloWzN83Z5Gyo7kk0hdaFVwrYLkE/nVB7htGJEsE+Fkb+pNX9V3vIpn4LpHuWiEnX7dP+i4Ts
Lh/luN56P1J9VDAUuBmylg4cV5ReOfqkW78Oh0bWaxPlyGPp+Hd2sO2GJJwSeHP0KYow7lFZ5HNi
XZSpDL/GzS60WmCXPV7/k5HNmUvFqOHBDGC5FREeXIINAqG6bgBpG6l00srWJEY1fON97RerAPJj
J41/smeQKeqW14g8SKmDprceq87ICzeA9Gzda3Q1Z6RiYFDx3Eu1rNKi2id5qXocHMcFRxYcXwo4
fL2VpxT+FQCAlXP4Jk0fn2IzdT+vkMCjzLaNS27hlW4rd71KOrz20fHuFByZ7fZegh5BHErwuGgY
+usROzvyuaaX9h9+2DoKisjSdI0eY12GdnR1Uj4gadjMo5TMgHCN+mvOTdUcYnisDr9qeB30YxGT
ti4pM1Z9UpFSBR4GAA5pIgr9EvtViYliB8C1Qlybdwqw1cfvZeYDmfZwUJeednSpxKQqKA42mY+2
HKYP0ERbVdZr+yyQMdf2jjFRsK9m2nSArGZ+95oLSRdH7QFiWQ5yUZwybLLhsVcIgWeU83gwUD9L
j5g7PXjquPj2UoxiHGvBeMjQxmWw5xuem8ZDrfW043m2jKI+R/PgqPrEhxonsb+ynJMlSagTImvd
zRyf4PrRcpgpzrpGjNQEMH4nSq8IHsTusH8CpVgCy4gpZa5GhOdALfnwYP3xpEUVbF0C7dG2/1WB
/S/THN65uXCk/JRK75tVvLU/lhkihnhy6xoa0ycSEwPOE13fZwjNNic0042C1U7x1ErQg+ySjgSX
QihBz3Z1HO1vBxnFdw8unfSFfGuY8MchIKp8A6d+NHRu12TczvBs9la/lKXe6ZNXPaTZEUYUsbgH
JABy+aX59QrsHeCev5FqdGsBcMMQ5FHLBiuoSanlSdp5Z1fAVDOUbYbG89Ub8g1ek++nwdlNv1gX
BhYwBhzID3OKw2erltvmJZN+KOPFzK35UeKBx1iruYrzYFoDTNuMllXX8fDguNaSP4Uc3TBbnB3h
i20Rutg1hXlR6/jWfVkJhWRZX7PylSYGPJnt9CrSTaT55UTVAxOmSZhBL2jo2YKDzQiSTIbytO2L
NeS5kjwdSNFt0xPAlTOmuFNIuipEqkjTJ6uhDyPqM659JTmtU35ZWNMu7WFUESHRwKkxwPV+FSyf
Rd2f2dRFGICZDMec0GjQl5r/v80OK+iNhmEWz44tn8GjGUNdeibGzkZzF/02jzXpQKS0SxpkWg35
uCl2oPoq8ykppQx5Ghq+GpJBeTHcBjHQ+PJVDGNw8zrS6xdFo2WU1h//RCPLNuOhdMDQ8WeK/hBQ
ntkEsbUES1d679UfyabXGfYve4TSBgUfb/2gm+oqpd7qZRTJXdfzKqNK10gdM+0TvEOUUK+3VkUV
Kyvw6ZlKc9g5a4XDKyYFxX4evsYqJ5LNlF5YkTMvkqikGKNQKNGsmPocs3jDD3g88X14L0jMTqFn
mgkguRYhCGn5E01hjgkhF0T45idRWeORicV516GqtWTw2VeOY3ugbOC80pJ+xo9HKAx/twIUlwSu
+XevwUIYxWpuG0ruDarkf1RBbmqvbe+Xv1FMd9usI3BF5/0iEjN6yE8Orh198IOjbbzBgxa3sSmv
20i2O9fWhS2xKbGvi8Qzhz/6ikVGYTHDdqSpBG3YdyJUsXA5mARI15g1ae6GPEWo19WUAfxgCEvx
aPYufB5FqcTJuC/DDOuwfSOsM0cxz9AOFpGMarboL2K18436yeFCGUV1QyCMQ9lqvRCFrvW01yfa
femQER9s7p86BisGtjjp1GpGiL4Pbfz9X5tLSGwyWVZHjDOkvYfT4UAmOrgKeGUG5u33+J99F4WZ
jtNGN+B1ODggBZXBPloBt6pqUSj+bzl1I7pS35vQgNI8gVS3+qnj3CLUywF6p01J6HuMvyD2zZTp
jilfnPoj21UskJTf3zpyeMSP1nWP3xxio8xbVcLWAvB7YxAygDie0FfoPI9pLxt/Q3Xn+rhfDwlR
xXqNWP0k+PeWU2f6Ur0lCiQlE2LUfLvUWnNXeC6E71VLYMrEtH3B8vmdiohDcNGmALmh01WniDpF
vU59NWwwchOmO5RJDiWIbI3qzbP4TBISqf6neNmXSfKXo34LLDEtgvLpLtxKKPf1PXr533Npeij4
t9rbFAtYHsjfVXLJzFmJb4YpUQqKZtxabzpyr25z0vmmFvw7Yms5bckn4wDC6YKAYcQQVyECAzew
RDvpzRXzKQ63BBdQbCZbcFeV994nmV75NeDFYCjKnfkzoXZs/JMvvxxg6TLOKPpPlkf+SuPWUr6K
/DXTdhMp2ogL/ydXN1IKTkkjVukI+ibqbLqirKV6tEk4yIPHvxdOT90Fu0pHyW9Axo5EWPeBFnff
6vPE+ShOXMa7frbvXDqWjB3YiBndurTnuytfgDopYg7XAE2JjvareOuXLzQhu4CEL5s6T9s6p+mt
g3lqXqljDhL0yUahbVBxtYZoUw3LoUqacNAtJPc2tJjfEwDgXuKTekkDhuxAqmyLyLDt2URjRxO4
5rK/bqcp1+6P+vphvnfS4wK/C3ps6SheqTXyMJ7J+TuG5FeIFnsVAZTy+cNKU6XwZviaEiDQgvdE
jivTQcl816BOSPI9q2A+l9xFxEDoweKfdwvemoPhGKNAO84wSOdokteavwgwXwbNahHJkfZgCD5A
73qjFwOQVWFw8WSBgiqWdcUPWZNIzsfJ0Jp2QAu05nSWkqGoX7TX6mZXEXMqmlO/CGKoyLZHi0Ew
VjYUHxiW3n6tHuYmtwy+atYCRTPyxkX4lU+x+ZZieVlzxDKPiqEt22VvexlWSVlJ592txykK/zh2
Ak7ulTxBL2IVb3jwA0dgJJ9C6ntCkeFpxn2NR0NIfXayMss4kCo8oHrDBl7SGsGxjenl+LqXr7oH
XYYTpTno/ysR2I/j9NFyI4rCCwMPKJT+6FblYdM/hwMHtQR8OmRsgPbR7AVkOREqRQZrH651w3Ec
UuYWk2VJRosAwY4lbiQOXjGlhkmZNPH1AwaNtgDXL7j68JGEaBYJxHxNtoF3OSy4hfZKevxGupgK
cZAU6GY5NqkzNrZLB/P59r/khjFZGL6D4l/PWQwfIEwnJ4Ltw3t+ESDFMRgqiAFnTsO61jcmD3IX
gI6InUe0wFtTZzvOgD0hITbLIfofn6ST3DqmdwzGmrdAxPPRZt6dM5n6Os1b5vrx8/29OeoiKLOG
5rOQdPJL4YrUKhnUO2vPvJtbhy2dSMu2EjKo24kwEvFVWw/1fplQq4jjSd0cyix+0kjLhWEkPbUJ
A4WebP4NJy/qHCdGxp6NnUuxzUv0FFbjvesytrbTg+qS/TaPs/2AkpQHSIDw72ZvkTYx/pYX0vNk
Ws8YyNgK9Yvuv8p3QwnmYifjGS29LJxnT6pFkaMmiZIQoU/5j4AlpgCCYytXRSQKS3eJg0BOrM4x
/2ejqlAWtwW9EKGE3SwirVavQjnmmpWnkxB0VHyl7IBP9Qy+uJqqa2+FuphQ2ofdIg9FSQCT4BMz
wSTxZ0u5v2pUh+J2/aMlTVTXfaM=
`pragma protect end_protected
