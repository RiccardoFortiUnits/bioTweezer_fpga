`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Tl4O7owCe27SjiaulSeF9/wp81UNoRqPu4Sq6rLDkN005083GRaW50nW5yUC2mYI
mqekE9FDJil7gpmMu6YOFUhZTS+zLRvoF4cSmleNYBxHy75rReVx/gyMTF2iirVk
VMb6vFz2jY4z8kp6RgtA92aZCdnw8jGduaAVCm6tSXU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8144)
Rlb6sWZ8+4nmHdGjETBzkwECvvRd3+pLeE/v+XWnRi7yUMjbk7pMJsMiyXrT09J1
wiIyPTzSN6VX43q9cZi96jyaS9YYBfNzSsBtbUu3J047yitDRCg0SG/PlPG8KY07
Wt3NQQ3Xmg7fVLBtWgw24nFZugPDOORvTFq7nol0e6pd9oBTLKLgauHb4QioGs6F
/gS7+hWCZbLvqaPUhOJj9ux1qsS/xSe0shRjBKb6StYFJx+W1n2Qh7tMas2Owc0H
m8tfRxMtmtO14YCLBIz76DtdEPv/J2JM7v3cF1D03O8I/rVANRJpZxPiWdn77PLf
LmFxuNZku4LguiGjZnN2VpPRYtcWkOHCvVhIL66L+bYDexcXkfKcdjP44m8f4Y2H
nIg/ZmwwiQWaNs4W8KgQugqrpBFMg8KqbES7mcyiC6I5FTgAyM+neAAPga4QqMDo
fM7F06oSHiJ7+My9VoVfpEjiSse/FpL/OA4gD00L8o/XHS9J1qC92xCYGliz6L5V
npwqYAKeYtkZZ4R7kU8m16pL+3snGfc+9u6JqxlLU0di7O8IrRd3OkqJWnsVdiGE
he229lJoomcVJmWreN9KGfi3p+N81XO0mj5RdguUNqStmbelnenYhye/qJq6y8Ol
NDTKI0UEwvFadEyPJ5qDG9FymFM6iD1MSpAYUm4rcD+ugsGMdHcQTDuxiTKJVVjY
hcI/JOnoofNzWohZlqgohozjrO+tZcuEVjh5eHMtNaUB5LQtvMle2gUoBfeqRpke
iYAzvTsySUIh9DBKpmUt40dOoPAllPUUGoFFS3SLIFYYyT+GujhrIaJfvZbEnoeI
IiBguZbJj3XEAg16M8QwglPRoUism5Z6nZ7zQwz9R2upZGRe5nTRlFoMsA6yBez+
3CD6NoUdPk4P1fGP3eSrnLzk+LPocy38E1XZGHk4Dl10PG+oSocAycIJM32XA1Cu
c+bpGgUYqM+2/pz9sTC42OagtBCzuOH4PLXDawGFLVsmXY9bgmZih1jRuwZFH/GP
40GN4y+txUpw+CyjjRTHEYgbX3Nqds4ijBHhZ9ZWp1UnL66MDpWL0dJw/Qz2+X53
aohammKjQsotfT+Ge6hjcCkKSwVorFCgld9fN9f1vuqB+eRUA6Jf9vzXoyrFyhri
V73xWrgsiwyzpyiJrzgLmU454l9J7LA0QJREs+39m9fMr1r3vjAZsc9x499UH2Pc
kJcRmm8/EbiEdWdOD9Gih48nhO6QgeWbVlAsg6NXGaa59LdsQfEksc4FoYO69piH
je39rz9WNMBgfJgA1si/yw/yz/+AYqXsuBC5r5AvBEgljlRp9OeuWv0CflctB6Ey
PuURPnvU4vSxcRn3k7HnbtyMFL0NuSt/35T6/B+OMAFPYjEr+bIssS8iRwSGIU3l
QPW3cfBUhBOR9WyRMvHCjz5y7tTpvCfxFV+IJ5ueKLPY+rHkHvbk2nzNH27nCnYY
xorSyow+xAphfcoLGusbAxD92GOoQ9kRfhBDvUnZwJx73tHp8agUw5GXthQnICcX
nLwNYSK7vMOot2Jv8d+7vxCgjw5IL9LVmpnOZcaZt56rPhLOpruIxK1hqvX1ch05
cCPVF32GYUcwwYjjgsGG18E3Kapy6DWY9jLZwTBr/JfiDCZHkLnSZ42/Fr1hKAGl
zkBSbdeZRag5hajhqK8hzOavApovCHBkV37R6AFIEZ6R9TYnatRRn37X7F2QWZW2
efaRT94nLbih6GnAcpEat7zRwq3SlTjSMgESWvi6R0KQnsV0m5+pjrEoECAyZWDg
2r+KGe5uQZmtaPsS1A9CJCYSom6m95ELWZ/Pj+6n7ladmIGiKP2K5VanK1kKuMR7
JiIVoOXgSoEB7zRhCeeaW7NtJX0YmejSNRT+4hZX8+sro+RiXHV746FMIhisr/vC
9dYXQefi5/9hmT7y6ipQ6MV63YqLVfzHL7cQbuUqMv8hfDd5N5tHwaWCAO3HjdkZ
QDwOzaGRW8JUEi/n5VAPea1GKZdybGcBm5LkXn+/SqCZoi/ZSmgNrgE6zeb+OvXl
UvR9CD2CPkMTIduksfQmLXVP2eoFIgG9dGFsKHctOGAwEspOGUhil+QUQHNViYPY
qHyUCWzAvYC7rO/Kjl1JaL071YfuviVIS+S4uk/+2hZPPtSUzIv+e0l7WmK9OQG0
t0EevzCzdxkWMeLKtPCjDPhRcHhxbuRrhXxkha+oUSk+C7j2D09qNZFTuJWTZ9PX
++v3u1wAUZbAOoi9qu9pfkgGzAvYYWO/jAj9AdU7yUpXq1fC6uwLRfOcjRorU/8B
EAeo/PBm7TiKjnkMZHCbT7OOm+QV7hV24OIInnAkg/ECX+awMNMfnsF4CAYQPdc5
4iQ5IxAta1MNbjPr1ckknkKV9v6+SRQ/mF+tPAVFc7O+/Ws+9rR263AhsdYkXAUu
TozjRBBdFSEebDnpYoVTGnGbKBubw/rehW86F6QK2zCPtleCPr7ALaN/dNl9ssTv
JFM8+znqgRhX9pHj0To6RucznjVhAO2snfm+nqLmofHZHStZcFHsdvIFHb8GhwWm
4ARf2cABLR4Pd1TR4rmtl36QUpYbiVXKFGTRJXpyvXyqQn3CElxszo2BmgW15B/m
xliRggR/KC92Tgw3HYdt1S296w9zH21+J5kjkcuI7vmYE3W1GfSy5L8zvPEtFccb
ZT5Nasy2CY3HW1mnhk5Mlo9iz8x82kIaFkRGphhFzeMka7fEBB/BOxcmElvsEDjG
ElnwpG93EpP5nIYXsoPN002p1HtaNglwQieCKXengYHJPuaPi7cDsO5qOiUKXVki
OYYVbE0jGrsEBRGa7pO/euA5KvsDIgfzHGfk04tuRXqMcMdWshw4UAitpOFDdrqL
Fa2+LVt3WYWL1aWifgTRfeRFfPnLclYZMZmX/RB1GQzdI0uyyg1ADTKE/fyxWBtk
LvLhe3lzIDR85l9+CLpYOjS2I+8Q25rO7eOoJ2IZO5sJlWueE3/NKQJkrp3S0UIf
8ILAaN889aP7slrEwo+sknzs2+FEy9b7YsywHUE6O7XLeXGAuNZv9DkoqxnU1q1Q
0RrOwaxha2g/IbIXrdSwcKB5hUJ5KsLbBkN5QpCxQBpe6XqzJ7ybQSqR8U1CkefR
aeg9oKi1y/vyL3jVdPeA4lVdpa+LvqtBjSlBpygr5eSZhuhjvPWT+27Jsh5JB/tC
uyOcKFto38CAZW328AW2ZEoCKZ2nRtnJFYK6N+l9PzyKvr2U9cx1OuhoEgsucBdr
tKOJ37qJoqaCEi/1hySDn0xQdhmq5AkuupyeX6LKaQL1fTQc1yEAQbfYn413EAAG
SbmzvMUvzo/ORzY5maew5rZZGj+nic5vHwsGAgZoV6bZ8HSdB0xD7CshYnl+31kg
Q1O8na2dbqRxL2ex1em3elUG5cGAr9eucIHAe8tBlb+IXMpxgIsvi64Eckl2maUu
eJ+3y2WH0wnALYbZK0jZFdV6eXSJMdc2FiCI7ltsfJQkJlY/DK+i9/cANzLGqQ04
Huw5tkK6EKir0HrdOYhNKfxaRr8HIeMoASZ82riEcHOZYweabdD0T9DJBOviF2I6
N1+rDARKmXSpl3Diii01F6PVhbxUPND5Volklk7sZg/C5ia/+/+xUfvCNwmpq4Mg
1Mp3g4F5H07G+RE3DLQMHn1yYcJzHKutnUISFdNqEa4cnWW6S7NIArYjuAJCDYdj
v8qEDBvXVBOWE8JZe4b1aB+cuppPqrO5z4J+2R03aE30a/3WUlKE/UxDdmRjCyUE
EvGx0ztN9hXAsJMIeA1Me9brqL1b4P5PZOZamxz8OOvCKNuIHkogWCXKcJvM9Pl9
OhgktpX0MItcwsiYfoPFLYBA5zw/WduvB43ZjkTDN+7Z/N0Czisp/y4Yjx95hvK9
Qr1Y1c00Dm6PWbw9ecqhhyD47aqb5gG5v57Nk9BoDM69IK3pJH93pxgiKVbz6dH9
066PsxvgMgrtPFBOipW7uFwmyBziLjjtUoChpbNCWAB0MD2xB5rzNUIoAi3XOZ6b
CcSZcyWPMF8y3iEohauF2SJlISTQJiefrEY9iN8HuHA1f/EuiAJ5BWoBYyYXt+03
hkLGBM4OCUJHmwM+7KrlHXtbvqx8xJYImvfjyXFig4RvFjdFFs8yZow/+7d7x6Yc
rVLwXtOW6qi4mRk5mFAMKcMTNaRIfKdnbqG33870puThFtMKlgQjolBIDQM0WGkD
wnIHlE003//w+aCGGWD8rcPHuBLmxaNUattQepBaN51iZAy09UAybOo2xkHuKiiP
Fraa1KnKEpFwriUfkilhbS/2s0IuSAo9hdbnSUKXJnk/6o/7232JgBszb2ltd9JA
NJO3Uqm5oanr0NowBc8AtMZ4UA95+pI5Y/ZEB3520qG6pqZR+XjEsnCsFFlLnWKU
lYr+/vRVdTOuvYPs9KK/QBgB3uNreje1VVLQ99R1WJTnpo8jjg/PqNa//t36btlC
h8yHdjIOKEmQQQKmxdiwBuf7hR3wM5DwErAqqACkegoUI2HkyMcg4Ddl6skogSvF
B+l1Q4wuRfPqS7/i7+XAGGY8L+AM5WUtWGOW7uocS9jxj9RE1PSEBr00ZEV3V6+B
HLtapy5IZgfU7ZBon/4WLErdJ/52ZcgPb7Bxz1sxXpgAOfT/hq2bfVA7vlpoBTEo
JE0lof+/OFm/d8+guIG/USnV8DeXkkINVjZpYV2YPm0VoKQTzMjez3D4DmbJJ213
bydO/wmZvlpOGGhrq3obbPqeZFa0Q32dw3pDF08tLh2VWw/Yysd7rI//mJd7X8Fn
NeD/VYrC9P1OR+h9XKx016yXEv6me+30r+95lHSj+B64x9yQVMm2VpPQ5/VxXOG1
YbvS5chrnn0Df283LqCAkUYp3CZPWpwe9HGwDbxjQFwrtgYek/eWT98bQZSzZjgz
kETQasy3YtpAYnyUjT0MwCaFxkFKznE7lpQGepjuu4707SLRnzeFQ9NIfw8UC/fJ
a5kHcKJ27SmpYUPzZPbWSmSJpXCQnaXM5WwO2GL6241F/hBBPTDIrk1xi9WJyqr9
avNbVP4Ct6EiZs8Mia8R0g4sv4bkC068YfGhIniePYWdKdeR0Y071j5d5piNSFQh
HkuV1jyVFC+lKYwPaOp7YOLGLKEA5ew5pM0GF0Kix/mEV602b+K6IvbUddrHl8Ww
KwOUrDuvKA+AceRgI4HNkJMaznDROPwXNLWnOIh1KnXb9YYdHzX0kP7ZUWHb6QLD
a6srjL5Z5CY0g3NXFr8RRADZ1TxSsvS3LQ/QN/0pgbLHZgUCOS3YgM6ElcC/ydZo
uHu4Q+SmR6/LqXCXM5rBzBqVSSMN6206kY5g8tLs8r9HHWy6UDebl23nhb5vM/Kd
rseeuCVAF/F95NtcE652Mko8A2Wo2S4K19qGlBsP/ofVR0M+ZhHfNJI24Wf7zz3w
hcBAwKD+t/wo9hRCHXlIrsi8k+tEa6XdyG8WSxdysSavsS+pAmJefICheorUn9qy
kmKY+cdrq2UyFCp1HtbhzcdpC3L0Ms/W9M9McoDpKuAklXsmwzU+49hpM5najb+h
e2MC/f5nGAetT2W/eE5Qq1vqZgZtO/Fuln7Bs+8vKfwPymGwUUgr+sVMVLN4qgMz
6JrI1hVQjWx6TqBjW9GEJd1naFq+L3jLf/6y2RsVKJVfLysi696xR+WkgY0asiOk
WxjJdt6fCPXVGVOVvpZY+xISJiz6A3kQBvb1v+nqCgC+RAlUzRtTqEGmaWAFt8jo
0iXPk273HggvuTBX8aeMJnMn05QlcIGj+NoqRo2mbox5rLu4UZjEquUQ1ueApUT9
VZOHm+0NimtCLPm/u7gS8JBtVI6/B/5A7aT67+4ou7Sawl4l86tpVYD6Q3/d1/z2
ozukpsQxYcI0L9l+D4wxo0P3aufUFxqFiaBEwyqAWWbFgk5JKbBEsxlgNZsc8Bzh
wrTp1VjLgEr2pmw2VsKMOZArwadFNTun/G5L5yByp0Z6e9H+c5gCf0+cPl8aQP4t
l2Z+Oo3R10Tz2qestN1HI+sceNT5SeUM/13ZYLM8EDxvCC4DBN9ooB4SfFFJXdab
ucMcCOi2vVF0YvLsqtnrPu8aNJCU32qm7qGC+7eYtCylVLIQZqD9oQa3aGpvcZFK
qThqcPsEM2e7lHJ81BkF7LEPkGOE7TcIo8h7Xha68SgvgCS1xENjLf57TIBqQTm5
IdxtB5r9og9QE6VMU8e9xbLZbKeKakX/qAMvqAOfFqNoT6K3IJ4osLKa2gvYdysk
kbGqtEnv7MM3E0asc0N9CFzafmQcmaEDNHeGofgu+lJ9EUb5mu0EanJe2RpBhg8v
luvDmfxQVvjlHghK5HDQCVawLx9zB/rCGV4c4utG4utekIeQJu5R9e5gDAxfYwnU
xWPkGzXTUhyIuqykkfC0xjPgOWwfaAoA4gEFNthRBi5UNnYnM8QvgdKhLc46eBUr
vihfWNSFblvZhGc04GCJAY7VqsaQU+xTiqu+VTvW0nuTHy5lbzZyfYb3JDDKkKsI
lEXFYwAPui4VUlgsKS29228YG7ji5iWEcIHCszf9yiUpIoMKknhQUMgzVFLiC6Us
ip5tajDFJWgA+WqJQNUFo/iBGy1nhP+j012rz+EjEUkaa2/MkgiDq9mGc0Oe/DSO
WmvVo6O6utDFvXHk2Qbt2VgFlUp7//QnCQg9PZgzTrShzKljniNkuy63q8rZT6/1
T1bIhLt3XgtPIXmQIE4XAHZLJ3A485IchsHPMinPh56DaIM6CHWGu1YQkXshjyUH
GFfMPNuhFtvcSvWoYMYNcEIhA/G5y6h44hrqSgccxh/mTrM8U8LOUEi0JIPA+tLX
xOMWHs1OZmX60Rp+FDCzb7fVLkdeZTylEWQwGOiqGjjECaLqFfVCEpRv3ewhr8yK
TCZop2bPlO8WfKpmCJRKSEZrn7GB/Qmjz2bv4b4XLkFhdiSeYa346AgF/GsQfmYN
28n/0L8Js2JUpECG++P+M0tYPtKEPYKzS3m6ioCaCoiYzwH8hEen+KCZF74c6SAV
IRx/qJQAG9j6rNO4Kj4txDmk1pemD71LR5PzHZtvkD/CeygeZeROJtzSyJrQID19
avEO/RKiCJis2VVWMsoqk0vtoVDZShMTp/yyAYSIufPjhELmz/nNHxMBy5bMv1Wg
QkY1/3EEt6JryNZ9g4Uoo1HwSBkpjFyG9PNBlxKQ2idN81ooGc6dOU0t8OkWlXAZ
giu608wtHjdne2imqGUmAC1/FUvEZgLpE/MakpvcjeYMnsLs/9/eEz/+nOFoJvSJ
uLI37LyFWZ9FaHnDRHi+oTKBzmu6kaj1dJk85Wb64FpLrZRkGJUi7GVAJDMwsfnh
9NFSsxkeee81zIoYrIms5sYnSoP1ZuVDh1sOouaaJWINIFtsLlKuyN60XIeSgzel
xaxEhurQmo56H9OkiseDJ+Tt4VMyx2UdjVMmOd+XE5oJq9Uke8ROU5p3aWRU3T67
+akoH4sIYSmaqYPN2jJN0mYfnK2O82/RihkF25mwYHZZ+u/PZjvPBuJ+4jbe00NY
+ejmE+NSrnuLLuBiNiWVOdJ6Qb4nviTW+VfhrlD4L1/QPxwwL3Icz1LLnYF+jWN9
03uBFW2DIdecTd+MM4tfhYKSIHKmiPXUZxjgX6//8yMKm1ZbHEEoqyWi0TkWj0H/
Ino2R8OTet4+Ua24qSheV2iWS7Z/8eyfkW2OoQqzJy6EqHqrr/yFTisLhPTke6bx
aQmB3LSu8G9C83Z0+TSe00mi6nOSLLRQrAYdeR46H+lxALNox7sLz3SOhEg0eTcs
AIaFRsmpwBq55NZlj4vBpOpscig1AZonKd+1cqK0pnQTYedzgEofpPUcsiQc1Oe2
m7ehi32dy5yQjjAiMt4tP04Cy6ipjQdsdtou8EhmsEbypZ7SxlcBJOfETnPfblbh
wiLptmWdv2lwDI/Jv2uzjelY1/qziwNRaVYTZiJDEQ0S2BPRWFG9qcg+EkTpJNia
NEQmK78kpsQX1fUsjprrLwTsguKX6vsgyA9+QFCchGNMF3Ma7f6pkfuTWzyWYNAI
okh35cqOtnudrHhkgyLiTxG84OL94bGzhltNMEZY3xh+rT+rjtAV7x3QdJWGn31y
nnCT0eY/x7b/DpKvI7wSyJRvckXlrKIfiKx8i4j4kL7UA+6kf+Y8f1QRowALsDXb
rX/fCfTGGZaBq014d4/Nur27JUYiMVBmmlMDWRqyWHbveDJDryPCWh22jvoSwETD
dk+KFU7wT8MaC+XbmrhO7u7jVSCjw4OzTO4gHHvyhWnLHfEqkY4OvcLahXEa5mWE
fQA9F9xoH9Z7rPGjK89/CefWnOmsfAfHcW1vL9VWQZu5Wk2wmWuAc8Wb51SmELDM
Q9jC/YHzfxeu3uGktChZDzmGU5gKY4UTfvqdGjxaUZx6X48jbF08NjBf9Soj0Mfm
uFTKe0bhPTLv5VcQs3m8FLCiGXwDLlpS0OHGbx8WxQbozz5BMvHwdZXZ4T0FQV7d
V1KBsroAYwFjqnCsqNcF97LihGIaGOT0n0uB2WCvH9xicvRCbn3GK081Dgfmnjcg
MPhxPubeiUAnqE1JW74va6aw1BrmQ8iaNFD4L7aoPCFyOZ4YipUlfIcXPjKxqSE8
xDW/eXvnOW7UQvM+HgIm6n6kxAETnLS7u+LPa8TM7AT9LmBbs21CFjmdLzexd9L9
7oJCH4Y+VDEShgQX2ebGGFJ5t10gIGonVm3bnRrO6MIsjWylOgoDvlTD1wvaXA2W
yDjIHuGyKfoT/xHW5e11FphShRhLLYigLzEnynUIK4OZV5xRgl6dwPTUSWUnsls0
YiyWrF0ww/aeMjT4x/bLBGABWh19G+ZgEe5nFHskQT0zfSoiSqQ7T89DAwwbFwIO
5UvciXu48qA/5sVVlrzxHp4KsrmweYz+RvN7E16EFF9JjIrSXU7ydAG1BOgzpOQR
wbzi4KYiVanjOze4IhfzAzSVlnem7cEznQGMiTI/M72khJS8FDnjny6j+jCgLT0t
v0XdoDysFkXJ+KvJb8BoMSgOZUWIPwsXbpeQ1cUqoxJi8djEY8z39rQ9XLf+yz8b
ti4FdfV9xzKXiWwmFajT4bLFYAiWSsSISOiF65dQY6UlHHeRqIkrL9G+t19qsiNo
5+H9EjSM+W2z8Jl+DF34A7HBuLrAY70Do88D0j+nSYgs5z6LiMNCqWMsFKjZEkD0
HIENMuY6AL+85RF4n42CAfcFSi0hGPpyvE2LMM6f7t5yihq6eB0k89D10ef3AdEC
tOj9ugrIIf87jlWopBVINh+w7c9/Q+BC/hHJpEIqNOzRp72UXS4hLiCrG9+Xw20l
XSEHj8mY59noCT836nO/mdLpGUoSdGQkkr3ulQAhaui/6QC9/G/+5xqCGLI0wqKK
tn2xsvDQCnz0jNVNOeELMRYDPj+HpRxqkMmWJb8r8DdBVi7j/9CBjFc+KBPwwsLD
qNjQLTlb/He2UuuVtkAwXHNHfOZ/CsMhD73KfoXs2nWQx6ZW56WQNSv/s8grQR0Q
NGBEOVis9d+wg2NiwToUfYGfiQVL8wPYaZrvbm2/uZ5yda2O7dxn7ke41vBzaBwp
NkRwJv05pGC7XNjYhpySlqr/mKGnn3p7LYWc6ewY1a7gsBJBXD+mN30IBoTwCxKI
JJioXjKIijI7sTMdNtaRtewYyDrVlYmUs583EriMOFBuGS6w6OMSHqWULLyyxJaB
LT5pPEBMmc1RllYO9xUq1Z+IdAGWWJIOp+R/ZA9NPNahPSG6wp/gFCpWMolqTpaD
60NsjYwrbMkctmYxEXn/dQOplC7elTpDtUqnBnITU9SY50f+icb9AZIOF1fYDxix
iq303BQYlSpKxcahAM+ol0ABmZqW6kuoXbZCd+U7SpuBi4UdIsRKKTeHUd4xNuuN
01BYfla7KmZcckFunteaXldYOG51B6YT9y6kpt/vxlSUhaFOZa72frfQNOCjdzP/
lIGxoAW3rrZzZsseTaCaZ2aPQUVjP8oT9qaKghDtTHoAKAvNJFDs+jmi04booCTC
3r5cx5e2xklpvdimn8QwD1QYJHgYDATQE7T3nWKjzSSslyH9/0aP0VcH4axoFdj/
vO+7gkVOlSDF+iIoyIcA5HflcqDpDdUeTO2430eXn3R77g2kwD5CWz4UtXXbWUtn
JF/hOjtMFs/P5z1AKkUbfiU8aEO5rQHv4kopwJ9HHmNRweMPVBehuqEGKcmeb3fR
C3XX53+Kko9VpAFwMI0hLaaecKgfQeUbEckr0rebHw3KCoiVn22G5CZGXpr9wfQH
7VksAjENlf/9kqal+fr/sPTyiGd95wX09Uw83w35pHohQQjTT6nBfhPZhT8WOxGh
h8a/j8SZ41SI6IjLs9Z0L8eKSPW7XRdyBVrSD8L6FNDx729BMuSZcZb1oqTSCIeO
pzZXUkyr7Hyip8hmv+t3Gi8EfEC+zI/fox5f6Z+WzptM/XnVF1tDiY3EYqH4HXy1
fbfnW+n5f4k6SgC0ZzkhyTL/ViqqSNbhfHNPFaov3g9sySyNCHH/q6H2homx3Yfh
Q3X/dwxt/4iWqaYJhBXZo2yRWr55oBZPP/BheUFJEo+cKiW7/ayImDD4r6afZBLw
8mZZxeJ7tcCX6uRf/QPmiDueuR3QkaAb+ufbE64Suk1dDCQdOCqP9GsAhuEmCsYn
h3ehRb9/YmE164p/6xgB9fKT0+dCjdjIdcUPYS8O8spoC4NlNpTqOMzyWuVuGW+1
skH59rNtUdjEpU4ijZgNJ34Zmm6XP2J2gfG31VZqz0QKG9H6oIcUyrOcPwmL7CML
DqN+aanPceQo/qHiQwOyIpDjyMKj/GMikO3Bkn56Agk=
`pragma protect end_protected
