// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
zhprFNzkIe2RFnZiYMn6vYtJ7NcTzcA8BzlYhF78DZB6GUcDz3e7Tfu3h9+Prnvofi4+by9AFO5o
nY8teT5S+fYSmI6HR37t7C6tyiFDb6vK5FZyRVhIGgWPWknHCquvlDsVQYkd5QGO6Lt9q8yBnzpo
LgCv1guATZuvG/Y9wLCVBEU/5rSTBMultL2wsLASkP5dJurOUVWw/fH+JEhUkSvmM/P2HjwBN0K/
qn76kuLmRSf82o9QvbiQnwVkCGFdhiNkNQvaNeVFTE3AKOWs0C8dvrsWcNVSwrPa5sNP3Jhl/oP4
tHcV7Cy7dcrFy83QRLqFHVK5/Mu/QlXhFIe1Tg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14000)
Kq4FLQUkACwRhQ/u46S0J8rsC6tCTiMWgJ+NFXAVlcyeQ77qVMwiqLV5dHUT0a+CvgNGL6bF9Kgy
BfazS3ITxy/1PupG1fKvZuMV+ohemwJkQLzceN33Ag9SE25OzcXFAk/xECZtOTGPAqglO3Wewm0D
RKhInAR5G61wdMGzTPhxY9VyOkLJL/jp+NCbb7Pw5qg1ojVpugLi3hq6yDJ1qZiUqOfzIAHPYyHf
ilJsUyhuzO2OOksW16nDstIQlgpdV8SqQGmW+ObBIZrjoM32ouNcZ22NU8xgzNYxx2k9xV0Kn/h4
UQz/lxwGHwjYU2Ub5vRkm4ibHUFLqOx1JtTjyYFwTHPsMuPvp4RXhRUuklvHDZgTukS8OFfukHX5
5HW9D0R2pMw9SdHJEoKwp5L5Ko1w3pEUBrJC8Nu1MqeSvHFFrl3K5B0VUHnzP4ZUVgF2qeWGBmVZ
nuh9R9JBG9MeR+wrqficQsWQx4weZNyQe+ICCAARw9+c6OkzfNJHBNsAp/VHzLq0k7Y3q4bWpPgR
+24pU+SRc+WkAo4EU1ZICipwxvC03TXfOv2cRHJ5VpWsGo94PwhdFM10jx9X58KLa1UIjkv8XODp
dpfKBqWaSQAdalNA+cokrIy00E0zfAfkuAxFVj4X4Zj6QD0UwW1SMqy+Kf6nC8s8vPO960l4rB4z
zrz4dqc+BuTU0lD0VtlNgbVkA2xhGqCYP0+QMlUrctOoa5/z7IECK7tygHriVZqJs4XqTu+s8hc/
xs/c6RNcYq5+lEwUByqR/QOgDuEnohijJHxeUUt9XP8zobhc3uvgAK1oIyzBsixX36ko229O4ij/
qE8MFuIvD9sPFH4CHK3G1tfht9YBuJ3ZQUr8/ueJibHRmITrO5yWxlT0tbTc3R3KQRkCN07Q6hB6
qHXTQo1vltP8MCyflCBeYLr+YvvusIBXsi59Lieq0MTTehmmj+8QLVRerFLKklZDdYNmLd2xh/y/
gnbjkmregesFx7FqB5lCWbDULj9PNCMRq5zTUa2N5BhGcpdqmTrKNPwFP1AR/Hm98wVhOTvMQAak
F8NQvI6ff0rkH4UohJfu0jhPDtfsx62Q2BKWNP+rWVsaGCiF1KPisBqbT8ksStrX01gwZAJTS5Hu
Z4VlwScrnfwp3IhQ3bha92gCtNUPM2D5JfYpksqpf9xYCB5pIbB4Limnx16jOdgUZYZLKTSnq2UJ
v/aGDrbW9CNshJ7CdVR1BjNuknHWij+gPr6lbtr2dJZQjpXtd/ISvh24ruNG5lvvWnjGIzDe6pk8
WzVVCCcHI4HGzWlMvrI5FJYmO7bU1Ai08efbM5gpSwpn4CDEt9eMMo61pebZm6xEwSnZp9L5D5IU
6CMO9RD0RPj8kD+UMfXPJ+fPP1m7UWSV7QhAcBXKMopX7wsEx2Gp25R4+v8b9aewIRWQElenTZfy
4p8I8vBiHt2dBPoxTLR5NbSfcVNtqqu12yncXRzLU95fcclZZMgxo7TEVCYso1BGJo4pa77CvlM8
6CkVOEgxWssvsVz/RGie89gnNF5AZNT6ZFqHja5xISPerbQdS2C1q9CxJBjEjwfHbeQqW/luz/0T
wNbeNesnQhmiLGpuf/khQ//9h6lrS6yYkVz/x+ahyTbTXWjGOzAut06t8soQL5RS4b9TZrGpLDar
9p9Ai+a+ONl0KP1w5WYr63hxQ5V9tm4Sz5jts9ArtfNuya4vZQD6TGg1emxQ0eRy9iANhsf4gt9L
ImVZdaT4jYCFT+2Bg6MVGACEoHCLo2SPbijyIbxtd63xsYSmDECfW3m9Yiqks1bTtTF9DnVOr7mX
cw1v5mFhI+Qyw4o9eCc68bOND7WlaBhTXtwqnEdwL+1DnqTXnDd2rPm3LxcW7If0+JgMpMLcagY2
O18O2iVs2ep+kopfn7PxJH7r7igICYk79QAoJoVNGiyA3S0eO671GEY8s9TPGpJx8ZXkpc/rmXNE
VmF8cOli7IlCD8v1ffr9GmsIC+8KLPW58XY+31Pn7mS7PHGlcuXuGDuzKOkeOOfaaO8an9Vk24cN
+m6SOYAH+pv9M0cL/Ji4ElzNzk/BL+gDrdvlINH76IHOf/Fb7NwY6yerF1q6ghkAXe4ohmwd51Sb
a5B0bxoukBHdL4/zN0ZLfc0VpJVlO7+IZSsLf4nEReIuzLefdWwJnqIQirTtqhEzqQsQBO0D0oNz
IxOvuobMOubyutJzS66bMsniJXQo/NATE/uYSuNE7tXg4NuCCKh7HCHSARrZ7m4TD42jrSjnUn18
C6gmEV8yBRMACWswYBPTRQvW9tcEf+sXZbF/N/Chvk1Pd2eQG1BAHsNie+obwfTpUuq260kXRSQr
b0z30MH8zn2+6427c7wDpVcZ4P3NZuKenXJtK1Y4FgdpS0vnC8CGyVlLbFylzyJ13PnuGrTIlj2L
y0C+KBYK0jgsA1uO8U62U5iL8Zdcq9fEUSHI3E7EYdWHhFcyJzBNA+6eN6E8oHsehQmoB44z5Acn
lCfmCp9TSES4qsDEfk2s0wH2k54WaP3wsfCIjF9x9KLlGLWrtEsbbJX6HwhRf+Y/mp7qOqV6HmPi
yLXw+u/as+fTC3R8PGs+g4Os4AGvCDDTqbR6KAKH5dPRcUPburudGHYwKI+yJ5UXwpkrLXm6liXI
KWmwtSvnFigS2BbqAGEJYH2FeD1BYfvCpwMKUIiKKIlFoNu60IqRUQl5lYm3OEe27l80sIHqdUja
7Gt2CrGDej/eIoJYQVOcc6KePMGOfXpKnGQKShUkaymVS5427e+BM4fozKgvzwY5VlKdChwgpHm0
LrdwZJ5+AMETqtFlGLCTZlG//dCOXGhU/NDoioc4nPhlPrQ6P4xs+U1WK5BOom91AADPbzGTBwBX
aD7Kzay0gEUxjX4Fd4a+b0bPAvmcFa2JFgOB/x8R/owoFeIvxCFfYSlS4qk4UBv29yRKjAkE9eja
WxCodEqn43Izo9GtzrNB36loHjAMW94KQ1L+/B1TjzG4JA+cYAxkHZkxm6WtBkT++abYpDLt0ifb
9r3LBGCTVzlqK1lyf60WDQNenUJLKK+zrT8eFJivA+ayqcadyHwo8z3og1lILCgyXPBr0upTV0WT
KHIeIjSt+oLbM3lywQlX9VDk5Vi6GsNng3lUsOd8/EZ74pib8wCdgBhXjjhVPIDspzqwjKDOgZ6b
pFPmqOJ6nCtGH7kObUr6PUWthlly42lFW8wWlyWeX9Te6mVrpWmmXoBgjcyuilc9P38hhZdoA7RR
q4zbRr7YRpKQXMTEdAmp4qWBb8J0HRzRhCkFfYEa+kdyQ3kQAR7IuGlq1Pnr0SiQzbEDSTJIFWVH
vurwILUT1Po0yrDQSvEydLIfUZBINllxouQCZPMUrlHgL/hhuCvE6vKRFnfjsHJm0S3ZnktUOfwV
IMa0d6FX1Of9lByNC4IdPujaDwIO1zNigB5m4GWInSOyy2xPs3g/nITh+zqYWNKX3Y01nmEcbPwB
p2H4R90umVpoULU5PF/PZ79swHi6SjCrRvYa4EqgnUnhn9ycf3kTknDrYXrf+TMWbl2Plj5n8JG9
3h5flQNtlO6yK99FGhBW/V5E9taVHTrXZ4HZpsWFNtL+d5h0WXq4bfV9OH0E+CjBsMuqTW260yYS
BonsuVHsNkn7XLqbgOpDCS1nw1c9vTcwtvX3+dN8qW72iP1wuK+//UganTJ3ULx2p7jX2TLrC7EU
XpgF9nOhE3qR6hbeyJTKEfJZjIJClH4AsZMyLtOvfkAnKsBXmIGg6IEEp8WA5iiILU/a0npm/3Xg
T7hAqA3+63sAU0E3hQt5ggburBPfaS9fK5SuUmVUMtBVen1q4N3DbAf1v50b9nnKC5LB/PKDlVyP
79FuGTW/cd+QlSOX8kLGqG8cNIvabn0UbIAudB6pdx2UydfBCM11HUHP/0GYeiPVnMlKQJY6TdT8
UsdmHwgn/MeuuKzvDmd25i/XtO6mlzmoxfVYyXjgZduPWktS6O8SgUf+4N4vZU90/rZXEuXXBtPd
cq9hG2rgNeoTnEia9r7tEEbf6habiWJOgvQ3EBIuRLz1xCnBUwtT/zHepwu/eOgC67TSiuCPEQS4
KNvNtcn1DQji3iKURkTe3LvxZP6gZxNQL38fPbXzsr85x+2S72ehD0dPK/zDl55Q0GqDfPNv86qK
59JINan6xgHx4PKWUqszukOkDn1Tx0Cs7UlElem4Sckw+pJyE438XQaq6zLepmAV9eJDvOKoigYJ
NJ683CgmIwCZOfcefvudyTg+D1CDh+6tW4rQRHJhHl0rxWQThRVNS5JlQHy1hF9Xsf2RiMVqs+EA
Bb9KcDhtVScbuZq4ybodDj9OxC2uUOOtaFE1j6mLG6ajgc5uM6SOzUiJltaKWAlpBQ9i0aKmAKzc
UW2kHJXBXB6JnIQxf0AMi4ZA7macjvAwkOrbg8+oUcW6xz1uRUL+g9lK2LFM5g2h2IWNiIT2FJII
iOh9KV6YQDqy6LVFgH/XYa+qamHP/CfSr05odqZm3pEtDlCZRzgDtaRv5RrWpYWRa12LmkPLGtrS
iUKtoZHzYnJFECL6RhbO59gHpevsenu5I1x8O8AZ83izxbY0P0JzW4OXGmAi3DkwiixZngOYGafU
Ib97r9puzf4DLDau3dWeqADnS3U95x2q/HDw4XWfNC9U18yaorr36UvOAOOEumoNKxEnxcch6WnS
FeQIDaT0yLduPCOJwrMlC19Ndc1RC/bd1W4+DNINHGidDnszczQnYwYz/eccfapvoZzdnv/HBcTZ
C0suhoidP/gBSGtBwiq+yykLdpICjrwznjUe953m+xQIMsCjsvb0GP7ciRA5It3hzYclUf7V17ME
nviGOcBv3gJs86f7f7wxly1tFU0LdnJ7pcZmIqAXL0UlIWo963z6WH67ND7dNK5EfKTuXppW/m5l
b/JXwCjdJQwOnlvrJx6ntIplIku7F8gLyEqj7A4FyarCc2xeHpzZv/MpHFMcxU9UJi5S7N4UzINI
i0UZhTaW0txdhmek0UU5YmUVe2Wo1s2EyrRpvqbfdfaL+lykxzlkiB0yswueidHHF8sV5DmN2JSl
26rWgzr5FrcpoLIlvrxh5IgXaRv5oBAc/qm1kfimspiQz0BPfXsn9Ex4wLU3DWgK22C21R63xoAF
O9elK5MS0Np8UC5UcWX3bjDqeRd91qShndJfLk21oAzZh+KTTBI/Nh/UJ5LAJy1J1Hrfi5OO6qjf
nK9R/cjmU2+agWzfwCLTABXQiws8SO7D2wtpI1+i3WPPCEsoYBbCpa5iayg3wc87OWhpKxohE8FM
aIe7XJCXr4Pwt8V/FGJMyjFb9Z4SekPSJJrZfk6nbPFnl5R8eDxTl6YtmFFva5p5Pgnu4kyFkAt2
b47sGzxoTdnXer3MswELxzIS8ZMFUN+3xgj142AqOCUqs24XZ6x1+HiENKubNej4ijBqf0fFli5A
Ay/BxiLwD1kd07b2o99d5sJ5Zf1eFcgBdl8L7uT9/bduOoC1ovoJDeM36UBrICy6K8Lu4zURms9o
7sg1myeYimMgR4jc/42veappZa8jWT0E6StT7ISnfCSsE9DA+3DBE/ufo5DDtFMg57sXp5MT+E7x
fp3KwAgSlAjrZCwPwWPhukM2TSeFOafQlFk8hTfma376/xYidtiSEtDY3IYQua4KDIJYN5dL7dGc
Soacqnzaq+F99Mhir+oHVEGQ/Q+UahIX+19/PmmN8uC2vW64i7a8DzetfSsTP8BxBNQ5vcNacy8k
KqUKn8ui+jwfTWF1AUjX9sPUdw8+tY/ezSdEcLgQwcVcBgZBoHdZ7L12+K7rxodKodPxUDC0qLfp
2lb/HNqCLpiZvO/TFVP3RDPUbzYmWZIkhlIJumC/ftxpgRz/W65h/ggXou4RetXoI/aQYmfh7/q8
96ai8WeqixRGvM47goIzGJLEcKZWOHjSETzHVyH04DOXObUdN4Pyoi+h1XIlZmQbd30Jl2DZL2TI
wgFHorzu6H3JIbTv4C3HvtoM23nBzZ8VqltRWTs4X4ulHLrn6KdMd0gBmNcDmX7/Pl2f8sasSf5K
uQKJsb2McVInOgFrRXmF2EaPCqkfcGsInLvLd3tHcsXK81ha8FOi9qCnrBIJx2ROEyS0xTtn9AtN
A1q5I1+xmjkHusA1re3ME3SY5BBuYZVYMf+ePNHk1pKiF1OrEvPNw5yT+0uitubEV+PfZfTPAXdi
sqWHzATckP5zToNlzIzR1n19BwYw0rThfe8I52jbKacVTi9tVvH359eD0HsyDhHX+FxakcCTHsQg
aOegt0mp2Xc827HXvpwYGXr64l39hNgTUvtsSUEydhllQ0nhPlIq2bt9eFtqqtkIDOkC5vC/y9k8
lcg0OXKi+NRyzlvxEYr1Bm6YzaRMj3rSx2VItql6l+djgKwHiUTYOXntPXjPfCniiKmUYd7vhoMM
ZfZOe42hE0ijCHlDGuEFJK5hJrLvnOFp7yINF9EgOLh1JbsyVvsvl9w1to6sVTbcOYY2PK4wq9N4
YczUF0zT7LPlu+2KtGiO2OT1kvuh1wmsE6vX8OAJJfx/e12ZFmwWVRvJKNbLKNL9xOZrb9ejT9jM
ND9F1Dzn9lJiIvErlOk5/pOiLHWiw1Y0l6ZrZl/S67Dy2gV++i9TdArt5qb5pUYFsYnQUK14ys8O
8a/MSpE/abZ1hfUnRC4IRdhrF3fooBZqB2nnde94OVIbscyEvXwF5TBDT326hiBSGKTzGqJr5CLs
QLljvFroBCZc16FC2k4SSgIV1YWCs1acvqthjtThmom20lO/lRrcyY8IQDZqjbwyvdDYif5dw3wI
o4bzx9HBBjKkqwddariSvpxftz2lzh3aOlhme5JqMukipXC0B84nGrXS3xiR2I+uNIz5WBpwcOGo
xq/S0MHOdg47U5aCNrtXawN4CDS4eowKrZdsGoZDuKvLQDUO4fe+HB0nrYS4P4yijChRbsW/LxiD
lPhVqiV27+hsmq3WXSGFc22rO1mVXN1JgjklXYUdNp3fKbN01JlMmDlElxOaVFyaN8aF1Gv+I4qM
d/aGBqDNDpg+erRlpzTg0E8FjQZ6XZSogMd9cuGCGdRiCX5WiXzlJKryjtVFuU8RgsOBJJ1hjvA6
q9Cxry0+9oesC7OiqztpaPm2cAxCpIyoCVumNqnasOrhFGAXRqah94Leb0lgxkeqCykM2FX+A08S
QDEu13fKzGVwq7FHgm3nYQOsKHk1D213A+TLg9MisakabQOo5uDwnlNvqcuJsipXf7DGTLcuDYP0
RQ6CE3vvN/Qm6551D3WojedqXTRjeCmd7d+cVrTaN/lokCsTrL4QWoQj6b2uiCdVZFo0CkzRlg7f
IblqDRTxPam4odM2RqmLWHYp/Rn6poxdpgHAyRMIaOYxQT7iPiT/WgwsfLcOdKOZHVQ7WqwcjIhi
RF90EA9tEu606VSTbX2cQB0wxWStH/zGE6ifllrXMmxdNmuhQR0NuGeWyCm1dhwEKPeOYo4s7l+M
T0alHA7R8oW5vsSchTNJ+r8irNU1NYkFcYCct5iNhrZ1EO74xXsujEbFNfDg3jeZPo6Mg+/zoI6A
1EUip3R5nM5qJWQofTSCJxhdF2qf04VmtjR9ZY5hk/ycbkeM8zwQHUVYy1DFLWt6QqQd6x9fHga+
48MPDm6H7ACxLEfSnhilZ5D2dl274eUZY16VCWX4wfp7W/YOrV/0dw/sII3awLACnFEIY4EtWFUD
rDgzbUx9MJgcL2UT8BZewDNeJk0AOqvbLX2+PkjNcFx1hUE2zwBzXvVuGAVWqCtie3X3YfbWO/ma
PTaivCRDFgihqu+/rcB4v1r5yD2lqxGCiIp5PAWHLPisil6AqN5UgxsKBFXuFtiV8D0dMci8R+5x
dg2NOpRtDea+YB4N7By+njpWr0pgFSEd/nzVffx+qF96fXS4uH5kG6jhEJL/5qEnFboLmqGxBvpw
16jBQmTk/sYyYDaKk35CvZr8fSugL415+SaluDu72z7SOcZRtfpJdDGy5E0DSlRbF+mXjubOZ/EY
6XZif84sohxjOfhHqmiFWThi1EFEvKTXThwbQ/O68OT+aGZVqD5TVBUHbZiI5yzCJCYsF/PpTTYc
h/cF8USlvsiZq8v66zrJY2Pbm/pV+Aezl2sSC9SpWvGardZFDztzvbjDtZT5IOHUiSKRBWjd++DK
TBW8Rnfzft43QwCGS46t24+Wr1x5aq4ty217wVVsNnGnFIiIXFriu8p1y7X2hIS9GjfN7qxa05WF
76DCfBjd9KtmjYk0WywzXdA9rUFeSXFOvWuzjnQVcQKNbCS6rVEi4ga0Yj/6BrdVgxHYH2aSM2OV
KNJDqjUO40pyFQ+Rgl1TvroJIq5tVT/tC4EIznigMUu8yU0hFLZp6apf/gndUSSswm1QKwsYZsGa
6nQwqu0G5PdhMVGoMFdAE+snThlQIydXUG3cpgk7rDVTDYFw+wUpmY0E/Tuvh8ZKFyygDTYtsiNW
18o3KxG/tntSBiAY1mG2fpKbBMgG6rXArd2hW+SceVdXaIzGjIUrPmLTZxNC+DQkJ9X8Mq8+99eI
z2pLEqbkYT9qTdOGINTwMM7L0NahPxrXpHyVAH1iEdyJ4wF1kIueAUp/PM8aGExZE+cdt3lM+QA8
d/UCdHWXaP1jytEr3vu6uiymdl6duzJ/bu//rf6dLK8+msKpXHNlIkugQQd3FEhI6toQTBtQTKvv
fKfiNQNHtXGOT7qCRRobhjro3zsctPFGjOp650qt0lxr6rVEbPLOl+QstzCPoFbd2jZo0RHn5dBA
rqCcCRV0qKJozw4DJKsTD+OsTxK06BBX5uaC35kl/kvo1u6S4g8VAz43P/giVxyS4+EpIXtXOx+2
S5e0Xy8M5UjRU9vQJbSw77zJPBslGv1hU4FrpoUeN2k/QJtLYwbSC85hrUe3yrDstZrdLOxJFOuy
hvewvhRW+cMvUrlSrpqioJHE4yr6RVlfHlhZq1aU9IyEMoFEUX7FpSqFLK0LaqSoa68iSQgpE7Fr
un2xDRfJwBIakq6biBl6NS/r+HJKHqLVXSRewvwMwwwG5TK7vKeEM6XNIQUgzm+rTUbfCLot95+b
iVnk/Dk3q5mAEDtMOBjrQvxMwuZeYdmKPUaoleEs8AbduSz4iVtcu3II00WByQ65dz6RT5MySEKu
BBGhc7tVQBc7wN3OUEHMSdLfOPYwoTXfq9zr0gfrf6WA9hWKDE/b6O9JD82uH2h8cxZeyauw6+3q
t5OZ81cQ2/bn7/KWo5nNpFSCZxHgaD1vsc1UoyoELlJSEe72fCnq8fhDhocyVk0ozruiJuf+qEp1
QS/hfKDfugnvpWMfaCovWn4TFaz/DSY7WX21V/SjPlqTqYdyUIbhTXDdpKqVZFgeOWaSY2v8dGZE
yI/f3XlG0RRAxfvJOXuwkwbLHpoazspE0HZbcbN5Zz85kIk3+xCUiHJu+gMqdDoXlHeiVaqZVKLG
6WN0lt/hdQtKTtE9znEewQIC4CChFoImI7s6toVDgnDRewtUDpmHxDukMDW7LkMih25whJbdI2sw
9Pahl5mXgU0f2He+eb76xR/d3utXU/QY3HEuCAEdgO7aUtMC3dqHaXEdIln5bgunG2DIBFyGxBbt
+2hGGUbhvEdpEMLGkxZ0g29YM1GMoZd9aPcTYUnqgW/h7ZIcH6juVQmku2byd2FP6MRB+tQO3fm7
et96d15nrXT5s8jch8kXRqELIWDktY0h5tlS40vpmpzpg0uUJBwiRowu/r+/ifBx1q31IRxy804M
YV6XQHdiXOozZPL7jQx/HwsAlirs349Z38pRXwnorrAFbm9ITtK1yHoaF9aJLYX9oyDEn549B0Uo
2PvfuitsiEMZz15aY/93ik0bPAw3wpseUOUzW1GXwEGw1cmnf4IdcB6su2wyCYiAPOwZ6Wd8gi+a
Awgj3xFysGmPVGEgdI/Unmpoq/yJ1HMsI/QCdKyQ2FWdFxy+QuhOzBjW/Gy/F+AszHh7T0l9I7hO
GQtiW98iNpU70myn/nkL9mcPUd8AqYq0+vsdvq5TNO/Q/uMewob/sMYRUe3nOljFeXUjOdusS+DM
tbYZXciLneVKgfcjJED2XZRg08PRg1kcH1oKHoJuh8eqEYGJyRHjlGblWd4xDLv5mSBuZYmkpOHc
m3LZkGxJwfAJ5BMbW1M1B+X0hvLwzM0iQ5Ibfah0FcEoyhSkh2y7VbZ6O6/lVXOIkkdZAfFvIh7W
/WEcixaVwdfpwis8KVmi8y+hf9BaVD3rKr4rYZh1QgXlBxkJZ/LgCWVlgw/nRtCLFDb9FlMdppzW
oFgvQ0Bm9NNyGqDzR4lgBKToq0dFJxkql0VCfyVZUJpJpPGllUUaWANn1YvVrgn2wSbAcKWSAip2
+Vwig58PzP9SU0NMQ95Z6xux9LMsTZqyjXy/TUpYMCEf3NBEy25s2bgCq8pZYUCD0vZE7Fkk5PE+
iPya6h1pN5hmecyXZmDte48GZmG75NFuETXkWW5ZTXJkdEWtNZwS7lsaSIHi6j5SzcvE345OF5Ko
9zhmWlEhvwIJlTPScs+vHVQL1cYJU1OcDFaEnjYcVcDum6oAxIXpah3PFfVCROve8vGRnJSa5hzK
sjTMrybWk63cBa5K8dVYVTX8ovp0wq9MN4JQv5XEQDUkFtNDDug71vbKLaw8nTAGSyCWB5/jJLR3
ecIyZD9z4zvXsX/uuy8QDCI2E0MUlOXRyyVqYaIrx56W1Z77jN2a9oq6hriiYIysHNWMVRiRuyi/
ePetexa74Kz2SYUSlyzi6hnx0gcsUOFEqDnkM0TisljhIvW7Ln+Fnhe1XhkRs91I+8n8jhRBqrp6
6w8VSY3ibYyGYv7tmQJsbCU1T+zdFcyvE+RiBs+ZfqVSzPOg3P3RulaSBKMOHCJO8/6qd5uNDNgB
/o20BwGuVPCrmzz6kOoCsnfpWCrpk7asWilVTsOrbCb8xwe9xmxS1KBWHF4m90fXGiyaPW5P0GXM
ioC5sqYS+BcDfD24wNOm53QQU/oEzmElfq0it2xn5i6Zbc1z9S/JmCINmnsPSPtFw4VFKta1WYku
YmQXbl8kEFEK6Mq03bZ/mIHEbo/ixaPqzajDOuRhv87SqF+cLxyfVxadHO4vqdUpv7iYCOa/NmVP
4XPgutXUXcEjrRIlMRd8bxZ6E+kF24i6qh8bOdQnTAxu4/jIIU/w93EWaoG+NSyFecIMvPv/6dLw
9VZrsEe2d27jD/p4gYAi9rhhTF2PEGOX9weOIQRPfUwyXJSusuHnR0OU9OC322yJz4rci2O75+hZ
13481xdGRmNm02fe2ygmRNaISFGY4lpn1DiX2lfL51iv8F13HGggRClBHiSw51KMKgRtBHVC0aCr
OFioEKEAyqu6bqWsjmQuotGtqA/KFPoQJ0DXimgEg+BGGPS9DXWB5o4KJISC3p0gAQoJgFGBxvPH
erWK0WgZHdCdVyujwyQgSEZKvnNUdywJ9fkX3nS56lH3hbQyewoly6GdziUUE6WM9NqaIJO4xPPJ
ealo2j08Tg9KVg76iKnNemaUc0LBHl3A/bpBbQ0PZl4s8xX9PMHdUXt16E8f7sDdT8nuHSYxWeZH
DAPWSyB0PH40CATS1wVOq15Jo65nwwAkduJRXRjWy8yGx639N/10MsMX/1iLm1U23tqivV5lWBV9
YScuKl4EWxZVbyJiXL8hDvoe3iPONsSvAX41m9Kd1YjlmeA8GmXBvK1ZioVdIHKaoj7HYEeDI1FQ
1PZ3a1r6s/5KiKykuLcO2zQdEMPfRkDtTetVQvCdkqZ1b/lXMoXgavQPEPvBKF+DoOSYXw8nxfJb
/ep4Pori+F7zBfO50+ajmZZFTseP5hwA+jY1l+V2e1hxt7sIOYpIqBbppypWgyP3Tggd/tKvuctR
HYQYfs6ue7bUIekW0ILimeD62I7rJgBweQrrovNvkLU0dJk2cJc9oJ6Wn9hPuZc1QTYBC2n9JHy4
Nt6RvLsw4/a85OZY5ISpR0mqSlvhPtbcQdrJJjXPnXFOrY0Ag31E2/tMmyUNhi52MNlPO+rHK4QZ
ahYfKjszY7AOMatPpWPieiubAXNFGFacTXBOfvwBxoVKjvE2gyrJrYIU7UVPyoSUfe7Jv4ubc2NX
tKpkQ7Jb2m/yUwQTNPyAGUSv7cyssateIQM2aTbmlJECT4EhgXxK9czKpy6Au+AfvFd4LMXhhBcN
jSmKIi5VS2nb+PezISnoKSt5qTcwsjIdCyGkScaBSCbmj6MDjhb2rwd2BgvBua/AAzMWwR7GZGQ8
S0JauwZoFPuPjUOIin2hvGpit3AkcxTeR6XYQ61DzwpWMqi2nqnyZhl/5YX+cjzamh8cWWfqdCNZ
lE1GhhEG+IHOoLZrdAbQNXfxmTLHf8Ads3LDn6CBOna9XSt7CjeOw5X6lGf6chMHVAhNBCFgGtpp
37VUAwCW/N9dkFIpzkKMyAgMvjWV6L/oCAqUN3pdRqSXyM/PPrLCSDyD40Q+XoxKqmpbLtWJp/5A
pKrIAuksmFmvXWUWZpnT2bKP3VCv6ILsx1SgX5+PqWOtekkS2fPFkg+I8cQyzL1Ch6+35LW9NXvz
lN21jwgzs0sth8RDr1cIEbrNzvOjg/O3IynuDDjs8yWsSfnvVshIpG++hAwysBdAYDKxeWhjwZ7R
aQHpRhE+qS3TsQ3SRQbLvus9MoOBEECFUAb21EgLEHV69nQl7KUG/W0KcAPUIYPca77uwunrO8GS
phtXL6yDlHjmvzNBtAb0EDVutjArErhlm3PiSy3/SVAhMbsncUL1cx+z/0jO+xVyqkbI1F/VcYxw
qpaV8BQsAJRquKcNGUl/jemyCqPS5OnW+bfO7P2Q4a4pES1Hkl5CM9dlQ4km9DUnepmmkJ81uoh4
AsTfCh1W7IIwuiMl+2OsyuUyEoj3vfu6hRu/9rFgF4WFlLqezYm/UPcdxSp0DIO2U/mOsily2gWx
GF0VcEx6A+WoG3rbMJwr857sbUjkx1gpKI1pg2+6Y20QJiFuN6nQGn9LNzab4NDdA8Pc4pl12tN8
6kmJxBuNN+QVi017siHhDjTOwutQM6qudUXDmJEndFZ4JfnPs4hTptKwNGSwgcorGQBY8qsQZ9Tz
cAWgDXLrG1a/scgSTVR6jnm1H29oUhrC0Fv/mkEN/LbJvHBI08CJMetccttCRXHVq75nILZrMlQH
l8FbIz/WkvIzV7jM1EVVuFYaSiwf5tnoYCHfKd/0nR5ilGGaL19kq37wx941uKjUtvZVaVGMrqO2
V48X8KdxBezuyvVUOrQotG0UwJ5Fn27b+Z2Ysl6cVY9oMqf4Q/GvxSqLb+md3ra5EOa0o+Niw4cU
lRYoYG4C/pyQdP2b0UkuDxq5huxZKZ+pAKlsbbGKIQ06wey33ZqjCwOngsHK6101INlz3FpSnQG8
P47gH8DXRXsHtL4KnmSUYkWN22vsRQ+Cu7I5AkrkCeBzm283x8KScdvR39ipzk4Vwlk+pNg7JXxA
3kGY5WPWZIOya/c9MEx3eIBlS6rbma7hf7NQN9+v73VNo4QDVLRFhepX7AmP+wWKKYIDICJPQ0xS
HBJW6ecgS+/CuipUwoPRdYjxxDOBdURJUwWjH9YcFOJ3femoDy3MP0lOEOavrfJC8sxxlGfTvcC4
DjLhZHGRy7GzouF75/jBqe10sIvjE7yLDCTR5dAyXwA3dzYLBXUhrpebKLzvqr4efBYZEXJrMP48
sYUfWez3XfVOTR5/NRBs91YRpY5uDHxH6uhOgGRP0rgbSFDoQqbmYQimUXMQ6BRywx9vSdgR8tI2
i5NHHeX1Zh4r2Rw+35RjHB8BCKDo2AyN+520u0DsJ55c3F5kgVP8OUtzwY21LKYYnr6lDZaiL7RT
0MPoT2hVhFGZtRiwTxY/XLHkiKbI9CdPkBjP6zg/nghxYJBYMCd2HmsnDruPTjaWyLkWo4G/EePW
u4TR/wkAhnelVJSb279etuAbkRAidY5Mvk5ZfewrI2OGPk6WsSHXfwHGGHKr1c7H9NAvLvPXhDLS
qtn5484zVsUILYqNKP3QRN2bbLAIt+1sDXfZKkQCKTCNYDkbcR8q2nNP/Umc9PFKLYNAF0xa7C9s
JZFfBD8Ss/ZaomM+6tfuo4kAXDQwFHFjZf3j3POeuqNG7acHHLCiNEXr9d2uye2F2s42kscSDV2R
9bkiXzHEl0GFzDD5cponJytF775AH1PtRqmIxSzPuwe0nsexDIVTIpW95po8rilJTp8CWUrkxdc7
PCkt5uaM5XiDX7GXW/xxsLK979X8RicaCd1xzpf04ZlhpN1M8eeZIniLhdUn9cplC1MOCjxka9bI
keiiI0moyf8/wGI0SIlJjJlq6KGzrc6gas/DchNZJ4DqrM6E3bSOl+pmBWsKIFIeO9kegoKeHekV
KbDpMfKYrVoInDFawd+rNPmoevi+NPMfIaFsD4DqTlSKrn5OEnGnua9u70PpuzM6nQRrYwwI0O4K
GfOIkicBMaXYsMDGx7QA30jcnsHlRmvJboHJU5Qle/B4EoiIBXMMtJxAqI8gKAcelF8tSnMAB4Mi
7WQ8Gjn6F7u+FE1+UWxjUZSWpJyyiIC89WSKqmfZ9Ly+8gwgpYEikmgra0OI0PmuZj6kMJd9Ig8j
AKCLLPMZpIg487F2X0fE9kJAjCxIw0ShwXjpAYFgHpqezTLRthzaMxL7H0nt+3VHqJ5VQlPCGvdq
HSL+QN1afKJ7tnHn9N0DqSBBmOfW69TtX0QHm1L3kDdHnG1w5MA8yAorx880W2AEMlvP3d9MbPWR
EaRqtfg4NuUONG3gPPM8QGnjz3nJEsCugMTMPoqfAzJ6OQmj+Y7+M8gxpTV2oh3oj1uT59eZHykA
S9Ae2OOCNIi5PAzBJL9lbFOhjBS7XsItDBSYtpptQCqBWqIt+w+hEYBh4YSLoX1m90IXbI2rGiS6
4xUthubDz1zdhnsD7YWbqvCD8gAYjYOgF04eKRoxSIUZrEQ9apIHxIr/kaYAQOBuziQp5dYPqnaM
P5sgkpiRkUZdFxMH4hL2nQ4gID6v7pz6G5VnC0rumpqPTTP7xkkwLqIxa3mqKPc04omjMYCGo5gL
fmCHcntiTqNyuwTPQXxwzuBTTrhN1UFFK3Ffa6wbDB2lgas/50l9xgNBqhBVDp6Mgn0qMsYuxf7x
2BIpZyGbLo/EqmZt3r8U7L7xYh+6c9klPLon3yF8sXsSYuAkiOT1Pp+IEDMXsDSZWkU8Mqamhx0g
h7oJJWVaw6Ahz4D60sBTChgNhMrUWGsF5iAJI3Lb/7SaSjdgck7M9McP6tgo5JBBFKu7g5u2kbCb
00HBOAQ9zpC0t8HrPp9rfr9EaLZkrYMO3zMs+4oiJS582Bp1TzDxCo7cXImPOEH4HZYnJ7/fRVtE
vS1PbF+vUikDcsNKIb2luywgReGuLgLFgcQV9iToPI3LqbNVBMT+dExpurw8wuA1cuQ4QUkfDzta
96hi7IQ+UcUAOF1PX5iyN1lOMIne+xBD+se3I6XJ9ZhZbVJMSWz3zb1LFJZaiKk4C8ZKVjiDgT8w
M2KcwzzF86oXbMjaa/5Ci9PLSTn+7XXTn7WAxUiG2h00SEK71xmIlWuo8f40U94uNqEOAGlHB+x5
ydR2eEYWqVP4OSmJSJYCd0yZ0tGUzA47NNFGaqNH3Bnk3oRw0lDy2s6Oe/+AP801Vqqs+Dviib2u
0QMcqN6lQgVk67lP7W/nNGqPLmxSjiKwLB0mj+S7UVuKjLiKUzUty9zWIyGFpf0TUpvMpjU528YU
Ggu3H/1V43P8UeQJD0RIbTYzzBPU2VFTFc8J1sBehauwTQrrwCJZI5b/9L5QIYmvH5J5zr4oytoI
y28ubcxCAYVN+zljHSQm+aMiG67ZIQGNIL/MN5WnhrnGnZ+ZheGYB1yZLgg/GN7qSlOLGjzy/u30
83zo2S49FiokbfUCWNm8dSrf1cPFCB7BLf1iPJFJTfSYrT5rDSpX4oR7UhOQ+UelF0KV5rLBPxOw
DxdevSDUmvzU9xKq7X9/bSnTUiv36/CMGwgJfsoWTZ6M2Yuz1us7CANsDLQ3Rv/YPYIsBM5fOVJB
pJ7W42a/kqkjQIt8Xyq+28OO0PgWz5jRR4ZtW4wPjREZHMbB2e0lluzqdtURU+Af2VGrHEGmG+f+
al8U3CLjDpBJ8uUxmoKSlqpkflZsztInYM7FZNo4fD48MsMbXHi2OTBkEv4VjTCCSMx84QWLHPRT
ZQI85L943LVG5WW5Mm6ilDmeL8oTtGIFoRxG+lLmLNC9yTFKkddYVTIa7xFzAhdyaD5qqAK+qYLB
2C4VNzP2BrhhnGXW1N/Bns7TtIdjauWmK9+en8fnAKjjn+zdUBzjtCYVobdTK788gdTjNl+0ihl3
5eH3dHDQqb3H/xoIjNLDqYdRNXJOiK7y+6c3Io4BgAZjW0EZo8BjYsQJTe47/uwCwj3SXcHZOxY6
A11uCI6mTPwPjsWTZmFnegWnF//3QW8lrtvhpW5yiDPJuQf3QgtIUt1UEdrh9viGC8mnburSaDVR
iCJUYsDzVxt9qMR6lph0trjFUs7x7W+KvOmAxADgKSXSdbgDOqiS0khMEfXzlCa8Y8H+oveLyqEv
SJTlgKvz18odsdpXsU0xL0Loyt0tzr70KRQHfxYS2In7IURcwVPhw4n9/Nh+CV40NjZO6nBm/nOs
Ogw+3U/oO16Uuqp/CZOxm2n0b+l8+hocZ+vfkbxh+A0YN6r1pKEzk7LLIPqXvfBi6VdOdm3PiAAO
9Mw2lsb2BmtnquSj9QgRFG55nm29jiTBrRDCDrmUlpOnKQnGGmbEalp1GGi1voJ/yFfQVHmiSYqs
rhFL7CMtjpCUPcD+OfRPHSBI2Ca7MU7E1t3sZc6fPAQHj+psDOFrPcwvMAx8qeevCtj+daRHQRbL
WU84bqh2XLt1xE+X3NtJK9Y8eIizNbc9AeZjnzGB2aRK29yBWBa3aSmUYdH8OwOFz3msSvkjAhZi
HsTz51NWzc3A5m2MZdP9RXsxt6LRbIhN5kK6Kpzo3bnsiqPyUs/w+IfD/3bHY3v8tZdaxrjDQJyy
OJDR84KFXK46mWbCnQCl1huBhu3sVorIXF/k4iIFA+Kt6njax/EpH6DHf1ck2Ocn/IASi+g5jfz5
SrFMEWdHsEJ7VIUYWTbknEtNuJX5WPUerp7W4RPsdf37uGckNiw8PwQt5kS9SmMP8Nic2qxG3bcg
41EWE7bVjWYwJZfhL3FYojVjwsrkocg2VFImqpirmhEWYzqk4nt8hF9w8qdKZDTZtQtk7i7i0OUx
p9FMPwXE8mGti3njZFTkQDR+Uvp4WCKK0OHi6ZrpHkxpJzwfy6WrxjK6uB3uDxl9GKpxZHvkOxYn
H4sQT5Q8bFwMv6HCVCkftJQQGPKkzFP9yherStCPhnVSRiBmK8LEw3S5c0TanJa7acU8rj6P8veM
vNc1sQ90EY9qyQaDcDdMjdqLP/92+h4EGlOoW3aOJXYJzo+chLfNJOeTT/pLggR+Y2oaMKnPx2y4
hjXWIjsiXVI6aQcYNjYLJ3gW/KKjVawM6iViZxYfT+JqE5k1UJ2Kb5Xz80Xt0s/siuLIc+kh8TGv
l6g5NIJo+Bzhyzfu/jecli2YabAl5LDkj+AAvM2pxbHzRPeZeKDEhC7fMFWARK10ndUQMt0y3zfA
C+4YkFElKPbf3eZPEITYyBewg+kDczLPZlXZTCH44Gtnf+w+CsXb3hmkvkJbMPdIiOZa+KkK4rpN
EOCGjiAsQAldj77vTXyj+z8IfOtv1w60OWh356ppJZOlhbtFNhMsNsfGAzRvinLbRpMddP4S5hHC
vYNVkUdJHK8y33RjOurj5fEk3oj2vdLNaIf5QxiKQC/gt3PGVIokYBHmEWcTK/zfj4CaBOZgNitA
OQXpAM6D1M4tgm0s0I7QivA83SuC2cyEyudN/oKzZMIS+3valGgW+hz9Qk309NuMw9X1ILfKLt7f
wPcogQyxnCwsc+0+k5ypvOlT8VN1YKaDyzOEmOQkA0HSE9kZxWon3k4CxS8MrJ44tJIRK+TRb/Lc
MdeuJuyjYnBpXSBtF0OmH10USjoZ42p36W0woR65aRRT4s4ddMstQLk45hTks6nG9/S7ogY0hEmr
uScv+EFwkrqVRtYtk0Q2+Afur4y+Gi6jXggAOHo2HFzBryLlBhkwbDZNtXODDboh37UkzQKzZo7n
JzncBD+rm1Z4/AfNYphHsEUkvm08YZTRRl3MDBZKBcw5W9mQ46VbwQ0R7y4jz3MMe5IRf7VfFcFa
DqMfnyMFdtbS8sTQdbKo/NeAqqKHdcAw3V0hd5FkroFh20Z5OXDW3ftzJQMyD36ilyPyo78CY1+u
GziJpad8UrhTVtoMGf/BnwEl/Sw1FhUNlHiJ1MM80UUW1ViWIOztDLPrrJuW7/t6orASU1IbJRNu
bjxRyerZLcJ1nCz5qMF7Ur6HPsw+Pwt1P6XpufIFAbFKOI8XUzi/+czZDN2/EHf2BMc7dDq1jvp1
TgTGM/2V/HqMJq14aNzvxz/J+zaev7jNacNXiYUKRI/qmoULT8r5yOoemKYNa+6xJH6M822tGZYt
0fGd/DlTHZroBCeA4NSU/EnrIM0KJEcKqcuVue+pBfCnuLY=
`pragma protect end_protected
