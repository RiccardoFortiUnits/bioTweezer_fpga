// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
UMRAXUBw3Syy3jQFl/N7jxUULGU0TtgJPU/JCvQsVxJ9lmQCnWj+Qce/GU8SYi1UrR8iwBYqv29y
UHEw3274yQ403+xgv3j7RYruxolj5U9iaMEgk3dHruS2DSP8aNdM/ZYaYpYXnrF8yW4GhHHdOooT
XWPa9JljEcsBf7uJb/p9psIyY2aq6yqBZCs3m7xcJndhEgte8kiNd65qB7AHIQvtU/6Y4WIXjP0+
KEQabxwhJPb6B6lth7IPDA3Taw3RNy/wENR2JiaH+i/cUBapqPqCJsXLowO9+LXqgsWwVaZ4qBGS
ApMweDNWCMWwrKJqUw/0ygv6W/H/nr/vmWCXyg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5760)
NF/rBWbFfMIw0c/DbkyB+UrooFJGSwZEGN2VN9ptZ+yb5ORUgscDmJULLAEEt7eUis5S12FdXvtj
Yq0WK+c9IYVnX/5ELd15Fe1xdoTNt5U5ypxFziii6uRZ4Wv0RIHsw6LZ8+fYNFx4ka8Nw+W1kI6y
rfLPV2xVx/S0QaN3PI/OaL/Vfh83C/rWs/o5Z0vC3YdfAWaoQpuQvavAW/7ENcjErhm8Psn3i0W4
ndaWrgb7y+356A0RN/iZEgfbFLNITyXu1Px5rNSkKCPnQ0cKkhSs+EMzDDmjk1rg+UzMFv5nhrTj
N5Y6YWC3zMtRAojsHAUD8XJSIK0Cy2QeQOsrdiM1U185SDJ6nZdnklM/GxTQ8WErNWRIgkgXSbBd
DTH5nMxVMRbN79X/b4NIiniULAEIAsqWJ6a45jZ9EyurXNjaOdkp9rE1MvkYH27HGuIyrJ5B3hW/
cyT5s80IPPsk6x1LV3Xr5kaRqeT594nVjXLE6EvyXGOXPhEEwwZBWDf/XgbH1W37Ajd5khRu+jxc
3Kzb0rr+wrKN2MURPa0yiCN4Rk1X4mOtAQtOzCLGC+lqi2G7Jqi8peyhAzXgNN2IQWu+RfujK3QC
gPIxZ36yAWZpMOitpqTtf568U9fdjzRhTtChI6kRZFZ+ZWl1AH4J97p+6+ToGhaHZAYpg1XYn6ge
8ll7arADGlVAKPEA44toPbAlWu3mN69D8pdVjtSaZKJVOWa6XU3hf5xDbNiOlXpadzkb9xIS56NS
OK+MUX5zgbCBYTh+0YQ3931zw8X/hPSj1v9LGHYrDRcrCdWgLjWpkO5kxyPGdIJ3qhFI93JoADfP
dbq5+GP9rW6VwqJa+BI19/QIMS7x/LmmnazaLSQ5l0bsY0o3rU6KXg8lSRrQcZFt9xWW9HrNnwzs
PGENKzHHjWZuv1x1o4xc2zFhlHVOax42QZ2FvV9wsXG2nGY6l75QbeinjYPhEwmwaMJO/d6seyce
FWGJaYKsp1AKEz3s4TmDf7mUkcH5pg+G1eG5G4APMNzyvGY4s/zjkwIq6DCNHNIbrH3akg4dxnBN
lEGW0qw4WWTJ2YV/ySOJhr41ugT4Loc382P98pDC+G+l9TxHJ0UQv5doE0hudvxE6QULJzj64vbV
2GhN1AHT6fdcrswl1hgbUshmx5o0zHHVUJr/Frgz9NPaHmkOm86Nbwa6c1AlS8SIhvRygwY0aJn5
5z97FP9teU80ju03cz4HhzCFFqYyCP+kOfc7XFFwhHs+zvqR0RtDg0gnotHHkxt3OnltdPlmGEGT
A5vfO2XwlVHS7/M00us06paqjo0wyylZ79orwyNJE793eAQhQmG7/dA9083stwla38tvaI/V9Xq5
F5dLMprfJqmf47IgyxMaE+85Exay+sFSI148qqm40hZjkazorwJRIjJZWnH0//cPVltY/DYnTa+Q
ZYwOlVDOMyPnjyywQ9trI3eASpxHCVJEkxCAsPTDZMLx/dZdt2Vzs59tnGM+kgAdRY/9HDGk87LA
dnQUb1oBlI0rIyF//vhhO9GJTTSNNp4wIPtQrhkwi9UZjBz2XXTqQJESs5ke2cz2NjuFeAlUYtny
341ISsMfMpZVne9RL3YfG48b5dBKmAU3nTl4XdgyWusmJQur96NDQ2ngwV0XaOXQsrS/058V6iNH
JebNdMUTt4m1zRvr+XVEtJO0/U9vXhv05EeRsKDs8+BLLRb9M+s+S5kYZ3XOnhDQ/UVrxQDQX4VA
dNcpV27vRDTVla0bq4RrM7LtvVAhJiGCbvzKCVlF9i/I6yhMP0iTi+U/v/OSWSryNOYMH1SPXMmD
ZhBSV5MdyIlKrxSgwEFVyhzyQoe631BIMzZEpAoBQPFvMXLu+vKorP/wJRXheEJEChlfWIDXMtr4
yVV2FmMS8cSQ83xu5sQlxZ6oo+/Sj4RhhuyqkAa99wI7XSZAnvdDKMzjz/mzL1AA+ZeCnEeDoT9h
cw3S4uU0LkrYiLIosbjI/6nkh+YMr3Y/cqeRMUqz0A5/f5xFbf2TLhmNgb5TZ5K5NRJfxY88Nmzb
A5AwjPcPKU+4dXsH62J84/SQ2itgo+VudBkxIQa9vimkkslY3cw9k/sm+iL6ECWp8gV0CYM4x8gL
k7xNY8s5xc/q9FJJ6Hu9bKPCXFNyrY+8FhfazRTpXRjdcbOKj0Gkl6qTy3BLeCYsuTfU3P5BYeUr
9b8dxt6E9dOf+aNLcWheuLCE/Bakv6sM3GfV6ZRxyPvgXXJVhIz9qO3GBpdSlzJP3zTEuUhuUpZS
d4VOd7yRKFIejW8KlYte/aHEwOO+HyKVZH0b1kFat4CKlpSfZiL9Qn21u/EeFMIPWknldkt48diX
EEhM73Wxx44zUq/Zh+Z/yqkAefZJcxJ7Px5OObYONXd09+QTLnQ4d87rR/wuxWSnUD5wl/WatPI6
Jrhw7dY3rfZCTkM0Je/lOmCdD2ZSswk0tsm8ukArujZHY9rWUkZKjUopdn8YsjcwwdgWMSnajh0J
fpz/M2N0BuHJDKLyirlo50Bpv41+hIfDlQxc06ZY1OxTJY11Nlk7YcIWj3EhiRKGhqiAcNpH44kS
Y6B0Vj+JRpaylez68chAzEANtftQDjKzzh6/ShHy4T8HT2Kic+RHSvh5fcvGf1spgjRonU3etaUx
cZmMJynZBbj35VuS5slPSUg6dgs7cHleh9+t+76TVlKuqJ4qKh4WR0hxpQEsr7otNCt3uUNoqd9R
BeidlT7MMAfJZ5x81yk4NRFQ4bcVrHMCUwTiKAxJCIwY5sfsnZfxBHov9YTLQ6J44ECzOEtnjg5E
cLnBhVKkJBGitqmD9vkR1jbHcNuZmYavF1634hmVKQUddP5QbtNfnouL5GwfL933QWeLy8d/padF
lC/EkVputA6edOZvYCs/46dEOUINKz4VMlrC4C7t8L4Hx5QQYW4umsgvyDCBTmtLakOO5sv+HWLR
Azfb77MkUQN7NFmr/AwBKn56GBiCHQScqycKqxTboxKoWdQJN+6BFAfGXizWGwASk8gl4Ch9q+In
ZGETRJMqiRUDAIRMTPyo2/qwf7xahH0RwuN5flAsC3+JYh9kdMcHb0XTSfoGEIsAud+CpuuPg41+
OQTNKcRS3VckZ+MD9/ZLspCDWufLLV2aVAvfJV3nM++lJsZiWubyFgRxXqe21Eww09mLilmcWdBO
X/zr6fBQ4W7YRDubJ3cm1Zo2wcHMwHEhLcKS8SVBydBtzfETutKxDJWnM+YrQ+wJAaPyNxrvA2Zc
BxnYOOaO3kBGAx5e30S9TbL9cmZDGhSUaowoG0hZ6m8WoNmdHF7vXXzYwWYoYat9ZmcTvBcA33v7
g/GiGITcv+uQ57WwSoAYVyzepjbJN+qm3LfbL/TiHIQ8hBYFKmHVbMhEloud4IqShEYKiGALhRyy
H5FgMNH06Y//Pw/cGgy4ltiM/ROUfzhaVAHYdIl7g2frogeKF2t5BpoF5gfnbn44JfqXXFhBwEI2
hdoh/kutWpVlx+v/nUq0n3GD4fEKSAGr2ll/db+HAOP5fmuwfyMXsUCFrpBHIUK17jgWLzRZXeLD
KEL/Tq6VzMZ7PmG9hAlHzcreX3HZC+WUDHd4KM111LQgdWtJzZZuj0L8uvTHUq5gWwq7B5vj/uz7
hjgC6rY/OKUgF4DgcackE66dfAFANWnJmVNGyF9X3UVmvaPprRLbpVXgDgWpVgTf7gafhbQ8/psG
CICL/9FKVC0GkiYgC0T+ACNxRNRBqVu0XkdYLchcCsSuLel+luyfbGcZPHCdYHmW0EwLJfq1co+k
X4qiKfhToEjbECJr0/D8dOMEBqSMU4h6t0ALFYwVC/OxrVIQcKcCtLErly9sw6nUhz/o4NwAot5M
3Y2FFzkKGDy3y7vHcD7tT6poum7tls071a6tdxoX2US09bE6ynSqe+y8mrr4Gg4bihUXgGwjWtzq
HQUP/wX3oPfQsexOwk/G9w1P6SK+YIqKKujl/E6Gb0aeVqpnQmAGrXx4CjX2LAZ9siIhzs9KvlTq
RNjFkpDOipyNIr/ij/YiIHo6K5r5ngnJSkM8aJ4R2mUecPi+/3UL9S4Kvxw2n200ONRi2whXnOJc
hxqIQT3LO9/m0yI855v8Ag3t9XZHjV5fQo7njgE4Wj7dkm405ZRVv17kpIvw97Wpv+yIqNz43Ncv
7rD1zQX5La1HUMQ0iljN0FutOCwHJxH42A41AuAakhycPzXHgMLw6I+xOVQ6lkfhsIEAbREQhPG5
prsv5JZru8Mv5BtAhK/I+OuBaEiqi+a0OdLamS3JxLB5BLgco+0asPRI+w+t4snNa0H3YghDONU0
dFtM4sFpCDsAZ/3q2xiiutYUKSSuyQbf4K46m/+gu+/+O2pz4KmBgdjn5VSCKGp4HG12CP6I+Qwc
sjy7PXn/bmVGCtQRf1ODHZHvIib3hL53WkBVifJZTGYHCfbjfSdbbNkkngzTNSnu/LTq+koJNMJ+
Yi/lzjFUiuU9XTRLgxS3dmGXKMGi6gRny7qLZ1skXMoY4Vvy+77bl+/CxWBLlaHr3Uzi/HvCBTy8
WC+fmNGITn+uo9lAZqfn2V+X/AOKiHvINa9wtErhcFN0wHnen5HnGy+sSLLO5x1LFPmz/B1LcRKa
LDcY6Dmm+x3VbMx8L8RisxAq4L4LNYgdaZZ74vm6H5+G81P+uAyWQNFDt8v6m0/m0Ur7zJkISOWt
7s6HHAxDu6z28FKiMCnn/nO+AO9O+ghMVDIlm66T1xSwUAXvudSVTb6XApGkGuQdtgZyIaIvVQ0A
KVpCEMQ4m8LP2ysj8qs2v5GoXYtZQISfSOPh32hgs8BiX5Qooowd/yOuwwm0SAI9dlDU69eXkbFp
kSVmddASQFoox/sEWn9jrRN79DBIlaPBtS90f7APmfywhICTfqBHVzFpC3Lw252BVkPi3h49nF2H
fewsF4aw8lBFhOV4kwWThBTEz3jjcBCl9l2cVHRUJ0A+hV51No4PGBqp4GKetgmUdF1inUnCBikk
94ceirYEJePvGs20TU9WGSAabx60Cimku/zJhJloJJv113ymdhDqaHfnhiWasqW6ckQ9R3cq1DQE
Tqbx1wb9cEcFxweflyEaLVN5tCd4O1DDk8PXcRUfk5uAQ8tC8ziRDyA1mlUa1lGZpR8UFqW7A5Tg
foGAXdlZV2VuKjmMBcLEy1QhZ3MBfdHyG8UtrXgWyfd8NR/mzVWxd8us8cPUtD8g5HG2awqQ2kyl
/geWXqGI9TTSWyloFG/jRXAHOUd3Go0ePuG+lfbR9Vv0X1GVZy19oL9ZuUAxFOUNmgwSXpXvJM6T
3EjcDapV9AaqcZo6B1Ot7BLvhPAlKM9/I4+2i0/4JMVzG/dKFMqaZqOKTKk51rE/1UMNAVsgx8mS
yrE5wegm+5jUo4Nn39D1zSsSgH3vTSwQTvVIcNjzThCuMYWLJrHoj26oEV+zgUfenEZZm2p5AyCq
3EBrIk24jgXlS5766XQWt6NTYZFEks+E8MY5Z7SoVOmvW1PZOsRO407xG8YXvdf4ndlnI/XN2wxF
HpmCW9QAk8lnPWiTNHjXOtXlTdsUrAMEF7cPsKYdzp2YK4VQxT+TylXea2VbVpk0vuhpbpSdMpfP
zRrYP2IC/Ientg6j/4r9xzM3zzkD2pV2lGnfNbjH/qzF2FyBVi2E6b7BV5JdRqGxwhYSbdnwqgpN
bhjNAPAalJRHixWkDq52SFUo4ZtcVKpUYhHpGzXUTflwJb8GjSZDKL8VMup32CiugFZiJbuZ6hLn
1n3jF0PEE/lmexXuUx+7EA0BtueQ8h4xHvosWbex/dTTI4B/uLjHcNHkMSygNN7AS1VxeYOC8AUr
2qtNM3srW6+eoDn4DJdVkziAT4q90kCJx3H9FC+O8k4OvvtU5MZFw0qbn46QNb1LsZO56kS+EIGm
R8RaufYAv5nF7XsRchVr+ChHgE6lBWGyfubn253x/gBm7xHaEEYF7aOTkaexnlbeTqg/v29R4Jmt
3QvO4lez0h6o2j7tQwIZPW1b2Gq9SfYBN4W/llCxkujdeOPGWKE9hmsStOhPVc3X8qxMrgzhPH0i
UHBniPrm1fRDKelNea8eowBMgILrbE6M+zs75UqxujaRG8byYfmURRP70FMCk1dEYQh4UmtuY67V
lKEEyV9GB15vTN+OqYtWFsQd1NP2w8Da4dNh8uy8jSm1Nwa1i6kVaC5IKrp/dUyLuOhKeCCaGvz2
eKx5HtCF+sJHGoc2kbnBT1Pk0ALp2bjrq3kn/QggX10Q/wjP4xRQwyKp3zeaVUZWhNilXOpXlsvg
rZwCJkCL0maOyq4v9/oUeVC/e1RD2YEAV2qBnzxeFQyfdC71obeYX5c/Wu1fX4VBNJA45MsK7rMG
g3Gxeo4WA6xAOA0rMwrg8vG4is8Ami6fo85L36XiWXFgdDEWNbaU/OPwCLMjeXLn+P//zczXHrtw
asXNqe3TVKtR07jEvmw1vsR8pzmVJ7Il5h0it0HqN+GZOyZDPar0NqyOgfBvUChj25ZqhJcV/e0h
tSOInnK/LyGhWDo++Ccr0RNgScJkIORaHbt1fwTUX8LXME+wosL9XVPAwbRK/VcH5SrdZQfpG8jq
qVtfzwsmKIdXT5TAddFh83+Mvb50SwLEqaOrtzmr2pwwKVfuBoRADFvbCgGosP9r2zEkhLOdrBFX
XMnNmPmeVtCzqPxnjzhc0IMb+MShOx0jlA4LAgGbMcS85HAekN7JLQEvs/5GjEhuRY7HlhIqsGaY
UZWXTv/5xy5Usj2uKZfnnTAdOiWA+LGnEWMrT4gTGfQxtj58H7WmDRtEj3Lni1WeHR9F55D6ktWo
NbmAQTCTVz92ULpjEUibE5Er4aQW3EozCEgSPWbvvF+ucUbgni1CxG2IhjGcNzec/3+z88O2tZN9
FNgn8ym08iRFYkQJDoOQZ1arDAF2LKHcXJyzLO4BIKBpdfNyECRzmk6TnHjM9vzcpLCdV2n1cup3
loTl1r3AjtMvAZ5THFIJaipxwc7qGUiIwFfyUFOYbIOOI6+zS5p+VRNMoj9Bs4dXhuN3A8iydT9g
/zCGIbSW/EdtBsCYHGRCMbzpKM3yO70coozBz/YCpSwCQq06gyj5nOzTCutFXOFCUqFRJNZMSwdz
yRrBUrRWXJckpiTq3RxwfE8ZDdlynwq6uHrrem5S3he0atsEPyjw2xF0IejE+TEkoHoap+imNolI
Do0px4Drp/u430Cw4/z3tf0LOShfZaMBqptDVP2GfDw5kHepA0vgUGsVEtcVou3CVlBsEQWZkuE5
rwi4XAV4GQ5P6Jidz/oWteVB9UYx8nmxIf5IrNhMdN1mnTm/nt2CUeZqu7AmCAEsjqUkEgkHcJyV
u+lh+P600Ps2J3QdbcdFmK+TUS7Sxo7lgbyFBcAwwYdIGY/S8t9jWds2r1/IpJuyDDiz2dZ2J+br
YvUxEU0ENDhUPMSlQd1A0oNneKkPrHwx9RH/oCDp+wxjzSc9Bd6OY4BpJ5jZmlLmQA2jH5V/zycQ
lathPpgV8F8A+OcbQGLw6WqNDLNwgz1YuIwvu+6CQCqzv4oQm5tWZyqFyBWAN0rWHiF74z8nC2ZM
VO6yWvhTGwgL6lgwbPNcuqPYDohEwZphPgKiUnPCZm8+6ME41YcpirG18LgyGNnMlbrMpLDapLC+
pCyJ
`pragma protect end_protected
