`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HZC1xkK9ACB9E0TP0BgdZ8drVzaTBRY14vA4HnWjTpW9Io1iD6Rx9LQInjdTD5Ew
TfXC/RtJz33MSP3gxGnXdY3EPa1h0VoAcmcYlSbfPTazAmw6NoC78sZ75QkMTpkb
272xYBSVBJJH0t3Mm/H/XM2aN2Yvg1VCJMlRlN3j9Vo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125456)
j+Md1mPd9VNG7z6YQARDZCcouGCwE6k7S9uybFFPUPf34OsHg04Kj4iveG9snDIs
BEeLednExmONdz2TNwbK9vs13VTMlBdMYOSp8ns2qKQvaNxytONLdvU6VAizI+0y
zQo973D7uX4qSfGxysyTXL5CVxuqjU3uNsMDCbB1+oa4I15NGdVn/Bk/xMwJaCTt
P/Osyrlz7ubnCABKs/+JVNneK6EI7JVC0K1BVv3tyTJCnt9AECyzxHxd/QhYbH9Q
OnjEWq3UYM0TrxEUn/pcJwa/YHurtbByN2dnwH9VcsvLfzuki0tRUPBwdJCSAkV3
khNvj7O9BbfBlTuVsCrBZR+EsZXzCYIgIDP2WXzsRKBF+lQKYbhbu3VWpUw7tcLa
SBXYCr9FeMBy6Sy/5k65iFuVNh2f57F/zYKXKYv2/6lBM/s/pWdTpHWELkx1tKdm
FPB5cXwbdJ7yt6QquWZzi6y6bTR1ekMrsyDXEJMuhKVCasBDuf78nkIbM4DqyTkl
CaKB1IWZBu5wr9BsPjTQmFWRxEFWk4Otlkz6FkbtPIPNxLZgmUd1XCBO//vKt3oN
W5IyaUMiKxy47v/XGT64Ri4PYT9hu7BRpHifd0L0Y6FXyhhoHrtezBj61PWbiQfN
rFAJ6W5HKSH6JzksHbvO3fNflcKJKC7d/4Ok2efCz0yWQAq4Kpw6DvYuobq2whgT
QORbCRZ1Kxf6AmQwf7ScnRqkEHvy9JcVCEmF289AysbAxM0Vdx+tlpqC/7/CMFan
bgAs75uPJ4YcsTthO6dgxU0BsnQ4apDjVlc7NcQ5xnkdUIV1faiN4Z1dNOg5XL8y
g6V5wieDGUj0N9PCp4Za9/lZxMPDtE7VQGeyJItz/kwOzEUOMZDL3ECcPSQpcIzy
sev8fYrtqRKl6L+lJ+u1PimCvVu+2gitXBUQltunRksTL+qktlZEDzbSNHcqFaFe
+DJdYbNiATEmVtVsqYFnAmREYwa/xVawHpNisRItdBJO9iwh9b2+aiaeGyR2GPYa
pPJKdj+B7RuNRciiYOoPlZG1SJ/UR9XNO5BSI6366J5DbGi0vXyxZMWZVitFsaf5
t20PhXNSYSke+6OzijblvM48IdjCoka2A6ejDlheIlZmh9hBSpS1f4j+56ZGYQS0
XQh+XAzMysM2cdMom7fqVKWgZj+5d46jXkmL4KI7WNbhEYoZBb7uGPOgnynDVxek
JfY0GdcwzEOxUYSTRvmuFNaL8frhzLo6IgJlfWoEpwRzDWi0AQEYDK1dKUPjtYXR
WlgZSQLiuI9URzXLl/6v+EsEKFI/pKbocxUyE0J8AZeMsttGtQkVThyKvfciGoK3
qVIjXSL1Fz3WED1DgzkRW8Ff+wPgG9VS9NdBrWpWrDWppeff3Es1HRUE/LDAIMhL
xaPHYSEDTKtzPcIyciXsxiCWCZQ+ZzmRnyvBZyu7cD877puNLxOqjDNu2ks4i9Su
eNK/A943nLjLttfgYxEJs5s/Inj7FIBoZaUmkERDeOUhH7X4UoPH1IbVjcUsspI5
A1HdZozLF9Y7QYEnwxK4qoiNi61eZRJKG0KCkC9ZpZtOgn55BBUgGc3JmVPbT4Wq
x4XWFxEYOe3jbLXL4GvAEo8bgJGNvSq/4ebtzrPuTWjXQ+dwOgIKSjm0xEpmbzHe
h7seOBx5anRVj13wzwa/JS+bDdBJCiSayHpphjUoJfR6RWYHsJDItxN6pFnUe8zK
sb0V/De1CISZpj5SN67g48dXJOaF/jNYCenzTNu/hSf/GT5w82/nD5Prw0QvZ0aI
sJ5gi0wQ45enyEWB5lH7vT5v4vBYbYjTGvQdT6cPggvaLyjfP6dsoyBu5sl6AFae
iLM82N0k5B0NBF2DduIo6dpzTNxvLaYN8CXiUAs2wYgNkTEKXUdnJAJ40rGs2Wy8
B6t6OWlHESTJIH0EXKrIla+Z2E6mA/VPichLlCM5Q23wxBvBQ2P+Sb+PsaHxe4oi
65VWoyvI+aFrqbY5DJJx+aobnl7Aw7OG41BIKfiuc1K6R3pi8xuVVZVIorv7pIi2
jwRMKv7tlgGOoI3TwyWGJSvMk5qSSiHTh+g4AYGajOWINojUTUZ39pmBiYYuGEot
M4yIn6maNrYaM+4TqIr5uyicfYtgF0beJN6qDXuiMNh7n4/9VvkKCSBcETktj+e0
D1e2ITRKrL51BD8Lqwl97EXvjFbppwtQMl/uYVn3cYI/y9VEDBERfgTvD7UaGOx7
DIWg0Rl8fMZIO8ZddzFz2QnHSethLy6MK5ScEtFCmva3FeyH1C0vKGXhJ3w+wHY+
AWqxQFV8FJH19Y3eBA60Akj7KIvR+O9FhFSweMO5zGu5djR0wyjqPXA27axfKLYX
jYL3dDi5OJI0+y+Ea3IlbbNbysQKijULwZCAL4i1V19dKCQsc2wYDe8x5wanW5xR
YGJ1j+aa8VlkfAd/5hGagn8ZpGvBBYIvWAUiqerq3LSH8pU2nmGGky/ODfagnZSb
XYE/D/dKZydfHvlqXgWEe8wyeGP7ty86P3SUqf8vyQF2c6weIRnUss1Vg7oKKprD
PXlAf1ua71Ly2/49+ShszEri4vIsHmNhEQfbdGcXVv/73jp5NMLt8oVPFLPbkten
lX/C4klqGIxspDOijvKDk9rx0NXI2nguJh/mQ5Bsf68ZUXrAW0TDr1a3t0KFYfEt
WxYGH/FcOipLXcHe0KomeZPFFZIc7J+NNXlXHzjxQb//AERHE2nzGHbJlLOM60Fc
Xqk9Th0mD8h8vueyjGGcjeEgfO1/vQEHji6HlyIzPGIvMjJQBFzdpxy8T6J2BXl1
dYziK4LwF09O80as/bqHUMM2TduEVMRevBD6xDGuGrYTVqjbr8Xkhzm057+xCbgT
vOQuTB8AzRdaN7wygQalC8oyT28E4AxqYiaau0OYVi8AjDQIi/4RjOTU0d21aT+J
NOVBj+zG6ii7Ndzn5A1fn3OKieiSLyksUNkrAFcufEReENk+Tg1g6XRZWnTT9F/x
mLLpFKQrdVyLsOL5B+H55nrr5Hxwi1neUZdTa5yd4jhQukJ6QuZYbE0CLfz11gXq
rYxVv1qO+/2kxUI9CCEyzDEHWstj33UCL5nIGPSk/fpGqqwkxZnv8sB1d39/GDkd
Z8x7JrJdisJ2dBlu8kq6yEYPbcguL4ZqgcqrUZ/abW5WY0gkXu1Eypa8JRwuTNpM
LA5w5QTdNq367yBRdEJ7GO4EQG4TtLdIWplcofDZC683+0pWEiietfgN7ZRYwCXB
tg4w0q110uJ6+At+k+4C+D6WG4v6xJZeXUR8GLCgwobYsXZehvYMQEIu+qvJnQq7
0X9NkTg+vFj4O51WL/kRwtD2MINe47cKNCJlq28bEmBvwbqGoUwEQ210Jk3GaKcN
bGdzcX3sA7Go8LBXSAASAFtv7Edgo0t6Hb/jZDnatokNefZYzBnhKJpRTDrwGfGN
iJfLfmi38pN2sx6aT25Udtgp+whSNO8pjtOxYkc606MevR4aSI9bOyK+ICox6eeJ
CCPj9woIu7ghfSxgYeKGU//SkHOLpFweE/D9sbtrdCj8agUBAOlgxHyLWlFz9poU
C9POgg8/uoEfA9yOhV34ETXKkBmz8RfpoXUBdU6OYa8O+3P1TLU7GF2yAThsg9jt
jN/vxhW3As7UUkUWoCG8DVuXSTC+O43mAb67DgTCZEguzFeBC7jciKhZux2a7hoy
eWOZ98i3iCPjGKKnI012AZKTiKXH35zoWT5Qf0EzpDatcHBx/k2u/YKY4Jfc6upw
5/2S1SHjB177H+cNN/8VIADqsXsVuUcQQ07I6zzPQJPGhuABRuKts9Y0vIQnjy+m
99/4aXsTcwvxkvcjh4WfA2amONsK+pC5ppUJDodX7JDlKXwC9lyOfhvBGeW9RhFE
OkMSqgjY5YkIoLsI6NQtKPzPixoYiNzt2JWNCfP2y2zEQ3XdaXP+DRQrQRwenA2W
3awK9fVcxhd03vxgFWZF1h8R95Iy+f+PPVvgswjHeDHconBVvbx6ZOk09QRizgs8
ZBJlya7jNZhPK50no0yn4Mqc1Z4rtnAUbzthHJAifbdbC6r8ccCU76BWOwDXsGam
D5CRPlXZ8t7SxSFBnch4LXS4Mxz/2vuXCJackqkuWF5g+Ec/uaKNf56vumk9/m2R
p5RpVgcbKR4+Y1i41SEDjvn+lldm1NPgUrEKuVCV2u2BKfs/oQsLbLEPmhVCjxzC
N2MkJ4Q+Woizzp43DBMsGAnnEAQS6R/eDpia5tmaOOQRgpFsF8CLvdr7CzYoaJtW
obdbP6U45n4Vh9BundbMaX6L8Yy+90ZER9TvewylNkeqm0mSshdAxksjEnNVBwbh
IPt7wPIUN9qLPKCN+VC/cojMtMxZEMOnSE7tzhGYJ98IdKVxCC8LdG8YctCb6V7v
tEaSjqZjLAB9piwaTKD4B/uPTxyvTSRt8F47oHSFn9K7vO052C3l7zHs9gxwTYkn
/oKp+g2JkurLYTE/gGQNbL1ZprGmGNThdC4mnFrsV/kVrwY/9HAa4zkTz4e0iTVV
V6Kt8cm4JIIWsd0cxaB0FG33LPN5refn8OgG+YsPBObUbK3YYi5zAi6dx7FXN3LH
ygErlazL8nkhMq1T/6fLWxvpu93AiYMp3CzNBJ2FUzH75EC5eBRNEevtsg/yxSXd
54XZdzmUctzajhCLFxMvFxVAxCDklvktWJo3RShhqmSC/MelSoY0EvXAJudihhjF
yZHhSjRMWR9acZ/SRGm6apoVoqSi2yjVBT2L9vwgtVp7/U2t6pCz7HcUngaGgEjL
OcVf0NlvjB1LRRgppUv5xwLjX8mT91+5W7nnjzn/aRSuyE6L4Y8aq8E3dCC1w+v7
pBe3mGsw8eapEJn7ZAcPi+XawPqa/DA611b1eULO6mEDySFYfno2dDB6f/CFTLMV
HdP33FqgP9DCE6oAbvkE8rH9scvNe2lWfoW4Hu7jRsMdv59OcMvinJspp8eCD4mD
XhbFGeNnr29KQbGjr7HqX2G4HzNjTLKGdOhR3boSoX6UCKsCNbBvLbcASyHHjWfm
dNoB0jRsew225Oz/EtCtr02aoQd4f+pepGsdU6NIUHonGr9EgJufAMO9pIzEf2dA
44N/Ed/8PghKFybNmuV/zn5vJAmw3O3M1qC/pmRyt2IJV9dnwyOmaadRG3LFyeEk
CFJ/0bKfMzUSGFGQItuI0/7gAYeIOGQYyk0V3TVmaywmcQp2XUvxGyBsR6Lr54TB
fT3TAn583UhXBvkf1+7jOI4pXBP1vyYy13+3HusPEtzMsxeU2OMyYF3euX8qKwOp
zcW07MT4ttn2OsSVkaOK9rkMdLgd9SNmivsF+9MjWnMLAGpy1nBxkgQMBpvWHuTp
xLQr1nStNjMC4cDoU9dUw3umxsuh/7h30yiwGLkSMy/lcvl1mV7GIMas2X6LMaED
sQeN57cNfHTrBByLv5dW2P+Icb7x2uoC1czhSaCND1Cu9arykYV5f4Lik9nMjW/G
4xqIxoAi6/3dD5ldZlCa+kvYLLQlLrxkHcGTLw0nH+swcVeqkfdEYmF90yHufv6c
260biUT1O/FEQG032ZC/0xRTtcM0Vjd0GEx6Liz++u4ryfKi0vKPLI05UrH0hGNe
48VRI0R37k10pBuisQ1DjCNLuOZeFbW3yUKNgGutdE0mE0rhjA2jRTozMCKsI5lo
ixpPWPdSAwNeD+R77mchkG8dP0SXU7z1j10YoKRDPRStVgm6aerxEQVvEvDfRUwA
JCBrZS5SV91A6+YVKK5WoJeo65DhDAoL5WA778HG9u1oFj0DB+nRt9lKTfjMyYvY
iGa/LoKkrLpu53+WatOSgSngFnoqz9MfMz4yB1A+/sqCVBkAYGXVASEN+OWgWbvt
pBreQEvSWAGH5Fj4v5y+lFX+DanPNb19P6CJJRLnyFpRXHjAbX1SSbFjk8n1v/hP
bMuJbQjQj4xwiNKOYwIPxMnzh4lDnRNhaZtZ0HeVSeGKL7DDwZgZTXGZ7ZyR4eLx
1y8vUMMO6eL0MFjcfAL5i691bag1hN9Y7g4+A53Ep5rvLVJJL7x50xnsMcEjY+45
rx85VzrFfuZ869oqm2jDNk8frGhULI1rjg135sSUSBSKHn6cjNoJ90VuJCuZwFuS
vKAEoNvBIxWj0mMQtTJvQYn5EmWp9GrhF7wp3Q0JOVDT5pFbhYeXVwCxADLPO1Ir
NPRqQeJdqgpBLiWivQccUK3fz1sfbXotH2iBd+h+rYb0iIRq22Ley7o5QxszFJQN
8VFlyE39+V3amJpvwwzraSli/zLdSRj8DieaFuh2z0++LsocQW/QZYs6mmhmQAEq
W64dhNhL88qXm+9iASzNAyJcy5KhYOLosAboRdE4fCFl3IukhOFlY7GYV43Mxx6k
OeGg4LzWCZ8pjsgDsdkT1nC+7bQhLjQydkD7sOWfg448ekfLWPeGuasNJjtZcMVQ
mDNkGuypCnu5lUEoIWKqXWrDqm9KMHOMfc8Z5HUeIZvaGz87Lo6Xi1qKTPsEKK4O
VwgIf/Y0iPkaYI9uAjErv7Qz/4ftNzFW8lOY4kc4gv59LHi5+9QD0iWWE3j+RAkv
FoBimJ7zp/2nclmNKkIqpmEpsEw9OozqX3JwAsPjVOeRqgpVHbenTGC44QCIZf6z
6YflU2Cha5PTgu7bNx+HUGk2Y14tlYR+mYnkZQlUg8HF1ZeuLt+IaNIOwZ3fF/GD
PeW3qtOdHoeFX1nJbopoZRjb3Vg6mM8iJtpIacAaE/CW+7NazIsNYVvzBXndaGld
G7FHh80hyeWnaKs/G7pJDftcaEszsT+jvaJ7qxpu7IONiRNeVNhXW+KseMISVHMW
OaqKpo7WfMVm6PGV6mGI+pielHtj1jrGVteP20YOVF6bTyT5AegFGBY7VG73M6O+
N7Zsp8LwTrfD8/BwZNVk6y0mLR2npbc437dyo8G4dWG2we1CWfg/1sdMZBjGNKhk
tzb121SVLXCsZrcQigkYGYlWeVZYoSScJk5KDd5VpIlwqgT3qQ4YHUEfEqin8Z9U
iHh0hPLxCiE4H+tqHVHsxVJj7GFaty/F84ri0a69aonBOMMr068m7UW/43kkpGpG
CK5fuMOUMNSVbcTBqXpODRq5NJpVGtN85C23zXZelZt3GEOcEF80lzdvsRuN4uuM
ntA5Ud6HlcIKKhDtCjTuh+uZcHXMubWKt7nLgpD/SRT3CTvPsbnqUEhBl01GvO/K
cBaRb+CtVEqki/WNEtZgthkf4SpDfzy11sxwiXgaDAAjo0RuIJQUqNfzfEi7iCfU
jgZXVZuVuBsIvxnYq7Rpxn0AyYujFZzt2gGQRidTmZ1hcqo+y9XD7gR/SJszlGeZ
N5qotqq+Vq5PnRX9myRiALY1KkUo0BLha0XmNo52IXZsop3gChEEm7S7cM6ozo6Y
nVIxJ8mPdqWkB2BgrrQw1tzZ4R5+XEtl1H8oikHans16Hcgp8oa7IpSKJ4+eZ9a8
I6mTf2gFZF5c7gfVbSubujuAvDl3ZWLMlBu1OX9UwHOkc1YlbiK0rB+SxbI1+5mU
QqYBfQnR4z0LR9lzh344vDo5EiROYgu3pBOnPWRRvuUIGX4bgn4ctRLuFhzC4Tzq
TNIz7H6+393fTrQ32y4m1Uy5noX+hRRI2/v59tIy49byH2mOjcShlNUx/ZUTMAFP
MAfBzU5we7Jx2yRHTdEp3hy++4/zd2AH6P4A9nYa7cn2bC+gJR6CIN/GF87gZ4vu
g5xCjWXe8Tu1+zYzDbr8ohX+VIA4V7T64tdSpFrKwM+sNa7fVaDROEbuwfV9MT8C
0+TSJxE56Qd69xx3OrHdXV9YKzNdBSGubFQ3kJNFrqz57tl1a620McaaO9ByHz26
KGRGaY7F71OoJVlP6uNmz3oh72lD3ooKGhCCvA74zuVKSKex9do1F3CeP6YEofLk
eBg0k6TYwjcNx4VlLaQAujkE2RYjJ4YbGPZxpvn9Uhjf4j907pQmqd/vCjMPP9+i
LvuuQIjDv0VKAKMo29gG7bYNVJSrYHh9ftHK1ecWCfYn8eT2HB4usyOFbCcFatqB
ST6xJn69GzdFJFgSqM0jakpZBcViqTxQUtm8IG5YV73vdm3oJNlzd/XFy+I2DfdK
FzYbl7+YA3YOer3tCXYwgXE3KKZR1p4AfViFZxYz1wtZKW/tHsw+M1B6qHGzBel/
krXgvR3mmVymrU4RJDK9hHhzgnjmEy6e9CDLGjzh7Ru/wteh6zxzd7gpd2prLcP2
h4l6yC/qGOZBwySv4BoWiESx3hyTtTnn57IulwI39Q2S6bO7OnuQKM+gUjUpCkph
bhSSh5R7hvPKf7P9HMaWHK/lRLyJcmXPPhOWj33nFO5n51g5k8RkVDRnnxfQirZ9
hbu/4F4EzmmqLaiayiYz9xTSsgiq8CRFf4jj3DXzUFI+yKJz6jKsqkMOwdXtpnIR
45Yi/Onbl+wftfJ5GVWTWSyvaOGRLUcbEigHDyEVZBk+UPkejlq9uT014Tz2VV6M
FfeEIgzb23mZQC39FcW7bSpyijuIM226QC80nhSsi2xvVaFPRK8iYcClz078n108
P0dJlL5WZD21nji6CfD6QUvlangeY2x8j5HO+oLP6L5oGJT2Q5uapku5AdrTkK9T
qvXqV3zHMtEHb2usRKQrO3CrL8uzW+PvHsOLltkse6kPWSxHDkpRkreCNQvB8asM
EC4DJXvoTr8f9U8A3mya412pqEcMdWpDHuzIOekDGDBEwhsAtT96IMgqJF09hYD7
WgmtKRzhSp0rRTVkCS+XCRAjhQAu9agoJUa5icphmr8hPmaS/i/AMdGzumTbnedP
rQGSoZw4JK3UvUNU9LuVeL0tTFaHEHl8Qph2tPhMg7Zra23+Mc2Kl4r21l94nIq1
aehgQT8JbTelqKwLyM8HRLZd4r5bckn/FwTloTyIaHnfOaaEvFpky7AJylDeDGCF
gf3teE6pJ5UIrIaTQWUIk+baro40kPs8YiTk4u+DnW3T8l4mcaEGr3mbGlitHrd+
4vzQR/2pyn0ZubGsMkN8F1zSgU6zaoyqB4l5ykKDR2IEDWblJhKvY6/E+mp4hxJ0
NPD8wDcniFX6vtpEQRFlpH4yvwfW6yMlQo9lRMLgrkyUyjv6Xl+RJSPgCOQpXDT3
ioQADSTiVjWe5AZbACB18i3zxSTeR98ikDD+nkNbddtZQ9WenWQRKt8EM3E/J9hQ
mEpdj+Gp47bjsjjbXYEIhWxQm/CNIQTgzmUEYEMtrwVdR0E4nHgrzCsZMQG9n22r
7aclvv1NJJsU9SGX3g42UUPAXfNc5FcXqabVWKVczmDo1n289olyw8DPmYUsvYFA
b6VvJkQnthdYoNbRUU0zxPLYSQJK9qgbwa9dmKNtzd8hD0HPWyHm+S/62cTC1gbF
XjqXzZNwnPteIW84vEXFpVOkssWG3KFyN9snhRoK9CH0SVlHkb3IBIVvIRy+MawT
QCt/iZo3R4FZSAb8Ltx6hIlMzilOytwTM1EYp318LIsB4NtWZPv5Xkrk1jeVYvVi
IbN4xYdck3UQBp1b3mURGGCCSJdZth4TC5P1QALtZNxjctJ19Ltmqu6qQ+DTDNMP
uhBfDjFjUHzSD1a2nFzMUEA7LAMPQ5bGLx/voh72yUpWkNL/dqZMbKeEdAeuqrdP
ckidTfEnPROc2Ga82kiG2GTlXHXHMqmlDL1WmUY3gpwkOArrM6yoRWgG7xufzN9A
aCIrtKTb5qFKQ3fhtN/syj/5yO435V9xEGcPPjzFhhnIkfTUEmSVLQLCtGUotv9i
A35WyzU3sCELlMiAWL5U3R94B2xV1Ng4RkMNedv5aYIU0YmEArv637q48oPdBSz+
fB3KDr073RJNhC8xTvbXNpNLTh41d77PZP4bTByksHcw1d0kfaXIWNv6vRF7zPoJ
Wfa+a3K9XZ7HDyTk59z56vZsYyC5KfqrJHdd5WpnXA1sb6Po0sFU+V+QxUqmCh2u
Gg/qg0GBzJ2zq/7aHLFcmXJJQxMXyId9PXEKg+OUt4yBW+HUper+6nzg0Objuy5u
9rJ4c3WFMaFkf4P9mzPUy5JA7fLM660lVt6u4CEPIayePGTDx2rKoGDMDMF6vh+7
EzGuruTQRVXoyAWUgUuwHxX4A9FkQ2AdvsWqRKsCmvRyLHXOZ3J7AIGaI/lflph1
pO3jRy5FNkp93A0Q29IRcYDgFaSk6l+worBI5eoWumsmu3ZPqBTcqUZ17HOrZ62i
5ba9DlFRv9NgQ0GQasGl5ybdrTyF7CyfKZSV5o038VenS8js3i+NKJ84fJ+wIkD+
c18mYxqLTtVtT5dHpV146/419E2royoqeNrCUgxt+kFBpJdVqgqOPFIfWtu3SeRg
QaA5Pxh3jmk6zRDoVL2AmJ64ch9RL+wS24LQiFKRn0kxdJReFugoSgi53cJ8pNTP
rb12DjizIaZDOlN8XYr57Sw96EjnRx56NpZIuWjkmiKDDtFi8EmfXPvu6LHTF3ye
h4hnsit3NM5lZ/lElfDR9H52d2N3wDBmaKPdtiWu2Gh876q2uVJuh9ZB7S+vB8Z9
WxHTA1XW5/UwC7Gla9YWHiUET9v/wsOJtllk0QZgZVj5c0/XBw2wbOERPRHADDtH
AI6PLXcvR/MzLPkUzX23bSUGjL3/1iiDyc20rxOT7Gg4+af6cUTefPpinkeZCczt
qaoo/UKClkdoVdLsYQgsyTMr3yZPzzpq6iXkS7ol4P7rVb4/U/mMGne/jRfE9DIA
8ndJWkWQmPxnbDbnW4jxmE/1D833hn0VbwwZIu7CZWvnp4TfRh6rEIr5Rcoq8upp
TOC0gUhZSnW8UK5Uz+W376ECCD0ygk3t7O3LavLF++Yt42sa3t2HnXZsj5Drwolh
LaFfma4zwJECfkjsGg7751kZ/mi4Urr9qW143I8GYrWV215Md2Bt3Xme2yrteVrh
GjGRAaYXVBJKbrJPMFs7OXbQBn/XBcZ9fyJZ8fIWzZQ1cg23cjhX14isHo2hQAHZ
FPyd2INFcc+OH4RlGDglW1+hFP/Pxjmo2PV0WyykY60XEn6S7U39+HP2zgA8Yb4a
NOOrMpSTvbRGpswHkxE2IPnO1Mb8ZrdFSP7gKvP7pk8GGZ9FCoGdtJ+Rtsd1E/rL
kLvMInTvZbisdm+/+v9/ZLvj7EA+/7RJD9ZE5jRkDeDoEEGcJ6MMkoOEu/Mfs3P0
NTpqcC1O2UbBBHk/Aa0cjrlPkch77t/SGlKnl54Lbb4DA2fSHaBYoLFy6U4vapit
02oHVmMS2bHrvWfCC98+5wqGrauEp1CO9ltcoN9Fj6Xn1VDPnxS4uNMoKRRZeUhY
z6x4FO0oq5DagfYDYw3z+Ua9u8IdhghtRebCM40jeNwBmPeBWf7nKKi1nxOzt1U7
Twizdh/gDGKQ1pPyw6FEn7sMudiTkbLgCB3GK/3K1n/TdA28MyRzbDkfSyf0qdPp
QWxcbPZ7+xkoAvKOHNX3Xn11lajrfsMN9OOHr9b4H2D/fJfQtUsa/auz9sTGGRCz
05KDVPSPijjI9E4hTg8ve97H50TxXr3wexqmyxciMKOmQfAmgF00CPmwLaR+APIK
g6Y2RI6jBtADSJi1o67XnbU34eJ1joC+T5KHSas2jG4hcvu909wZnuqquU0+jdws
IOqDpF0SeS0YGnQzCO/kWUNt411qFRLL9oOdCRvJLmA9cKEBqERV/BGMH+ProNro
3+p4+kce5r//4poa/eHoVXdFyXdeygxJIRadeMJyiOL6+IMgRAEZRW1MdoW+4Dg5
z9xOtaFitCuB4YqTq1Sw4Rs9e6OiaMMeB8u/9Dv0IrEYGEFIMVH9658x1LVJ3HZm
goEVWTQsu2E19JvFRBMNdxrTfpBWRQIcFCwdPrXGwmIj721l1ZHTrNUkwYUCnGiq
K2Iqd+BHvzxvPWFenZjk1I3Y6pPuYYMibTdzOAv8oqxVACrn2prRpt+Z80wanPUt
NIJMEpy2di5C1B5xBOwnKiJpKAKrude2FK8Y/yLXkTpnlTk64PmfkOOI+kuGG5ex
6qXw7XVIBnr8HPKtN0yoqj7jA8cRXIZnE2OIpU46k+Z7CgbgsB4BGA4oR5c0/vj+
hEvrj5s8FaqE1PQcOfm8HWPEidBZaaWSTlinskaPTkZrAFjdVK0ivoYp/ZYHxZwB
A97QDpbcuqDAKO4TCeQ8wEBTn3jFpMFTWAwph3mLvFQbTkcs3hW5EQAAt2tFbRpo
IRxQgPAe566H21kWzN7U91Uj+Bd885DbVEjbZUgTVH8c/yGEF327xxgTsG1XRswE
lQP/+K4682MHP6WdG5ZZTMDhMx1ooeHIemzd1NOJ485qedXxMxdvFJ/3bPwK4Jom
GqeVyeSDNMt3dsoMzgPp30fLoTbz/EcerdWLSbSiKFRInpCKxQ+1uulbl4L6MmzN
Ltcifv4r5jwqTqpGfTuaCQ9xAe5m0rN4rsN8ibzjsVd3Fqs9eIckPnv+DSnX9BbL
WKEmGHjWhCKB88bEUzPol8g+UJ+mvA/9J537ZoJayazcldZOQ2w+Gkh99brvJQVi
JK3R43lmPoP7LPZavaoefsf6W/ot+RZNmeuKBQLlM/IJR/YfDxPsfCXO51Js3wq4
azNhHKSe/cxY1aTb2KeFSxl6N08xbyOnRZRVJqDsj39vubYC1pQImwv6U07QO7bt
VPFre+ThyOFmkmS6asfIokFcAQofs54YUYAfcrOc60tu41uq27CzT+2py/ZmXv34
Qo42q5Oeq4J5xzDxYvAJG01ypRyP22zBxOZivirPBq6dQHMNGZL+Xp6wCiG8bVUm
jGM2tWeXEQHe3cOCfsBqbtgOxpNE2Yc+i8vzE7s9QujrW6HXpDrNg/cpWuPvujT4
SCIZCHqdkiaSCPlXPytMY7KEHcZZsU0ToyBhfwuc1XlCRqBo8y8E4jALUXDQxOr9
RHDDmpZpHdP41EP3eXiBGr9zGSKJzqmV+MSeYczvKSuC+NR7vDbjWiozuGN/Ilaf
hTFsdcOdLBEg6uzXlLvdn+xNzVLYetUUOm8V2sXCbE36ctVrDai1g3gmg3TQhDRg
uQ+Qqm4fYimPejsSmgZEJHiuio/JavXagzQA+//sHSJp8mrZHN0WFeZVKg00HNSu
6Xlx9xEW/yDfuTybO7A3LZT8I9DIa2nUvAGsp/dD3t8D9pcOeuulMS/ZR4gtK7na
NNBwwVdEdsYNqvW2t4u10iA/gRKud4P8Xq9IAihPQoNNlfoCgKdSMdnd92zE355x
nksYKVYdnoIHVXzF+WyqddWv00rq0UlWu3xVnqGTfMUGcs2BTUhBdV0R77kXlIM/
ZuxSwHoa51/rPi/Z/0WLs+70NmuoJ9YYTZfNwCxjkkTotOcKjUW/jlAJhQumMUwG
gdEE3gMaWyqeVkPKnqoQor3V7rKtCE/tgAWIEy1ewG+Hafu+dDYJFtZHqlfyNe51
YwO6XM8UJFrxFc/+2hnBc033p6nhfu3aHg+WYRMEPeXgpfbKnQ1/2tjnLZTJKJJL
QUNAYiECwAisMhABdO3vqJwcGyRaDkHa8y5jOhfMbpIi4Q3a9g6wO3xT3AheCZ+W
FaLVvexeg4uHCd7MQchk2CMaExo8HKlFp5GaUko01U0RUrig+GoBUeUnFuZnXRYd
AIARg3oxDfEuBQk5vm4jC6vaGoT7uA/4VrjazZH3uU0hmJL8o0gXGLvNnyCB+KLQ
KPcEf+4kwwO6B0ZLFms/LkPXJ+tqnT482xOnwx9UcceNLdlJ74kB78JDRcxIQSNZ
pzetaZgjBHnARXTMcTbW4P2pt25Haq1EPW9/nQCA3lIzDYN8zJQmoSpoX/GzyERR
6GrYy6HlZWME3y29grUu6uzCGksN2YcN3AzhsAlYXJRSZzogn9FC8W0wuUD/ovrJ
KY1aGZxyVky43Z5tHTbzSdGQatEUCrH6TPjBZHGpcRKugr9koA6XTDWbt662aHir
L27Xni541W7XDRcqQKjmtg7MQJXuckb7ysqy32xZCjGEZca5NCm4ysuaMJWhyZOS
nkxftt5woAYJyPd3XAS6ETgfNoMNnuG7EFk9rsjo+CdpdRoqBXVBi686+B0YqtSf
AnSl9wKG4U9ilh4/QIH+UyCZmRlwtcmv8VtZd4yKF2w2Jo/eU1D8n+X9QcXodlee
Pn4GkN+A7O/wI/mraQG11YidT00tbiYJJfJKS0ZDH0SRneph1ByZZWp1QA6H5xDW
BFZMIOajXzW2+p0F6/SZEIlTGE3iu8yXWb7bkwpy6ko4LMzAoulRRAXy0Bpkby37
xyF3PViQlNt2aSxky2QIFiI1NaWHKWgF6CIZJXaiK1kLUWsXMoutWTPkbTq1J/iQ
Lwax7FM+PfGB2mIv3djBaYjvrnldVaERyUyryOH398zBtAwCJfoal5j5z/zm8TE5
cWe6f7gMQW+O52IkYdNkpV61GmWXI07h3yph0wTJUHpLdNQpumVoVQ/QhN7TO57s
5XhAEi8rEzrJslrKmaUM44Nlqm3dHzBRrhaACGG3YqZOuh+/fm5S2mJG7cqIrjWZ
x4llLXl4swkV+cQ1eOP+UYyqyQBRbcew/PBj8QNHg5sEPfvf90XHoCy1Cnn0K+He
G0GpdiS1XKfLA20Mbvw90Rat95h9Ku10y71a5LciG3xo0UN3nBqR/PLfqAtM8LBk
OdAezIxk6pLdO+YWrtit8YInauvTzQgEmflWb+RSk6VieonGfFr4+VhogiGmmkVg
5vjE7oYGLw/hbSdKKm3sG7wSi/mXL55WV9XY1a/69k9YrOxuIwsVOsNdOYlYIppP
bbffDzVkgVULOmXVY4mHVBBteL99UHG8b/BBJ31j0wqQZ9ABYA6JvqV2n8nCRERY
Gs0Kpx57DMx+7u17mPI9sKvPgdYfx9EogbM/C7Hvjv0XxiVEswZjgNIuHCRE0krd
0rsJamc81AVPnSbu5LPp92M8AQfvfFJ81Mbe2t3MS87IMadH20MJPv4W4O8SPNzY
b+lCOwwN48sNWwFkRSiSEkkT/CoMy6zw0OVVeYKXuh0GqzgMUbHot2AvabNadkCs
tymRKOlrJvaHis2DvR5XPHo9kw3pClsyHNhW3/gQr1Rg/Opf7rjo04Qz4I2omdXP
pq6UyUBnAM3zEstP5o7MmyKcV8BbjAaSTMF8bXrffpcgJz2dxfO8xkEqqLYRnJkY
oMWEkaIve4eJjdnMD+hmNVTLAf9yEQWFoVI4vAcrp0cO3jFnGR3QN7GUDhOaEBKU
XwZs9IGeiakDeiFoQG9pFy4RMI11HQTNGbW1QYFt8LNkyWv9hU2G8GYsrFceAhE9
fsv2tF4uXzoJYA2YXXpvRFp5DUQHZXKxtAjdO2sszOjwjMTnkY2PBnz5j0WWd37x
zTNJMgmr17b9RhQizzBxg9g6BPAgWwtJZzafZxmxp0KRmb/DFWR2emLstCulCYB2
lqgwyQeSk6yiEgwqfhf3VtuJtXVYbuhVDKWqX8tFKKAWf4noEjmYdBMxpomPg4Yp
/aCKrqSbmPPUGis0KZmWYNek7n7hSO/YQLxG0jQ5Hom3vj+mDJU6aw3j66oJ75Bz
eF5lQlCsLiKl933WoKaxZyd7m3HQKYGL+oXgXwoYw5nA4lzf9t2goDgEl4WKpyGB
egvBLSPyR5kOQvUpLiQuhA1ELYxBLWLiYzyNlmxJZRUfs4Bup3lqhB+YVlPWiay+
VZF40tDoz0W47XiD4YgaU2mZMTh9BbAU8rnH3KZKB+gxtBgMpEf07OWC8eLqmM18
rr4FdilISptlCkAUfKMPQxTJePujYrHY7r5kgUz7nbqx1COWJDIMgV/TfBK7+s88
t20nHz4Z8Moc8kKAyUxi3JMW1tJVMi/HidSAFoLxnNDIV85uk4Mzb31055ewmwXY
d9jq6iueFXETabwInhOIQ4eDA6u7ikRDVVGW1kg4uW6cEcpAg9ODEXg56fsh9W32
8KSvJ3D5cgL6tVFvG9cXx7bWt0r0B2fWRaaYLR/6KllqGoRbDMV/KMB2JokwGelQ
CkZ1cI3h1XX/cG+V7YuRsnEWUba2w6+hAIbwECLEWZn7XdKOkL6G/zmo1kvKv+ib
doBPcD2f6P+S9FsrjB85pwYXKafSH4zoD23T0jqq/sePVvCImoJeP3br0iBqOyw/
FuEDCIoJIsGhppLPs3KRTSJDvqrjcbp/tmThOdykOK6np13UdDqTVGmrVfnHtEui
a+L97yBw5nuUn4Q3huAyDA10fMu3wYgGH+5KzS+MLnafImQOloPHwnpleKABYB6S
71lvaVb9P4u3d5kgckqODzfLogfiqlFBqbLkk0Wj/Gjov5LJUdDE8r6Z/Smnzpbs
gP2Krptg1AyQ+WXsvoAVMc+qrHwUlOiWjswh8m8WXTjRB1Q5wHhCSHdzS0x8K7FR
4eqtzbMZPxlLZ+XH3QrFxcNogiTPwKFcoZDpIDIci/sWY/NurUAQXlJuSyQg6v40
bCAl5/0wBf/I7xHZ/kz/lkrg/d/3NkfKWzgWl1x9uP8UzpxbHeqc+WQWj38x98fl
9R5v6U0IrrkNCJhttw+jrq1wd3Jf2c4ndN85XiPLKp/pcGv4BhzjnrWf8Dpsqf0V
A3wfZWdQwKZ7E9rVCJaD6bqjuY05Wyelmg5ly8cAtlH9ihxppZkFWqUcnWXuiWdT
oZ2aXH0rm5RbNQcxyGIJcWw8K2r1HExpTbOAmdbrBG1yKfFdHtu7AB4DuG7tpVEq
QG5DgM84veDMBpj7lRl5gC4TVmryj3h65UjmBAVFUgz5ShE0GwNlLpf3qEIBkZON
afiBW1VjxPy1ZjjdbpxgjbCgirBXmWcqH54RsKA2fKCHASX+EJQXKvzGOSdkI/O3
43g8qo40wmFoDCfs3W2L0N/yUUhEFSMpekGnMYrv7Tl6DFEj3R3se6LC17QP9ceq
oCuEYHKx4pkArxpixFprFqIAOEpYN05yxzyJwqZIQ9oLvT86TcV5qiCtmpP/Mkqp
k9g+NxZg3UxoRKV1YvTn5IWHj3KVNIi6hP7lnikIgYrx8fOLkX6VtqJ9MweVSrGk
X1F56+944j08hTgYvyeeoedUOdcNhFkNV4jsHNjC0yKotO89P5yLINK/9nevo4qt
A1Cl/mLh4cwBlAUL06o05u71dQFpRiCskpWzQ991Qzq8n0ntg1L2Ca0Mr2V0j0kf
ufH5rdwWraNcBNK62wWORCCQ1Fj6FWa7cJdAdzHRKFlkYGMnP+A3rmbDs4FVgI5I
KSBWzo3rFUzW4NAx+BZlViAY6UevuHac5yKb5omvCHApdKJGWkzSUkmU+oWwe+BL
kkOUdjl5QQhU8EZFais5jICZH2T1IHsJqekM8TECS7L9aVg+cTLcHTB0Jsp/lxGY
LkS/p3z2yNHk/KAGhO6slCzzYN0RV7Sr6YaiXmkM612zIFkHgRuoAM5ODOSYuExr
Us/XcCj6g9QHyoFPss9BtrVhQzPz1ZcJrNd+6yMOx+EF0erhZrwYybgtkwOXH5ac
tqFkNHIqVnIycnCb2zcbsz9ULC586bnJAEnrMBuMtMuekY+LcWo5UiUP2vJYrPWv
2YdK9gLVAyo1VpuzwG3jwso/gx4NfAOSExMkVTbV7TC0Tnifufdy88nfrLhS09gh
fc0Qbq2E+GyeUqy891braLugYI/DIgh5FiPHWIIySjMbcjNbriM7rxNkoVfDAoNW
sOTBe6/akU5OkiLo1ebUBNIGIYzyonnmP81lTXYplUN3khs54dlUc3oZSX/PkP+/
MBTodFMkdg8DvzFlOZaaVkb/IINIe+1NtAn+AP/2CAI5HWZBeSkJJIoPT7BMIkcO
x67ktQEKaLb0i67/moCDlTMbRQW6T9ge9UyB2WRFR0uf5NHExdbieELsjP3xWBUy
jxcN4kHrc4y4DA9jyMLzdAybU/vfu0uZydzEEcfJnPnCWapMJgwpdk4zn58P30EX
eSrj232ZzO8xgWeICSx1CYi8S7KwFJPcT2EdmB0JJpaYS/xniK/K8Nisq75wC451
FBs/2svF1CIrtqnMl/VIkI8OSRVS+P2Oye5v5UluusvmLAT+zzGD/nGYchVew9D2
/vvuQ+IM3EtqsdsQAmHJyPrSnopaKEPrNws11khtH3/r7QnqyanRMuNZb9Zcxpvt
mbGGa0XGuXhMo3S0iNnZ6NtVIYtwY7SiUgZ8Rv4sK5n9O1J/n4HOWijToniD+NmU
njo8LBO481C7YkaLjfmW+ODzbn0hbxOgPhR5fwK11cencDZO0XfJ5EfGq9zqBk33
yUfgvs0htu+lquEnB3U2jPjiAXxKBPDUyXkCwwp2thl96RbkLX0cMPJ1t7p8rCor
DeGdmIwFkO9QTGJRdLv1esmbkFz11YkwbUccF3ctkO1shCu/zX5TVta4XbkyyEuy
wgd8yxA4FuJID3ZrAYC2TnBC5JHqhjYTGivE7HsGM60d2qXUF7YtYneQ2al/4kBI
Agm0Lok19Xny4EbY/gRIEbLlrtwXemiP+3Yq8Es+PZH8ZfFQPUiRiU+k6mG3IIV1
2NxzXhtz+fmrWbDXj0QnmFIRkzy5Pr6oIICvaE0+uVvo1iBYomtCeH2v5qSzUfJI
iO1HeuaQRlyo6/Ne0c2gutuRmPfaFYmdletXIS6ihDwXirW/boSByIYLZ2I/LOpZ
ZMd+wlzCbxHOUN6MRx6Ey3Zgu+FUIH3tjr0CIGQmYmerB5SeRmUZspbzyDUWsvEv
qvCiEe5fGTwJ3tBlYWIFzMMsAvFd7doOExrwY3qgI1eSF26CdCk4yaXIOc9B2s6K
NWQD8Tnz3Dbms/k1eq3MgKz2bJ7i1hNI8I4JFN1xpUUkT3HEiCrGVS8y8x9Ian5i
xPzY//jMS2FiT3hrf+QC1V5c6Ph6JKtYNz0nvk6cr9I+TatBu+qfQMLUIn5Uzp6z
4ljjb228CYxVFo1JC9Q1SYp4Wqrwm9Et5YITgrK589wAU3xFiU6JsjA+7OPn4sch
HoM2IEk9OxA2STbwHVwIPGFnFDYv25gsILhOVgEOUMEoTs0Rwn11ujAka3jM7QOn
mVYGHBwSPADiUTrSlE4Svaco35FYH1QlJXiiPmzXdv+7Qq8wmGX5yOyp5UyhIYv9
FG/Pw6ZKBBy6QJEUfT7prjxPj1xEYKCgqhc+bqojMj0ep2VojCGWz5V8S/3fTCBQ
v+CKIRV2Gzx0iwIjcOaSlvHsSZF3PWVHFQOmwmOFFtAxeThvYxe0iJx7QdHIjgik
l0OGFsHAePM/DZaPeRLYuNc6ntrtVzSoXmov9AvM1VZUUarxi5votg3KNLZlM1wa
+G2wyUrc4pKrlYpXN5/0agy7WucDs/4N6ZL21BoTh8E/Lr+NYpbpJT9MH9b0C0Tl
tdNYpJnDdrI+eyfhtSHX6/SyNzP5iTfcyymaa04JEaKO/gowZbzD8/snQ8l95sC6
rUXfhpnsojV0x4tHhASt5hrtOg1WqroE/rnpAbeHP7Mz0D+mAwL0VXEpK8025Txj
WbLrpHCgRpOKdCRW96PxCh+2AgZeOnekhlP46FFascM/DQR1rkg+fPPHnncyK22v
xHoyQ1kPKwCYdDIeqLV1LvlPs34rGskFtLq64k5ymHXh+CbFH0gKtsvb7AG5xwx/
LyMk7fxWGFf0mjOCcXlv8cZwJfPTIUbuWdOLqiiQbj89RfcwJK9GhvkowtG3Esuj
cmhmBfK2zAcT6XPdCRB9WsTXSuEEOj0LryjIhHk0uRfw/sNRGaDnptbeAjEfF6OU
6iDsukDVfE7gPKXKnZ+GoY96LEvpzuLPKTvsF4NPFksqnk808DWY6xM3aiQyqI/+
mNTti1l5PPQdpMMrSWAVlqfjAzMEcO2F2nlSuId0/n8KD/s/XmyAa0M7tdM9Vnmr
PHxGUdRL1o37Fny35XQvqGqY5HnvhvfECyqnOrMog4sIRY/7RjI0rWfONRuah2pC
4zlQos4LsBcZ3eiNq9BfBCCtEvBfxAGB13qCJHnGOC027KY/LzNnrWCHwTIr+mC9
CG5dP3/BgBg/o/h+XM9uEEnHknNOUgZ7Hg0QMWYfu1O0+9Zzz+9y4q5LnRHao3L3
3LdnbGulnMXxr5Tu3C8FIGSjkxZoUsDagrLXHSP5rIiASOwZz87nEwc+dLOjz7Sc
MpYI5EyHmG6u6tLdP1NChe9UcRVY/k1rDQGgHXvxksd91VZoLmYNvM0C3yHP8Eqz
tWNY8hq45n1/ho7Ez/pi3c065QCVBTX2fwP6m9GrTmQrnfPsPAi4NbLCdJbAIvH+
BhobJzVI2mnFzwng/LkBktAW+ePrhbAeB5QqKKjZCmG3iaxf4mmwibSRIsmqAWex
xTCDz4YelnI2PY65Zd77Wm+5QztQ4Liit51pu7w5TcOdFG8VESp2egvp5t3re3+W
/Z0czRNM24aRJLRGYF4rxn8tMhqH5j+a03GjHWWLQdRrKCd73Xn+91tBsegLQ77z
6L71ch9g4omTE9vbVl9XKi/rjQmyq2gkz3B6U+TzchWeJqzHOc0SDKbb11/NIBqP
DHZuw1Vh9Y7f8se8Dw+K+/K6USyBvx2x01q2qcT4LsdWQB3z8RyxopMmoawhlZJe
vuuWQXQEajT7VGXDch+QiGZK2XR4Mfx5nfRHgRzuPNRTf23VAIx5eVUdoZxBsv7L
5KLNkH4B0nA6YVKOjVoG0uVEutJSV6BAdybdGFT4Jyt/URSIiG7gXYPiY9Si4A5y
0NUfE0tpBfm4l9CAcGXt+yky+mKTWa0ryKA1MqCqnCBJ8qCV8qAad34ksN8sGm+Y
qIaEIsvJ3hlhJsMvvwS/bZphe2RYooWslpBAF9t1ckvz5xyPWc4n5DaYvSiU1Z2i
XAtAS20g0y4uhzS80+faRrSy2f9CxSixdI3fM3v76QEdIoUoA42P9Rv+QMNkXa4N
yPHoN6qoIOu42A4dyePfFqG0NbHUb32wBqkXcc6Z74mWhR9hRj2GpzJVuhhjWCHL
pXo5ZgfVxttSoOhrMlTfwBNgJeJyEHlUfO4oIAiKjS+P3ecEGb7+OiOyhfp96Va1
d6Cq1qz58fdBUUNcqSwen5IkZq/RfbEpbxVjS80NyIWcVxHZkvdqD/9T3F4pCxWe
49HlnDOaTTAzvfwOQ3uPIarUlsp3icBa/uD4pw1p9O9BbJV4hd1DGnhG0AXaPICC
jSnhskRRW61umQ2cmiAFJDdKz+lJcYuE1w1ZFCGaa932QQ77COHAiRV0P+0biJOu
DO6ZSfSqahBmYRgzz6YTFyOD3UcsxUZ5KYw6888XMZyeL4d9/0sXAkRHG3Cfch21
RQzIJK3XunVjtMpaNvPaUGdcdqH6pUg12oNgThe5YwW1+zymd0GwHAzn+fBw4jHR
vjj+k2UQUAOJhPj7Wz137HKWVDuqhzf7HLSobLEoA5416UadSX2aiRDCipRaOeuI
ba8eCyKHAFuqlrFaqX1E+UHfEAr77cEbBgCZmRNHwQt90yocVbADaUitePTmIpQl
1SMDxRdixzK+uoThJhntb3+0ixU/WS7Z3rnZ4LIAd6rKQDtgMorsQEziH3/k8X+K
bjPm6cfrTR6WB6aIX6jFTp9QFNLktPdOushtjslFFnqU0xvfVftCfXE4dQzlryqI
M18gop5eb6Pl2p8LZEn76T+1EXQ8FqSGWW/95f7ejGZ7eeAjEBiXkzN+2/aoJn5W
fdDTaxE6mv4Qd1zTj1ghBIoVLHrRzhGydYOjZHlee8OJMYxui3dpiQ3GV+SUb0NF
KLkFYcepT5Cu51c7x/k0EAfZ/NF+G36MAb6tubyV19zozR6m4CbWY2hUWnk9v9Bi
LpmSFWdaJlSytA/Mt/uaq6raQvKFNkgD24sbz7CFB9qcRlYeTU0n8VUTdAlaeIqJ
Ba28lK49jYEUzoCfFINBH+tdNHFmai0oxxrWay7yMt9CimmgYmmdff5fjICRKzfF
nhZ20qdIzKZSnCNXEu7GxJ3W98q1hSqWoNNNqrM4k1e6ehTQhZZAofBGYyM+mdp8
NIjwts7EL4NLh2V01pjhmEzHMSQetQVbP0yyYTmKaT/QgQxeq5dlSO5/VZ1iNBlR
KS05evLY95gRlO7DcTMNl4VLHksCuT+4HR19KPh6/HezDyaG915KtQnV3OUtRgME
xpmhC9uZgFRPadeUVyUnO0BzNP1jjANSoibNVFXKvWEhAwV6vNpKgt18A7IYbtQr
aevbHJnFQ27mveGVMbfVRSCLtpLkC8nwriezTEP7H3xzek0TKNLKRQp74dLvlFwl
MQpf6P/SVQWx9OwwiDBaQka8itJLaOUgOsVW1djQMifihEfQLKu2gtYF+S+JuAL+
GsCYsY7aL5WNs5kmwPPsSnj6xo1XwEgjYWVZcPP7xCgbTuBJW2GpjZrjOG1s4HZU
xCsU0w2/1pphBFW9//UYXCntIv0FQK9A6BlQA2Zmf0cvUt3YmoJHaoa3nsgtbKOu
0uWfptXqx2dmNJSSYRc9em6UAkG/c2gymTujuKRcmMU8Nhb+lIAdkGwj3rbCucxw
51OhCs7MIh+Zbru3TfRFe3ADNwaFEQ3nUSSd83ite+uhLt4zM3c5QDuT0E+q/fxE
wPItv2sRg8Rxn0d51fcPPcoi72Z+Uvg0JpVP70WWTFQPANr47Lhr7uABkRdooqLd
0lXUcJRL/f0RE4ua1ybYPza55ze01+YPw9O1KcPyBalLK8dqZI8JShf+D5BoxaJe
VwdJ/BV19KuT1j5pyK/Y8Ho+6gnLs5egTiazamOgN2IGR1xFhqceTabKPzTfx8Ww
IDqVxtqP4gpzX5Ql+BlxgPgA2fR6FNTWoTc3LcwBNo4bYDpGagb8tdQlKRiF9OE1
XsJPjgrKg3oGxALnkKAvF2JlS+etHIc7VPtd3dyeAoTC8hs2w96s7lrCDZluQfmp
D/1SvXfN9av3XKUbcFc3rdIWFrQe8GlyR/lW2wXCja2TFIS+JfIjFWh60bQiKVta
I5Ru8izZfGpEXA/RANQGXCQkkRDDujAJa6Pek9224KkX3bK2tNkfgaBx1S7Q6CTQ
S6pSGOaKFdpHS5zB36Zn3LxvPLyWZ1ahrFnMTiNbVHi8m7raI/+kxfxUqI+/AkaC
sPNbyHrOkuOAgV2NxVPmbZUU6W1ufDMx+GyqtZIBSzudtMfFGlRzn3RlNPJi770v
nE7zAPyPqQ4xy5hyXFFC8kLsNOL++VyH/puYPRwAh6zCV446AmW0rM9sK/FB++AX
bIgms/vr5nEHxuO1tYQz5AG/TJnQL2ap0T3Q2LXjz8nL9O2TAHBbyMcA4pK8HFAA
eJnP8aIO8PprKstnvHvn5YoLUI52Yg+toP0EyeyobO6VEyQX2Erk0iUFTBfsDCW4
yhi5W1ok8qpqYpmY2jcIhOAgGeQi/Z/7hArskbyd3wV1nIG+aoYsazGVlVwEUe9Y
g4a67NdxIoBt+3y48W20k/KSHb0/P0WoA4fchlEKLYeadDyyB/DTFDSZuhuLNIaI
7AWdds52JHPdg6vLKIPzzqzN9jaMO5U0YJ+781bJIRZWxgVHrmHmwcPipvVv2K6g
Ng5L0B1qXsNSDGHWqME7FyqLcgR/3vTHq1xWY5FtuaqRPmVG2Kld3sDCJUo+CTu7
MiFuhcoiTD5WvTScGbMX274kDXGcFCixhpxtRDcc9Tuq8hicixYtsYLc5khnNfC/
Lr/akFmboL2pRFqy8MWlOea9nEwZira0Vno7YXPdWslfqiE93ciVzbCnC0S2cFva
Fo4QZYn4IZRwuxCnODQ2oqkSlpFFOQ2durairYJ0IvOz7S7hoaFZIVGhcvGbQQdn
rM5AjmiiRX4ITdL2PykNWFYjBTSd17gotlUmbUFlZbCStnOrj5ZI/+GGcJ2BfBPY
u5LKmqRhkwqrrYOCfq63DwBMWuuyNI+dQwJ2NLNp3wfj9Y4QZkQ9xxQ3cwOVRpee
IaoxbWG4KUItqWwMrnifDyQ2I27LGLPplvCdo1nvUkZqKPP9uCT9YOLe1rni1A2f
hPa3hGMENAVm9l8nPB+dhKQFKm4Xm3LhjpN/ylBb6cENoIUpHQfZQXOUDmlW9n+g
LVmsnF1VcsNJe0ZilGmRHM8Fun0d7nxbAsAuBoWAsh7FnriSHwcdQiijBwd9PfSo
tXlsTu58T2Kpnp9pw1ehL0Xy1kU+EuaTBUCpPYGwWxRWwGql9jymZz5Hj4tj+Fe1
FB3i4PxqjFA4C7Bl34CaeF2YkMTd3qplbh5CqN8RqAsIdVfHJ8F+bE87QCtMmH4i
dzqXghyBPVsKzYpRRMvo6s6P4lswh14rSggFQYg1WMJED5LHC97/KuJfu3CVLK4q
dmWzkLTIhn0Z71RBIWdtu2YIDlIE+ExNmRo5UBBKHnPemYv0xRBg2s6kxnj+8zHO
3yXhGByHmZMyPA2IUgLzvCZlAdppAZTviD9LCLbuPQMMoMbDR2Aj80Jrl9dOqh2Y
vfkegvWDUJYMYWCEWeA6jj5fMBossA30SixPO7gIoYpz82cFX+mbc8QtT9NEfYCX
qHb1amXOIV1pwjetPB8PuvjV6Wf3Fm8xrS3rN4fyzOHDc/zI84MJ2U385/EIuBEM
Lcr46Wri1E/yi7vUoMOqwytjay2NZxnXBF/b+whCC1KI3sk0za6iTSA9dsLfFauN
iPqaMAV6WS5ShKumqlELCD6crNtRT41kqweroMwT2SnFhbuqweICPNYn997juJ7b
gMGThRGkArKdqS5BxBkSaO5ymoKYznLelXhRcYH8I2uKQPaspwhefq1CwPmAowq+
pioQxn88KJp3x6Oaa6QhuQqbwDwFG0rlTxKQhruyO+gCJzXXQ0hs03zAdv+Pi5a+
O/xnO9S2joK36HA9NXNTOZT6z0Cbu6T0OVZv/YN1uLY2ZH3gGQji9cHuMPTHJZMp
F18K8B015QYyN6VCHSSYaobCwYGcE4sFeUsxE2r5ZcHjBx4m7fwg08XI/J05yPKR
N4Yh5ZG3cp2+tJNDpKfignZYY3WY4bZF+kX+CHhB8GFoymY9XZGXSJkMd5SfkzNX
6yXNzhiCu5jmiWShUlIJZbKWSHWkTJDG1so7wCkrksb86cuSuA82CEpLRdlhke7M
usS/b+wHfV1Clr0v7niJ+0uqmVdjIIFCmbzUuer/BVeIvnrt05f7H0eB3sfmfSWM
FEHaRghFGEHp97BqVkkK2PSaztrFzERA0SR6dfebF5Pn8RmnSVleiVpYomothW1H
WzD9YZzS5neGXXfTHdWV9TJoaE6rnEEkTo8pCKRIsghvdX0nSfib51yQd/7sKHRh
r7fYvJZkFaYs88M1LF0jQYt81ZxtPEGjHSAAiKz6Ilm0g/bZlyVJjWFTEl0l0CMg
4ZQU5a4ipsJppbXFAHNu6z+RkzbYLTYnsxKZsk9bvlbdoNv6Au4OfF8esUZAgX5L
V3EPZdVePClE9sn/vJUHjaywtxE7Lt/cbVbF15NlqRwF4mqSGDidxpC7LePDHxKQ
NxZziOWExO2dyFHjiGneqbrBJg+g9i6iCaaLJOYhbBLk8msfgwiXZn67NCqWpZGz
v2180/UvA7gl+CEeKOmX5MfYVLxOMQG57ls+5fxTIA5KGVhDM683cz82Ky/YsM4I
DnZXZJO3iavSr7ow3p9KEUT9BTyRNkwlqMQGe+IkiwYWYbFaiF9s1D0CarrFfaKC
98eEAV2w+426AhyWyilZyaDV1uM+r7xY6KxhxDFDijaVLsITCRltJYqn1lysgfHk
JpMnt+2M+nSgS3WpI4vZRQ4K8kX7wrqNNZf8qAb7VTVKV1anz8GJMOb1SZwa4SwA
rN0PREuLbkLyeiX0W44lai7bhiRW/Cku9cZcRZfI5ZYY/KsaS495lPwHlW7rNyir
kWMExbKJi7gsiLTra02Z1NGHmniO7YD1MsS23H0R6OQB4CxwvmHHKuOGLFkLaSCE
U5gPFiWAzgkwrb1C34JomAf3LQPyVmx7utI33fReah2RZNpu1WsykzmaTh0nx+6K
8P/pKA60pZrFXP8cfspIMQjreOPgP7mCX97cwIA1PaKTagDcS8rhtsFDxGetKl2i
M1Yx0HH63SfjetuFinriCDdplMeama5aO7h/xzpXuSnQAgQ5a7+xg0TQ3jPGCP5E
jm5SiUrmOOif3KOyRVyEvMdTvvvDItX3hD7mVk+96X4+JrUDUMqUSUomqsjnFdc3
vFQHPpjF9jY3S8okoafWjBhjg14oKsW8N+NwOuBwTLyUsLPqERMbAM7Laes9qOwd
cveImmCyX+A/7qApa7OQqHA5shKREVwFhs/IYi1XVuflE+PQ8UmvQXB8qVQ5Hwe4
nDlkUaswdo9tnJqqF0Fj22PvZD6TuRCt48Mpr+1ADwTv1WiMFbpRfrF3nqiMlH/g
okfhQsyCsNZu2bl9Kbz/XKN58bmefM2RNSvpnK7/Iiq09E+fse4dMpg/KqWGOe15
D679MrvYL9EwspCIAJQb8f46mrjlTwaXegUlZFXnASSqAQL1CLQ89rnNSB+qPANu
c1wyuH2s4+efHL0aEkdITlRmKmyitBjPjzAC6swDgrMvSCgTqpN2FMQ0DSrjxCJv
6nlah1sTDsHg9+QWCUtzbiKTeWvOz4VwNG7DBOYwH3pyh1nCH+Y9dczrsQhfLe5A
nbDXb7WBvNzQo6BcCxQiiQMVRJoFetuclmpEu4qn29x8wL1au1FK9fMMl7Z6VfMr
3ZK4LxZCYg5ztoTUr/0J2aJgFmn38qrPBff9Qsab0eAHTPrjvUAAxDiUUA8ah6yt
qRkYxixWkC4k0h7U+XFJn8LZ4aibAd+u4aOcIUGs0LRY1SZ2VmAE5X8kve+4CYpC
m9bDdGMZGM645dvqlNUTGTzRgyZFYWBhCqjpzuoKPpob1DnSphvdkxqtjrFVHcvR
RkLIYWQGYZcSkqjnRlnIgGqQ54RCN4wMzhGk0nuorivIPI9cw7JZ+O8dwHk3WyrB
OX06dN8A1xSDHpGNzg+BqfTbhCHcxyTZ+wNaZFus3yGm8MG2UsCb0vovMkXUx4sm
H6uj84UjXVqbUfqd//bOiOQ7XV/Ud+gUj5dx1HpCEz3NQAAZfHN0gwthmaLaKK6F
Orl+RwNB/JGaa0+pbnMMnl1uFEU0Y1zKQrbNESSI1O4tzWS6tOtiUKH9bYlQ2X2I
U9hQh+k/nG1P/qX13vo9eNCFeNcSYE1v7cZbFoecK/bEjl/KukB4aOtpX1vBqFqU
t9HyzPYxMXLMAHnPNpGuM/UYJzy9b1Zq0nYnX6T0eRpqYPI46hWD1jrKaKfkuczd
2MNMPjcB/2SjKBw0Sh14hYd1bn50mYfGE6mD8mHHv5pcWme2XHUOpMeD3u6hMR0x
JVTpmJkMPQb3wBp6rzAqYjhqZiigyCL+igN3b5yAqi8Ys/HsBjixculRLHFvG1u1
v+Es/Sk6U7TQ0x3IDc/tG9jrgZUSbl8p9L6fGTQVS6/mTOS/EcRQCI0q/prZPrI7
/JHfS3adKIDNXI3AFCZvXUV1YS0aueS7ZTgcx2QBhNnjH5HZHkU/CxvoaRuT2EFT
TIiEfU1kpbmBHjdB/W7eQcn4TmfKaT2ZbPfmY7fc+JkS+HOfPkdtgJazLe3RvCcx
Ixu55SVRA1h0mXKT+TaJDQ6WSiRhprCwwJfqsCqC15/cxuMP40FF488QK+afenAs
UwA5jhyQwPC70mr6XLC2WOxkkkq9Tteie+QAWo3iXYto9BNSABFx+jjnbdjUvOu9
Fvl1E4oskFy5JijCvgZooDA/rYpAXCW4kw648C0gNIzWg4TteShb29U4CYQv/bHM
csRebbUZTeRI8b4EYZF7g7XBs/YCZZBpraxZaXynfRfTczTg5XLEg1Od/RPHtx7V
Xe+oFfigrxRvno24TdisnfM+k9jIMX4i6/H0eQdd2+zQlc8kbQtmg3NIQsAm/pxB
7RmU2EPtt17RcsDFuHv+i5b/JB1qlUZzFnijCjMpBzCT3rQU4fb9PItQOcs8Q8nw
BAO6PF4kAJh2N7N19/Lj6wbBiOe1PbRrNz9wM4J5MrjcFcc/smj3NYzWje34URhF
K6BMKelOEPX8LsWFdxaNYDZuMsalwzkhuSzmdGQcl7b119Cm5QwsTPbqW/pabcm2
78Xak1FvcSS2cneP8gu9QWs2rcU3eHivYtMKJO4kNByelPtYx6kCH4LcDd5QQ5AM
nR7USOT4B8CR1y1lwGCpR+hApmlAyXK1gch+tk7rA1xHDlvLXSj/5ye2EAxdNp1E
b40+GmqxGrxulJIXI2u6PUkYiIZursHxggdnjv9UdNz0AFQf6sG3ObYYp9TgsBuW
hc6K9lr1ZnrQcY1jwnNT5t01B92e/To1mMYpSQgnC1CF3zVXCfVfZlRFoNH9jjF0
EHQpJk3F5cFutWawhYpILHCsu2I38Np3mwD9vWgZ9QBPvsPE0BkEgZo/Dzih1S9p
0k++F99HcxTT02SLAVVd8UVboHvHEns65oEJP+5LAG3JzjhiaoWHaYLg2OQNUdJi
P0anA67yNS8+fMkA+saoz0eQ1kH7L/xtUgrG0PpnC38TRDJvEohdvvCpnOL1FxWr
pxu2hr3fm3h8ZFBGeNaps5uqsaAaPKaFqPddB7bW10o9+n7j9YYkHW1HcuNZtsz9
66OiyPeDfqU16TEa4XIvcp3JDjWYdEoXkwS/Y9qFROF2+XDSw//PKvFkt/+GKXm8
TyvrgN9+3+98fp69eQC7ZlN3MjnWjmWkrAub47Opt6OSybz5Iuvas/EknJnOuoMj
8fQZGwJx1kG/agqKPZo+7pNqX0ODaMpax6oWQjP3mjWYA8ZJkMv12sbKDWyf8f95
7Se1F/WLcMULiqly/IW77P8mdzzcAq8611vNxg78/kmup1OjTTvocCn7LgcyVDjp
x3vVbQUxr9483zS7asC+s4K1tk1ElLiQgdNm8ER0MTU8a4Ln6Dq5WHPGgewB/pEg
PFNqZ/xV3LEAf9/zst01sybGOC6+sGpF6ANJ85Dw4O0xu9PC7POFSHVG3mSJIb25
10+fP9yNwCNJwpx8pob1FzgmqQHp8VD7NRdxTz6BVHmCjexOkOs4tf53nTpkPvF2
uBTN7nMxjFCeoF2ExPl5aqm1v9tJ2dVzQZY1lPjOo03g7j/aWNjxG2oRz+mxG42x
XdIG3DCvrukv95OWAB3zqw+fnpWdHwRoOcs+7tuDFPH/s+ob1zXpBQvU35e7H6xu
+MceCmN1f8+N26oVsRV9eCv3hDyc/mHfhgkQDeJK26N7kP9VxBL5BP6hsiX/ZyYm
TA0C/0UICph1ThFcyt6RYrdRXmLGAJVB9vV8OZB0yQcMltrtjnRLTVeLUuOhcOtg
AF173vVPmZJu+KyO5N/dE9fudq0LuWsX7INQeKiGCT/g0dghMG4KdKCXYg4tI8fY
XxFIF5A529rMOzuy11Nqm93OqZi9yJTuO2OodL8hmAqdEaHCIbAAwig9DyDNUUAa
uDt9HxP4LiDOPAvunfUX0H2SRsMg93UtcJ3+jDkw2pYfL4urycnghaokVfbSQJA7
mMW9Hs2BmFojaPsLviwFoeDyUq1gRm2LoWen3zf3/APs8hfWOH6BqeXMG/dwFgJB
8DjO3mEXW9+8oFubHXkM+lvDuJeeEyD2qRHSnzh5iLgmVPNDRRnuS5fgfVYGjl3R
vet/iSl32ZggMEE43dvmijCOXu0PyWxhEH5mwkZpHkfYyQSrbLi5ve7K36/+Byjv
7uffBuzPNH+0P2F/4nDBD5B9jhKpVGv4SdRFRrqmaM8/XHkM23bpEkQOOc4tbd8z
QGYJ35CbDdDz5lwOAj0uoHuPHM3cJ7jzKZz5EBmZwHNrAvJ8KJjjxfvNVg4waVJh
/2t0zqkjg7wS/bUg3TSxLgPMTuIPtH5rSpwLMJsSQbNIHHQFYaE9dJmY8YeUUwgj
xAEa3aYiVyzCdrhEwLt6HPb9fvB4i6xMH5P1+7WUETimxVTh/l4n3Yaimz3U0NpC
FMnF48SVG+GhwwLr9rpsrDMO982cPDKprRdwCf2Mkt6JS1hh7Xf5qx/SFSfixibo
3UOrs0XNe9LAaXoXAWcJ1un00wQycHyV+pz12Cxi1UiyW1upzssy/wdOacUCcbit
a3IZbofZ4sjglTmrGowJJHhJc/pZI0mxnBqA7ig+m41w3xLFxrNv+N8+BggiUTBq
KnG2eXnKwf5QQOk54kiEu5Lzg5AHk3s1/s6ezoLhFjoPzaWv7zj5U+WXatu9knip
QOkKv4zu/DM7OQjTQ9+tA8Q2prNcAfMJB4HYrxbWF2vO1oTlOcKkhMQHOkA/ncJG
iCFE4E4BNbN1DV5zpiiHD1mWDooZkAqpl7SElxifkdcyIxFZ/CZaTRdNZKvNcixJ
rSa2BnG/6HIikxPsMooGq+St+u2YoL3nTjpnPrITSxFbw0h/QP+O69aMJUsDhqA6
DzkEUoZDkvE1w9Lf/fWtSK3XlHOU1N78LWjdBhUCYzjvZsSse7+ub3P1iHXkqs6U
ORa7QkDq5+Ms5J7Jr35DInQRdhxCcWYn7QsBvncLrIHhwhlOGMejC+afxFcv9Jtd
3lTB08wgX0sVrEZBO+QeZtCvQeHRCaRD5chGL3sC9HKjk6IU3zm7p3QbHC4FGbCN
tlz9ek2kCqVmKxAYUrH4LotmegTx3SUBfS8lZaWRPR5snrv/SrXMDNI/5xTENvx8
0nEng7tu/Xbc+rT0Va2rTgoyCtiogVJjMLHRgGb+pXndVuwJxyQtHgUr4+1QUAWU
nFnBiniarg+EnAbFKrxUMWtlPDQjpDasSQctbLJp3kZWa4KyCQKW8x6BJ91Sr1gL
PuRsuAZF2Fr1eNvkfVSDwYTaJt4LdiKaxajPlZr2qibc2M15BCylXjTZHBtzpWbP
FWjd+vqzHQ2OAo5joVG/V1UIji2JpnrwpkaBP7o4HHs5WiA8xoBiIwwm3DOhIkUo
+9ayoNrqebETbChONRBluf4NnT3h8M7VIQNHLelfIxVfTz3in3bvTHyt5PgDP2WX
+tlTbCgi/ywZL8frsL8gQMYzKmUxoNGrYUMoPuQ5RZlABzbEQgfXBs7vduB+GmE+
ic1louje3CtPxjaT8cs2DWDs8RTxpeKNBWBEIj0cQiqbcawpjWGC0ryxzxp34o3o
z0hzo5mSwo3Pu0mu6dKdxo2NDsJDLYO4Cdut4Lh3EGc849xNr3EEuYlxiehr09kF
RMq32idm1YNQzHdcfpm3PhUjDLRRLzksB53Nozoy2y/vpfU8TUsWESZ2tSkF8HrC
HPVO/DcxtpR5zOVp9D7P38Z1AzzqS5kdOFTLtO2HDpEsz+ZTfj7mnUEeqU3j7TFd
k+JRC+zhRYU9FITU/Cp/10cJeFKNbv7bVFeTOJmabzzzm8kjIeJzJOPAZPNcU97R
TV6B9JApa5haQAz/PgnguJ6d5f89SYJZe1Is9CG7yDGLngoHG4bzN5Es1s+i/Bnn
QZ7FiAUc+ye8elSgjk5V/H9srx5yQyV0W9zbPvf94e5JxUn32Ve95V2lbK2kxAMT
c1FCVFWeFCM9vSpi7TpX+M8QU3TdfglpbtYlR88hFnUiQdZrD4GENTseYzj45lMD
hm8jiz2deRFh6Ak786uEJRKyUd3lBm8kqvmG/DkzhNK2YPLPBvZlQ31q8PcMVNiY
mhYYvy/XBGpa72p6WCce8NErdoZAoNQLQJnustkbjHBdEKbSPxGo12L7yTCLb7RB
Qhw6TPk/FNizIAWB12QQJlcew6SvsK3M7g2HoRafo8osrS/Vp9HrykZW3+0NK3DP
O8KO2felvEebUP/aiwD3SyO3IqcaMSttsufAf22yh2SO3E7Pb68zLufAeeF73L3Y
PFFp/uxAUl2qygY6jzkAcKtVSwhBwSbeFgv+1ijRuKQc04NlwO4FnJF0t/HBZmHD
a2ZVdMJFFOi0qtfBI+pAzbfCW+d9VvEdF1h5wft693yiV5hTQ0+Xjxt1N7AqDUe8
TWUGKRWpP14ydWSynOV7nlhnE1uUVNlmUSj7Lsg+/zdSmok34j+8xHhf3FCP18RW
wWm4shIlcIaL+xsN+UUaS6mX6vbN5QP/oitIkdgWHDrOuaeTFPq2iaZD2uXtZZo0
78kZLFg0fy5/6iIvVSZ3i3CcZRSGiWpQaOHEd4eJn813GYczv6XVn1T3Y0Gjl91e
B06loWnvOVEj1n4TAyFLsjqPX+c8GQUsVSiP5OEX1vwQIneMghRFeCW+Jie/xrmu
9F8UHbX8nsJu23hAX+yraUBvH9FldDSGx9GwArt9akGWWLCNWzLjqf2vras/wGcC
5Kfdo7oLyo4Jc2wenB7vosTD5BFDxBrtVv7FLrQ5m4w+JI6LdDzSE8FmRtF2SvO0
ZK/ooUZLob+DiYmcVy6zn910Txk7jb5BrDveJEiMjFZruZZQy+l3/xbyiQDoOMQJ
UChmXXUgFGRU4db5rku/7qW+9J25iVIOrvV/HN9vjlRmOjO75+qZlFlcpnuK3l5W
nMhsiBOR+a4BYGNmS14+KMMPM1nbAyB7+dzgGXiDE/S9RrK6O3uDiIHWHaDUcNxJ
b0F+bXK40druKBCLq5+xbR2eD9N+rr4yLUkkMBZGGk8vglyv0ldP40hhNjPqTqyi
/A937o4ZkZoHWkINWXLBPcAXzU4PSstVhAfSRejlD5drHuNoutsSDCjm1idyXBST
AvIR+1U7U+oTitXM7CBk5g9FLDpS+GjTUTBw1iEIrzXHlS/JhpYJy3UeE6kaFC39
XBFBahtPh65ssdGbReoMXyxRk3vEwpVmdYxhD+NnzZCqk9U4dJWHvrJMb5Xh/Mr0
x8N/XgFEWDsZb7TiKY59gelubmdHfpF8R4YzlwYrYB/RYZ6lyaxcTvsnkU8Q+TqG
HdAjjzr7lvQphX5KnOJMJOt5v5bT9HW6VmA8QHTBV3yyiyu4Y+7MoSobbYfbmEwW
aQ6BZ+VCrvdz/u3oO0RR38eFWzSdBeBvTHUY+o05YYZ+e4PN5vuTLeKZf2CAJzAO
/clRZdzw9Tx8jWd9BF9NGca9ju3UvB/TOHXLcGMMGtdKU1WbFOASxm8KUuKVwWQh
LIHig2DceZgzfNr7e9nivFonE1xruodTmUimH5DLSa1JwgeElOj7Zxcfv4SdgWTx
8gXl8lK9mbgM/XKP+r80O5zETtZ3M7nv/tEjiokHsr/Lpc9OuxBeAr0ocHtYWgcX
ljgB8wmtCVWsKmnWgT7p2NMUw5KBL7U5Hsbf8LJf6ar8hpQBkg0CD1rZFfkFNMw4
pPRqoUzUIky/0BOHY60/0XF2GeWpXZ2dSox6F1Uu9RisAFiv23XZ4udoI9z57wV9
O72H9BC5ISyHWap2gZpfJ7KDDloHuONgShV9UxFM63dbC/K7cMzIhwcIyE/ErKHF
E60GSz4OFA9XbyFO8nywcZzd5z2RJRGHEDGAkSEe6gvSz+IvnNDerBjFIyuZH0Xc
N5eCckgPPQ9em34DODwQeYF1XGTIXY6eCBz1+EgRPU+d9bXYslzjZUxRJrTgZwLs
b8m4bAFmUHw2aEBPxuWmBudVrzkgBxhVXc4nCHgGaiJZuW4OyZ6YPrsDQysjV6He
Q+co6xcYyoYiA3c5HdSxGvtSWNIr/0b3FKn0Bng/gsBYqbHVVBH5kOR0hmcEkcUg
TQKK2rvqSXVbOdFFZzPHWRDkoPa2hN75X8mzAgQSFmamYqRRx/mg7yRjCIcj9qdZ
8S9brh9Zrtdp28rsFj2sJiiujWsqZk2+KsZvxbualQXGCyRT6yTM/zxr4gO+CM6o
8X86y8nG5tLIm+EW2ErwwkP99NVpnlMjCElYOyR53ScRysFUd1RTVOjTFzt5ewzH
Uo2GzBmzzTHKj1po0kZLC67GrMpdEEvwM1J1+8lxNsnJSLL7wlzN12T+hFxixyOe
JK1o93d7YHR0XYxx2N22uY+6uca8oXdGBtC/fyoVR576n+VJ+hlJ4V6gpEssRI0u
t5qrZsCh+/WxHURbCAtG25/sj2LNKCvWiyjdJ14ah5SCzPRiv2y/cwmQ6SHUxBwg
kiS9OWnWpFGsbSRPWmmQ2I6ifJspWRNtqnk7Z+SJQN24iKGtnkbbIjg9SfCdqolQ
6sHcZojQ/j/+n7HjiEyJPdAL0wf+mtpclRfmJQ/e7Anb32UkHNQnXXzpDmRZRDiC
JWY1BJ/sO8EMk9pIBsMpgxChZVWZ71eV/bdy/HAXG4CM0OFOQ3Q5Vga3WthYzEi4
nSwOMCf6foHHfJZt45i6knqvR5yll9ozb9GiTcV1S2MIyKeC2ybpUX0h8Mrm4wLl
kLN1AqZkrTuaLhpczLJys+GWHAi+k7WsHV02ywYnJuFvlliMtAur6QCocuTw9w81
ohN4v6dEZNBJChQ1CTddCom1zwOanYuxYUEyIkxPmR9OiHe5m7yJ4oW7PpbG7Dv6
Ayc+kuSFpGTrZT+7qrD1UnWgZqK90BnF+8NHwjT7QJnOh61huiwCDwyxnHpnZD+J
WgFSQP0jnY65HxVFGyw8TuXgCvfllDe2hYMggBoB9pJXeqWd/h/z45AXc6SpAKDQ
m8yypdyK3QnyeiFJjD8wwcQooI26g6Ey9Bq6uoH7/y5lM5eTWzbkUBXAqs+Vxpcn
z2NLBVcnPDlpF/vAZ7QTWDV52DvLzTUDmWCPfr4gzmc3LMQYgR7KWd5q+WM7IdtB
YCoNSwK5wT0bZccVWqDcMbXaqax6u6LyqjmCFpM6qB/wIIr+pXFiahNj8lVHiSNo
1FCpHQqxMLvBZnFG5QgEzYRyOYS1A5dXUHGYu8X/IBevi/VQjAiML4nitoPLvUSg
M12numEJLE8I58NdeZ8nCGXHB5Ba7bYKAfgGAMxM9c0vWWuEvL6uJtSeVv48A31Q
Q+3GxLWRsL3sTlfXDTxF6qHsWIpbC2ick5x0oeI7xfUXrddEGJ3NYyMZ+KeS7sAu
py8H01oMKcFhIsSyKdfBNNd7Jd8bT0x7afzQZT3Cg/qE26Nd64W3a8MZec3axT7/
Muaq6DKYxgU39pfEKnkO2Gf8HvWrwO1WJhX9kXEAkYKt3On+/M8V2hEQnsXqXrUf
nfmom3i6vJkUI2kIFuMv3CWmHagjSDyCFOcvc920wLR+M0eNIlddeybb9Pn3wHj+
429pEeo3fGZsxheRFUUGGN4nCYA6kMNsIE+ztK+AMd4zoakTvaD+lU0ysycoNfdk
dk9CJn/MndVdf7SrcMcc1ctH1x9bwcvgPnF8tuCnrhT9Qt9ZZ7eOx1AxzZp7WR6i
qc20KVP+NnniGzuZ/qELvPWyKoBB1rxCozVMpwX7Tk76Sn3DFadEdSO+Hv/Xzcs2
tIXdC4t4u/jrRv6m/ENiG0FRAa2IThD+jp8Q2TpLFdpXvb4pBGsRHWHUE33LSKP6
9E8YQgvrpcU8ljdJUxqkruYQCz+N44t/4W6V52VjTuypBBizimdQ6FNkdSaGiWkE
WZj9D1F2kZ3hgP9DucUkcsfW74KEZeUCSUjQKWcXyYxFuG+PHXVISfTHZi1mrFOm
pHsK509YVD5N9gRsItQ+tGmGbpj64CZpNZixR4Q0H52En8EljyOE9+REIrTycLUz
VqbSs7fX6K8XHiFmNHmJFMcQvCwuJ5hkpqcKKKmarMRPH/6Lh+e9b6MSSPBa2C5H
GWHHHw8G99UcvIM0Z13+VwjcN6jfZRtjk+Mpj4lq5X1eukzBGRuKQeMX33wk6hOD
BEZMgFGSvTlUIZTKoWbFyJ+VjNVZZoVlFL98PE5Mzt9Kl5FA4TSwAqQin+5sM8Zp
iEVbdftlxQz75rk7H7TnB3hAdUz4ZPeZKFFn8PO/Lke+WYXQ7r6BTVmdvaAa7Dlb
y+VnkunRHn2QtP0/zsAvqHjnfFk1IYWjs9XrsBm5YOU2IyZfNiCrH2M51JdFEOOq
bPU6g7jgVkkM4kyGHsbKvyCCo22JUrE78apcLc7CC4xIGDdYTs++XAPAIG8ekHy3
/Pm+LlF4zgMElusT9wnqRsiDPNZ7sr2yOhP+AMl4PN4JF2nG5Q1mFiKWudEKPTir
sittanK+cEfk9KzGWGDT7raNsUcdXZBLGqwtdi2jKDWt6+hOduhzWOZRbK/+jpKW
S6+w9S+0ZTyllXsrqZ5FeQ9sWnN3s/3yM4HBgeiQ+0PBWQJqWVgxvBLQawtNmJ0j
9R2fvbFe3uCnSN00XWxvyd3kvT3a0JxnV+IaUb35M/hwNRgemz7OSTrtrCL4u15u
KZUM51C5yv86ycANuaPnOBiP/zoi2h4Qmyt6QlP7S0FW6dBbuoskAHpfyRPvy7Zi
tX87RG28uWO42akoy6riLyr5zgeeqSc6LjBsi6kgfoIvHceuR+xmLE4CdaXI9Y/s
JCS+saxAbT+EdabsdRQ6/MPqSOV+5LE1uH9Wif4AqhQnQtpDB/nI4undmzMGE04E
/SFgyS5lP4rjJ7kv6yQwDLY+kCLW4CG6YsOut0k1gBntsx6TMwZqgUQ136FrdtOP
XzPXxvxTXK6A+h+GYvWTZWILntlCdGxBM1JysaL0roPIqD3JTGS0r+Cd+6rxP0tl
Dmay24h8CD8YF7//TJ7iSyhayGoXOdrj9fvIcBOXJbomRGDLSfu11XCj/DFSnmE5
GomFCJ5gvVRKMgW63uTEeLdRdnOQZ6Pcl/pZo2qa7upKNeoaCPtsN+MewPu1qnLJ
CJBosze9rg6k6TOXuLaPEelYal8wyWhwxYw6m3dNdlzzaQ68ljoAL1RRXH7mLM/X
MCqF7KWUiEp7gDzA5xzXhgW8VDNYqIliEfpbyzQ+pI7sUULzMaoxf6Wc90o9+Amv
OZETX0WzuqWzKMgLUpTUJcUfoBarCguRHXf5i7K7BUfvTYLji2vNPWvXGCsP/gaV
GeH5kn5Rf/okdg9P38FXWkpbkzIxjXexV4U6CDSkpVGom1BDgJNHarxOGWqhq9jE
dR2E5wg3NAgwxvPVLG5LY2CUKnaLcwj+pUQ8IwYUZ0REpVYyIax0rDNr08HXMELa
wkrqEQwqjHNG0nKoEmTomLTfF/vnBYPoTC9vH1R6eO6PkT592Ng4Pjao5F4mHPC9
ghfJRXGSsed4AES9QeFMDULhUHune+47Ts+vaZ+yGECbH4WmG8ISVU16gx11j8nf
+8bphNEHsBnddC/y5FTZV+Zfw2AKIWnMrJHjvedJ8LBgMLZk/3WGhwyXg9M6Nr7j
6JQoV9xb2zu1PGLT5v6uQufz5/THWpuf8hU6WjlBj+Bfyfg9eEXwI+A0W4Oa6CET
H9t4RiL3+VYAc1oTFa8SUKd5LBGmSTerkileifyPys1UGVCGUgY7/bU1lh7fFMmj
0t/SOL8BdHejG319hW0gIFRCZFbwp8WwoJ511rYjB7l7/bq3ZUxg+dRB9Mg801gM
ammibsUSfXfIN9NQD4mLEaEhg1XDikek3Uw4Viybcj3gX6+w0oSCPfaxIpD26/ZT
LjMnulTZk2/CxMrRDXIfsTtXefRMP5Jsy23mx0Y9u8wZWeAVbttcJgVTyLDedzZF
enOyx6pQ2gX2iK9KBJLP1N3aE3ZkeHEsn3XQmar8X355MB2cvAKJNomVRe32zjKm
x6cCSP54hNfPYdbO6rbXGRsApgvNqETKh/nlj2bPgBcwpL4NQB4NskjUivNKy5r1
3UsxhBd+qzzncuozAIjSmA795YSE1kcZDTPruybk+I/nlsvvCE896rzitx+sLraW
isL86wW6crayMVEYkzOUg19UdX3JgUnVNOclJjg7E7I7t1rfLBqjUc5Na7ZH3MTN
OMDGKKeVH6gz7am08kCmLDLnr3GIWTO3w78cYL4h1+pQnl8nHpK5KqVK/QGZOqbl
5VMkGXLDtU8Ge4y9m2LwV2Q8MkEdicKc8cjvLWXtTpJxdzKvy48bBR9QooOOTGw8
LmC4y3J5zwkJYueRilB+TYR92t+ALDfxBEuvGJ0nz6prG7k7dvZojvM3CbXx5MLT
ttCAeUmH4d4NMK/Q0q7ZbTd+GiJaLrOAN7MXEl9xmsFF6aEtUeNRBFf56WgF6vLa
RCkPT9Ef/te5CjL21JTorUyVJiIymz0PQR6xWWzohb5QCHoHM0zGwTQFXp/qQAkd
0Oj8oGXanmwocnIOBK6Rnf239kQlMIw+rjVdGYhGt/tt2/4aN1rWESjSpYCu3weG
wSB7gtLporKyh3U7sDXWPERBFsKBRPczdQ0Czqt5vv3xCnsv3hJsKqoocKlLYXcB
GQC4pCMAMSELhE9KSztly4uGIaM+Eg912PcjPPUH5mOtII0Jo5/kXdfM6EpZchGK
VrMLjW145naZidvlk7qi0LyWgiMDQYNQApyCI25aWYJgJXb3ijvG1DLfufcHE/ac
YeTEupf4wruwb1b8Hhawf2hywFItgTSlrREpY077HnYJDHKJv3RCWVhvuZCUqCAP
LRANRJPrebfU+BWZwGKgMukiNFMFG8ZOk7VCSWNZUhlr3B+jxGTfeEcAvWhX1kb6
lG2jdLvJQk4F8bqIs2soZq1maT7oA5SgJcXMmS02CogImotman8tcJe92OzdfhvI
FqDWvuUvKbnTppWKc6+I83DZRXW7Xs+QuesMXbLkLRChUR4sS4PqCkl53DBKU2xh
/10rAJA725O8ZzVcBG+f7VHGVPAcf/Bfboe4yAFHxWUYSyePVRVTQ67Xic+lrQpQ
OoEKk+2dLgPPCSjnXaNyZEILLiFROH2crRgqAw+PVMC0BZcpyAdfoZm+Uxt68qDe
MZ9bQbdQy73aTs42W08uPExOTkwZFaH4Iha+jppODYCKRGxypWacIm2U/rOCn4xX
Jlvn1ZU4nhyW4FLdMPjn8v4qGOPx14fwNvvUvXVQykBMVmMh/n5aXNwW5i8UE3xB
DwEDHQmAWdvqXdbjf/CN7KDZz9JU6c0kiKPhq//K3A+w39iD3gCb1B8IRWaYWBI4
qoFjKI+3pV0y4UHFNTAgbSyJeo1U6Hkod/Kuoy7Koz9peYKVqUDd0HPpxhnhCHIY
oVm3cnL2j4nXnTiAVm855prackUwZILp+0LHZenUQmIn5Ss1TYXtkXULTN7lBXHG
yrGmKzaiC6TL96iT6Ntu7uo4CjDFjcWXpSVrcU88XyXXBr8WR5K4/V3unJbUnfJW
goW1lzmdiDBNnaJtKkn8F6BXARNzzw/k3Uv++bR1tkUO6v6UVB7x2NyRE8GGIP/8
Wwym+TW4Pq0liJs8aJYCbu7O7bMDoB6Tgrkil6/n8pIASym7ItnFG7H0oUyRg5I5
Z3iTQWwsVundPUhTcncm+TorySvAOeqALqI1TcMrjwkfwOhUYnGiOQdG0BHCF9Ns
W/OTgocO+pdhkvqaY5uy8Ey7GG0847D9NPei7W6SI+MAvr3R6CoshZgbj+skswZN
JsWglc28pKOMugoTpEs7RIiZmCjFj9VunNGR6YHcmEUf9IDqhWpraVe3M1+vl6UZ
g/lYevfAIcqulbD4MmoTePj6lgIJnUTogCTdspexpF2WwgBX/B5yOYCKsOjN8SSt
xXpMRYbt6q3pX+JqRWIwrip9XtC7+6QX1h9/oe9dDjtRwvFGB5LsG+tmwhpCkAiP
pcCHaBzkahiatVViahEE5xSmJ1TbBZx+KBenzepnZCr/kDMzbimrg0o17c6LbxY8
EmHxS1qYZhh9f0AStQ4ADuLy/L0LNz4OtffJISeveH1bHNat9oQFmRH55jCufQr0
/ZxKyHwnxkTYX0z0yahpLbYg/SzrXUYlZgVM7Ef2NQozxPLwSUIkzhV8rCEzs+jk
pb4zHLaO9XoYfk/HJ4ERdpYEjuAWO+tGxfEZpoX8Zuxwjz7QyoHTBVX0dnqPdogv
DyuX5WWnmuVlMlr34r3hgBSxiFQny1icV/YV5XDt+zQRK6wFWeO4hDutv99aMrWb
InwGjteswNyY+cHiPjyVXTbXsYbcmVciCP08TJMJG2+BjPVOLhLDb16jZCV26OKa
NhgS1nRopWfxq2JgrQED0ghsy57QJftTWfDLUAooSdbR+X0Sj5xlHPXiBEGkRCUd
1zKEWvuo3Bf+dPXuGYjyRI2X6Wdj5CilTm2HWonkGqkDZ0OVwuCDG8fW1itVKnli
/zroaFwI8oKmp/YsPdcYiEwQU/TQpPpVqKqd876BOUeF7bA/CUTyUFlgYKM8zyDa
gFfl4jOgYjXpwr9PaRYX6CUdspEJwQ6PScxsQrE9LgLj9EaNBX7NQE6ZPJ+qwJxK
OETKR247Ao6Z6/41gQXsC5oucDr3qyRpFN6L8IAgnMTvNnplnCekp2ENH+YtZjTO
92h66jOy2mrDqMw0tR1Y/VpA9+KAep+gF1ucmPy9HAWAdhiZoVojGlGcL5p0Yh0l
vJUx5w4FYCa/Ce2E8dn/mwaOTjTmMZSvKMnKmXbUmKjzny+u/4EBgU5h37Gx7R6/
RgjpYuVgT/zd4RpA91Jb1THVVrTf5nfTAtLBRrFhNGsouNQMPnhwSPwF0BYeBCMO
8X1j4bo0WCQ/IDqEjqS1LrSTTJyihzJJJ2KTIDBPv2zyIHOfe3C4tz2tfjh7Z7pn
fSZgim781DkJz6hICu8zEkZ4pvLxZrWS0viM/XhihnvRMFjEsC+WWEw9B7SKxVwD
uldcEaKpeV/NAF6Z/K813U5/Zh3eoBjh1VQdSdhAnBccGkgeg0uCjhULTtrWGkAu
Q758I03xBsjAZgwKXyXEXUZzGcUJJ0MTIgPwig6+xfpIIU5vaqN00U0Hgewbu0Dl
gNPv+94Zy5rD+2laiyAPQHUVs/y8XovlY5afYZspJclLMlXiqynunzXRqSZ80SeQ
djImrJ9XF58xFIa+/liePs0fpDOsOBn8s5K9UWbvgFboP+cTkTRGYRhjkfPIy69j
xOD3LjgSlrmhTju/qIsPwA0Sk7yN3QetC8LEcSfYrxLc0vwL4bvtdsLIhUmWM0mU
Fnhp2slpqtByOvL/z6A1GQqSvqkdfG4DNJtZwclIBJIiWrgSbw6KP5eKnWXGvX7V
G/+aJilS1DWRzVAmdz1CueNPvI9J/9rbe6fuhJ1iHBPJo4ZoyVfKurOK3UvbKTw5
QsjU9P2EWqSDNRu2Bz4RHEyCzqNZu+go3JDmxH46LyUdzGH9gYz13VT3x3aLgNgI
W7M2RjXrhr/gF9yx/R8gi/cMXV2sgALd33FWkgXmea18qHjwNgnGo0nxh6BzgBAO
hv37Xf1Rk4HrnYyn+ekoaP+qNInovrLAQLMRMhA7gBrVugJSFNQiLG4TuRIKDPnE
CPhTEa7/fMirM/Vk/Nap90qNToQCeu35P9dx599gxmeE1DjY2w/hi0hIV/ec5D9Q
Qm64v4SA/iXO7+7zBfYW2MU0CgcSqg4X7BmHRnZgBe+pqUmmVH38uD/7A9NYj/cL
syC19xz0mQDRvDWic2ZF6YeyvKkQAOSvSCRn46GWbbDLLTDISVtuztr42B3gijKP
chwOdAUzXJao9y8u6/EKL/hzB2BLX/TCTRbnx2orWq7ZvcjI3zCUMffc0JdE+u5R
Mdt59mWMnYV3ttz0+JtI0K7+wD71Q4+uUODLPIV8bEVGrQBgOIcIftwJc0Sr0aFs
tG5+jA9mi4jW+Iz6NQZPe6WOOTyvJ8LzOtd8+B7dtd71f9abCLvbIgkfGYWXzkOB
qO64DVHce2WnkNk/MoBe4XreQ6WcL9tIG9lMKzGDyQf6IIIChoFqU1BKnUFjfohS
/+FMwkqeVJpHUuFOqCqbLogKxYCkp4MLkEBFwvKf2h/B/BsvtdZGTdFh3MdjjtzV
m2HLXRN5XkyvzH6xMb/6jNbMoRq20V4Vn247cslM+P0My6fCY0YG1kMXmhQ/oVFo
D80CIrEumA81BoRI/8/V7PszQYqGeRI1HYJF1OXwZ16k58wYhe3e+ql3sEi1MpsL
vpGTcyfNbcGZeqkxDRgfLuNALAYIOcv6Aa24w8B4bGP3qwubNApvTvvUS8CH68jO
gb5/23pD70MwEzOvlUPVcf7Hv6ZHq3gRtLfXKMj7Q5Mx0oA8fDjtwYPenAr/yfFp
eq8us44U3vtelVIgGk6sSB/x+pZiYIEozfY4g3zeFe/xhsGF+umGrlxuoMpY/yqn
pYnCJwB70GgzJYUjTBPIsqZGcEchx7KbfWfblk48rKSoU0BA3KChZ6/Ldp6z9O3g
6bb+FdouvM5po5yOwzF0mxhu5+r6jon/BkPmgtjOMyL5jlJ7AE/hWrGGyUN4DPoN
XdcYVPTKamuCO6I8tsD9z8vyKsCNu0s1Df4004jmaGX9p5fZcTUXjFNzKRyOwPNQ
jJt5yUPV6jYAGdVEcuumAFPwAnTFWyzdSWSrKgAhvQqOUTuCVV9tJexf8CJ9L1Lo
GSRRto8+hKSoq6VZI44meuHfuFWJNc/YhHEg0wimKHn9UxKlYJp7576QsM6pUKMb
v89bqn38a5l6I65YtUEw/CODhJ92bnAtTVHMen6lZfcOn6xCybrhYje52n7cRI2I
zlP9nFoSt3+jtlcOhu1HcXOqdP9xaRxXns8/PK35K/XaVOfALA7pFaLIGvNhORya
Oy1gGNt3GMMWgM5Qi8x447zjniai73iVq+l2m0+e25mc0s7QhY/diZ+CseKlIHI8
aob5FHe5my1Ol6jxEM4SFNWjhY6ub/yjDKUd7eipMVaCme3/uTeILlCw9VSI5Rm4
eatKJL9lgsrecDqbm29w//ievXb+aAz0VGVYy+FysnSRSyN59mwr7utL7ycoh1Iq
RIuQT7JrV7M9oSfiV7tw5uAO5nlC2zIUt2W2Q0A3jEl7tOjiF4BAEQXAV10vXsZy
xmUPXaDoyicjXOSAEkZAklt8VY3Cwewd0c07s//rjHg1AWiyuLeP+/x9TdZQgaD4
HMJe3zeD6rM65uSKwsWkGBUw59HDQmxT/OXQH+gqdyV8Cak1FhpK/WcrVD/NOp6y
T8kn0eF5BtsBsgHO33NB4DzKQWynhcXrF+vmtvMpGVXgKXR2P/p8UCX6YPOwzeQS
mz4pkfIFsObZRi+yPde26Ampl/5hRFVMNLkotrC1U3u2Ix+ep1fFjcOHI8vHrU/i
jEl2iKI2tg2uX2EBaFAX19+eTz6nFnP/XfGA8Hn15JpW29MI5oJ8QccdGqDvM+Bh
ngwKS0i2b1UxixFaCLmRcLwJORr/EP3A3rMrPiUo9+oouAIeMQDJHgUoNR3+X65g
wtZSM5jPgXAk+KEfCmd9dX7nWb6X6PWUTllBri0tzwZrjJ3UBcUq8vJlRGdIY+9e
n8tCGmjwQbB2BmWBt0CiNGLWyxENKL4ITnFMuv7Qn40ZE4hgHbsk5euRfErvUwsS
eBdWwv5NzA7NfzvT4nF8x2gCrqmUgifXPgWGwNcC6+GZaXB62WbvhVR3Q6C5luhs
xsU81Q20YA4ZsyEDRp3KhxcQaYcwV1/pdKKE7VG3OV4rPYTZiaNktXdQweRnlB0G
yxwAZIYxgGqAbtLomRIh8Z2MGNJldiLU+971GxOyIkWoIyBEje6LWXcNdvIoqF0V
ILlJ//FftU+OcCVUN7YFh9QODRjazkeGafi2l6rT7aW9N+IpHgnbqj1qhWTckfS0
PHXYlmj9xxu19J2fL3wSBIyG2DzGC4zfBtq6xoFBkPRPGer2ryFIOnNC2lpIfJB2
55FUcbd8y6itOCy3seFLflstdSAbZ2AlTmRmIBiAF9p9ZzAdh46O4QNgZ1Lh0AU+
YHtuGsNgiYhNyAyMQ2tmwnXwFO82G/prlPRAhhT6nrfRdFHULTYZZjJRbePzkKgB
iO4Y2ULF3OM7izTWXT+tKz3s6kvzaRMpMQEww0tOCeJmkcDm0/5JkPPSnHV1MpGJ
Tk2nRTcNE+QQAxKEA6zEdsGEpR8shI05tbaviXZ7uzA9p8L22YORXV0UNFrskdQ6
++hkSyXunF5DnmnOHyYiakg/2vpA02w74tymnsCEg8mJnx6rdgivl/W9AxXb4xAF
RmyM69MMvSGX3KL/gICCgF5sXHfx2Hz0/LwK8DQAf3O0iAb6AmO04mc6RDakz78u
gHVI8eMIDcLVgQZBS0IyPFI6Us8pU0H7iv684ACaom58Rvrhk0ZHZSI0kI/q4/Od
UuoigStDYJmgwL7Cuj4R7XVBUW5GqDEqSdzEwv/HCetN0Twl4eQGjd17VoAUbcYc
H5CewBZoYlpwnX6WAIvLyRUQbLHJdqjt3Mz4WnszBK17Frsk3DB6lABpSf7KbVBM
qyGFbxljvpTvOLJwAPPKplxR1AarEAc8As76938EHUYF9VYcKsQm8qV2A+k9llKy
I2nX+y6GN+VRTfZ96fb0ygc0EKLiKv4K+uciDq11lXs7pxe56cxTErDlDXmwktXc
UT4ZrXDNijvDkP9SIB8rxAQwkCRi0O7B/yBWscdtkkFI1ZZyYGJxxZy8yUrKDjOR
4v3zWWap7YMncu0s7uTjOxv5t8grycX4BOjDmciRxlPNrmAUq762zxtndb64cdTY
249jQF3jCUKApHNMNBN2vxzZVTqSn7b7rTYqogTkJdd8Q3Ufjc0Tvj5fvhFjsFzx
qy2Di4ti5MoF8cI5kney6SVSNlvOuC/gskHMIqxGNecrrm7Q8+y+noZUKFE1VcXX
+zrSo+C3/fP28hJfoGfciLEpSxRxI/EjeItpMAMJw0ljoT4G5IMQAsnFgi47VC/d
q2l1fw517Nl6GF/6tXC7R5BKNEdm1n51VV5NOgGj3cJe2g4RM6cN7NZNPJZYEPG8
Xoixy8j06HQL3GBq0I081r4BQQ7BMzBkLfOWIzYeohjq/1nHdVzbeitlVM81n0+B
ZZTHAd4zdYcvOEQST9ofKkU0/5q7AvdUSFLPhqADdghgLoaixqFdHjDm1+hCzHFq
V2YsnfKEprW9mrGDb/TOjmL+Dni11Hz/88/pl6SpOItL96ELzdBvWfNxiEqbnAYx
Bu7vyx/j2cjEhxZGMsWHLKhkaBYmfqCqdgs/CnAWsuvxdc/CbYcs+X3KLUXiF4p5
3SvZaI/50Xe0PwlML1+me7k6L+fFrKRhFGsz//qo/xLEgvnjF47jstdITP8HSNrd
NF7HdmKzdhAAmwm1DBG9gfeY/lTSpMWPpmF/t+eEpXmgvrItbIIKCoknnVmwrkl4
iiakR2/L5SeIVciSDq8GhhWB+RCjXwh6j2h11cGy9pjWBKdHpB8xBrKBxkoqJobo
Hez7rNo4rXU/b1rsb3qQgzgCY4knXNaDQT/ayp/haLEdyx1ikxovGhPLnyPcNECf
BjftMjlVwGUXXx7nqhJr75o32WDi7BHeHmar2iV6Gw6aAZZVI822MAwFyPw/G7tz
TyxiRZJXOaMNdzZpVEB0F9BgyX0yrktjmRBk8BqYJBpAmDY1Pje+IXPJ9xKYzu+w
qnAq0H/6BdR21lIj11pfb7S8XUPUyVU4JPneSn+V4G9qammxMmjSzsNPYAGEoZIz
CfN9McMbYC/5p9R5huW7iOIusiF1QXOsbEM0yMHDaUOkzuwdFzouagtMw1EPLfD+
lkArEitt9kqNfrtFmT6mltHgPS++fvDJqljkqpIqW6clsNLh0//1AZprh2+/8eNr
N71DRtErpddivWTvr0pX0cykshjnJa2bau/34KsHSl4bHEhIJ0ev2DtFGqIkzXXh
SflLNSFTqCCpr5Y+krG8F4KTarcWG9DqxcuqjLXdhw4GYdsUi4LqnIN2aRaN6cq4
u69DaUIPwMKs2a84LYwbanoKcM8Aa3Fe5lq0UxP+TOOq54HLE1g7SVcmNawqUmP3
i4RdNX9i/K4UWieJW/72OleAQhkZXcpxiEIo3D+zqYsvCC4uvGqQCww5zKGJvvK8
qeknUKXIud1NQn+JqoWqEMMkzNqNPADyAsOEXNEuOmB3vbc5AjexuhPDLahBQCUk
iANSkN0EB/dWBM/n6SWWwCNW8UQCSyxb3vbDnZ+pY9Jo7Rng/N6lW4wxO/nfwUNk
JCtyjBQ1GNRaqL6WJ4ASua6b0hmIKdkCKCKDtEYR3ZRqsanFN+vD1DMUzBOwSPRE
1wnBo/zb62slX1GrVOQRtg41loIOqseUJIXN9UDD6yXeBtRCXhG0HjX1MefGniFS
G6z2CJuKNDEuqpL8aWMprjaPUN7jStZV9I5N4lwMltFyit9Wo4r5d6WTBPtu5rlz
TmvzVAWGfKLHKfUa15zPVucnYOC1rukdbXeGAWw8CWJ+zANG36cEeRwDLDKPQcjL
CCGomGX9DV1QYYhbPyUXRB64pmN41PV9MqO9V+1PKzUIZ/hSLGAcodKsubNMllZ2
cIZxybC/lc9YDqOCe5KBM2uftxqR23ShHnKRXPBiramcz5w+oEefIFQMu1AyYDS9
HCZNM8IKvnd51fvqX7/i5U1rv/fLNrCH/nX91lZAqsgz4OcchZfHH5YDUgQyj+bW
1MN7rM1MFhJBeniC5dNrbMIbOaneIbUlexR0LBgk9kUG+5wFVWzzp9Z0a84/B6DQ
9W+q/qhG8TK2cOC0dTEuxOWpQlGo+9/UTy1I5aCLL/M/vhbQu/PeblNs3k6lqQ4D
aCFHGGvUIXg5BelQio/mqxpRDiYAk9NFJQHYgfftHIOQJ0jZMRbzrLdFCzP2DKz9
UD7+OsX0ShMRww32eR26uXtpfIPNj/OVOA61Ou8Rheh8xE25tK9m1+pYj5wUw1ba
gAFpbi4voHMUjDkV2HOEznD/8yQDFoH7Jmxm/nOS3oYAovx1EbfUAieAEvtzlD6V
ltqgR0cct+RRvWrR17N1Gs3TyyLqm3StlSxq14b4hS4Ma0FffyY2tcbuz9/iaVPk
hchExw1vWzyL9hrzM3lpnslDrOElof4YZTVGSvhipXM0RWdIv3+DJ42Qp0/n6Uuh
iWK/7aMc8neOe7/Ix218Hb0KYSzU2YTC913JRIKwCIun9s+bowfKyZOpfoGBH3Mc
y2UjuVLFtXhdkMMS1nfsVa7lDtlKNVmXNtFW5b9e8gAJVkQZrpKSvInp2djnI2tc
ow3Ngsh4c7vHCodWQYzPZQQv+aUmWO3kF/RAZBYA/yU6CclRiQJISys1tGx/vpKT
A61gON/ZNsA2RMbNQKPW4nU0REkRY9HsZEadDAXaYBLLGuA1efcQZzFSgW0zoeUP
ClX/S1RiyhqKLpanFE0vUrEOX2BBN8OTbAdneXU9Rq4tQ+QO1JykVOPssXnySxBq
zOUDscCMbsKGlO6WTZTqsOoPRJ93mj9+tg3eMZ4Ni7rkkE3/HEtm6pI2/OBDYveh
ixm+J+5ZDTgs+kJfJDc6aJKHHHp4sd3fNMQkGuYI2zo9rhuen9uY2pNh3zsWhvRY
77VAAgEI/GUFSbPdZscYlZBl7Z77Nbz6oYlJwaMGmx1ABwX8ZWxZ/B2Rbkych73h
09j6No3V+BiPoVq8+n+x5dtsFVcvjTYyLdY1SkT7Y9l63Pj9zKnQTHcnV1+JeRya
bCsQ2GV/eDf61XBN+Jv9cWUo5JRwoVYK2HSrgCdpgiQdO3OsdO2GYlNlgDdaCJpl
yjqD3jgrFoOBMWok5o86zdzBCffcetlg0140s9YxlofmMGW60oKO3Ux0O0CH8OIz
1DYFRwIjm20IPXoPUcBzy//Wc2Rb+R2FEkrpj3qJ4oUQbsty3jbomIHjQk7PGA2y
aTqNZY4QXYvUtagJUYMHBYBqgFt2i3K+/3719f2MeCHDcB/pOehzBWGO/BNYT0y7
+rqS0StQZJ0+W64+zUkyUinjp+hXSls+2DF6rldmlUndCYDk2p0+YyAu+NNaShok
GBCmznQ2WQf4vfNMaY7f5Ga95CacUI3IVCZD3lWOJIPG59vpGRWux8R7c+9vmJj1
eRhWCyaOga3STrJr/pyHJ2S8SxQ8aoN1iXfEca39VmPuYN35WF+uHbniNxZ66S0h
JLb3befrStOq3CVeHsDXhj5c6YAX3Wb2DT5rCPrqLphB+M25AAjeRD/J45HX/aAM
8TV7bEZBtnPUi49r59ORglHYPFm/8ld6w02fIbH6jGJ1JGM75eUJfJbuFLkijsk/
vxnxwzR7PF/RHMNGRVe+DId+v5LCvo6UKtmLpS3JsKFk1Lw6x1XxnExOoQ7vhEDL
fFnP1uHbAdEvKs3DQO1Zax47P2BxOlT82qpys2X9JroBtUOTD/gqKsSS1ycpnN01
YgOo7t7n5l4r02C8l0R78rIRqA6lJNTLOek7cUZKD1UeTwGoH4uwD2a0MnvzXO3H
h882GE2DsvYgH4oodZfQAd1c7zwBAYpUAlF9Pdt1AU5djQeR4zCCrQOYO0wBO0FS
mNMplzk4nxfZzelGkXdukSMlYM92AIVTGiEbhzVjAYp1wmq1Z9lEgJJUR2uhwCu1
LQpJu+4Ln0wdXs44jEPzteyOtXmFsnLroIdcw7Ktb89Bfaz5CIMCGdAFErJG/mX8
g1KSkQve/LidNgI7iXKuJWO/BY94gw9yLMMoysCbt0wBK8QRI6p4YJ5R93+Rni5v
JrOlWKQndyAF2g4Gb+yPfQET3nu5CoDJjQrS2CrhTrPiW02uiry3M/l/k34wCPj6
MN/wLcXfw9vIIv3WRduLFW1PyOO6s99O0pe7eBH8Pl3Ur4CKddWiILtzb3X29sC2
KiUDlBgu+0+FBqWFcUgz+gfdzy0ugvbcmLloDAIYEdbfgHO4qdplnUDrsRj7zkrH
G2vqhyr6C0zbMkwTLxaKcykanWtYpfz9pLTp2oej4OTk7bdMovY57XnI6HKnggbz
Z4Rv+TAirLced8bakMJ8rSjcceAl/HTNg6ssNOqbVVuO0B4BWdwc7zv/BPb9St6w
yaVo623NrgaN3t2oZ4h2x4BxnPUzVAHY/7BHQ8YnCRudPzYxf5dUwgKmqiZLtKxk
QfDgiz5x3DIW7ZUqCu3G3tpCPJQan468HaqWO3/VSV51DjxC9uusLBOX31CZYZzq
lzF46Dc2fG1n8lnCYZdlFKczq9XhVRJZsLMg3fZvDNnhY5zEuShS6+kToGQsv9Lv
nZ8DiRwM2/yctL4uA8PospJ8L8W+Qti2Bm7a4HMJHG2p68Kwas5ikovbXjzXnFc8
CL8hxCaHohWATAvjfisYclKq+aqIY5YX9tirojE9dtGL9uoadlwuEC41rzq6GPap
3RL/5kEFXhYJPirK0Yvn12YhyZ//mFRugVd7I4+n1etG/cEerM8UM3bONDiFwL2K
X+44mZFRHSqxR4lROCLKeZwW/BVO/OC5kZS/m79Ge1xpiLvxAfVjJDzMtDbIIN59
UEKhgx93hSgIkRta85tSvggf8sNMyrRu/12NW3PQfzF9CsvJQdaMf4yKa1Zq3uXz
lFoflLVhPTZbp+p56FoyRzZBRr6GG4qmEhvsYnHFHgOzX704k9fQXRo7RFV+pWhX
tBCHkO3UKXHLk9OXVv3g1av30MHvrBiZtLYYENO2K9CPAaN+fTpzqqL8NW8eUaPa
0uC6F5tcgwswVaFaVq69XKl4naiO5BdiScWK/WcfgJgMRiStJlJZBMxWvjJ2Km/E
D7g10PiyEmUwocfSc2Qqn/GPICYOFjp0hJVBxSKGpVdr1c1MUqcD6xqifzuBV4Zk
bEdUfapqjCz6dG2c/U3hyrX7/B9E36DCmkWjqkNymJNjUbAy7FWK0lEChYGn04YN
hjiIkXsDLcZ6etKuRMEmCTnzQggMumB9hud8GkiCNZp6f6muuwI+kM7yOAwr5gHo
bauda85N4E4Aq6AoNUpRhOzl0hSz8fH3p5/NaRB9gmVS+c7+vml3RhZptKkcNYXb
5lVrUchboq/8CXNbK6eTiR7RgGHBJqZv/g9oF2TU7RFLj9XRAiPwE4zJCEZTobfx
lCC7V5ef1e/zJpNGOtheRvxvg3Mky/Zz3p8BiCk5ZDKrXJ4ppLEsWATPlE2csyI5
1quVfwAyBO4AExyBPqwdAFuXInqOSHAFl/e06SO1MFwPNxzZKAS3TTIZgdzxPxWs
ynew9xFw5xMhJuuOSSL1xzCAIGE1AlSc8c6M0kRGyrO1EL/IKX8dlFWEffccuUNR
D6HgyoQ9dUtrHrXsUyLFXl8SvMWovTh6K+cDQJtiECdG8QYBWCF7EUQf4Ut/EUiI
6huGaB60HrAFvlJ5aosSczMezJviMMSbxqLO77WoFVNQzEY81+6MtZCMAOtj7GmF
12RkB/1ZNPgbcKLEpEh62IuZrU79LMvicA2OR1Wvb1n/i25NiWCP7WLjJ1ziJsuB
pJ9dywAv4PhLKcTmYbMLBJl2anVuRnSlP4b7OJExdKyKVkc5cig/1U0R+qp0ewcm
Ppsq88CnTLnfBBoq9mFpvSrgKpg3JK4b+q+EgsOsj7g54TNTQF/9Ckug0vBMN3i6
hJQyh6OFP/+rpwmCGHetrG8PniwZ2MK+mRC3NiBtAkLitnqxARkviVIykhD9WvXy
XtdpsIajbn5trdP3uj3YAVa8hJl85HvvOktRB7e44jwX/1pf8CuH2zIhRL+llM4W
1UpLyjCZ9spsOKCJkT6MrUn0mgy2nOngX7C2DYQLqPZwLMJ1dMBHtNYGrvKnr/Hd
SkXjtOPYAFTDnV+X57C7IqpY6Fl3ZU4vt8LvMJeQ2GoF0JjLEeUo/TaCeR2A3xPu
IVTpTKlTjn1OO9kWuC9EChmBDWyGH75WYrHpB3ghv6kHuALhq6otFk+yegi1HZkQ
4R8VK/kT2rjNH83zkl1/GWBOuADjKsdtAVlDsZvJAm33DP5PQKQ7ePhWCfR68yqq
/z1NQfuaPvp+bysHHERW1Qb8O6DpSQS4/9VIJ+FH386WFo9Rxi6e/jiB0ble7+0t
2Tl+TEH+tNdd9DizUG1UPsBDQ7W6e1/roElHTrnkAKcYCx3ZuRBonYM45AWQ2ve8
bBWxwHtSVIj7hhEXhrshA3u5bflseyn4+Dc9jJPXPXg+8rCVZl45NAJFQiQWZWfJ
IgbS3N0N1GLvLD1vtAn+l/OXIAk31YCQbyUiwkhMSZgvIMTu1I8XN3s4NToHCoOc
GFFoqiu/c4oJ1ulQXYEqxqOMcRadunoTTrk/zm6BsmIpdEzhWrISes6CCyb8sfXq
a2qmVbVW7BaICe5ybJtM1bxMMHyTiPN4DDrFOCQcTVzk7e3hkdRCgSuq7e3Yqr2z
cDn3dCtBFBDlZh0OSOSfPV8Dm0xppqN5hU2Cb0MoEbzh5kYy/FKySPxbyCXeJeJK
7NNGY+YvD8LzWJFIdpSF5Fqbj7pIwFvT/lDGGQxiwqttdk4actgYGHMvUKu7p33/
g44xE2q9oRAlLw835qRL1AuZeQJcegSGTYfB2KUAZbg5rRICxRrupgRK5Q+d7558
HPGnhxSgeYjpmV5CuhD5k2+OO9zqMvq648ugpgeFqdQ/w4EDX3UBiBA/OR8VrR7W
bQplX7Vfqis0TCto18AMUKKMlJ1EoyvPBZ57h/Uo/NUZeTes/Y+PyQ/6ssRzhTA5
kAwMQjzE1t+NNnuFAh2K1vPP8GWmA6nWlfjxzNxZ0qpwhWsDwQUuqgkT2YyOxpNA
YC0dL26mVu/vUhHzA99cxHJ4u2RyjY/lm+6u8N8DQr9/zq+NFQ6qNI8FPpt8SQQU
46jwAg1Iy5py5nX9mGKqpz71XNtSLLw8UMXc38k58jUXBKLbKo/IpAx8GykHni/H
Tjkq5Lvy+6jKXqzUhUFZFNfwQrELp/d1jB+5F0EX+lsak2JgcuQA48hOPY1Lndfa
512vsETBVWbvPCDL+uaejhqYrSCaFklaape+Q6dWTHCkj7WDID4L6t7uPFs6Slfg
ZVSIHDN7+awUIJpX8VMOhWdsOC8x9lPNv0DP6JP8OYeDKMfqMmFUZTxKEBNxvEko
JKZB6tLM9SULLYViGS8FX1lQNd4juZ/uIQ224M3HFqUDmJnrSy0ivmeUqJhQ0ScJ
slBecaGAhrhose/lymQCUQzLXByBqcKCSbwY48qFDXTgdX0GI7+8NMB+gOXL2uEA
kd8B4ZJWYayRNQNvQdA8y1ayekICUj8qUmNbprcW6vtDn8vcd2AMFANtyAq9wp6C
qrka2SGXAR1+yMsRtviow8ma88VvwHQ6lpTpET4Jt8heqXtKEwq27Tr3R595dqR5
SJ9dz4btvGLCGPvhamL4sWXS/57p2ZJOqNM9ggDQ4OqN7QLUkpnj93FvSYG42S2h
0txa7+BE9s3uWL8F3tvAd2CjINVcSW70MHCw3VR3dssWy3h/Ct25EnoYRM1HvmBn
hnNFhcWuqFiE8BirE145/pU9iw5Q6hq9ugyG0gYuo0u9Q87aE3clpKlMzTEZPaL/
nAhgENpizgElpJXLgnZc973LFeK39G2FAkjsydsJF4S1OFScn0woJPCVDHJd220Q
uGJsc1HaNOjpqUdHc8Xq8HHUcL9RH1h2MWajQUjkB0EVSII+8J2aY3v/UCkQIS9p
TzF1wUQqtyw8pKQSBhC8gMDKuApRW+vcpnkT1wU+lE8iqRsgrouXPSWW5MxqKG38
vNktLimZgIDp3gtc1gZVZ46EhTvMUKbTuZQsMgCRfStu3WY13ubO2iJ6460SSQBM
FPtssjO/ath+phrIpLKhFAZHQBB8Wqe5msJ0eN1PqK83eD0HlfrMN9pPdk1f+BcR
IFuP03KUmuq/H8XDW9y959fcZlQ5uCGo6J6yJVb4oC+ZV9Uvg5AMtGcserx1lD1K
rWTUPoJ5zLE1mqIAuWqb8hfI+CyjpmB17kLb9iaWjtGPyBbu1FDfh8+HnE2e7FB4
sk9ZrpfxcKIR7Ir9radro5d4CnWgOVhHVh7jQoN4cZgokcVvQ9TD1mrjpHdHB9Kz
gsXDV6M4C0FLlLIlrLNTEvCDhOgEbrPbPCd7LHRxP5LxRDp7E7BW7fypvzfCjZL0
tTUaXADr32LeZ4pNeIk6iuGYOKcpXsdJCsFyQakYOXTHZgV+NbKFsax8YicqoWLx
YxWbFf+M0tAQN5IfB28mdUA7o1hGu8cXdcnkd2WeRG/EcloIrJfWPqM/Js2Znf97
wKldwfm9XwrmlNyQmn6cZr+mx3sm+YcMMYIgLZNBbAaHtju7rnY3VmoRKdnTbsoC
B1IEmbZNhzIABmjWjxkG4ZkSLJ5yyojDDZ7tHd3S61sWESgT5xPqvWKkDe5o1iZ4
qRubCEZWQiH1n/VEpG0WmVfhnOMQvLld0JOmHp1+NeG4mSnMNgkArLb9bvfJ332s
dtckoWXpJeR7kZX95Xv9XMh8WTKk0H5QhYdsAwQhWRgFHqMuiDfzi3CW1xBzEPaM
+KlE+0lp2KEzqpUxWjgPp8OZFFJexGc+Rjh+NBDYvkDeRySfm7T3hz6A4ESU7jH5
F1/iflG6Ag2Pe0RMzrnOGcWwoJGl0iyPjFBlVjiwzGoapdb0/KhAlVknXOMdBRfq
AYHSh1RgyqvwKS3THCgoXhR4vl2hIjMTBePNqSzdhGkJnO7kgLm6/P8wKJGslVqv
5/RZqJUi5OJXCu9vJFC/ShMRAyqliSg8AedZAv/5JDtSUJl6mdixiDwItNZOmdE2
CHUQ0LqoBpyLv2JpkLYdmrd/4BhHnyhnd/GnMdZvk7ljWK5GI9CqEax5qsnZOpFy
6qeQXW3d9Y9RNkZxzLsOdSvv8oDdTCHejOVI8KCRrsaSZINZRu8Pau/+lLP4Sb+3
ldl3c/CW+13sIk0G+BVjL/3l4RMr8G5FIaoHoKD5zhmv33jEcAsTtkjUcigaO9Uf
ihMn9LmNmzxu73jrGURB0siuL6k+E1nYIfcPiy96pUOY9L/CEoSxOWXLOPDpBFhn
rBYuqeBXgxft062yml8/ESaUNzwOiGTCnGfbEb1u2Vk/cX9tWSFZSeCWYQ5Aje5h
BlGOfJlcMkyPribvT/dmRTtKH+LldWACbO9ujVPdIVROcW9Fzji6/XVmgxx7tcZr
jqU0pyEe2wBcasIrRsCBl2kbmal5MrpzHXFhH0T+5R8Ot0gsdH1mgjX/yBVEomta
EeiuQHPEEmFtMUVF/AmW/raXZwZE6doR69ygRoGHBqp/Vg9Fo5d48qy94mn5OCYY
2PPAtBdtbiQzgv9kuRx5h3KRmODCpq+Rn8FBIVRCz6XicOi3boaJHgNZUvMsysuY
3YgZ9ViOceCNccq7p/g15T4HYJ+7ZUCU1l3voHaoG9mMcRoGMjP/rtK9AbD4klro
8FM3s3AaK6AiDW16bl6GDVQW/C0hADO30hJ7O/V3hTl1l89pHNAzB7r+DDkqv72s
KG1si33EzxhBx6I7G85CknSVx588or3u8pO2PFNK0FLP9waYHL1254vH+HSvI2RX
fU9zfN5gXWv+WG/fUsW5i1y11HzmU+ZZiNgLpi/fJ4S8lqTiiw6t16Mv2knNhncO
V8QtGrQpCKHJ3wVFf8bT4i6pIohtT3NGBh+m/JVX2D+dQp+LehZuL0YeS57V/992
4DC2YxXTzEYA3iXBR10EfFPg0vHjjlz6Rh5YPmKhSFCRnYCf35uK8i1xtL6y4EAc
xCrdX86l9lYFTA3GnxYpoeIyHEDs8mSnxABRC7R/zRlkk5S1XHzo6L2qmvIuNLDZ
W+TvZOhQJsTPXE2SbxVS4pHdjN1T24QW93qcA++vQbjrLog/vYUq03Xcv1WuV66n
AzSrdRVaWYWYG/R29bSCl8veF35xcUj5gT+0axXWgm+mbuQSKeYpNa3YwsnmsD6V
TttuD/izB4gfA3Fjcc0tBoZCZ2pEv3IughOBFW//bnsuO45rqzm633tY/M3cKlRM
7+hTX8wONJUOiMrtXUmZNyI/Oyzj9/HYImLDoOdENm/2O1TnUKOjsJbC7Kpc+HHV
3sFLkkqYyWHtVm3/H15a2mSiiVf55XP9VKgZKuc18VJuZzAx9REEYplszVNAbu+O
ff8PA7KUhUJGPChxn/h5Pe4CAThByGYt/gf2ZbR5UOXCYFAgEy+k58/+iF/FfbgP
3DZvxVXNVqYkzktgz8K+gmcvb7lEwAQO+gELx9cUnZomYkzpu51MgOI1yLH68lqF
rDVoZGyp47YCEQJ++GTjGuixD0b5ltVu82wF8ApQBPLvZAxyoB5E7yFmVJSMuSTY
u5i0VLBYH+UHU18Sa9CzP+/OgzXm2NLJgUSaQhgZ/dmtCWju/ce1nBuIcLO01yPn
IIUhSPb1n/CIVvt+YZbJYXZsqIJNUhLSpQJ8nlJ4h3XlEVqADRP+MEvRO6Bh14gH
vO6+ck5j61D9tPVxOoYpBv3iA0jsKvAXeyA9EVpm78r79SZKkhbOHnoSrCvxIkHb
H4qyGgrHfgSYddmqqDRpp1jNzGlU5k0w8XhFXXXhsB+hXjLA+NqhKH83QMA4boNc
Ne0eQTauGfmReTE2YuVzf0qPUlDmZYzqlmcpcX+WrdpS01UaZ5hpcGwgW2pjW325
zN64vdFSgtYX91OpEVT/3B5/ZW/MSAxedl6H4zVorH3ZJo8atcJ79/cUDsUlPEik
uadBmWKitNhV9K1j4DHP92oO5ajVQW7N9Yqkr9E+F7tj1qdyJmXQa+c4RmNIMGst
ceG1Q1QkQlFxB0NWBv+3Ho7iCf0L9D3cgw5WLd4/CqGHw5Rme3tP/+pXeIh1nMJM
ClyINxjFOM7mJFJEirYTkom05Q9nIjT+K6TmNsq5W/a4RS7Sx0IW+EzPdoJ0lJON
oKIcIIGLdGqBYxv8uCPIRzc/BH0DKz88nkaab+3RYdY9hT3m9bhUMRLf1l6cvHvf
nLXFnn8BO4FVdOpi56NxmVXRe62Ur9a6khqvdvUGd9Wh7XKaKDJSuRt0b8EGHUxC
qIpMQYKOPadE3E++WBCQKcqd7rIt+oDXqVZcRaNyLnLMZchByxkyFdUida6HzZWU
ANxfTU+vxDdsKEOxCrtDoEZX3xCpsKL/NUcqYlfNKgh/eYVQGUnhCt5xao5+PUaN
DzWDbGaRa0SV1fX7MgNyc87PcCX79+uudIwfg6WCH8CXXN8X0mNtT0MYOfJQ/Nlu
mD4oDCOAHnkYJdLxBA4ig/vWt593yPRA/gTi7jEc6M1F6/PKY9vgiFME578a3eaW
i3gs9MAMVqjL6Gsv/nDxAVgrdBjk3195UK2miY24pv3zRg9vRFW9wYlcwhe8MnY1
8JVLBqLcwDOtEyZqHiTHq2YAL2r1wEiNbhYGi0yFygmORBaKzKD2A4Jk06GjqaRP
cT+8WtGBxadKuvd4UymXik43qEBt/9vavHJ9dOUPEcruJ+Xh26fuBnWWgbqczhbM
zPK+wNLnqI2Yrr1jd440EKVyjyuT/D/+tibls0ygNlyfbBa+ibLRGHefkE+/znAz
m1CJFmRLm9hJoMLKqKk8iN2vemCa73Ej98SCLh0SDNlb33wsXv5PyYBJaNl033E2
CgAlDnuY7y6XTPunPwR8jh9x8m1lStEy9rbzZppnKJMqTEsBtCegA+tpFFkDjAv3
i59yJ20uU/lseTLUyIJl7yVOgbAYdTRvqxFd5gUvNtX7p/U0zRXYFi3zWczXXNH0
lvB9UjW6HNTSXz/+ElRKhT4YzImU+utjm7/UXg9HxE2e/9pbqd+RgcIcQ5mC1LPn
eETd50kk3R44Tij81e6zqKLMzfomTXBjWWiRcExIEW3adyYMYNKBhzdiBHbnF+07
4i/fbSIRMUeSRR3tLNSE2rFN4e+vqWP4+xv1JE2oANtJAaj2U3z1L5Q1437Eif45
MMQoKJxDpycJvpwu+E9vLxPkFnbmGuXe6jh118iIR1ZkZwfHs4Kpug0k4t73Zvlp
acp2HNSTDMC4VZJBvzfPs7Czj5Crq8WrQpu5IJt/rDypEzNRyICRsREEUTbb9KO2
vKqpS9ezCaMq9g+YXV9+8KmhC1S/TSngIqwVqKXmdK08+z6LbFbeBNTPqx6tBh3P
osys6AweawVTx9qWI/Z5R2HbZEAkHH3YeYjFhuL9IhhZvYT79q3+0kL4+d0fArVj
p4iiJiJCXKO2QkX0VC0WMtrZXBAdw+viSssI5FH/F2eACaD0cXuQ8+l8IZzFJPqf
hsrkE9bg146BSgh5Gokv7RNGc7jtoeg9Ks36pMoLJ/oPjcmoh8yhCXHRMGXyQU0F
5x+I8Om1mzGGaCP64P5pyo/pMY0N7AEQu0Q0c/lDkcoet/qqI055WDmHyJgWjFei
Jk/DBEmnKqIQtCr3YCmnhA+4Drx+bl0DUDLM5luvV4P+hnBzvBxpVmYFDIS/7rJB
nEuEVNpaJaeWsgLYxfZD9BMdPAmtIbUMe3fJRjvvrBVpf/1hWBMhoSdjEwI5W4x+
RTlAqX/5CqZU4xEY69wb19P3yqrW+PoDjKIw/a/TWKA/BRnHkic65gH6HsYcO3yt
oq16ZQtPrugEgkd9VRgRaDLS1Lu1mlsdNEraOYWfozivkmNejg/Ypz02R6o27Tpv
zbM82+8PV5KaANoeH2yWAlpOJDd5F3mLmDgAbx6tMLU97ewEYMkhZPccTKWpAKmD
Lg0dqtHLwnqmO3eiRNW0EWgQLeW9TIhziqaM8j9hIV/15TGAKaJAC2gn41LaOPcP
5+RMdNy8y9xc2MZa0IlhFS0GjIE8872WDzuq9/BkdhTu2PNl8QSc6GL+//8J4585
fCC7DtLOCsQ2HBQQsL/cFcy/ab+Fv4gMc/GTGS5iGCyD0yn9wBySXRZSMunfg9CG
rp8PE5Ay5yGBdfkA5oHHDnZDCENi4Lt642ldJd91BSxGDqmN/X9CsshO5MT9qCdU
BiBIwdfjJK7D6bm5Q1sxE/t6IGB7oNE6dgdnNT7lyEjbu8a9UAn4nGg8Uf3klAVn
nArFWmcPq10uBXjAF03/yAASEJVoA9HRGCJCM/fkEThXEZ/GOtlXT4L325ItiNxN
FEKrrEiJ9A3HAOr3H9OrhdgHiMQ7xsrq9EDEFhvg3hjH8u3JZcwPYe9kh8qcBZR1
0ZELdtgWUAPyyS6k1uNGOnsMJYcpcfAJb5h6Ni0XLDJMKkjXZ7BLr7LyedL2LvRJ
dEi8gRpeehKcrv9jhIZzR9A4lJ/k0KSrdRoHpzEmDGK1gfC/vtrNJQLnuohWuHld
a6rFNLInG+nI5sqOjY+BMK7hd1fCam1linOKSkITcZCLOE/da2O5uv4iiPJ2pBe6
Cj+DpijnDV7Wbv7ZO2yU+5KEQOpOZxzglh3Jb9F+duKPMe/cWNBL/fhSsB2+c0qH
VzS+GCU18AA6yB3tstHMHGiLHiNHgOKBP7zVvGnSW4/MbX7mvVLhm/OR8m2DTWFs
zumVT5OMDjFV5fZsaF7IX5NZ2yMgMJudCV1FLgm9CalqSSMlO2JTDEHMTju7d71D
ZNVUuiZnHd27oleSd8x4fz/TOFSyPwFHgHIOt4ZFl8+P+hU/kTMb/6z5n+LGRgMc
aQZF5HHO09iXkDkxyd4fkNRc2dl0UYuzMPwODp1N1XfVmEkZUVlJZPSpFVfozl3m
V25njS/sl5fzQHqVc4wH5N7TtW4onmqjBDzea75FANprMpZFYSxB21Szv4YDsD1y
Ohl6fnd9jxxCsO/t+AqWuJueos4ImqgKPIr1K4g2bZe54e+uB/LxincXzxRPmA1r
oZFRFkkwAu309ryUpzAdpDq6qZgqFxcC6j5Fh2BiCXZ57yVR8/xuouVYsBnwjmFO
0BvImVbhYawzp3/yZcyFsQ3Q3JyClQMPDC+W9Ro88MiJ3HTg7yzgHdXQ4OQAzW3g
ylWDP/yzvhVC2WbxHvV5MYUwrNn9bCgwrDLTZTd352WHqy/08VR98Z99uM5vcz5e
6U6KXobMZzalOgvEpYOOSS1731INdsUaZOOkPBa39C8PuWCBJOpGKryhro3752E6
DScPKy4p85TUWxazRMNrWwEUHBtj97J4sCxkQSl4Uw1JlW4HTvXMaAZ+KmXgGjf2
FrFW/OrjqHjv+WvfyZxz+ZkVcGMuY2xR/UCUC16l9cHlIF3Qz2LIne3rhNFhb0Aj
xDGij8abW14fpk4TGLiWX1sKLmgFTCxdKkeM1vUFUpNIk930UIQILRSoqaeUv1SE
/vbrr0BEM1ypIUiIN21lQZ12akKlfFoDEtdiiEYlgvfu5urblD0/HZGDfhHU5LIQ
NoX7cV6oHPOpNyhxhI9GgUD/8PvCZszy5SdtwDH3lQJ+pNUUc/XfZ0SpEswthjfB
AAh8nwbKigDCaYFPx012TNkn++h2UOGhwtJZuKRKDCDazuoanwIQU/7OIo3hkSaR
t0THYCrLDM+NuhImEQxro6A0prdx1kCoNZGDKNXPz3zPXnICamMwofiYqPGItNfS
4MEEvLH9Q9NA9Ss5xA7OhqJPGl/m9gfMOTGMuKMNqkCH3uU5Yl887xgMgfE5ZHXu
BAswzl4y1Itodvdz8HtGpWrmTiALi9hA3kAo5Fwys49U9/tc78wq+KH5oXNZmX8I
4pp7u6S9KGDTLITzhP+54TCF0mXGSb/VHyn0hLjOKzv2Tkf+5GFPyf3lftCwNDWa
FWF9F8eG52oN9fwi8NSfraYc0cnz3Z0/bwB8iONvtdFjyPaA6LD3keRq+UATfiRn
OmZdWr39rY4qSFKHIdm5dUB9anxurhl1tbQZ+nQrVNlXDyBMsmqIwp5KhIMxl2MD
DInAmNo8zBLmVozmtKhMNNRizl/5HNQGcvcmOokVIGecxqzs+rBbyPurDADSVNn8
433YMpsuDNE9hDYM9UfrHACnthuR9Rk4PqYYKYz9zEb/ivaeOftbvZGUlUgZCo8N
JowW/DF53RK6VCWG2bYslRyG6VUEozL7tYJlzDVpMsd9DNU2oU43/oT4pIdhCS5e
rWO0oVE4q/I6dU6nKcnONDx3oUPabzMsVa2dfjGg8pr7zuzgzpX9NdguRYXpHMuN
+VnJhnOlmFG5e5UkX3Lj4AywT6AuvryI4JXK710Xd8YSrPxTH0RmTr8b04ofJS25
DZggU8ZNgbXkF+f0EGh+sgDBGoVVWZ9dRmJT2GvZIPDRIUA5DPIiX8/5/0/wNhOc
8ZsQGfvcxmjmHdfrIfl1We7j/pn6Onzg0QyrxOAe1IWum7pFjO+qM3Sd2e74FLIC
sfLwbkgNkfkCfHNkDL1SdmaImEO9QwV/PM9ZrmJwtPJ9aCHXLBM2GtQG4fH1xDQ7
ShYgGuvM5i0HmfUIZsE9tQy4nfpQJOYaNXdHbdbq5ExKnLByZrDOYdVtyZRQSngn
GpctYQgedlYwrzS028mFAqk8Ql9Yg6YJnkCZoTP21N8Yzm6e/WYt3uEypOhIv07X
Rw3yKfNMgPL9F93eai7FiYHY/9uO4IoMNsTf4/QntXpCI+dfrFfJWwgFaq2oAFQE
qqvVRzpzziR4S1Jcv0S/9YNgJuGBSafyshG9sD4uN2gol95iWjHcXE95U3B1GVQM
hYoK0I8kBHhsOpzK7lG31JowNxDbmnsYv9xRzHCgFewlgJ/O3AnHl0TmXqGhwv4X
0ROR+giZ3Hm7+AErDFUe3A8c+xaMZfLDEcYVvUmo4cNZpSiqIyHC754c3rFfOYca
nJnhP5O/Lf+bFpB8NjYa7Wh0N3ak8/B+E8vuTKRyn1HGz9IFxSsATjswCQvciSjh
nKdlV6BlX+hBP9pGUIA2F+HMP+Du5uuP52mPF8m9TkjBWFe4SmzVlNPYIdnc+Q9+
evLBGKArSKZVcboEDmwQgFmICDcwP4X0TekgXviLdgJO4zmfi6d5j6vuSu9jyQz/
HoeSkRJXAym+mSrvwmEpElx/ehE2fRblQmcZZE18DY9ZNlD27x67ayBHg24cnfka
qTXxaVR/33bda9wPbv8Vt7mryP/9/nsZfWoMInOOJX9bQn8D1hTsY+vPfFFgX4H+
E9ARGtbTjyWm9VkmZ2F892B5g7FR2aMZPXm8riwy+6eYHPhnu8wBd316KpHvaPbM
fnzeJvIsjqVy6pCo9jHvJ7TOdMPQpmSHUJ7FzG316SGEzRtXvwsUheZm2J9LrakJ
wHR6LL6TQ+OSbwNmhLv9QI66pBmfBQ4N2COH47Dbdnh4NvEPJtZ26UL8oKJvUduo
0Ox9s979U1YP0dkV10x7If8x3PGaYFhyM914r81oKmhnqbf4u8PaRf8zcTkkFFn3
RQjlPNAaedjCLAQVoDTA55Yq59K8MZC2pRNOALGnFVzfnAqeGwyO3AsN20ZNf686
VjyPDNdk8SamFQyKXMby96RFOn7nFrPKaVOP+YflVAHFLVFdx2UdW9cllWiukvbB
tHdwKy6JAz7YNnFCbpLvIL1AZGnX4N30N2OUpyLI15l1c41QNSOOREtTC3LYRSQW
j4DoYZFio/yLMWxldhhPwmQL7AhhT4t4XjmY1FFUe6jdTjeGZhXq/wF3+/+ThJop
ENViMOPJ1XKNh0B9Fx/vR/sLwlQv+oxO6MEnYmQt7G2gC3gwBflLYrH9K+npkzvG
kR7pch91A6mMHotW1i77BwKrKfcfpmmA4oMQwOw5jE5xZf705gT/x9SBgkJ0HSgf
0rHQszrpNld+DPqCS1MplQTAFIDku4U7su1Kncq0yIzSw8E8oKUa/e3/tneTYt/u
Fe6Xyw8292CgO6HM2hdNRkscaSC3Am/9/cE11DZJZK40lG+MjqoQOTcA2p/ZHa6O
YcVLoXJ5Rb76nLDPaN1ZydRVyXVQrphLWju+S7qsQJVwLa5O/yrWrzjTPniXSaKT
PWskVA5VHvpcOIuF0n6c/8sR8ZiumX9Bt+ePkApJ/xYxCQCEw5BDnKU7IrMgyBjW
NKtg/IOYsCE85k9cdSPkXR5BiL+JQkpJdTWRyMpf9xmMhacEP69W2NWaRM/EKRFJ
7whQu0rvBBAfgPFnxIXJrYajN4Mo2ap/vWIj2lsIOly5HFp82102+PEougA+0xPt
8aNbrKP1oi7F5/+iXkGwO7CYgRlcO7Bsjp6KImYLqjPxWWRBDign9YWFPXqYX+bW
OxncawhsDt/B1ev4i/KvdAkq8mFg6P+AIvMup15MXh0MtIB0KoT1+DyIqaHuo1an
MYBZl5ukpy89Tp4JcDkZzhw2g/hEhZWBHdQuqwBWG/OyyqhZxfML/SgoW2N+jM2F
JSJa2pFrv++2yNz1ZzJRQD7L4hK85GU2+VGxkPQLF5DAoNMhDoP6H9k9RLW0JCtL
0w6MmPCL4qUbby1FkuEbys12URhAnqIagbG5sedhpKrwnFXq9cvregH2jgvnjVLY
pxV6qdzgswsqOItXgOYAAY+gZZmhDsH5vA/p+BcO3SzPETatVdyceuB9XiuX9nxq
57xAWtUfhGs/uykzXD2c/jqELqIgGStyHYkEYDJ82jtbQAZdHEPx6bFbTTG1hfpY
1e9D6AJHPsMVXtlKmcQyvgzbNfi1nXLwgceSjJZ/Y+wE1QWuOGns8/nLdQnvqyRr
KLLrSkhYj7yBhnaGub+S0i+JjXGUynO+b7zNYdjn8Z/78van/koLdbWdCf903Rvk
b7ZfBC+o/AryZs/vOJbQk6NCxCiya5tNybi0KIlP65lL7MD3/4pxaB5ZXpVMpLxo
y+jqApsSaSVgJpEj6jzFwNTthVIzRagG077xkYdd5cdej3bWlOob8Bj8f1DDOKmm
JBmoongJ0sAdbO9luxLgYZovM1NgNY8NDBxd+3AWflZlASgNIwEt8pve3E/FZquB
cSGstJWSrY+5MBHbknwZLHZm01uJi7rj7j7I1aCy8vBJAhfWs5z5g7SztBV5Jznz
xAcmNg6UkpDDF9HhtPBlXMpMCUSIgzqOmPpqxBsEMsen5d0BGXSIwjiNoTzzvYv5
DPAJL5iH0LuJwgCnMvbqBCYTQzlvdogbQyRVm5LntAC9xU3lrqrTStKcPP+fSc/m
Q8y3WXzwMJcOLGoEl0OpmJvy2Z1yGfouGmEXF4Be9JfxV3ZqT7tq+arxFyRBwZ1X
1mf/PprwAGKm/Ehotj2hJRF1MyIbhRWPH9B3jcZ+M5pWqbCHL95wj6sffO8KJ4CE
MLgfcLLvWY3c++fL1TZeT3GXNfrC/7puxUHJStfXefW2FPwKs3h6LMUaTREaRoN0
wpanlX+5sziHwYN/xhmW75F3mmKKIQ51YnIHa9RyIXwtd7J/fduQrfmj3SJXLqz1
zOi7eo17BQHx+dDvYCfuI3OKxgOjr104a0XZpBjb9fUhGXq7JwNF3Aqnfj4RZhuk
gzxlOVviTsgCmk6jGPD3oczYmIs7eN8SszsVtp/k0mxuw7eLjONmOJhdbyGtexLu
8vCLE+MntE+mb3pWs/tXnNBe/ctDvIHCJnR4xWlRSACbxNL2ofCJxduwpoBT5nxO
mGCgiVToziFi55cGHx9Kc0QzaG6IXOMN5ATTjBBmbXr24K77wLOaT3Ydc+CLZFQg
1dYtIryY6G+K7PH6frQyc64/tnhPv0266VSPPzry/SiC5g6guy8dhOiLhecyU194
EgI4uuVXjB4PZ6IYdR7zY5jBr0VE9kWZg4XAv2l/YMyb3WidMxnRu1J5ls6WNhdL
iNN2c6M9A9LyapmK7JI/qVb1iNoa2JpvlB/570PfMoa6O77ntuYN5jLWJLAlnD3w
Qh7uAMq2LuBBxzbx5OHtP41alZplkB1Ql2e+GdBiqEGBQyVsaE7BKEvoSr7/hcaK
NC5pPyjBTYKrDjzfiVagWiOaXNwU97T8ZfI5tS4AcqNQmFUzRUrKy6r5t1Fe72Vh
eFrg4lQngIHNvHkrQvT1jLUFFZrChluVPQUIzkYl5j5mp9p6SVoYPYoSh8Jsy4Em
duiZWB9WPvYHeSjKaveRd5zyQlSBlRH3ZIPlbr4GYlN/KrnhHSQ1kYRg+2H9zRrm
HgUBCx+5c9cseTms0gQZNEZRFsLBTBeJKzIMFSa7PEkTu4L3q3Vcm2hpwVcwGiGd
v2cY+n+73rFKAE9hTbbzciSlLCtLyZ/XeL+pgR6vWNAdetZxHjTE0PF6KYzB7srn
/1/JsckMtx1Hq7SzmYN5yH4Hrpg4h9vjctd27LpMWv0VCAZu7eJNFCtZSfNq4rwc
uYNlPu1xf1XqfnWbBvfmpVmk20ffQOgrZCVwlFhH+KxRpTWKgjcKApCHN/0cAlqX
2ggTK3C82CkibCoOqAJ5zUUCF+QfPqMZFVROzP0vMeLGM+ENEKP1KfSUUJVrMLe4
I1FxYyG5BhAZfggKpzgzww2W941j0FNrwggBNyBaMnK/GvGB2kqVkWEGJR6tneQJ
NCx+ILBFa+R/wcXhMGmNt6W30o64qcFdx+t2M8ILVHAFG+mbj+5D/MCqMjEDlfy0
JVwYB+UQoszxTCzOte8VwSu5Jz8O416WodN8h9QefZmlkvReolp5zYizjXlMilPw
zWUXUt2P4Hb1hGnGUbMbXjjAViQfswhWHLlBuSL6MuyS6eh1UAHUxMhxT1wtemcI
fPxUofIkgXmAdFMj4WsBrYgk34hCB4+zhUYAkcJbht4TnS7jmNr7FPlFlVEtL8hA
Km+OYBNj9/Fw/eEPsxB1I8/4AavD5Mn1xuRQdsOXY0VihILfs5GtbgOxH6H3c3Us
erAlh/Hhpc+u+xfqc2NiKf313kmQo1Z7o0WGhuO+eJ8ZvOx2CvnDrzE6JDNAAouy
qH3X1JrIaAfr8GKkj8Q7aaHuVFx5BYwxrHfZ9Yo3qilzQEeXe2cLx0HtoULWBOC5
nkx3D/161A9m1+JmdFpyrqUh/UtY0Boga9WhW+zEYVUK8PKN83tddUsAJNQ8XICZ
KbpVOh6tN/zV6SgRk9CNNLgJeluvBSLm4r8tILd+pSJGf17B8YgOLWqVS/R0oYxt
MybcVs3/zh4wj1ixJVHRLC6caHxFsm+01uMkArJsA1Ed2MT2ZkgYOOZKyFk+80ER
f2VdjZ/p53MDPiDrqVCyO2yQPAspe3csZvZpWk3RFnPvM43HM6O2QkiFpMyyDaZN
k2rVZdcOGQ2yjT150luM96zZxhKGPI+IFiRWX+tfO/A1nDnyBwtwncxb7P7y3JAC
bRKIsQTi06WKvxHwAgN3z898TVDJC2tjYCHAxZwpuKnSnJluBqR1n8V13TVqBsKU
izhYYBGscg536giTW1Ba8HdR7+g68TcoUaBhNyBQmfccN2RMMUYKQ5cB+bZySPIQ
+kNbW0LVZXjwJRmA8BDQi5owr4tAKpSix28n2KAYjsSuFyerCBwF96T9qKMcGmuH
Z8h1IRWiKQE7C7Aw2xbz/in9K55kcjAWV8rxoIAkxcdruJOdQU5Fu3hCMyX0bn18
SUIZsAvq7dc4v6yj4j5g1JAiYFaDEiNcqsacE8HKXYZD/r8y/qn2nq9WgPL6/3LV
sn9ISrFsoM0LnOJ3ofh4ndCyPXdcwtjJnLVATIFlsiYEciJjxRvTAUn70we9ug6x
HC9XLBNBWeQRoiro+fYdPSqRwjzxzVxOs/x6VkExJ3MB/ONR5lIGrmH3jrPPgVyQ
agKO3MGnsyMLJ4vSethwn1gRbDJwMCzG9PMYGfWcSTH7dw8dK4m//ZY7Rasykond
m6IIO27RG477LBa6naFPMtTb26vTDjuOTby6FkbJXtzZxY30JD/rh19URocJndUk
6sIL9HjH7zy7/Xhkmcw6w89hLZ1yBcSgeCQJ1YHeCBQ92Qz906U/rUeos9xto+Ab
6ujYw6iP5sspeNhz61Yx0fRo/AX995zfFPNYy7qFnR+mpTa/4tyTwc6UAn+MxJtj
LlgT7hI1BUPWMyIU3Bm6h4L3m94A9OUs4H9YLljUMHU/W8J9z2RV7XWgwqIfw+H7
duDV/iGVmv/qp7Vwn4mrknd1u0+sFV3wcu7KFzKNrI2YkGl1VMCQJIX7DayYTht0
gCRfoN6UgAbtRUvwGZ6s+BeBrLx58LsA4howtwIJmPcGSYeB29jM2h0IDa/CiX+0
vty2V4ZvZvh0oMMIYiKYhS2xHi4uUjdBRcRqEqBBfnR3lUP4WHWhFPmMF/x08XFb
Ts8OqBAt2BUDHQxRErrHB2lI3WY2/bKIW/6gRdDpvTQKtyVTUi2QXrAuteQVvEId
2ryq3X3yWc4KYvLLyPKmBkHjmCQaSwrWTTs/2ydZXbNxjVcDgvrTR01nu327chO4
SAK1nhVuA4AxDmBkSeVPNicZGzHSk3XfvJH/0PAAKz0A2B3QXdav718+IbyLqiEc
VUlaiA72ptHFvgp50BLlgN8u0JL9tO904yN6u3P+oADhh8E0EwL6rMHargoH4FYK
DfcPEtJiqfZvuMSWP97VnZChDOd69oHy2GGNG0gTdCxAWLhUta+HD63YSeLtlmlT
ozXct2cQKzWXjmPQGAaB2d8125i8Rj9/x8FwXFZX8V3pXkkdRHSTBpqNjQTdtfgQ
PM4u4KX293aOPSmnlGUz670IFQa+iZT8RELua0SL9qo5yuHlGjK1L7I0ih8rP28A
MIaLgOe08IABfzVf6XqyTIpJtzxix8y4LUdDTa0G2ZTIy4NIRCCD2mh5LGaCR7kX
aGOxdpuR449xW8Do5EsOuPS43nqKe8ltCZcAUHuArH7bedYyjDkdDSWX/Dmq/nKG
vxImIGx52tPp+HI+Azau8lYNAkXbjItygXJ5Mlusr71OOqx29U5duSR3ixkJZ6Rc
YaI2nv+8E1dQXNZ9auWK8V+D9JiGdGiLbEnHKDU00wU/2Cu1dBsGMpKWRLxITaiB
xIykEIGAVA8apdzs9YwQIEqJtFnvtD5X7w6AxjJ960LEbJu0Ds8XGfU6UFVbhoCZ
JceQhMUNuzLaMNW69bKu8ixZjuJoEJF6iLwgRKrj6Id2mjEDV0NtSqha8Bo50/md
IfaaP+CeRmdqZzgk3HVjSfeVklWfDwuPAjJqOCcAHkJQdjoPlW0R6YjQXWL+9pGD
xXt4y1CjGMFNMr6USReMNzUp5u2+aChBeLQygucXW+RpT/+5TyQPO6WyF6T6ph7a
CvgAKkzzs22KBWeweu86uS6WNKfJAxKQcAcfyiQvAjnCbLpauwPnDwYAyhOQviw1
KB+Wbflp5v7gtWx3lWrhCkoS+iU4ODxeBzeouv5ST5zox8g5MDzE8YXkYPadk3B1
D6QtpXDxSH6WMfMikVxH/GsGCIk4k8sL4lgq7kMt3oJblGU7qYnWxNcXBZBVT87s
aUbcBfRh7gqPjBeBKlBif7vkmsyN8e7OFO9u9pyrv36b8zZuNwAYUjQ5OZ3Ic3Fj
hORSUUVgvX6mwaHcwhwBbfNiez6nUPdeZQG/PWoXj5e/vqF6tZ2VA6Fec7uMEKpj
T65cqV5Iqin5dZSFyJpAdjEizhe7D5LzKNd0B1vHXWOLUdXns1G6L+i+9a79s9lO
PFNrAnWIli/L9eklyfhfp4OIPVKvFqeVg/kHaJac9/esXrnThwRaZaoZoY3bQiZh
h3Q4Lq311b+NTKKELSktT5VuYP56PqWXISEETg4CaKYe5Q7VXUAcSRbCLGpWvTa0
10c/X4UoJ0/PuLJnYy8hqVXzkBKPBvTnho94JPvRWWMcKAFc5BkWKYCSLElxbgmv
E2SOu26GuOaV1YMvcTn657J5b+HQKG3/mkmcy9pMUDqhjtPQlS+fzk7LgcqPKOMj
6x441ZvmNvFPdDgl6NSJ4DYkxG3gCuHIE0vMf5GjRW4s50bAayOY8eVpsjUIp/tq
Fpl8CAx/2H9QuZIznqyafQ2WZNZFuFaTCow2iIe5qQ3r34v3IvrJ9D1ainTw1A5S
wTEijQQfh/VQlOgaIZEWyFQyzs6oNQEQaxnzpnBx9wMzjdoGPNI6XYyoeQ4gwO08
JrIq83n1ePnyOcKcAAjYBlVXAdnXTxFTj4BwjlNYSo5sVYyfavhOZj6yzg4eDAHr
vMouC5HZtLL11Fc9mIMaZXKLSWVb5lpw9e3FDeYVJYI6Ubhnjgr/GC+Lreg27/+3
Nm79U/des9AzzXpzU14zxfR2GHvPfbVxQQYhi4no5ui12K2k+tiJ7f6U6FGZ54If
qVJBaIsQm/sJHw1qLqbiIia4am0uz7HJ6xywZEek7W6vgOZxdnae2CYapZJS7P84
+PcUB4Er+mwtPdvTCg9aeJGBLuUJKw7dieRmSbW3b/e5MOpN7TxCjJXCwPeZ19UL
DzlyU4MMaJJLwXX5/w61+qDNancXmaG9+v4eUseGaK9RZm/kwhP0fIrMLJ/Rpp4P
BtzuligY3TI+Rp/r4DAw+cGDxmXD3JsQQwb0JNnxXVeLWl38uPmuvuf3q3N2fnY7
b9fX4lhjsxabeXds0ChFx5mhC93OKLbsmSxeZhcpsi//Kvgb1VwjD00x4zkzJOOf
lBORkmrGNVLgEUqLERggHx5uugHhCvryxTOkwvPXrWtlLG3QkQhhHGL6eRriPXqy
YfPAegW8JcBtLN76HppTqL5cXcLay5+wIT8NIzVmKeWMI9/BTybJUWYoNkM2g/2p
yA52JX7F75kchsE10KCDZsokbkjdDzRjNDMzEKymFPp9ZtrBJkmaNm8FVZOicMRa
MFxZkJE5boeofV/V0nnqEMxQhJ2MLHISsazxZ7+BPEvxOORBJB4U1J2vRQxmz4mD
b9zrFfTF4S61jQPwhv0rvIMvocf+dbC1IJBWW2yF4E8FBTrSzE8JvPxEJdzFb77Y
y/bi0tlB+4PmnptbibsZgn5tu86dLA/lSSN/fao/L6xhR8dzYkbWIRJXYx7KXg+h
9C+MNuucgt5Iaypzg7hleqjOn2wM1wkR4gwEs45iy8QNDuhcnRW/8NNjIAcbG1jx
1Hnqt71xhMcuiEinTjzYmP2ZQnTPlduR3Qb915hfJtIoSwS4OWtMjHGYTMnENnqR
lSTVihxDdUMggUCS+ACP56cbNiC+3lgw5ohoXyWy5JBGKtcy/9q+Mmh6P75/nlzO
lYxrBmA1v81yOshlUOhX3F9eyth4eoNWPZY+BevztQNoI1fLIbrgti4ONW6M/o4d
2gOdN92Qdf9sA75upM1HOZhxu0c3QD6N+Gvgy+24zx//yJ/jizPDYlff+jaW8l6N
qABPyaEUrvLFgD+ccn+cv5RbVeAFkDYEd2s6rUL/+aeQeA5gCrKHmX2mw01v+g6B
zuC89JtGhIK5QGW6RQAlldz+gPCUUUN4YzSPe3jXR/g50ooEMzSJ3nwDq/+rHu+j
kLiGkbrLq3uGJO0BXYvZ/v5JFTKOdF3rKIN8HPqWGNDZXN9fIE2PVrrRn7BxUE5u
QwT+itzv3kSTyLQlDWa+Onwh+I4k2i2ivAim8LrOrbaUQ1kE+Hr6wFV1xB8SOvfI
/FZF9pxlrP7BmakJvU5yYdnMb9Ux/utw1QviSvYpqc2CRGt/y2Nd4bfM1lXPvLv3
EcHDw8e8yv+vQFRzLxVAc86oKabtjjc+EcxeiOvYy+UZNVbDlkXE7iZxba/Xsj0I
ZQzxh4otIAuKJTGoGA6q06w5lMf5iUmTVA4SZFkLG9ilprp0WIbjPTHGAb6K0K8d
9t4FWrUqwvhyfzqVSZcfygEnc96nkJVW93JXbmLJMkvikWUlnGiZzSshCC4V0Dqy
TFg10uMcT7Xgnhy55fqsfAhhufy9eY5p0idcidXlptF9Ql1EKFRnmqU0e0aZhS1y
YZvr5LDQydzQ3DzA/3Gs4yvKwStSfiTxFdNqyk3Q7ymjo9U1uC11FnwgZa2BjbVT
jmvkmMFo3oBHSpImZcHb2bYB8o90Cr23rlGQQvLdBhM8W9pQtv0c7Xd0L+C5NQ/z
QVJR0qCsaBPWySbxdbkNwXErl3h4BmC1jJRZdPmfO+oo1RPU6QEFb5NWle2tAGk9
D7Mjl8i/ACBVv0NC3gHecZS2wudvs8kz65mzVJDWtnFWFmJV1JjNWGmdrtKmsqnT
i/qxYhNzXjiWA4hrJAEmvqK5pUd2k7472s41fIP1HC9nsTgPHTCxOueKrQLkMT0u
Y7XUHg46vUopYT4FUOd6d2Nz6RJk+qUiswozaBasKdyD9W6wQUfFFFDJk+7LNfrj
9s+SUwH3OpfLtT6zP4n+syj5uisDAIH8zQIII7UR+qir/s8+rgkzRl8z90Ep+y7e
6TqlfMXQUy/PO4oc4PBTEhsVU+oZIJ0zVFUA0kVRxpcppxfKZj3Q4gFKZwEf2huL
SrRdMvgX0SO7scHBwje3GPGACKXW51+im0wgP3iEYJb/9pBjCCrpvYjq7c+hXhpb
tRuNpGgRnemKtnzp4ljIeALxXwI2BUgJ6ZDd5/dLvykHiaeKtRr3g3HJO5HeLYbj
2TOEyUBBn7XV0bb7ohLPmDjd54Oer/LTisaH4MbX1PsLGZM2JD202gEay8OlpmcP
vRWKIqgnMq1jCZaOsNA18ftLV3NIJh2b2H+7pFKyxnxpQVKqJmg3GWmqWdSO4mUE
LBQeiy2Al7cWRi33CF7e8p3qlf7rGfz3QJAwlb0IOdmRz6VzlEKzgf9g92YvrUZV
RU3tznoHcwP2kmKDTQfuEMoy/qOxhQG1oUBiEJXVfa/H0lIXASy7//Btt91a/fob
HWsd7t6PwEdLC8ZOvSecDfvbryB89eQmul9Wh6BOcgPZhDOq6qdHRO9tfGoycFKE
GiIHDsENquk2VejCT/iDTFvYGcwArGQPCooqasnsRHdr+Y1itki9Y33rtvTnEtZp
YV+9Ep5oqCjNm4AftT9cG6NOqz+CC5WyqzPg+fQmYcTrilNWxB1AT1VppELYeque
DanH3EUpqOdii/3ldzavczONyfXQZksy+l5/7Em63DjeupYjQeLlaz8ffZ67H4vY
h1ApKFFuNIy3DAU3WExvTl7gl67umU0mCF+TElwp/hBv0Sw5OOEACoKjjOe6w16I
JENEm/ktzlVRA1vbp2jQfZf15nUJ3ILauxykm+YCpX11kAKrsj95R5bybEKm1sCU
ORVk+RJZYxak+1IKVIZN00G7w+WRxASQeN7QpJsWQitItS/x6AybD8bWRBpJjevr
rSeFZUdKirIAy5D/+PS5T3ObNy6BSQDtjMsCDBuQ69YfHa0RelHIKdYzw+BcARqa
kWrxav9AKeAQqzFBUIrTcKVMAXo+z6ZQiQ/Js7l1WHF2jbuS298f4satFxlmqaz3
6uKv9HUKTuuOjCfgGid2f521SF2ef3qxk5YYIcfot5mOlLusk1FkOnANRle6/ZYy
xOas290d5p7haMNBI+yRNtC1zz8CRhz7xXhOleXv97Wa+F+kclPcxqbBizD8YOes
9DBgwRh4VddZq2oA4y4ec8hevT4T4t3BUgFRByjhaHo8g3564oWvSJmUKwyQ1Yim
fVmQVJxoeXdSFPwr9lXlGPRkB85CcedKGU0/dcYZ290ZvL9YwOkeBFy9EotWU7R7
dENv6fxarObvGgKpRilBmaoLxq1VXSmLa8R9oRSoyYOPTdTPVYaLgwuN4TlSh67J
f5g9Un6bA2e5O3icW3OSxM/9gCXxcpeCZI0MoxohBa/1m/t+2vx5vL7Z5/HqO6iD
jkD3aTtePa79zAZDUaPSDWDzHk5Q8D5YAaBO1T3IjlBMEeB6RNlGTKnYARSbAsvy
CWp7034+gRcogBjie/Nu98GMJ9lUFprDxnI4kC5sauCd+ugUHcsk2DVlIsqnZCuV
JBBZonj+A9Lj+gIRp0sS9heTjPDUWYIW8pXcuswMcy0XdYI1BGnnbbKa+SBukwkR
NSX0nz3Jc2DH6YI77is3dn6pWmLNOk3WlHbEqECNtkmCzqdH+5RH6Xi90/TB0vnb
dbIn97C78WCKStJJnmGM66WEMrFDOVkQSdjgIhxCw1WUCWJReDr8X/4CCpF7gslX
P/LsqJTMuWVfKP2hdR/aq9jST2BHj+z3LnPviIF5bPVAVhVAEKdvVi3RHyNZQwkh
oemNe/C9KRtvXsdG937j6URcN2+fEuzC0Z9eFO8nheDuEdtR4+ft7WpSQ9HbzyRt
jI7M3oFScuaHSD39SuQfnp8xLmddN5iuxXOZubqZHAkGzdSm47iG5JXSWdPcd66V
s8HI5lnN46f2O4WZMDoQxS+4LpcOGRMnU06znlH39EcEhTuCnXUtggkGpDbRhD2i
/X7ooypgEppgxQ08juw9Ep+6xyFU3DJgvxEXpiLblycAlae615TsdJKXAXRFb9lY
FRgYd8rcPSWaM7QyaKVydQDNIVGcL/jdspS9DSul10MZC1Ip9nwMeJ0PX/YJZqZF
8tOIwwMLDgSII+oSUATqbWmsliqCyDYy61oT68tRMTLbsdT53cjVbJzzo7Qqwp45
81XBfgp1/++uaH9ngY7eYC/WstFaOWvhcV2/7kJg4j8EYxWJGCME92HSKLY0nDab
U4mJIw3c0wFuMbHG10i9YzeYnDgrEb/xf1yRXxBZXtzE9Dv1+18BY2hLqWVTcp9F
G/F40d88bUlXlmHPU1TV+FpryFSts3lgH18aTQ0+iCMf8oa/Se1IZrOdP5r/dJOI
6rsBOl16B2NGOGGhdJPBsW6CsFIOa14bg6r1F1SjAYheMMRLein0V6yzioRg/H4I
uXHqVpLOdqVKD4zQGOONVRAi8AbHcnbnDUeIBsZHVrnPdVCNF73h/CDyp070N5Ln
oL7+taLg40c1oSHuDHC1M/NzJwhgNtugsp2AmACmgvOnSyAEfvYpOviXrAodeVXs
jBYbTBicE8Y9lu4U+yAgHSUHcGUKvfRws/kwbl1vKGEV5shy2oAH+1T7oaQR6spC
k0duVpjnG3K6J1Ym6NCtEcHW2kB0U3yweYaW5bxt8VMMF01UQqaEk3tDKPpJMYx4
Fb7PAjeRuxg76xtpSxreE3pEjgvYNE7hXskdVHmKijWFzB0DZqLvXI8uGy6Nab28
qIuUKshV7oZhJ0hRwIp9LYzQOIkNZSDt+egPaX+/SC77964+TbKL6+tRgLv6/kgu
/PMna/EEFUfJKolx5/vOI9OeN9C7R1mNmDJAe5J8YF8oxiY7gy/N2iK5CY45kmSC
Ffd6g7K1FAka58XoFhGYBNOq8bnIUWpIN3YMbNaVn+fhipv9Q4VS5OA5ALCmBmwE
rPIEMYB00J4kKvGutGel8KZGD7adrwYE04bIsA9wU3yZaUwXzrPAC7VoXu2UbfTQ
uNgF0CiMh7/oJEUhGvS33kltG5znQ5cgu124E6G6Zc4MlbxhE6MgawFhCmwYfKMP
U7pJ3Eq0XawWUGnt8UhXQnN6Ebj1yJauImpdmjJwA+DQ6aXAEHzHv3lefDcb/aeW
phRyKsqLoGYgxA75FDYea2TevfCbEKBUJsUCWV7keVh4focyHxG3anK/ueg0BS7G
zH4rsEqFIZFsHINnjs+2SV/vTRgXLMJpXC6gJO+c+4Ghz/hd1NfBlOCIBPtx2x1Z
G3mHZASoRv0hrhNSvMj6kZ7+6yx85BEcrSgOosL/1fZHX9m5b0w+yMRvocSSgDoA
fvN1Ts+2fuGQ7+XCMwqG1jIOsqP57lMyxREPWjAo3hXJqb/xUuC0DI+3dhDDUg6J
wpsRuK91rxPl+gUdBn0N0+2BdBfeP5y8aTZqcOV7GgviZmVz0uVx3MRNlJRpTNeh
EKuQKncESZ+vO/fW1be4C4CkXljX/T9niBzfHZ5zUsn2Lp40jAZvnsW9J9VFtaPn
wITmvTsC254XK4OcZx553kaqLpV+dP5LPe/15oif++UOOw3oVL1aKZJmTPrFy5dx
DsM+/IQSVzhEzXld/2fFiWTwBuCmbp2LhdTLAYaFdDPhBFjtFzzIqsL412D4R+yg
9cfoPGpKzEVz5yZWQLnzy1eNKOMyPJSBZVv3X+SMHDRIBSTuWME3ll99ZqlDgjAd
Td+HgKkH2O95SVaOVkxzP/SiZGSMPixqbOE2AcpOy2UTzDicpXqOuts/flJzzxiC
LBuN//RujnkvKxOqgHZXk+PvxQ7JQ1g3Ki288pl5Mc8nxjYbzVjr7Q28ksi3OVL1
wH9LOLicet8x3Rlr4oxSbGSf7swGKPEN8vuZysYegF/i3EZETOTJp1OU3vq5RdJm
DNG+J9xZTXYVxO6zTN8iY5kwbDRuzygRd5n598FpWkHQLZGX1pklKozRkPPT5qri
+yrA5NYA5/aQT7wjR3Mu3sFPHfBogRNF/RVKbb6wTLGsfy/MXzyuUkBR5f12eQBq
m5bh39QBw1IV4YJQgOo5GnOflncXq+NhzxkCcdo7BF6SNb8F6BCZ+Tw78H5NRCFr
Nd0+OieBHRDSUHjxyKEMjziJ5WqU33yuRJE1ccTNlVK1Ii7/0biEV+ZBDJhDZoru
uRUiLDY8VOyQdHXwCk/TJJ+sr3bIqW7ctOtNcovAvQOyju6QdsyU4+aWz0e58llC
L04J/TgjAuZ78imTieUCTfMWTtX0jiFtkevfEaF8c5gcG9KtQJZcdR52KZFq6r51
hoI3kNw+1rqYhsAvP/VJF+pSFpjlMj+Uw9rvC2HCdam7JFiOhy71VEq7JLTAedK/
G3vhh9Bg5mf/Bn35jceHx8qD9p4tlUNTAHMKOqh/249DUjRdecjaOvMBs0HFcRbk
ktQUUZGAWL5R+I7s18blMfTrk9jmPtmYK448fHrJopQITuMtT/JGYD4gorVKP/RX
T87RrTJEIBlKopGEzXkYtUgBS9FKrOoznJOk8Kx80Zc/qnib9J8Rm2LAF2zc+Cvx
ImgSjoYUuHmVeLteTPUVA1gMRJratVr7EZANuOSPZP+XKHGmzcm3RuB2/AAcnU/q
XMYbP7PqxmSg/zkBZiR5nXGyNfqbuks/TyP4hJpfGEkM5+rvyalCJ8n8trmnROi9
ox4dO0Nj0GucK0zgGQwf8+I4wQNNdOYMLgRGZxyUeQIpA8ZAgyumgAPwIlW/a6Vm
mncpCJ+wHZID0g79VDy12jC88s5D5m7MUpcz/dnXlWefE+lzvnG2old6N2U8SCid
uN3JWwd+iQWGKF1tMGNtEl/22U3CuVeLqE2wRMbbVEAl0go3VIlnwoUA/SgxQHI9
xvb15Ngf0Uqe7DC/EZpBYGmDDgItGcLeiLn8paCccucUJaBN2zu8BE6wDENP1JxP
IQrEMPRljQkyaxL/wPw85XEDYlXUPKt01Kb3g+y2gUtqL53KnkZaaUJGt7ksPmC6
cO2NFmLlQhNWD+uOXY45+9DrF42L1t5GeAV5x623WpkHRWeNVnROrlzkAIfYxSgh
LrIiq7Ch2mKKIJXPVRLxmAKMnDMt78uuKBBF/JWsy1BybUlRMOiEJ43YIE6aZOIK
ucZ0kelPK9sDMrLnPhkK7NMnmtgT/xgofzv/PVFifsRx28Zy3bVbZdUIOiN45Vxo
lOfNtpIYXP0b5b/xGxec3cjeQlDl4Y6+o7JPk+d2Sfwtnk6xm6zlwwlV74rHPDQZ
t4j2bMJ3r74JM5rvDCX8ufLjNrfg5nuw3VMdcYUulmt1Z6jAHYiVwJOUA8P4/LQj
KQ1uk1TER2/oC4dTTc5RTknzhkRLUud0LC9ghp42Jjg9XQCm04i2POjKuvKczsQ8
KRPHAwi1JrlECYZtDCO0G77o/Z83j6zZl75s0ddlcGFGci9E1camCiUieU2mXhDu
Xe91VOPh08cmLTiIUCfVU5ZR610r7NS8kE8lb5GP2xRWUVgQiGUvodeErrB+XImH
CRf/AS/E+bx8SJTysUnHc5xaFtZLyIMfGOwD+mcQiTEn+q2OBDtJm0aTWHe6NFMt
sgbiNmjf7vjDglGf54O9DbVv/hR8yhPZ0qcPdFqpEEqIA05S7KY89lgimOJZO9eH
6FhODUQH0hBO/ChwbpxOwHlVJ/qUPI6vqhlBg4ZKtZTwkNfF77PrIc8RQxb1DgyD
9GEMNauvmM+zKszv6IonjF7tgjGuXYyRGt5guWCPg01xBI0Yku+Xuyx6AnXoA7xb
y5sjqr9x6H7ob7ukIhr3wXcdSGlwnfBC0O0SvPW38lmHKQVQsTLEj8OQWd4ksxRO
NK+QCZICiI/643cV2MYxraEyK2e+khru1+LMCuvaWJgsvNi6JwexH4fXThK/dypu
EGu2R2lqOi2QmZhO/ij0dOjQ9oIpjZvlqlbzR79Xsbs7n/FOyhgoaGADe66zMw+h
/WzVevVgu9kaUHeWBCLlyiSDLFUYdBR2PNfIrtYzaiiGpVKjl8LGa90Pg1GO+J1p
S7A3zxSpT6DeKGLaOfhmY/0/5CsXLmxQsfWYzCMb+KKWRrYuiRIdnLoHyJDQOw3q
0f/pg5NbdFgqb6/IRE02VoOyz+d0N0zjA1uSv9nNNECF58m8emKCUibIkcTzjxdX
NkkNeW1b6zMICm/6GyH1uKJ1S4OpplAYqt328eQ9Osm16FsF8PKjtnK7eVRYUmGG
Gi+zmb534pE/SliaXvnDf5ogHSfPlg5vdYcZdt6vOPHtMd+RrqPwGOB/46wWrjHi
5HRhtVa7FT6oTwPCwQ3upTS0RAOrEWSbl21qCGHGozS93ycA9BtZs/NfUDF+yLp7
c8u6r6r6yFUOibZ9gfrOQqQJKOwUSu7+pavc5tWgaDDIG/cjOqmI6yFHQWWC6QRZ
NcgUo+TKokKno9811dCGlJAJJL5PzSGtqlPtDjE8+BVL5UvMf4t1DFKjBsIbD5hX
s1B4HVdwTs4MOsr7JJAoJINXcJtORP1+z6WOxPTU+tRNgHBdRbQfgPPNe5smxSa2
ghxYi6TP8OioGpFen/kDDZRSxKO8INLwzYptzGzDebqROBpdBOHq+P/ksWLN7mUy
PiM8CcSfu4EdDRxKHucVdyG7k92JxHGyKGI73SGzrSi9QybXbURka3yCVtnFFsyU
feiLcJPMLtmwlWBytQEe9uWrU4oE9GvIzYjeRjVho8c63+WC34afioXi8VTnwYRq
DMENH3c1VA1sVTsl3MamDrOPcmlyQzQH2LtQG6vJ3fwrjttcjW2pnL+/yBr3a1gd
AN2nnDYcVPhROiEfb9brO0j4ZtopM3hqXgvLzqnifIC7UmfNzeVKYZyD0CmfhLeA
bq01PonYLqoF6rKU8VtmwaZhWyi+t6XVqJeV6dLaJQ47aW5Yvy/hYW45UmI1yCmY
DY7zdspiHqWnj/UjlrGX6fOHgpo3dUXYKGrwaKNS1gEPl2QaeTKUSg/JfOLdixQ8
RwVCRQ01hDywxo/khWLNZvPHJvGoTFiAoYHLQbhZWfn1ZDwLudyvDv/V3xQ4Fbbs
BCaIeVEVOSvPdqwqbDbN+DGVF4A1wOVrR99nnlXTKd1KlECQ/8RirY0C4hwW6fUk
Y9XR00i5MbS1giPOkjEc0n7OpTjSVfvN9ye4cPr6kKJImAfQ9dGRXrCpOHpghTz4
ZUW8BKPevTw3+SOn4QhxHS1B2t/V6osYup3/y7R8TKyXOWMWwGwtUtRxguauQaob
6lfLLbhxOHhAmpcVMiWnE9G6YbL72QDd4Z0h9PIsmfOsjYIJ6+Bp3usilP9TSj8F
vd+QJUKJpz4XbDgOKzKuKwg8ZmUt2XQtGGxL1P64Nb0k+ncZkpGj+OO//F6eqFAp
+NL1EKNce0AWBrgqgtbauSIdTY5Flha6XI/QAR4sBHcW9INLkIwv2zawM117yHpf
a7WnWRV5BMnGEPy4c0oU/iUUbpDSq0yO+R0nubM8QCCY214lU+RCLoRAGCcTIpzw
PleJawXPrTVXg3PEV4hexDepCu602/T5Hqkihna+aTpCxqe6BQ63/Xq3ddYox3Z4
JL9lrUhwpqKSXyvF+anPzBvC3gLQ/cFZ1dE5QURspzxZddy+sCA6/dQ+oltlt82f
/Kw2kJ7rC4k6v2H8OLTo+C38Cm2xK/wkkjGOqUikbxMRYZx+M6He60Hy3aw4lnc6
jZHIU4kIqyzHaVyJA8bEhY1O2mU65ZmP2OpEn5G+NAK9CrxrBiMob6NV/ARWmEEt
rlsbQcKO+v/LmAJiSs5eDFluIGuG2BseZ+fo1agpkA4sMCYyz/wAq3X8gQ5B8aje
Wc+EvH6DTX8UTANs5i7QCGz8JoHagfdgGLer6hf7Heloko6SGtqnll5li99XlK5+
lodxTf2vCnD2P888XsP0gnXeShqqk+wZDZLQpxr3Fw8nnewKVBfoWCqkcnrPH7cj
x7Ey9ga4fHHjLoE3LQnLhOZCllOfel75/xWR3u2IPpM57FQzSrmswTbB+egdn0sw
YqNoi29WohIif7fuWkkUrmQF69TMh+KiVnTu/rm5WcJ0dLJvzJ1RL0WZ4Y8VVtXO
YoiI0HZpv4oi98KFPvI2ZCPUUVGMxBO19zAFgb2cmD8Ky4CbPR1k9a8T4V1zsYdX
fRGHvizV4DGkgMyWbLfD1dJy5HwAyYCmYsy/pBapyOYJmt5QLmK9rZk63dAhYRV5
vZMdbZnGQJxzL0H+bKgdZ69WL97pEZo2ljqx8l8Iry5n9LuvjFAAsThv0yxOl/R8
mrdMZ0sHtF0r2jgd845G9r0gITJSLKvTrNxfL/6xHKHH8q6Q4Fk4c2pCJZz4R6QA
+aLgSmYXJRbTSL9q97mx0z5Vnk3pQoLiyW+CAgGljhwahLFALL+nDQZU02lRxZ/j
oy8SwMjHXmS0Aq+o36tnJni31ZgwnkWEQ9ByhOozdJZ0vpRynFee4M3jLmUmQAHT
Atq6kLQeRVpNu9z1G8wVGg6Nmp8iWmvrpqw8PHc6LQJf5jGzIqFQmRODACl9qnve
TqBtqeaiadGuFykroQUhKBsGxAiw1V0ifDlwKcf8BzvyN0/Ua/IaPyp5U3r4jwpB
N6foPEpefpANcIYVIZYr3TJNIKLKwCNVie59Vz+5tlBfN9aAjvBIn6F91iUwzooy
R+Q+Ij2w4FfB+yqmGheWsuZR3tlmQQrDpO0CZOf38C1q3pgFY22KNrTqQgn+kfQV
A02RWR7P64Omu/ey7jQd6ZM64OjHUPodvmbJ0IXKi0qjz1HQIx+OigH1S8oNF9ow
IFqInN0+0ih7R8GYfGc/GGCY+69RI8p6MyGON68tfoXZZQNrpED6K8Vgi6yQpJu+
CLB14PW8G61SXQ7/gg98EdhpkvMnxhVa+sHtEOaVGbWjmeGS4vj7LSS6sDF+OvAW
9ngMJKojsDZWoMHOulXn9FdY3lGltqBR+3t2FEG0P/pNqjNnSoKN6K77Yg/SpVI6
KtdeaFIgUKPFT+Zg6kWXep63lg0tR5XqrPlUivXakCT3ntNlbbJ4HqOJcbS7WBVr
ei5xzJ3pCCCFvn0BLs0Dwvx/Btx6uFPGe7Eh/0jzSjyFiJEg1stBh42GYY6Df9N8
+CmDV3+dGKUDVo/qSBL0zahdnu4/tiItREhZAdQiWw+4qlH5B8Yqq5PxTSTMuMib
HTtChF4oRxiF70Z1D9RNRDsAGwvAKgJoXSZjDABJ2RRO2TPaRHQ2fiOq7VJqzFnE
hnrkq4Lbng/QCx3OKk/1ux8NG45FQVcJVp3PX1bsASC5jKgFCSxQeb56AxmRi2T5
Z3Qn6NlwpUF+vysmI7wjGzIr2oVBTRP2vDalHlwbNX4dwxpfW3gXus+1K0+ABSMN
j2JIdpYy55xYH5AItmlQejM71hAn/iaamsRNf1SdlkAfM+iQgAhcN8eUzGSjKAD+
rysEYqr4b+BYITv+ryo6ec6ph7nD+sQdwrj6867obOv34bVTf/5vbCczyG+WPaJX
FiV+PfK4LvHx6wywHI07nf5sithejR6QAdziWpBqXXHGG8oOpxfd3O72JERNmtmP
7FkbvH5lrRKzACPDaG4NvNb7x+njyr8fnRRc5img7bZnJsq2asJIu0CCnMfecUXH
Ljmtqd4OzMD0uvwnzNmpLOA3GZ+3v3Jg+4QAHpc+xg6HCEeDTJ3yx9LMOp3mvgmV
1ZI8cnlz/ii86dwYlzpB1KmMt34xgBt5JRy3P1eFcV4zD+JjheJSqOWxoU6ZkhWc
00EkX6YYnBaE4GF39t8vwEk27Uex63z59WBg4GaFLW9yhasaKpMkOJjmoGXdYA4u
tQRoN4D5xAYQ4dF+aT/uIK+JUeQcwhXb37nBNVD41xR/klSHpEkSCvbMJbeIIQkd
zMqt29NQvayiBTlXMPpn3BK9PWhfqvxv+Y9l55/pPxPUSND7cbbUlDd8W3td5Ebo
n4CiHxxqhqJbhRp/biPl+cohRaEscyc/g3HZO0jbW5ow75dYZXN3AlOw/s6l3rrt
S+aMhmRzfrnCOeLbpBF8W6FQZtG81cpNvuAhL7Ec0AzER5L2+IaYsb0/yN5vrSIx
FdTh/1dingQjtJMW9imd1KDA4jYBB18hS+ReKI+MQnhZA8JlPET0OMgHEaR/Dq8h
7bsVERQMQEaEo2E3OnGGfN/s1H/qmIEqY3tEV67Pm0nuyZmnSEJnrdkXS7AgOeaM
Ce9IF2D0mRYM3hLXZ4Dzsh9KFWz4DQqfYB/dDwAJCC5JmfkH1q28H6kfGiF/oKfz
mOHjPgPlbFVn12Ae5mJnObPTpNeBIT7x1t7jzKXgxvCUs2Ph6eaK5XcO1FQYBw+T
z5dQlywoododS5wmZnhgPHpAsxeKfk14pfLQ/aGeVFub4BvO0pEwJ+sja6yfDUyB
UbmRjVWmmBz20y3pCCKmbmQD9pE5K6ZH6AZMisZGjjKCg6sru8GTXAkdyEj5KjPl
bUaD4+w6ZqTSLwvF7HyFfsdYo51wDwqropBdfxS0FRSetbBogfByh6yNuSWiS6Z3
OvyWC0shYRm2sNhyjUUQnHd3NV0+mCtHOvTbwZGhZ4BRcpu3XIOPCou0b64bWrlJ
ocY+a8ww4Gfu5FMehgBdmSryGd5RU0SGL5lCy3S20pZpt0q5lY+6dvCIyD+9KDI/
mVzuus22eE1zdDTFilZl5X2RrtKI8jCLSj85VIbxWRuuupah8Mqga+Otfd0ysgKX
4y0wYEECXrXoxvg6DLNu+Tzt4bEux6e+kMkvJ/QtCwy06wBRL17ut6/7nHD/nxI9
DkySI3bDmDT5q5r4cDMzvhnp7TAXx27b1fC+cQd5Z7ga4kiWN85HCEFbaFPmm/vq
p4O9fLYt5fSLOBfQ2bYlcjwbFpRbemWEjxE8JDgi8+jrgW9cwejgkGt2O9jm+ktu
l8GhfQvb2A14dNK63lUPDngZZjjyHw6Dqf66IPMDwpL3gsYJUz9wTDROJkKh6LZ7
w6KrRe+vzQpZHaq0ECQkQR9ay1wPcFHVY5me8yI0jld92fTv7fcP6Y6+Ophb+dj2
Y93R+6rT0JYpqdxuaQid5nnsFM0bOAAPLyUaMpJ+bYRJXeJU5IuhpUxnrxjWdwey
8onQp1u1KVq85CtQGCM0BTPzUItiue/+w1ABow8gHivXSfV4lyx+6jqUGHHzncRH
GNUyYs8E/84a8cvK3MmPUkGRFD6N1cVCPw+mrrFQQIVIp2jOiyfIpvRL5buFz+GA
IzP5ISmkQnwZxU+U1xmdnhW7BImkPTUrwZVg3WgM6daNqy7AS6yi0MzEIT4uJBdi
3q08gDJdWF/ewyFA7d5EZPJTJl/MiMp0a6QpgQOlxFPdwkFApkG5hohhMrVMNeYl
8K391KSbICj7Y2CeyJb7VYrTGjurhvSPA/VdBUF3OOfXmTFH9NZ0S3CqWvylyZI5
T+fB8VBsqg3Ish57w+4PiQjHhyjIoA/YWcDl7+oQ2YJFYj3zsgUGsXzFqs7B2Bnv
YkEhDdfBz2tQcj9lorzw/dxIC0c22ap/lpYgYa5nt9r0HUFptv8V+AmLaNpbhVin
IMkUjFVVU+e8W0ZD/pv90cLdrqZcfuRR2PEzQyRA4lgu3fbJ6evxGGBeSXHECsYF
MvCWxi8qoMYj9jY3LZhtPzoxa00M4FGbma5CzRQ98ePUPKTWdrTgbywqyHtdDa21
mnfG5EByL8ARxG5PR8JjPdmSfG9WyGjn07aamG4NgxvTJzMitbzQ7yNOmjlHdciP
3gOzTpaAGLpLPS26GxhxS+OonUma2XAOET1KChH8xJd/V6AAwAOFwC3/0AWjmDoG
NOwmNyx4jL0MZoAxT2MZWxYdAzm7dUt0eAzmgCt3pkIRwgGftzA27zFBwr1EcAjI
a5C2rxYXoxKFDNDXPOuYIGUSEcM6//roS/KNaWwIIkP1w6JKLjv09O9rBclAe2pX
821Avby0xdYakJnHwkpjYcedT5sbBWyhjoLCL1z/TI1gZeJYwR9dE5FRXS7UvSQt
LRo1qspG4HRLiGYKMbZ+SAObpHaDlqv00l6UgeawtWKkk8npAmWlMj+vrSpYj+az
n+UcxR75MbrDxpLJrl3pOJA3kf/mWYoIzHco12CwdrFMdTo+UA3zpxf7aCCdEguP
Gdu426TShVwBjZdNzXMTgtxcbr9CVc0HG6AtQq2/vf7PAnE4LU9me4347NSkj+qM
GBnYZltkQQnPk7VO5POCg02mIouJj3kUjAlkzkzHpAR9HtZiY0ok4RiIm33adBJF
pwa5Eu1NsRRdHcdZYnndUuaXK6BEfCu7l1vzInutLB6CTSNQqYAQxUXRYfvsaIC3
BZbRJBYfGNn+xvycgQSEEJFe1WKSS00jLpd5Tmq6RXPek0Z/tTW/Po9EoPLmp7Sd
509KzicjxyojSsH5D69wE2z/VdNFqzGAcGqsBiSjjqvtpPX4B4hjjEUltFV3YL3G
WW8WuGF2ctSlvYrCDQ6jXzF+eoRHBaJ72YsqIwTVHAj1sjyif78IRMfPDLgpw6K5
Miqlq87PCSmx0XlUX+8cjPJt9uxorfgrBxiFtafVvRgQmBYWp0AZl8kvc85nVeaa
DKDetOk/9gCeVmF92IkgGhhdVWkUvn+3U/u+qUbzE/gByQmQPUI/2mcVwR57wOqu
zLeyjARxQsQYdRLHqkavb9aLjI+vaXCwBVswRt307z7npbrLM20TL4Gkp8eh0o05
n6rVlD5CzNC4OofQlkYx+cYOp/se00SoJuCC68sKKlQu5821X7YSRsQ8CBu5UF/O
S4i6toqxZ6IAIj1dUmGhvfZjWJTyh02tc5SfEE186NzWvpRMrZ6hS12ZmhsfsdG1
ifRdJ6Pp/5svJ9jvb6wTGYvix4gZ5s1coTGGjmtgF0DcZwJhqlhJyx1pEw1EwHka
pc9yceF3ANPo7qDDPv7wKvCT8PJBH0SSzgu0Czj51Vo9JEM4pwyv2z9RrY4YfGQh
n37VKDvpE+3o89snE4pheS9xwP1ethEWJ1PUDZzjeemxvCe+S1uruG9Up3bXcSlr
zGT66px5+E6te37uqn38JSAnF48Ij+YNYXZ3VGZLgZpTM7PKuozKORbGfZrKpe3+
BQkXDYCJ8gv7NhpGnpEEeKQjd7SNWaE9m+XQua+p9s9CMcXo54NgAfn3L64lSiHi
0Td4CNjqtev09T/rMD1BJbGtZ2ctvrCUFbE7ySi+qV4Jaj6k+/Axren0Jm3f0Q0/
zRYHppZJ/csM+Yx5zJOPuD5r00nXushy2RbP1xOOKRlqniYfNIfhoir+gP1pFeTr
0rTNNt4cgjTkj0upHijT0PIky0KH2NJIEzBPKpJ2ukeect8wso1l7V1dSkSwdXQ6
T53P4dMkD5TK98hv2cQdeYaNsNn1x7Z+Ap505QgOzuICitWYmjiiZtHmS5qu3B14
0AEWCqEALnBgja7mN47AU0NgF08Ezhf9dmUtEcsqITuiPBhrQ3zMeNQu9WbfFDiV
yNLvcYc6eVbh57aZPA6VrfDh6i7ZRwFPyo47bAdc/41N8uFUayeSlZkUEaqJEzmF
K0xjkHuheYwF126F3Uc8gV6XfdhsdEyOmhgP05+/ji/gxI6OEhsY0YEezeg/eAvl
C9+/GQv8rbxQElCmZwwRerObfXnybypYkUnuoNhm34SsOCvsBNYiK9NvDGOawCHm
evgOhRK0WvT8nvF6xkqFHDt9CmsTC9g4LFBkJVC4ufo2Dbkmv/8IdiF2mCDnS9gI
9q0vGrGXMmri7fSzR4Ox/6Sjo4ZjX6mBnRhddsj0VwKpCyFxaOC80Q7pqlXEiqDu
sCuh8GVp7S/Dx2t2TyYLHtMhWm/D/U+NLqDVaPVxeN8nDWF3RLIgcf4CcKYT6OO+
zSBWMZVI8r24hm68JFK0iDqSwhbP1yY9N5zUcfhCwrcwcoC5IF29EFvcibf61vKs
CBDSl0biRXVn7bnRwmTWuWThGhz3A++6jKhNRUzKNzZ5Sy8yG2puqWDw/iEHGNSn
8FlC54CZI45Gy01k6/eIv6+z+amymsWQ/CTz6Z/LjjtCExIT5rqhEWWy3RtYxuda
YbMjfTqZcyGMdZiKzdkO7+CCaBCO2/9W7ph/zBFigigPC2Xy9ylOvRnn4UYvlNxR
es2+PbaZOxSzkhO3O0iqgeA5gsN8DggGrZ/1WGDsQX5246DKGY9ZWsRbyJgFuyMM
V6WVpN+5edU83+OPzLdz6i/dDnWKEbpsEXTBgh7iLwbX8foOfBfw3IyjKcuZeOgf
yK4tHxKjoC4nVr680fXwNSbxceh0q2WRZSd+Q0aFUdxYgo7yohQwkL0BbBXP+t+Y
gS7Rt4UFmNyGFHRupUUNw5IyNCR4DAZcLveKLSfeANzNp3xqLcttdU41OV17Zg2I
6cjP45ySyAAtxSoszirz8GBQ9zOGwiV31xhGNu+zq2HkE+F8lYZnNOeJ8ZtW9gV0
/NnhwnJGzWCwNpSARWVYTNXKN0f5jBbD91Kauads8RwxHsV3wBmnJ36LDoc4u4sL
vxS/ieZ9qWYzro62fr1oSBTuUJtFifQ4N7+mQgZaxgu0Ey1025ldZdTN7NDt2XdM
9/VTHWzHiL45OVBKjrp3wutyJr1jdCno1THstjalOHoiYn2dcFOMH3W/OuEs2esK
9zs8t2sHhBCR40Jc7KyuRK23XugAtXyoc00Q17fWcLK201snmqU2rHBThNeuf16a
QnfU40GUJ2xt/eiKr0I2mRdRi5gvVOTkLrYy0gn/9oGGidWSt3b9gOYloZbN1jfl
eo39vX6oEyXPael741NjvOWm7EmyQ6gP7E57rayeJXL1m+eRzyWe8qnTxnYsvWnO
yVZnbJpC9bASp3QqyfhsA9wzgkFb3XUTz+uA1DsBa8+30EZ6T2MM3WpqjF/azkCe
UAOshg9nzbglvq8xsuyx6p9Z4tLmARRJt5A5SU4j+NyLXED6LIRYETnpqTvKIIQ9
ETWCsz1VJ39ga5WAM4RGT5NZ3g+NDL0cZ4Zq3XpX9qWfq4dBRNl6Yiog4up4SH6T
g4sv+q79u4h/7s+N25by7pjFM8q/qj4DTtox81TLudlEzvsTXrZIlk/ukJtVpyvb
HNN/+zpBRZjqhAHWpS0eh0DANk+3WYSFlmTk3d9p85erSnkwX5PEFqlMrUWsXkDT
1yIjPe5eOXeh+7EjC+5s7JqNiAeeuzz3qcv6pB0i26kDr+0zEsvyGj6YdfBF0S1a
G6NVUoenniJ+b7/fs02iVz9egA8noV8xNzI7UYK3oqCJOPisshBvuK3DwJqrupbh
55v4Ea56xY+GPkFzzmMSiB7fFloWz3ZvexXxeHtN6HEWJ6bbW1//GnXpFZ14u3Qs
gRRcDVxfGXlI2yFHFR2m2UP3Hx+JNZbbuVsiOVn0iF83H6G10kagQKTakeHLbOfm
MCV17yenlwZGFiUh+xxdw/ZDhlKPSuT8IaZR3k0Vd88rTYRJjimdPVgOtvr9ALQW
jEdAlKkapiynYuTUssEJ/Oj633Cq3Ip3y3bMN/ezOHLf3+OqfOe+HJvuCjA6ZRA9
rpPL8su9zRi2+EBwtafpEb6OLPSRq6tLWap9WpQoy70hxnpouRQRcoryfSysfJQr
0CMty4goZNnfQjMeul4tdamc1dr/Yr36d59oP86eZoeRaw0GD5GSn67hJytRPKJC
i5P2/7S2oxkR9jDia2wHR4y/2O4IYo4W3ybr15xtXnm070lGtlgIlKPEjikq4HjW
gxzdFGaPhoxVVTQ++sl9ubNXyptaWFHdLyZbfl0WxWPWsPg5d9aozZ6stnOSSY0S
n4ZFuPqraWY5viFvkv5VJ9uV4C53By4FyFo7YJcGVXkRJNjcpN0xmmmEyAg1MSSV
Om8DnOGwVLZF3iA6eV+/EgdqA9AYb1jSsFT9CnOUaWQ02hZ2e16noXpX3DxeLnE8
cRAwIBdDHkNZOXZAqeu25ifPZM+9sTywR1ZBm5LUdbfa4HqI9Fd4sKDZFAFTDqsy
luKZbcAfkO8NV1CvnmkuM8kJmNSTBvgpr4yV1C2q2+ARGvtprBA5znNS6dhXFsxh
uKNVPdbUgpNVySEvRfYZL50g+IK2r+UHjWN6gHqC6TKOJnkD0S7Q1x4QYY0OtS1F
WsvyM10IqguJUgwNitBaMfoVxs2dOHwyH09EAvcihVPD8PvdjB019owPNDzPe4Qn
XrtV/Yp1cw5IBOLn8EIiPxmmtNi8WDIXwvDBPs2PqkhjADStDvuq7QQZ4dyDVuUk
yj0Gerye3zsX5tvfmj8+eF1ChDKELYBz8Olu6ipXYJyz+aQRMqxkIBe3E5ilpouX
4IrlsmDtcfbD7tDTljZJy85nod7Yor7H4GIa1WnNFU9nn530I0Jp6bMzlrg6P+62
D2gPGo1Nj8NaaHjuGJwagXoNbRD64sxw+0KSdHicGK5Ny1hkPJI40LdF0x/2mrQ0
F6nVh0sFBHdV1GzDwyBS5GjzPNbEQSX/TGabtqzXXTbS6zeujF15OGSM6qSoZV7u
ELMfZCdm0Cz9aCcdjGFPTVZUywlhBInXi8vyIeRm8TlxLQ4GBlKVD1e8WjwM8SI7
1BsrcNnDv3z1dfxl5w8SggBkhY3MjyhKSefS/YkxNut+yy/TksnC+tpefxS1TSnU
jD4mOatL6bGgg3MnyGH9OeGKIFxRThN+dWtKawy7qrXysBE+YmrC9aS+xbxk5B6J
u9RQQADqdwxasVIzCRbJuMgtnY/f530OHFAqVvq5JY7RQOcgBobKYWcJzRHc9r/S
ok8w9nOL6PyodWt3+CFJCdCHj2cLByJUQrxsX/1bi0yI9UeEx3dKGOyDInneeaoz
hDGjXZNNVXZl4v5BCJVegyPPIqR7s0wmDxsE1s71ENB/91YJlMhRXCV/+d96AJ1E
Biv0OJVRWIbT8YAEy+JAqkMGNfrezktT3CfX/S9bYvFkBp4jVPO0jWTqM2ctevf2
WU23uznhM2rLZ4pgAeigd/rPV4Lc5v/g5xiexOZKI+m3ksiOB4t5/TCrLF8cLd5X
FID2R84wflA8Lg+nC/JpmLoRisNVOe2PNbiPM67jVY+TRukd1v4+8JKNqljdiM+Y
j/d6Pw0BBQrtdUuj9FrVw6BqFqtPV0Sh+oEmGGp53/HUxZS3stlt8TpBLIcDvRor
xRXiuVXLKaUPyhVEwn2R0snhd3pC6U7yaj5yvtE8lRgV847lSb+0zukXRZ9IJqgv
gKzo/trqbmY+Mi1StytmDB+MOkHKdgPkypP5vQqjfqUQ5hY0roGnpkdCrPabRJB6
2Xgvj6jSY6p/Bue8J4o+4lcQjUdQg1Z0y8vHcQ0qA8fqG580khzutlrqWd94D5tB
yeVs6ouMIOTRAc5o7ceyOldKB1TFtmy1hEZqiWXI+WS0x25bAPj3X/3fRuWglqHt
t4S6hFpneNNZVB2Vfn870CvK1tQZ4X4JgbigZ7Ga2hNTm+udcbTgkwCXODEwdqMs
2h9Qs2ex+NfTLUVoQ6SCa74wsauVXKynN5XI4N09airVtW6kLpM4j9mQE3wyrIpS
BSDf6U3ZUuaY65oS178rD9pSYk1S4VZZj1hj2KKMEUBlNwQ5o9R6uxuekFENaaKU
rledzgmC2Q6XGPENsFxv8cg9SF/fbYf61/Hx9NthvJUt351cgVB4VU6mpCMgRCiF
4JeWoH6A5wKB46VOW7Qgj0Es9Zpowlrf3YGraa3FbV78uvxDW4L3BGjJn842P1eb
YLzPz+JAHH7aXW/5kd0j5sT8ti/2L3kMlF8hedDLkBN3RKblhXcANzVqr6YEG1ar
iejtgMva59vVJbvmcsqt6o4FuW4CIDW+Ji0AxnfV+uV+st4KJta5O0BaInnNhLc3
TyOBC2ZIufyHaIthmfJMBPbqVPOnLGb2xcUzv67izR0hi5rPCTJWc1V9kQ5OFJc1
RHNdVmYUJONIjX+bEZVKvYs4N+l0+ZiA0tAgXi5IHZS9zLHksTU0qtu5OXiWo2f4
NPGbYrZ2nLTqbxSIQBFp0rCribI2C1limV9McxgqFvPf1hLxHnnpeLuDHAez5ILH
ZDM9Us9SyrVDTVaXglgsOiDDJcV/s6p+ca8t1ruMEPSJnlViNZS1tneKeZNMOJOi
IFZHwmU6rZzO4ltRqh0y4AG12enK2gipeEhtaZTgFozR4eoKUZ0w7QolrymJV85W
+D3zdR2feHTGFUJiL+EmtLWbfAcmnVAK+J82u+AT/gn5TlmAgG32Jlfmo0RBFEWS
a4jbGF/aT7QoWWqWLAuZ+9GSKA7sCT36XkpJcxmdexnAwjRjibEC7p1b9F9dmBYr
Y1m/yaXjNTpq+ghTDj5TdJye52Dfs6QNXg6oR/bLNEQELOhkroPFP0ye7UnQghfo
PU5vs9IJ8EOtqh+k+DgpaSjr/o4KoQ6pqExzRvoV9LUAztWA9SlNENhj6FcFUmAV
eo4Vm0yRrcVldKeIuzLjrLU5O4EWBBZZ7I0X2PlZPbwk6QS5a14KhtAs/gwzLYE6
QmMpULFR+CCxh1e0sMOsz2RXfv/j18lwEF/tM2krkAfsDeomD6KwUs88IgS9GMOk
RJikvVAR4TzptgJM3QZwzOBp5mjx6pPl7N2erPKvR81yz7T/AzzqZrQFrYiESrsy
BrjbgPqrv33+b8JoG2lq+Evr9Err7Amlv3VyDBB1l/AES2a6/ZHv9fruAjZtKe4d
EixSCnlcKU77lOfkO23RgdM4e8/ihUsqisnbnYQojJPO8ATigjJynwqryO8+k7tx
Q5Ma09te5Y874gKD03l1h7aeiwN39sAPCt30L2b9+HBx7vz1YJ0WWAv6fOCPRqun
kLR2NLxnypQofysO031/8Hyn5f8h4Hm5DShsQWIXtMN3pUqCy8bpQYy5nkKuwkXG
bq4vKWVjNsOsFLQLjYbGyFhBkamlbIzQphvvM796SliM7dYvYhPsdKykd//1FpGO
I+m0hvEHn8TeWW/nqXRPRTVWycCwq2TRhCUtmbNMDC5ur6lSPi9EVzIZcFm9jjPP
Ub43RzSUCNF5mE7RoHiLWMgUHL61JtmMMWA2bje4L/X6iSXiqEJXtY1M5E5wxQx/
ySTejHxtteTog4hH1fsx3MwCRbhmZENb1z/d/vIzsuE7Gi+/wTmozZdGA953Kwb2
bI2mP1aPhMvWpt+qfF1MC7JHKyTNLMhyNIfyEVLzjV0heI5LptReNdHFauSv1PjQ
Q9pVsUTVIcYiXc03mlL5FNM/Zz99Ig4LKtyrGTVJd61bHyj8oVKfDv7ruSb7pPur
9jNvyi8R5jC7c2uBtUggXOUEIqvuOCY/PTgXqzHh161SXRdpZMu9bQz/GLv3tev0
NW3PdpSDpeE9IJNxCM29ZvN5MkFQWuZ9fLZF1eUy6L+8ApWB5mzyr+4djU9u72TL
c0ogBAVyACrtZaxfgEU74OuYT2KXZDbzkrdKTZEJ/0RHCvNerMT47go+z+Fm7T06
T/nu2kfUfOTwML5xBuue6yVNv1zPU3tSdg4PqD5gg3d3hjkSTspBI3Ai/IyFJnN4
IvWJeHS/imPZlEsAqbQHgFae2qe3Nng61SCpdKx3gr4Tr9jpwd/LQwhCfgdFNuoO
6IQ+4HN/bQoMFFaMFsslsohYtxKlZczPJnYOid9RnnusrMVFVJSkbtfo3Afox/tX
+DCCc2GR86GTrH787/14bxtHHSBU2WZjuXFeX+B2qUPG4jS8UFIk0VTHYIOLDMs6
u56Aj8sTWnVZNnaqt13+C1fhlM4V5CMXbaeuAOd6GAzazMWYKSKuhjRsXi4/VGTc
HoZw+CRLOdgguRzBfqh5fvClKDr3jtkBEJJqKxfwj2QRkxvGgTt595D6OrKSbT7D
btKzxeDJE5uJA2Vve3wcuJqYJ83CohZYVeQ8Pvh9EKYqNSikrbH5mryGym31R+Cb
DqZoiB/9q3d4p7nb0CZk1QOuxFVWIEOGCq5BySvqjWZEIZlAS344L8DPlk9+PCn3
qF+uSah1ptpn8QO+bt5zebw7a04xW27ijsEjUJ6RHZAHsr+e0C0Cldqsmcyi3uxR
AN7L0DxNPYnZHwiRLMAKjFjGgw0fowhpWNSMBKKqESGVRFCZv5XsM1exsKlxOZWh
WaqyJmmChkxrpGMV3d5aXUG1wayaSAlELVqraLo+EruNbHuR02NzKuJsjNwVcddF
ARjwhb975398qA3qhyRWbep4c9X/90mEN86lawfzrZI0z2ImrBvlBNuPvQDrQ1xp
GPD0twnk62QhjbiD0/UrLn19IpOjaIBJc3/Z1hEVzYC338EQy5qUWHggVGZmAgZF
nnTTIwYJCplietMmKrdvXyhT4PVT0BREBGMD3K9YFviriihMu71gK93PPeJUxvAC
7IDSdUWldbVxZxeOvwEd+Tfux5j9YVYFZ0cl+ieu/V8V6I0S3WrXp+7q7dx3P6Kg
MSlbNn8as8XiUpqjTMec0p2P/5gMkLmB0WhPhT7zuTLFSxR6Z2VjXVoT8beWUzfC
5jKPAIG7bmFbXsuAIyvoD3RohW61hCmUwiWBGT9/bt3iO4tg/0jiV3vcCgrBBjh9
z1nC24npfyetTemYJ7ClRFpc9mhdn9kDqImi1PZNVbTRjiL8iHlBADV47/7BfXik
IN4v6zrolrqGSOg0wnJEYYiYaG5BHqihvgr1TgEJVnm0mJfZ+lwApuwOWxBPLToO
GmDLaftxKnKwbx7msKZHKTd/l/vYbif+oCqIJAVL+oFXwk1dHXxUdoZQIq0Jr0Qz
92YTElhkqXMndZa+7p6gBMiETVRyX9LN/bP42woY4ncxW8QBafICmSd4n+67jU1x
jSl1qAn6LfpbhhLGWmv7XI4g9vE0obOdwVcO+2mKMClyRFwOfh1Eup3EvQMg2Kg/
jl/0N7vmgxH7CXVuYqPr/Orwd8WpZaFw+zst0O/z6erS75F7HcfN1tN03E04FTeG
92BLsR9FlLjwOBJ2Bj8JLyfC8qIi8P9/diRf7FpBxkF3vXJN//ewqlEs7WF7tLaI
ReFKtB6iUXJHmMgw/yTr5z7h1pfUflDmN5dkIzo3KurdEvio8dbFMaubjvT2bPHz
vQGLpMZrskt80uiQ06t6kZ5Am6wMbUJdGa7n9tSwKHCgiS7cF7fUiNj2ufm9I3JU
Gfentpf7KZfOwrUdx0XjUNyEFt2LmLRwcfOI22eA86XysuuK3JSpZ13hTqhHfOss
M3oe768/Np5D/8ARDdjWybiwTfN8wvtZbWfL90lB+47BfTPd4RL3kzyT605zi3dI
ge7lRbLMM6V7/lt92gzPwdUGFou5fvXMTGju4szVg09YyK2ErXaRjoiSRbgbazB0
T0mdpRUG6MpFTpnY7HOcCvG9FJmciEXf/APAhy8scAgkns9F0x4ky3KkVBikzLz6
8tTfa1Q8Ji4OQY3pja5HbiJ5TC9Sg+WaO8VVjH1wZm9H5zJQO1J5mrciWhEDH0jk
dMbNC4oXrEXcN9BvrmhQziJcsBktw01drcnMNjSX28qClptcGNLKbpjFBe89R+2C
Zh/1KGocV3BXYoO+siZrMzogVcMQDxNySf2EASkWwEWCoIL/X/hIbddnGo6d7sH9
hcmOIIyCHPNxxGPZEYs+xk4OvKGheZHdeGEphUxQTOybYAuLp0REdTy9quwpX1nS
wp5s5k1tNsUIe+K+evFZ9KXsrV7tnMVQhyYzgPJUkEm6ZT+VvM3De7FoHrTyOCvU
H2k+Z59GKIgkpI7lw795U0msn1NCDMtyD6ewqxGFSPF6s35r8J/AV+jUiZbvZVGD
ky7lMmQAtf/FvbBtf2AHmSQ9IIPFvQ96isDxnnMQ+mKD/Mkl8yHI6ZdkhL1rYkUx
UFpw8wL3BWYTCwRxNWZDaTXTZcC5TMJLKo6/l04ffQMACkPahgYghBJT9JOVo0FG
R7SxoDLVXtHkXU97Ue0l9A+gTwucfKRAhQvxEvLPK53Is7NUfTCiiFfVnaz1oKg3
4xkogm80YA+150V+gFPygsGbF5krH+6hYzO2TG8wI8B0GjeKWURu5PCUa7m+ARnp
1XKzYlgQ5KjgaKdJWsNRRt0WGPgTh/p7Xsh321y3OfhLvhibXmGiQmENmiLSSTwT
UNC9v2B9rbAr8iBONk2j5QBJRr9r7BFb9dai2QzdI1gIsWpeQpzHcTLdMP/vaPsB
Zd98AWY/mhkI53FJ4MiySs2PhdWRN4r1Z+70cKRGUi0vgAd8JvONLBHlSSL6UIGh
hmNewr2EzauBBUxEEBAb9Abq6uGL96xUZ++iF1TiquYGyDlw0JRwbY1hxM5MRO3U
D+C13jUoB9ON4VbiGoPS8pWyQQvXOy/v6n5YahlZszbTPjGrxvp9h5JAlbTCUTJb
5mhS35LGD4qrcYDtRSi5FaC4jz2qb/liaB9b++s9zfIhjLxZl+khFhwe7rnSRTPI
lKsSF0fsWBLzZmNtk7IPDgh0PIqU+zVQjuTziFhMqXm/ajsgp3zecZKfR9Ros7MZ
YBYiHyqKwNi+O0rQdU3pbJnGSyJN7l5TxxvpBUI112s9mDQePGmypIfPlayduHLX
wwc7wasXRLNUhu1TzEVUgT9sFBSqgVbVC3hgoMaCmmESycg5k3sUyYT6x0PyBlN8
n8WU0D7FtqbgfflYm+56EUduyQm8vB5Gzcewc4sK1QACSddmbgC0q27kg9y+YSH0
hz4n1hzTg3yJ1Ukqd74WMv6ukgOXzTK2q5O223CQ1LPQgKtfzHUBjPETTPJwHn57
R4tlxAdugv8hj9GfyV3f6lQAZ4z+X05FkCvosYvk7AjqFjxZL4UC5YESN8VSjK3o
WvtlUa5SXpKIe8qoXwu1ViYwvvfBH2h/HvJjieThfORK01jmolw4EoMab1/MQspl
9N7W7MsaVYUee5i6DexHm7La2CTMlqIyN8PpkF6MC4eCARJ86s+QMuPaF/odElA0
uOEnMJ4/a5h7t0Nu5AiJZ6n+q5Ejpch6OP7EcIDTMOGwJyLyc+IVg2yJfKTnqboB
uON2ZMlGwWvN5kvuYvHHOlvbNF1Pu4/GGylBlQDW6PzO6w4KP0LtiIzK92abiFfe
SVeze+2vH0rz7dmyvLhn/mM5uz5zdf4ZFehc7VoSc8XodH1xCmqZXHW5pzkxZcG3
1y9KC1SgKYhCPyADRILb6TTAAK51+kOSPp/3jispHHYoQYPewTCpnbqf+rdWcMOL
KlbiZyI0bCGwd+cIHd9kT3+Zduph/F0+7xPGiZ7nLEvZhg+Knwm/4H2GjFtlE2rL
KiSnvx7PNHgiE2WPn9V9NgoiQianN0kc8YnIJ+1fbJsvyuYQzOi3Bp/+HBOAvTiZ
WFhqoigZTD9zlxnORAXTdl0vfb4unPaWebF3wzuDUWhn+L9enwJFER5q0TXe/hjS
I9Uf5NUY3cp0IM3B8YAVgxuAbQ1E9Bd2trXSRjkAIotEd6t5zJRBU7q5kQmRXUhz
+duZWbHcB5v/cXLjhjcE53NWsbiy/U2l6BgkwhGHtXzIaG09J7ZlCzAEU1sdN+Fx
VvnEfAURr2Ka69HkcMePwxowHZixD4GqD/PwGc/B5xs0z8YZkUm86TnsB4GNRjjs
Px4yuR1yZzaWeiovweWrwCkO/KUxIIW6XU3IeJdA8ZCtxJ8oRK4MFaKWsVTaYyeG
zBeXo48AOrwE4715wn9ezcxxnjM/iceHvHFFEUSovu4QZrQu1YLZ7itM8k9AC0iv
4Hsr8RCGQdgpZuQ28EfFgNaVLRPUoZJ7IqohEMb+ikmF9oApZUZkL1jKEjHc+ATj
FdwFryce1yHihooEwNpJ/+FSpCArQ9w9SJrYBGKYsMRnYdpFmHt+2u7C8zIHixhG
9P2GRxcRptTN+o0M4iqJ+BNriJ2qOFg0eFY1ni0lEsmpXiFYHYtAmVyEzSAG0Wm8
TV89j5SLOIgxuWU7F4jhAnhtdbqVVFeVQV+oDupQRIXu3l/5vYXMqhMPX3iBAoeE
Wne0kH5dYkDzCJT9MbiW3sDy2wLIQaGVI4OlVZcmJrlCo/ao9vrcSc6k0vqcFgcg
9Xf5CohAzfSb+3sFcpyQN04FArjDCjVMgMV9P0tKVBW+4toRwYjOolU4td9kEBfF
q7TRcZDMYKzey+p9OK0RoO8ywM3tLwOrV5YMjE31Df21IDPzfW6IkR9gs0D/dr7d
+tk1oUrfpU4cl/5Nacn4IlkrlgKHNEaSRB3tRgTGwycBvblpPcSzM4Ew0gd7yphY
o2RIwoomIncreJapmNaVLTMPbTeJPvaaGFsjNdYqWTU21ulX91DNIllVKvzWW1pV
VWNcVj8Xs7Dvpyzx2BbQcp8wFO77fDh11NmhPui3GBAsCjrQXqGHnanbpT0UuszB
ebDWUv8G74UbN6mQb2hqwp7oFSg50KIXv53LguOqlIkxHvCTs0Zl3dE6Y7T29Jh8
vDk0eWmJ6wClRoAJcnRu8mD4u0ZiyhlkBD6nyHukzwUWe2CKnQg6F1k360hkE8pC
Pn2kbnfxFQ3n2zT8Iayt60AMdtK2dvWLnokNjLrFZhmSmhdT66m6Mcv5dlxmQNae
OCFutkcilK4eSZbJEgh/AgJoQh145SM04n6S1FuMev931ACHBFbHVL+KotRAEp4T
xKiC4DPRMa2hzXYpY6KKiaQ+/mlZzmU9o00fJhAXWCTzqhK/dYz3logpnpyqAR6q
JRRj9mFZhSRBFw4Vn3qGFwOW+QfizfMxi98VxuHHH46dlfnp+emY5jkAmLOZLtOY
adcc/2Z1pUwH2+oVmIF2ZeSyLBGIdmctm4E5HdrBu+SFnHOAowbSqa79TBgK/2mJ
IheyMRtRCkxY14nH8tw1tbOaICwZSLebEI162oDk39lZrSmKclfNanqRlV3qPpFW
eZn9s5poPHcAUXlIkluvodWy539l6346WO1Hh7CLyRnUK3mnZaJl3ldwOK3BdMk7
W7f7FLfTF0JI6DbqW3OSeCCGolfHTk5kLzYb53xv41kPhgRHA1adbWlozPvly9nW
eSSYk23Y4uBwoVOVZ4QE+uAMJB9m5BWabMjIur/kLnyaKiYyEbxVylc4Nvsi1q+7
fHUkDYRyPn+ClUUY+jJcNfeRWya5nRSG4F8RCjez5RmkXZI0qFnOXqySBUnkuVUW
VbuXpmnFmfEXBnAtQq6YipoElwbJRmWKo2jCAZsIg30ALHErg3RYiMASnokF94yb
4WVRf1Y+uKXNtZ/CFJtPfUtH4D9swEJhzdBB+ukMg5zjx0YYxaUEKhKD8U2j+F6C
Z3eMi3m9bcm3iAWYD4aBHrm7s5dabCs5VQ6BAbYPmlwsztagxOP62y3wTm8Xr4Uj
KMxxOlbQ0CiXcsyJHT8mqiPtOmBSCv8nN+/0RQtRV5lwCXtr4Zz1A/3xy+z/AARP
pKsR9aUzeRI7jdMcEn1VZCDzrnZwdY27ukYn4Eve0V+nV31Xe4Q9YtK2sx4Jb0QT
2chPnuKdGgTmpZ8xUkYNthPav931VaqxDm9sgMxTWnFgBDAyAAUVWIkqOArnJfRg
9gf456N4arLai9FIWErnO7i+LlPlGnr2qnfaOub4Aq2VfaKOU+RIaWuJsJMiORf+
C+m9PNJxub7STvgIVlGbohJtidjNC18zxLgjm975gMH+6BygHTEKJT5wdBSddmBr
HY12juDCFfIhiPF1LmxR52FKdukGbtXfB6IhlZIN8b8dFOudIgz1yVUNeRtIAELZ
KjYAsbz5fmLh8tq71oKoqoeQqaWRQutr9QUBg2ZoYD9iyxyUJwaQMTQFsy9ZYKy5
mFbvdPPJ4lfEbOKVHIdBqnNvIxxVseC8xpK0iuga/Y4XsuZyZ8zlFUqPeiJNFpLv
xLSCxG4lS0D9i7UuNw8J7nj6SSB7g2vPUhoxCj5IaieexQzFixLIlPTcOE8hx3rK
7dyBa3fPDXuNlfKCPKTi6qX9R4W/CDdSUdMeCcDiDTngXmliACyDdq0tHz1zVBJL
tG0tB8LF+1TvHnCu1I2WgR30jWLtEGk3uz/o1SWKutvoSPNNkDcrDZ3N0wwlKZ80
+Q/0U2ZOGhP6rb5JnYk/GTqH8dvHVsexpjfefeRWqn+P/CQdBwWasM51fma3fngG
l9n24n1SsZXVFrhmJi/yw0CdKnmxz6vzyYkc5Uoxm+8nrWWK4VyBmg2B1Rq1mcP5
gXdR3AS1vXy17YUujn0vhHt0BLHnO6VGm4yed9uV9mGns+ElT3Zq/Gdkx2lu6vkb
4xre/zhF8b5vDGdfnGcZktaugQfrTmZMG8B4AMWa/wJ+RO+LHMTUg4q2xNuEF7i+
LlwKBMo1+opCH49nXywCDziAGJzyZtNra1RHiCtLwj8+CPEFZVcpG4gStAr19gD3
a6jzrg/BQEqBlgWqpbg8okmQqASGA9m+0iJ488EzRhd+qkJBSLBruilmuReU6/c+
HoZOAl2758dOHOxxjzCaRFf5cUqCxBtHau5tnjzsyy9gZqxmd6PkoeKfPe3hlTpt
BxBgAqXTNU3k6qE41mNBOp2dS+HVmrAKYf4ayh2hfUHpn08EGFX7+FF2KmH0By2P
h354ig76z35VoJmrPbzTg1XrTHuxWghTox2OAQF+MIGrsviMVrZe5oHXUTj8NHEw
Mz12n+fCqkx8fElIXn8hvab8DXd46iJl6B8HpyhF+1Ck+NlTBhVJwvRt4IlkD++F
o7NxLJ3CbiKffMAHgdd2TRENZ/SLEmZw09gGC6LwPx9KaWykOkq57cCBS2wKk+wp
FJsCEFXwEgcGXSgwwhzZLjPjPwaqo2Nk4QiMkUTISbIsqgXP0Dhw8KV9e/hRD020
Rm+hUcrHKezbnljwKnyj7HYge0FfT+J40Z9m+67Of/N6s9yMTr+wZVSjq3Cjuo8M
FKR52+NitIl5IgFID02WThSpMGxx+7sdyd1IAnawsmogBtT1DjZ0VKnO4eCFVovB
u6XWqUtym/UWomUoqYHYcD/DJXiACJ/FEcgSAflEW4fWPpwDfExYwxWSMno8DqSF
V0Tru3pkY8xLH6e4Fs3JQy1YWunDRZLV2SpcHpWnyVfDDfGyN8SAiYmQ/sAoCE1N
NXkXunAvhKU/H3KHGqX8jk5tKDsBuD7ue3ooSK2pcjP1ga3bF4Vu3RVgL8ZzOhPI
bu7iOLGYYGKjiqA5ZOpiZc8c8xO17g337MUjizr/CJi8GvonBjT3jAlL8wB1piQn
KJWaO12RSnF24F+C3FGYtSfKOlr96BGpDpC0HXACjw/u9bPvPrWSEAzdBlbo+CgJ
okX3i0WsP/Iq9SUJ0G6vkir65cxIEpSe7fPWWqoePNPJt6UmPcaDTXOHy8h79yuf
zriwUA9vN1H/WWz4tDSOPFLScR81qNa/9gGnECaxWdo+c4NRPBx7l7OgQU5unzmr
TqNscxuaNnjhOevikjP1T9ieXQLzOQDW5Rof2qJx+SWUW57LXs9sQRorQmjCgNK9
VQtAwaPysTlu1EjcnsOs24OoF2Ofd8hI8ZIfArIrVF1D00jaVc5DbIeTu7lJL3Yu
eGDyMKdJPdCdjp/O9F5oKVRQY7GJO7r/IbRpiN2xfQOGPb1ND6FfxY1nw4/zzd95
8d6xlStLxrg/Dn8NZC6nP+8kUF7qpf92POREO9t0tMRj4ZnMAgSkLcKGBBHigO8h
oHnsnaJkH6axmtvqTcr9m6NJlOMBYC9kv03v+ypdwXEm+rAQuqc1atIzeprRx3j8
jLdpVGgE0OjTxb4XVgoEdoWFG98aB9s0pAFK1JrA1cGqMQ8H5oZe8pQFVT0mvoQC
tGx3gYGfWdI1xbFXtNHE9NselFkGk7Suo97rFK3o/cmROCPrRzgbDgzfWvO4sPDO
wGUEvzYjl/3pmilqbJN2WNvIj4Qyikc9aXqLIRXa0JHAzx/ObQp6rLMvx2Ft4lbi
53iOi52tXn6cQDo+wpBK5gu3e4lXzcYUSDE3cCOQ94p0EeZkHuu4WkQQJtnjiWnq
kd5JlGeOqWQ+3Bf7bePsOueochL1ZE272U9qhb/4Lbarosfo4EqoyX9maU1EEh8d
yGKtWomYx28+Yfncqqq0NzkAiI4CtUnkW/H3plmCzDLJ2yE2iO66dZaYlSJm5cJz
OpovHJ9kymifqy1Pwgy6JKU1S6av+Zt8AaI5fDdbr6+Ak3Mnbhl0lSZt2U1DXr9w
St0WGsT5mzkQAVb9NjKpOzll+Js8uleid2bgMx+mCzJp4vmW/im65xcTmyL3cE5c
eudib9Vopuz4rZ+1RNstXyQRfYYcmSJZDrPqF5lB71Pm5KlLU1mmOse0LkdtODmk
ISZEpAGOZF9aWtc2XlshgN+8+n+6wHxfQuSLtLK0P+5iD3clMB+Dy0eGF8lx1703
cXLQXjzUTmgEuiWmMy8E0NpGkR6ueeHI50cYiBlxb9nK1Gq1qBpSm0WvzkLPZftH
mrtnw7qgXWHzq0dMRZrdlmZucWqV1OrUV6USpRTFmMPfVkwBQYA5ajzoR9ksvJzV
M0PHc3A/VA2WpTvY9FLyVOxzZ3G/279wx+NKPQwXRhqTro5e2J7dnnGGcB2eCmvk
3UKTpanQJQnq75qwAryA+zQhWfJ1Otq5sM1psnqGvtzt4b8MjFgKyVujz27/T7Qy
n9vfe3UKhsDMO9jfiJZyKNXtrZPXzpCjhBZrY7WyiNy/8VEtIPbiTGHqngpBC143
nv6OW4BM4Njo3gaomSUyI5kM8ySwGDtlHSxr/MdYAmMZ1RE5wTLGwxqErbj3iHwx
6TwdRQVLAI3z6l6PpPFz0OZO2rEgl0IEBh72twsX7reYMR/Xet/hrZqZF5uzuEZJ
M7hMacL1PJsZulA9xiFKQfqLO91xgj/2eBoFB9akulj17RP3yFxiNixATdCR9fYW
GNya24+SFsr4yIysnfYN54bxjr62iP3v2tsqI48lLosup2Aaxef1WaaK0qbRk2pr
mKwwZN9tXzb1Er3oOS8PYC0BPmqd37ArfOeeAuKlZuuAX9B9lJRcmu5ONqjkcCFn
yoAqxgZBa7soxIXTwZ6mzKkMQ6wO2E3nEJqBssYAr4Zy9QCYncBM/n+3xGmqrVy/
GzrMVT1RkziZ6JrjhiKPTlzeKtLFReFwsG9Uijdx96Xjh/6vzWGhjeD60XXxHIWM
tNpQn0IKsyPQ47CrYG6RL8Xuz2OFipcgsNP/Lx5FZaomlUh4GGCqeznSHv7ktzdg
RuASICODSbnFFnLyyKejeiHtFxCM043up6BwdyIBXNGHmei0Ws/1dpa3fsC9DTon
WBh4ncOXnruse0SAMTCTay+FpL/2WVgGfzdFKN9tetcdL5iSiSRUxe0MeUwe56wp
5tq/oG9/8fqPPk9WgGSgXTN/aybSaGbCXviJHdnshr0DYSqPU8VVUftb+26AJpSs
YK6jtDVCTkoP4ONsbYhJ34/js+7oiUaPzkksPcZrG0yL/7LI+7pfnfWrPfIZOAkc
TJ7ac4AHWIpVoS2NiIYJzPDa0DNNQpnelqVRIkgKoSHpht3KnDBHq3at71Wvajuj
6jq8oTwmuutupmqsGnIrM8/4eViECvWwptfarbVZdPKHtP1MTfCmaKTesMbp1Q06
0HaVWqCiD4wOW9FreAKOS1yAaNIW6tUkut6vHuPGe/Q8fyi8tvIO5PcCchxfy1he
ezsma3VZThmRdEvkah4RDT0xicKcqFA8kLp6EDAJYd80tmC3ZX6hiZq3BdO2TiWV
iH7CQN0XMdt9HgipULUuvtjQv5/7tYZynQI3Na9auQDKJGplkA1uyLmQY/clnZVs
85DsP5IcM6UzyAGjLqadCAYelMiZiLbw7fA6h8uXefLxBzHD9jAu885zCqsvFT0f
XD3LxWeqVdflUOKsxcZENLe7mwdpn4UZFpXLzGn0P82fec/61H4XMNBWk9YFC75y
Zf5Hs5e23pqN6CfXuF5+spR21X3gMFceqNk6B5WPJpJO1iF3RD0apnFhUVpjOFY9
guzgIFcliMOWpNiDM2p4yhHDcSQbyBMsuNPIGrB78GHGrpXpXp2eP1d4OTwpFE8v
9ErWeBBlGQezLQcucJfdczERv+1n/SPH3hyWc7RkNLJs9I/rY2cLishpjd5ItK6a
S+OpbPeB7/Dor2084ClWLkrLcGOD3ZcPw8GwBDzSt9j6+Ucfazwhkzmj59R2BIBg
D8WDyj7NSql8gAKESS8lZzC6CG6KWYPIvMW4+/g69zEmlGNhQidOp21QH46ftav1
rVY0nEnYuZYqhuuGdgg3hq/IptAl//29Mvh+HxWv7vlz/ahUMyy7c8PcONZiAvEm
UkrgerGOSazxAU1j6qZ9olRqeF8GROTmh4WcyuHflr+I5GG7BqupVrU1yBzE4Yft
6exa1A7qB2yJXr+lloFzOIW8x+xHgd6L9TAkEXrrEv5TYi4zRLN9BYwS6Y+fzYEj
7ytFJ8A0iCiU0uJ/gtI6c5VG+RjZo5/ykfy11s5A3rZnFYHIGWpKoammE6p4W/yc
kOaTgFG2M7vTEwKY9RbboSxz2JY7Xq47gu59df+dngifjQXnvLQvPTARLZ58jF3N
AIv0wOdFMnWG+38vlJS42sSvV9Qk5OT2r4THM2xR+D+BLg6MiyElKzS6jgmBJ3YV
n4Zocgg5k7Nwarj0EZ6yRVohemmmkENDoAfNA1xZjk0G5wZFbwV18LSWrEsvIlPa
jNlEPH2fQPnANHPnoOWqTElLKAY6zhcMw2dcuvRZJNGVt1oun1vZpI2V8l51wKvW
czVlunPflI6E3VFSo69IAHBzyCtYOwGwW+P+4C6lutvfrmuIqctc4nCxdApXxM01
i9+QQIDTupN9Q2BEeP2Y9T0v4fWmBgALnUnCPjGxnydXg353tHn7Is31rDHP3+oD
ze8ZctntOHELexr2xTUZEFgkXVlFqyrxqaTnao0e/TXBa3CIq91JweYwm/Rdtgik
jXA4DTd1Y5DBFXaXF87HmbtSWJf5K5eRlzTgQRTFDSZzIVVaLs05nEHVgtlpnZmB
O4qfizVRH8og8aJhcIsmFlL9WfpLeXePUxV0jCAgu4c5cQwje3DfwXClNylZy6N7
pTMzUY2rOkgAHPqAtN1XXrWfCEk/B1x493K1C7bj1RO026ZYcXwASc3vKPZIvVAB
MCOFexF4ZPQMbjrJg53Na07lJJFCOmmZzKQOmEUpJ5oBQF4hnt5RgsXnLrgPEJzl
Gmh1z2NBz1LqY9MBmmnpn21mJ82gNzbxZhvk975aS372Kujrx/1ebZK0SD0bD9y7
f6tRrYToq0CCXIMCluZ/mi1/7DnoPmWw943l3qlN+CKiwsuKdXn01m0yrqAvDr5I
V/vo8l1W99CeMNgqxWp5sviBJunNNKmyPUlY60V6Alji2Sa1r0Zey5qmFisgZiHM
0AEoLM7nuahz9VBSoeavl56vdYR/xjyFU10RcCiNbLNpmkmNYcC4RStVQko8Yde8
7imTqLasI/xs3pGk+yLhxVbqeNckUoXyMEX/iJ1QvGRRoWVNUZTmX0/ohsQ0+aqh
nBzonHqMUCw9gRh7y4VM6W8tTVDfPgIO2qL88tPXSNXTfj7EjDYQ5yfep4LKQ+NT
24CR6+X3gW9HiicrQKTzOl6vfjTttq9abEH1KJiE0/iQ7wHHo+4Blr7JJZIEi7Uq
SnUMNJ4ryEFi7sytRm62GKi6MewIXvPthY66WtWv8GCrIDA/mVt4zqlAK0kvByAE
a/ilPjdQUawirh/PKVpnJqIhRHRHtfVGwgOBMruQ4wyq+LIIW3xc+DSONFf+JOdF
iArUnO++RJkwQNwimQgvIu8GbzEJzxvTU8NZqQdBwAWdUiSaOGRbQTNTohCOB3Lx
YlevQXIP0MQj7gaOrzHR0kRinICoEnMZ87Olpds7Y8ALxaBEQJ8Puf40kGctcvw1
yLMfLiGOjHuguxI57COT7zXyk5spg7sE50GOMUvlW4bk53P1IV7aHxjwqCPQimte
mIOAeO4PH/xg0qOqJNFd2UJ6CzwlWN/w5c+B6hDvNSjnaWbumuFb9ibU1UdlLe0+
VjeHiz5+2WoZivMITsYPGRNyqeXVerIoFpOP70duAfZI80QkFU7sKaStjXhRQjq3
r1WmgJy9i45Rb/saakyj2uQ7wQE6dFRGDzSdHW+EovlgoAsNUqUWnr14hjJtjpjc
JXwlad1+0PUrTBPTosG2H4EVLAAgejFEtFcvwgX5o5eLxetkhEE6CLBi79BuBa6W
lcTARFCflkJcugRQ67SBGW0cWiHLGcG6PycHp8Kd6t72GlDXTyagV00uf6AtJIqy
3Vfwm4AnbkAyKnfM0IZJGwUOCiFFDZqPsFVMRqxMqGrLlv+BAxywtLvLy9txanmT
ejFgrpURGFlTZE7wORK3lbVMWPBTa4qSgi+xBvNw/bE1rnqw/+DNQ25j1YbIS35N
0VDNtNDtpuPvlSelytMQKCBQXMypKrBCAXqOaJ7NhXH1wZi1h9fL3kLqNwuvlh15
A/doc41cl0h/iMgIAbjFI4WhofbpU0JfilTDP4Ayg29FeERao2psi+K15c2bfIpx
uvkGKg25slideshkF2aDR++s9Fri+WRnCG2nQNByv8E8fbkykKR9+yAf4bVjggbW
9KlTB70nG6zfnHtrjvfus7EqZOc6mzftfeYeRZH8SJ3URKTGIFZTVT/eH+xLmHhS
XXf99eJyQ4YvuIEHzquFf7msw8vGQ137M+ENgjenETLZWhF/hQogejpWQvUO+VOx
vAcVQen1hSfFcSOAfg/npMutPvydFG+MRqn7mNQGDWgN955YWmlwx8lF1uqP0QWz
Ls/GdYgoZX9eKTdzDhAwcFAoNusTg+QgQXMmIShkMT9E4tILw+eDBkbKE/O9/G+6
BqItsSn2SYUUGqjUAASFULvWN0SDNuQd1k/qkV2i7V9nQlFsX+6vV2Y5bggpQV1i
0ySRaVX8Di8mM9Ek21r0rDQQKPvi+14Io1cVN/MPW74DjuvKIuiZ8ajok3N4NOpD
FvSl/2g+XpmZHeereuE6RNEODxeuuKhW5MSMDsc79KZb3QAx5PvSqk7XfTPHaBS7
K8iHVcHNddhDmMVIT+62UF758Rm+F2FS6UBQWOftLzzs1NwjGhKqloEiJl5hz6Jh
DdgZE4wrQzpdENXFzb4VUOZXXqiqKJSn3V/Zia+3t6z2eWVmhdksxtwK5cU1flcF
d81wbNY41D4j3lwTooHJENlF1xasXUMYTYgevfxvbBFmwIDOjQLfnZjL/IkxxKQE
OtWOj4NNkFRe6CTD1HUqRej8M792i76980dBnY0D3/slDFb6qeanyA6HxWNA+rqt
fMWQTeIlsjjnlCFqa7J5a5fljJq6kv+XNevuhuc9o5tyM+tCKgt6cZRDfcH3oGIJ
vbnm5TDjq8ZtH41Ug8tjsV7+RwawOPd7WpOOVAiqbL1ZtPD1i6PFOdV81PwgJmGU
NDVsCPDdqfGWaXZLiKanmaIA1gPt0KnyutraZonButNqT41PHYnnjkjUHStKcgRF
mgmb+drPmlOqzIwLX/T5h14OFGLgypQI39j26GjminnhchyI554GinIEo/b2LFta
ofCD73ySuK/jRdwPBv2DtrKs+XH68ccJcALz9DiV3wsS+qqAazWe8JjpGxEYSyjJ
0kW++wUKQMgN4mD0sGMeTuDrWA/21Kn1pLdt+TNUOnAX2W6S1Ic1X7vGLjnOGjVZ
nhFZPVMlBC3iiTUJr4FowAGBk6pNdcFveYZ3zN2ipZ46L7ruIwUk6j93cNLSDeyD
67jbAq16MeWbZbaR/N4ERvbF51oqbaPxDbC/yGqE3HbgcKtTpO8bV4YUWeXOn10v
D9ov87gmGH722DAYF9W9xpGnxwc9Xt6itM8Zn/joEuURkMbNlLWz1fBAqabRrnrw
q5sqrCMcevw7sXr2vm+rxVw4eckNm4b3CC0BTOXvFUoZCKRAmoZyQjHwX2FIyCnP
qyUT6PqWEHeH3ALVn0cQ/FOQNwR74vBIIYn2pZLwr5ANNEK9fV9IQMIbNYAyh2Fa
fm/SwRdynrT8YOPa1suD3gOg91X7FF0tx1PG0oB8MnUeNz7Cq7/4N+1Cb5b13r3l
fQ1DJqYeJguwEYOqw0QBc4Mj4M81zvHhtOrNlgx+GPh1UWMvHKdOA3W3NpfLq0yr
yFMNLTg2g6yzi6GJD7Aa9sCsDFs9oudLvF8ms5kozeyV3CfHoOJv6C300bQrG7zA
ABA1bjCXzrvJY1PXj5KaP/TRKDET7nczuet30yciuRQczBnhiZjbJXHRIoa8rLdB
UwZKyTY80AoC6AqTbpUgnLvTQ093R4nZ/BiDDcRXggN4h/CSWIG/OSxGYW2gY1IE
cXicNP6EIdcg+mpTvWCuOjRrqG2Tt/9+I5PHDQyM4TeXEnLpEvN+lC5iS5mXQxIh
SVafGCZCEgws4RS4hVwNB+Vukn7ZsMv9AQa5GBQRgMYxnslZF5g0tb1jceE2O5e8
XLoI9XBwf1a9vmSDkwzCGqdpNEtC1I7rPCWl918L0whcMUj26581SprvMd0Q69BQ
5HVQhL87q57t3zsqUh8lyQcNqG6JsHxnUp2cjgbSWljopI0yMU6V87r5GyoI5XD4
axbnx4ZRf7AJSWM/IxrfiJfbrKqOJpCgR6Oo0Eep5Kmj5kv5WT8KKBSS4mgfTWT6
fRReeK4XMmIYYPXRgjX/5IFABsghigKYIifmx5rEuqa2rpGA/sN6HRr4oZyU06Cf
zfqGw06K5q2jTjwaQwPQm6Kbw8y2wuI7k7jv7ul5CfaYVSReAScagIHCIsJswLEV
uJluarqrkmHB4eMm+dqUN6jRyDKPeo2ARGMrmtopUzxhhV2nVEuC62KpCXZkfL58
xfkNTtRTWMhkW4ezfGkgczTHMBGOOtTCuqaTLHhYVBzRGy75Ne7Bkp2d50aZwyru
InkVuzWG20oGiiJnobi+t/bbpBvP2wC+kuRvlCYB1X1xqj/vVuyZv8r0FTiRezXX
x6L03q8Jq7jiIyFB8Un3uecWGbi3W4tesZdtScoxXpLV/w2AnufcjSHeSFlHQjCY
Fbot0LVKvcr5R3OVE15ETF6tn0RyIOOOJnpHx795wi1GJ4tx89AyACQY/ZAacnpL
ZjPFQ5QOggZ/Z29sdm8xyPU86RQZVCHtx0ZhSIUjPwWrnYsrBIei5JHZkAYfhsW+
5YRvTg66cxSQhvccRD5agf63YkuzKgX1jU+7Yoff8h48lygDVuTDR21ppSfMRHrg
OJsgt5u1Gb4j4AP4FcHOXQJ7CAo6KBC7jC6tXzDFI//XD6QtLFyonCqJb+EJXSuJ
9eYqR9BJ6NGymugY2nhzs5RiHeCCeLB7ichgQ2YoAKYN8bQSf4NXEzNzGbxPaUxV
Bez4QUkpqEQJ2SIO06wgg/9tJ2sCLIJ3mIfX08ds12C/Tq8i6EetCV5biN52UOAT
jqcIMW5sLANePOfK+h4SuSiGZOE/GLPIcC6WQE00c7Mm/+I/M8jwgxj1XNkahZ+M
vebXWzDKhrGbhYilA2yxgd9u97StT+caqH9mxunVBk8hvcPE/hRkTjvbzB9f6O7Y
torGIz54zky5cL6usXo4ppXO/Xcs5ya/p6WAZn6tO/VwFPhYetmzAXc0Sjk29jZh
egtso/CCx3tmYwtRo2R16ra2fCW5uf4+8YmX7jR3vhyRw79n/XAzfcTQ+5ly0HvB
TtlYRLEmvFxvNCJbReCXUN0DwfxqMzpwOzDh48WOYXRCJT/ZFJLh8qGbFjlyv36F
hyZbYsxQ4dZjtPARln3rV5bbDn2qBYCjFxw937AXnjDKQXA5lVGZX1D68Lr4MpTL
Im9Zi1udQbnvmQZcya4PN4YXkul5ywH9kK96gzcn9f+DKowwN2olFDTYMAMs8GmX
fq0XlIKZGCReffnTM9fk5/RPev2xiBsJJLIbFxKyIHO4lMp+gulhGfehKCyydHMZ
qpKpjtKRRpIIjwNE3tZzdsrQmbCf5E9sP2lCjTFBpD4Cm9MQYLVMY6LRRMqxrdne
FljpvYrTc6dRv+fas29ByeHHJ5w91i2yEZzIQOlg6plmJoOYOr3uC0HqAW+BVOg9
j0Q+wzVc9TG715qrZ+aGiqDnX1FqtCdsEi8ywdjDddBBhZnYxZJUyjdhsO1Vq0v7
ZOXgTNbozbIM/koMEJeDoK+mxDd+2Dvp5gb8sbM1r5p2+VT+ANhfozAi+9Bs7+XI
y39VSUO/esehoPFjWDsyPEPrCaFRXPODyVEmhYzYgrhW7ym4VxrFADnhDrLbU9oQ
DeV5HbIMpc4d1t23vajR2ZpCcd8VJwt+UkXFCYa1zJ4s92vb3qBSvYBTduWCO8Tj
oa7I652EWs38Z5aq30db/da/gweTnF1+nT+QDooVclt+U5WmJ5VC41gYu/NwPZkI
/pLQypVnHTKxKVeGdTV12tXAuEHyptShBdMWiSPQXoXsdw+YcswKkXgF423lsuMw
9uFr2/Gc8Kykhr9XKqEKVIc/wg26E+EnM6EMNh8HbIYVGIQrWpZQo+rZI3O4sN1P
FJXb5/ex3/KYNWblWWs7b4ifxtcGzp6ZFq9usSOX0p3MxjF9lglWZDt/C2C6V22S
Gdci0eP0548eShUEvEGTC0PXeIyRi52JEs83FYIWZKNHBqzMSYoEH+gJRFpKBRyP
tL4C/0m4nNUUXJ53MKgfOxTa/4V4EF6NHLN+bsMeEtjx3co1hDPEt4Ns55aj9sRx
U0bKOmZm9QVR0MqNIykxSD1MTBx6OCcn24ZOCR6m8mSltwMbbtBnozrfMgGgxnVr
oRtlU5nnJAv0aV8k3yNxKwqWl+1xU1oBreY/oKBE9zT+rstsBX5z1/J/jvRf7G1F
0NjJXEh9oZI/kVKybu9ZaRdFYRT1pHgwDigDaRB4OJiVmNp3FMWdmnAqhvEJOl2r
lfe6CApCLq0A3x9M+4Xwts8pU0KSQSw387k68/itBTP+SWcCcaOg0q70MbFB14xD
2u5wOV3tZXDQ+vkeDDZCXgSNhfKyPvlxcH6T+QoLJ8pumJBEu9LT2WSsKcp/3xBS
FP0JdP+UZ0edTs7w4J1ORU8mj1UYyUjh6vTIUdgeFVc7v5g0ADZ0cqVO58+OGSpx
sK5WtxFUnjWHUu/NUcj2hjKyzaEzCx/wIVv+H3WZYEIvSmp3qKrCEAi+Dd4FVdpZ
sEhKvEnqWvVjTpN8bPEyD7vu4DTzhND8ciHDawbvzQsT0qNQwH6DZpRi4Q20Ean1
Acn6Ys0blc9d4/DiKuGsUYYxY6vQFzJMik42CSVggORjRtODybyA3z7RXE/9unb3
a5BxxoYBpTkXF16ATJPLF2n6fnGWkKWadIyYuDAmVKH84Od2FpekcRF4Rn9v+DJG
cUqJE2rv2fqqQV58PaZTx1TeWilUtpcaXg19fK1FRz3epoy0wGSwlv5BcPsQ/QvX
aDeB59Xyn0ghmglEJZIws3js7Wm7PzdvUAkNGhRIpmkPELrII3tVK6DDnjhpzCfr
IUMWkUg4SPMtKFJUZaGuYZAVTlUbuQcVbsso5fUoY3QOswk5hnUEN7fPekYIGuBZ
uX3XlrQdBa8Dw5SpDFQv7AN9Mn2F7dLXlH7WoGMNA3OwWA85vMe4kOI6i8K2ueYp
npHrSfP1ZzbWUGwD0tuhVwQRFtQTN2IY+eSsqUWssgj/vo5+QUPUOWRTxqMp5Wft
HZ8npOLOpHAoIeE+R03WqSDpWBTuqDGkzF1xqzQzrDfZkdI7C1dE2F0Dx3wOSJVr
2ftQ+KWZJ5Fv3r2RHlirgb6BABdL8L1Dun9Bey89WwtckNvgV9yQNzdUHy8cTdY/
X2TGGQt5Ic+sLLxSH/LIgb0sdpHCl6s4clObD+gEPmc7cTFbehQKfs6BtZFCJ93R
vAKfX6E4RGuPKwA/f/qDgbziVBmU6Bh2jdCcSkGQr19u1Im6MLM1SlyWxprZtV8B
JU78jvL79hbuhKhELDAQUvSpMfbC3vlHqHvoKCk/n1jRrUR226ygv/pYicFkKQ2T
jUYQE6OuLC2fdPbxIJCEPhiw7rVqCNfMarPu1hqNwXl/ppxgiOoiMJxWPUntQq8l
cFjQ/VjaXH9/ijDStG60bI8scCXiFbDa+dWzypucYE93FHqwlQFmeUQ+kI+gy8a0
cRPOSJSUjvReCbCFN0Letm+KZk2agbYBtWc67O5nGCeKsRLpiiIY0J1ZP6LDiheY
vKLhwictBLZEiRSKNER5ZDDOMKlK7VFNsUsFLs5TnUOPFMDBBEfMnl7H2sw2uQuC
KqrTGvHaiKzDKeLVDQU/su4kR1pHnBgDb9GhE0vsTn+zbtISV1uxgD/fMmi0eU8A
IJFmblRNZOqPXTDTaVhPFe9QcNFnJdJ2O5PyUlTP66Xk3I15Si/br8vqAXQo+6g6
KBlfdHJyMk9RRZdrRujYAClf0smPudTjE2eZzx8lwGpL4X9KRO9ydW3plqFouD74
YGkMcpwbnjriTi/AI2vULD9Hl6sc0Z54jObbOPW9jmSFi8EbT+ZxJ3KiS5sqqgD4
oXml7duemMjXdgz9ZjrZTwaP1EvrQKMmrZ86iQRiwua9gFfHfn2ceGRZLk8Fv8mU
GoCPySeh4v0wD7JPTe5LDN7vMWnk6TpyC4bf2F1oU4P6mDvNyATvByJAf6zfBAHL
a+alV5tWEWLAlmK9iwmSw+/8Xdv0Es+9RHrr4OAJWXLwLlRRex5jsrfBZ+9Wec8R
eyUyPtU0jK9uuim9Ew76bJwPWW8UnbqtjmeMd5SMRvSH9rzi8O3UpkyvA9OFPL28
kboruED2r+KjnpiiJSF8tqamgKTIHYToNsD4cq0jyX8TWlMfZGJrisgD2FzXN2yH
ZEWpUOUjrANY6E7q2UJSOKoMD3lOdrZvo8ru/S5sixpJzpeamyd+zE/srpMv9uhb
auAWOm+RpbyG/YR5aAXQcSsajd5W9MMFjuvFaoPJHWlIW1IPj6tBo8ubbNa8GEk5
ipSXdR53K4I74FpgrghH0XwahZii0n3QMZcsoALekeCjDRIcT6MYZWuizrTzGi+3
8eRf8hQBTGa8FL1CgaxfW8S6m0HlFpIcRvPg1Cn0ZfCr5dQPuHjgi8mvtHqcAmmV
VSkqOMCrP09vH62HGnVBmyieKY/Ob18Jko9EVn44i1WFNCOg6MGyAZRWqnpwEyho
al1+LqPwZqd3NvM8T69EWIqQffuYALK62zxwJ5aHadXp6IEAH/rmWu+nxyCK1xX+
O9G/GsElfRT8QcLxjLKFaDuNcLs1GGOWOuGRquuOtM4udZ7N2nN4Tvyv9NmDVG0L
Kd52bD+s0wfqkE9VMK41bvp6DJG71MDVAFOClGFf30QkZOnVpApWosK15lafqlmp
MhdpTKsSDezuxHd6IKr0OsSTtcYFgAMi+s7OEhr0WntEbhTKgwVCpiTmAyWLPBou
G0I/op7NRn4ydBW58MZ7mjoWT7I+qXM+eYZy04ydJa/2TczROudSuiwP/0iOfUDA
NoOL1nDKdX3TbYMj5bQkimtv4pdcuqPvepKY862ae3lH1yXEl2DhzXt23iwT22b8
3vmPF/PLWIAVCrR2kZuitQUvTHiNISRh7u7jKeaDGaokZGm2pfz/fzjkfO08wby5
mR8NaMUaqTFOeWJrGEgvV1KbfrKOhAIOvVfYJu3/0T9GNMnIdKBS4m4hsXUgt4jq
QVrCN2Mu53JRO/1EA4d/MaGXE6TU53L1K6MMs7vabgWReZCjp1q32NGewwoIVFFM
q80JlLCbP/GUF84LKTtKkjusWWrjLXvyYmkE/zOGiIHealXu1Buldd4xalpDVT/E
LyqvUurHjIUBOc/pfcHlJ8GoWswZnm8N/337S28l6+wyOY4A2AeQefjgm0py+oWz
WZA3qXvCQXMZI/pVny0TU0J5vKXZd7h3OrHsoIiyq/FJ2e3Px0hVptlRw1dwhjdQ
YO9/KWOt8jo0aLnxZKK+8SRTzI51MFeHaD5M+ZshcIuX2h8gzZPSiMZo5YCHXlv9
6FUzllLWjjA3VkZ66OPFbaXlXrPNDUKgtn+3pNF14j9/08m0fOmcHGB/LFYREw9C
TkpC6nzHDT4uBkfv8zGF/VHbVUB4iinDRK3DiBcxYZ5/XlUCUXh0W8Kulflvwc/3
8ka8qGmO1UqK+V6mbAIZsAu5FMBPDKYZApuyl4IbhslNZ5vP564SbIcliNz8iSoJ
v/kiew0H5f2HJsh2+//zEP8z5LWJLQBMeJ3ski/euFVn4BXbUNlxwx4ptSyYgAQx
h5ck+5n5p/2K9Ml91nsRzt5XVoZHZjHA+Dsvrs74nspgemFOJc1RuhzpPfdYkmSH
21LxqQYYQppEQsHEHZBqMC0iaWmWINwW6vPgtK4X4oImS2guNJU82O4bxJBv7FY3
GwaFEwJcPa1O1NlgJ7yFvEYqe2xegj6ki3woYuD4KUg6N0wnXZby1/XKpFPNGzC8
RpNkaDSYHXXLhv01xkDrUyMene8UapUuJQkgk5HXvK6VzaiQ1as1kXEaI4HQg7BF
koyL1rQ/DtQwSL1quROb/fusTlc+036+G26rHv9XK1WHAtO/SbJnCwoyw38hoEDT
4CjrwWgC+5XpDOcIhb/Fc/RkwsozqCkEtK6qVJljk72ImOyBOWGafWb2ldCCKWW5
ho0vuoZ9sDF+wUNtdfvMzPHPN4YBT/gyO66lxCnRr6uQAcgJCQ+C4ngNUoi1BnXo
bOdv9GRlOaCrPe0EUIQyVXZT/T2MSzLbzFg+LrBZlrrfAdGCEIOvxdl4xlcJpu+f
ZlYSAFT6IgIrOQgmrhcRk6+z6ztlKoYeQGPPJYxow8uMnPnaaCGeT+m0u8RO5AO8
0VPOAAiRmDMViL5IOothDUPkYkucNQpP6JE38utUxdjtwCft6mPlxcZ+omBLQu4d
nFeZMjHxkuAkDBg6IR5PUK/tFC+6Q3SQ6KV9AoK0Blanv07vji8Vew5APOoM/xg7
PTwOG80Kt9upBZ4oBLhErx81WM84c6f0nVifmPsJ+CQ138gplPHuuaUhJ02P9U+Y
V4thyIZ6A8R8hmmGBE+bLKU9PANMELL2a5fFzLg5z6LmDUA8zbejg1USfuZjV2PY
c2Wc8z4GXUub/IOK5gBzNL9dQyb5K250x8hfLHGSdnTM9Gqsw4dOUog8QOO7Ncvt
s2ZTdLFJfinDAQW9I6sqWG4MOJ5zBMBI4BOuWuGaBYSTzOrTdf4GTX9h0nBYoAfg
Wx6swAm6VGEmHik3vFypkqS5q6HMyk9fNrn4aph051XWkAZl10xX+UW7MX6UJ35j
oLTomO8hhfUVC5d84dnYtNeWZ70laaDeH9BLiUIPzUCspWhr7xTqx95Ouj+ako0L
bHAf5LWLe5q/SZyvAeIHLcaOLmOm+fOwPk0IF7UF+UlXNjxp5QpEQkmDYZRQThR0
goMMvsTkdJ76BlTOGTSeCzPm2T8EaR4U0er5WdP9U5E+7Dj6GHUNpJ9h8blD3jl6
bGR7apwtPKr7EuSOkMWej3B6RJ2mryMh8MpzpZG3ivMRFtRKFuwN1NB5bSN/XyHM
R97w08ZMpX/dFgyJ6IN6Kd8k4+/znETYsiCpcyRBC4KlTAZXmlsweeHsY6l5O3Nm
eMwHNZASL2KBmt47ylMjBpZWJrs1rMyTWmhmlxaSMO6MUB78BVBz0l6L6JLktWu7
V6/HoTYDcmnOFaQL0tQNhfNJdJNA0KSvPI8sHmBoBKyQsNHC9V57OohDEpS9FsEs
+hFtzGp7LnXzJw3Ez5WzBqBOQhEIi4V9JJe7gJ7exZqLuTYu6mYSfkejnKcMxO9S
M1i+ajE3akBjk9Yt5cc+9UpR4T5839+5YKbhqbBqazP4rmHg2/OCuTs8vh3e3THj
fCUfImYkR+rHRUDPcftuKMkJfxsLrmLmK8ho2K4S51QP7XxQzWp2UEgyAwTl7gBE
aEV/rFjPejC7Em3lEB1pxnumbM7SYV9w9v5KxKWWey7dsWfvPQjBPF8f9/Kph8bu
g/gQqajmJXZtsnuKZiFDPe7l6vWq1PHIdvjlHlcVUUlU+HrK0YVvBxi26MzHYZnt
sSLxMVMBpMfqV16E2ib80kKh8/j/Tg8DmEi4jfql9Vz8ydhaEQKh7gWyVuwsohCI
l+sYoSg7rCX6bsg217eVsmb1cA1d9APLSVxo1o9icRQVxcrlaqRcZ8w3r/RaSUgw
hnyLJEiyuDgDifPmXDxGRuO9l3VU0w+r4udrw5WXCHZ+HtwsBo10mZiWPP/xWwdG
AvtBqpNQCG/LNzNLOVwVALJsFqmiJ5h9x+pKbyODc7sxwXHYlbkxxcymr2iSPDYb
9mtkDz2a80zW449jedwGyvkA1d8dx0uTqZ1G5rlzasjWdirC8Cb2mBtTkbh/iE/Z
gTBA35FC8j61QK5m4udtLUooYvk02g1HzQ7v6vFCB5fMhe2T2VJwPABhOVvGoXR8
Vp6oFywVERlcx6FKfq1e7hoqtBJXDVtu/fGX7UZoSIUi13xzH4z5P7ph4Jz6LuiI
13Q8PRg10IhNjv24+WEUVQfUuYx018YS777fQa9bz3KiYAfSWNg+rTvrIOdrtJwf
6TqNsKs1gR/EBVgOswSqfkYLuqzzaRhVOIknGPTWiEwk1aw8ORhqX0K9SnOEv8H1
HXMwm2p8BwgYwHgS6QgzYnVlFA3wpQ7un47k/BUngUeVvZhariYUeX59hdyE2vkr
XRzCGfn8cdI4wT2uRvqLmUiqXwMBGQwYUMT4f9q0wd4y4yvQaL2JnlBTro/9pBx9
wvjZ7Uq+J6tOnWKo6HPPMKmA57tiQOkejX5LOf19okpDaPAxJmWXM/dsbeznI9JL
Q/P8k2Gf0A2rJLwO//xSyaG7JYb9PK2ky/Rt/S9VIoL7scICJWp2+jzu/EJ3xaJU
ni/LyxgBdjYMtD+lp6hS3wu5TJz3pOOm0a7ObtfTGAQ5kQUz5heF5H3+2vVzuAOS
wMAglUJhjscIk//O69sW+CiWT52WDwLqbppZKdiO1ta8+v4kdoA2bDk2rPFX3lia
5x2MniEciyhLvPK52BvnvJsQvJVM+LU7XzcUKbZV0bggmW6L3WSgJwYFxcJvZe6E
8URn68ypbHrgNlcoj9KDO/D/Gf/ONctveYPVBRpGuQRFz5IVLT0hlKhfFVw0U1ue
quqUEuS7QWzDN0uoId+pbZHkAWy+ynp3sgjljMWO6gTZLpzImz7B2GMWSlwcbjnE
wmtjWneEZ2N2K134S0H5gV3rZk5Ly/nvuvBPKjynjb3c+hmCLjmpZUIyLJ5wpN+m
k+VCOBKx4rZNuH43bbKQjpqa/KvKk/mXTyIfzgTnDcq4YX8J3WAQJPY90mzh6t9I
qqvZBk+35prkvCE/lcxOpQQ9UwKekjyZeip6zwGsUp+S82o91GzBCPU6V5aZVZI0
Fpf0OOYEc+r29VP86Z7V5roax/qGjWAQ0F4/Rf/6alYEVWERafpQKaZSCKARjQ4W
ct76YTS74pgsYr+2uCqF1GYjKkYt1TZfFFQnZE+iJ/l3RzLS7wRY+kwbFYE9DIjy
AD0jy+NDcmPUqHW/wCcpygfk8PKsX94qlOcT87ydFZXXFq70CI8L60tR4aIjLyDk
+BjaRipUrsH8C3vwEnjeh3g21VyOw3lZPwF/4VBrjrkaWAFKjXszUHd4bEJij7sA
Vq/hceZ292s6r4KAGsZFMwp4Xup9LQrsCGv9xyVeztRQVY2OxS/ARV7jq7efyMCv
sbZbeOCMZGCW6MLdXiqh3sNytqxopvHrxZaXEhbS7GPrma6yTgFgsX17pxRxIkRO
fiSUvk7WjAbB3clvFewCxh6k9gjklDgl7f2F82I0SDDh0ULGRSmRGKRHEKOHBLPy
7UcNvHAH8vozBazVcKKkKR2tlIjA3U2e8oxaBHqLbr80Ylo0l3KD4tl0CKQedqxm
5rDNOu1ATueDCVaufTU5iZ8zDhpavVCk7ya2IIPU1dkP4tHm0PMqJoQff4m7ivV4
v+P+e/j2v/v6h5Omu7+JbSZDuYqh06GHAJ6/6zZwmhWMFDIaQYF1qM541i+AgoyY
VkGTjYbxgdFKmPpYT9AwofNLLy08j6SIJWLTDUcYsGMeiNVQzCQF7VR0gPjGtveb
JcpgI7ND7xEVELyHVJ7+QCpXx7bi963akK7rRlLZ3+Zq6L223OZRJmjEL+QJOUHk
JBsUXU9UR6vpzVMzgQPaM7PmK4lyklALNsQA52igQx/Cp0awz+1oTBoRK02G42fT
TQY2s22ZIWH8iwWmSyz5YCjWdhWVupg4jB2CGBGIgboQGf2FHFriUo34/pHt6npe
V9Q7URfSDBaCfISgb+pBcJDYxXRN+yt/zspNTSKQeCJqbI7Gr2g0+FC45SD34/b+
wwvnDS96AxhhPohSPGMQ9M0PX6XblVhnCtoYtqDY0RCVGj1XDGUkkj0/6np4UUsW
3R30ayTDLwXS+Ooo/u2dVune4WAcbXTmvFcOZcyYXtVBYBgsVp4YIPnIwq/5uNOz
7c8ubUCR1aRu2PQxmZevILzNYOCDdmdMGnqd+uv8evyZVxAUClQuZyFK6R9HZ/9a
DFWLDPEDjs/blztPfL0k5BkjgnWznJBx6+eeRcr72plxho4MBrgm6/cVEK2IH/yh
H1A2ag5flymoIaGzfytYcwxuhBcYSp3EAH0DoBaOC9lNKmzp98pGwnSNn6jgx40a
oICAv6XLaaGyaP/RGtMmSwGC4rJOMIMYVQquTuxUY2Of4iva6jUkCn8y0XLuAw93
vvdh3Eb1wMy2tFeKyMtxN4MyRZUzPhKSq24Dh5TMBDnaz1aFka1KNq1wJqcAGibc
f41znYncLf+5AMPu9t0rw42Kal2FgF0xc3cIR8bD5vNk4Z2jeZ9vpldJUG4LmOR/
D3NT1frtU73hVT//b4+BXb4qKABD665LWyDV0kr9TZs5G7xwM9ncMx5nWnPTh6ef
XWhWfTvxaem32xxKF7MHNCWI9h8CAIGFGKCm+jWUQflF9e6r1eiB7p9lW/LpDVba
K5ZFiJa7kxtgWgnY19ZwOTr8EHl74NOZ9k44C6+ToIqIUQLSb2O5AMS4srOU2pMX
+0TJPHlEeS8Su/TBvyY0GwKooHlwvCr1TTJZ1iF4nukW89xCYtmoVTOeqs9acfoU
jRIWjVWzc0WFFKUwDHtBLo9iBanRnUNXomvW+SvNZJ1CfHsNRIIlvfm2f+C9yiJ6
7jAjKoEuHzvwm0rQVfLI80dwBu/ovZMm2uDq64q016gMRXP6c/2pHkDijuLQFzSw
phHo3GhgOm81EyQg/NAgO1KNCLJWXDrxjenDHcQw4tpSYMmClZgIUH8rpGvtnrhY
PPWoxOTcsBIwFY34Ee4XIHsEW64TGUFS6uzfP5s9BBHdZG0bayKB7ZTGJDYNvA1i
tqx965wtQvFGAB5g91zXGJm/coYgnl3/7FGX5mnas4a2xA8kfuJSO7BkwzyGez2j
meFABrX4xpyG4y88nWUpSin1MO22WGBpJQdo/VYKNVHa1NFYgXAY3gVHtSOknbVx
lrzsqRQ1ya2qBN4e/GmIuIheGWw0ASDuyqYnNHEh1Nk8/nNDaZCDm4e/efGdkWS9
qLYR6VGsuFmoYmsS039aJPPGfJw/p1uKMNpRIvnjUuH6wn+mTLO6TmkvTDdHIA7D
Nl25DvgkvHLXAjfDLHZBcrimN6HuN1wKoyycC65C1RHvj1tfRw9UB/6OOi1hTLWa
hfoNy9OKTymzy8hiVs8nQ9Gl2Cb9/eNIdWzgzwJ4mGOZTLrDPFbWl/lW6vyxVKhC
7D88NOR52TY8Ht/qWGwCzJIsS1iIeT0IE9o+C8egmxxwrUydTyq9evwK/WhdKzWt
u7DxCTBe9dwa9YUse/rwK12ME/FPfnnTeNQPMlqnWgPwxF03yb0fdcgA6gxdqSB5
7EvRk40OKDspQ/Fy+6wd40c3o2RX5ab0IM4CfI0kBwbSXz7waQ3afDRvoPfAMs9n
/9CqON7qpYASVV6Ep8Sq2Qw0ovIGvrtjOMJmSmkC9+Sb/qUauHiFDvvRgbvGxkUq
pH7HOLtgzSNEHUuUOyHojcj+DWBSsBOXF+sx8ILmZ446YfDDvhdoJiB4ktPaXvVz
5U16lk/9afzG56NYkhA3c4D+EQWyBa2UXw06CoOu7cmbvkubBEBW4hF91P6r5/6d
rFS6MCvvNJAUYsqufkH0fFzexoVrq7Zhk6W7osdknd1ysFa9/jPn8pvXxaBhHOeh
epRTxttpvcEH4Y+b2zwdrDEWkmQfqvD6ffgDCWbUo1dBNBBIwVUogPs3y17BAb0c
eLwmMh37n2F+muuGNyRhLGNUGdhFmJhBsRW7EnHk98r/+HEdaICnFyK9AUCNS/N+
py/QcYksg4OqHMIaMrQfR+ZkJSC5onCBTVjXsLGwKcLC1JHSmuM/brUKO+Upl/Hu
ezSkh4ulCJBf77Brhp0IovbTuZQ4zXhpY0RC5o6RtbAikTLhqyNSohnb9kM8Vx6Z
zk+QQbFZ5yVhS1tLtL6DDizy4jtEWcFHBZPtnc/6C053dKbLQaJHDrxyt/KWLLRg
bbOud/raFy0gcK5Fo1jKuylDsSVzw2Ho81wHgzK+bBsy4DC2igNaTkbj0BMqBj8l
QVe4gvnbwn0x2DXDzBwG69BCgVzINq5a3ekrmuFTrs1YZdTDHLECnfMkgBBPrKiw
zaid4O6v7YUlIdOjBog4odZG4jZrgGi71ifpeqZSZko+uGmAdJulua5lkJKMOaFL
go9YKrJq0veg8/fAJhuGb6Dff5mvLqwpWRQj/jWstzkHOT/h8GbQ+L7Clp6apJx4
qrL/4xcJbI+9uzgzKg3WqZafKPUP0WCpY0pFzH7WGInMSQ04w7eQUxShgt4jxL5o
LkGJF1woP4HXv1UG75KoVOoqmaMwGIgeRnIbx88eIQI511qUzOx/+ihqGydeuP4Z
q3XKKrciE47D3bqKojfviktwX2z+U6UYTR8cMGfjKo4YEMJnmLa1HqVTVP4uqOw/
vswxfgu9GEFzzBvvMWwqTvDv9Yas69DpPfq4KfxotH1N8HCLeceghzUuItL9phmC
F8RX+dnfDdNrcHLtrKVdNIxlAev6csgsSNy7LKrRFFc6gxFus0sex0wh5mOnA+Uz
yPL9cLLWjFYwQDSFduSCmfoGRrWfl56OqztDv4nVOACGsuSIOFWnWbBCMzE/pcGM
IFp20JxH2NRkRikYPrCsOn2OV7QnSzPlO1S+7yDLkMRBGbdcwCI+LaOXnWbvicNV
RNXWnP0HGZb6/dTtwrsnhsDxKi3IBzxog4KRDsjtbEiPwQVFzaBQNN7eHIEdaUhY
G59CmHZKHV7D5a7UuB8jBG6LciKoicGmhbL/MdA5CwTDU79a/l6eFGKzH/zZ9tm8
5JOoeoEsbeQNplEoahvcHfx1B6oR+TC+JSO1MgHoZ79n7m+HsD0M6vsUHs8iZ3PN
o5WoXPWjG0wlmnKojBE45TeFUm32XsmiEYYosVzyXHcVbKdrFUPL2a30Q2HV1FIg
0dNwdbWQcGf/WxUz8nuhLgdbDQ43P2HDuX0CllrUbYTNIYgjbwVGAFAOzVWFJ0ae
Zz1wRKhbcI4S4qeJJzZ0e9S2MQHJbMQefxatMjHBS2WnYRqRqaKq4y3KosYc4AmU
hsFLXU+JTmC7B+27kCTKwSpPc4U4Hu6A8qZ+bQmly3uyxHthp4kFBStlWM+gGqCW
MIcwJyuLyujyDhaO7g7A/h0E8iIbBPfo3lAetwqNRfzVQiM540FZLNw+2KCBkmMx
V/l8gsTjS5tbf2U5ax+LOxWLOOKH1QcgV1XBA2kaB/RS3O66R7mE6OkUZjhIfg1q
DlExZVFJsYxi30OF+kLPzKMO4FIhZKvrJrGx1qFptn8xRQLeFbUddd5Zc3oMvZqI
ZDYGEzPCivH1h5ihCFMlc0CKYhSniQvnou8mrDPEFc8siA61+gtZlLE9YzroiOnl
/EBB464TA/kmJFOq/iWOlwPPTA5HPNMzTw0OUyrRY4s3l7h3um9P/1omWzNP7fHB
0hbx8oMSHG0WEuIyQ9UHNf3/0ihoC4gl8pxE7c2RaOKKXEjhBSjW9Zut1LuD0ZzZ
b0pCI4QSpk/hSSr2nAGWXilr/ZGUfqXLCreBBRP/rNzmcjwvfc5LvR6wNptsuZfl
J7D2rGXffUWGdNdfJbzUA/SEnnorCbX5DQWSzdn1bvnKwxfO650K19CV6jpEoK9F
awWSBw7P84KAU2USsAJvHuZpq1Y8rV78Ayva3m2gklygmqbw2f6PS3E6kaikWCGO
sg7vfB5d62f4pxKrWmcrMfzD+4QqeW6V9hPzB2AVbMA2swZHBCzhJJvAFBS1drTm
+hrWwQ3gSF0fDXm1QFM2W1bbEPgvlpjX20CAD5JUghGq9ya0hCtlZSOXEsUoAGLv
VdWIFg3DiKD1dFzTfchBGd38qGIp+U3Ih7SVUWKKD+8mWA27lDCdqYUgPE0y5Mv4
csK2BCm61Oa7RoD9MQ5GiQPPZyBUYOXLHkCJpYlNtpy69yupasIlGEvjPy0jRYQb
ASlzlaSaVi3adPN2Z/eXho7cNTURe6hpKyeZu8N5OlNwbbD3ZwcQQDY/lQ58umeo
lDeBUOXNX1I1o01TyWv7Gb8IqVnDTJAaK8VX86zXgNSmiAIZXqtI4L79QRrou6aU
K3oKhowAWVdEuGNhWoarABMU4xIuSQdnPlOzgcMvsBa7V0huJer0WlsrL87if9mZ
V4EQGY2GY3QZN/qZEsQG/pWVM+kIm3wsJlQMbF+pbizTtZ5pX3uv7dIlzwoYjiH/
Yu8kqwuyxNoEvIkILv/IPHsKpeTuMmctiPwev3QhWWxmFJRjJJN5cGfW1Ww+JBdw
9lfZXRrY/JelqE/NdezZRMm19uFGF67uMAcdhDYj2K9Nm9p64fgV4fcm1mpEev9Z
WiAyGAgZnI94PegPcMYnUfZ4TV9PS1NTVsyXGfcTfR8tbrPWZlrYzaSPUyiHEA3q
Cd0uLCsZUYe+hkFbVlor2QjC3F6qNMKuDTYV1GicVOVahGFcbc8t0PUDDFT8h3fA
7vcZuziu/gDh3b64bNZY+JzPusgX2oaLBE/RSztopcDVZfjOK6oHqWQy2iVLzip9
K6J+Zu/qdWp13XtlHkTgL3iIxCVjFtMSYyq7uPhpvQhWOK3n33DJvIgBt9j50F9O
Ha4b4DMEcO6oFyQktoLkUJ7BmIovQae9tC8ZlkPpJ2NUU7wnsRQbbzwEdGm0JQSJ
juYWjUkIxvjwt33M540BKi2ECKfQpqcAgqcZa8WCPjUmySeJAhsZ5mtddbCkkyAS
y2Uw2itJ2F8ms/G1M1Trd099HiQu8yzix3qjSW6MzBlBIgK51TpHkBXkZOr87RUI
8i/7vAdUk7lIgCscVjf+/fVMK+G6DMsruvw4Brui7CR3ICNXLiEHooth0DauU8ZW
xXOD/tQbPMJiAkQOoF+gtYkYjDPVS7sWsKBbOdCOq26D6NZXM78npmSv+HVaAqHE
/c83ubG9YN327H3+T79XKkJO387jVFZAfi14oa4rnVx4xGgtqgEaZLcOxKr+/vUG
K/5fCij6mzfvjeLnz3kYF+8vpSpKSjwzDHUTsKWdMUpt95TYBkTlsLHYQWSt1AdP
fb2hnqmTJRhpAtD6CJH3ApcKj3vydPQr3fZ1xzFkqdADeiVvPZh+kdJ11L98bBPM
Z2atyDWlTAcOlAXCUQ7NfPLtUEYHTSXLRUu09cZI5Q7TtTqADlPv3qAfAKZSsJHg
yg34HJA7o7HaaR+pb1s6aDR6zZPubZob/Ad4RILN5iYa9jYSLtv64yljoGirmLGW
jll6Iovx/ZnZqg11XjM897T57winLHWoZfF7leveRo4gCuxryCufFm7dy7MmM6KM
TnCjkTziKukOf/OQjAP2r7EdVfcUW3+Fv3nH1lFnlg+J7WzF2TdFrmDeY7k3pesT
xIZrShT9x1YiB7KZcXyf5EhLZu9qTnRRchE3PagLPDMCoA4Z/UFGhUgEzDvjWsSE
Kxvw212Xy/DvE7kdC7cEDelrNwAhD2icDeOZt8ZoYfTqEErxGZA2oFUaXhObXso3
XWJHXXk3jvwc64saSSdc8h76ZrQ2+dCRihr2kICx2ytaecqoRlC0Rit0QJ64N4gn
yhTot4FKlS9AIz99l6GELchUQueVKcM2iOdzBlRmuBYEDPLZ1uspPLmorwefZIV5
5kqBHMlyFr8CTyoi5TF1zACRbh7s2oT1Ob4410+rIJ0SSARg1c++URpGSaMUBZ+i
WibwCE114YSAmIuhSMvUg5BGtWPN2/o0xac/04YaJ/9zfstkW7d3CLDZXhlm1hmN
a58tZer+koyg4BX7m+zwPOPCjpk8sy/vI4glTl4bTfGErczjDuvGS3N9E76GNpJ7
TymvHAp6nqfLm4IvhNUncPvxi9IKyWwrikx6r/M294xkjJBzR1Wvk96rp9jFTTCU
r7lQtuCvx0UeM5BoTHZzDwKvib6EGoD39vcnVTnzIukPhUt2BsLNVcWCFj9vV4xK
2W7bcBQDPIS8phVzBxKneDQUv2Z9AaJtbxs0HEjP8iMKB8PxvkLB77qrqFl77EqN
eLApywzkZibjj/ml7CtT2ldaOlMx8s2ZMUyCG7G+M2BBW7n3iHHkEqyHDC1NZdG2
k70l4qFQHJS2cc3SKmmDCnbkHmPIyG3LJgp69danCvtDllDreujmJTOftHj/DJgX
57MQmxYEnOVRaXalXxxGK6Cjo0Crx6NLiO+tqOmtQt2jfgs92uD3kcz2rfUQgw5H
1+4FZbvbOhaXKIO8KoKyOtRGw+NkyhLUcEkmVzvXKu5lG2DpWNfq7PKySKGRjG3Y
beY5q9LKBzHcOybTSjjqqw4DSmZc0VP4mG9JelzDOc+NFBEcrNVT/UwJvAWAx8Y1
QcC34XffsHNHUfq2eJs7L2q6FLoT2NZdyjlRhQaNMfgSIwNNQ+GHIl8N94kINbY4
HgP3fImCrKAfc2rENmo70NkVKhMJP9LswymemIR61+FYVxn9mRAw/P5xt69C4R5d
YSYQlWbchhvJCA/2JzT5c4j8rrCCLqBX3auJfwwpQ4I+uxpeBa1ytBcfZJQ+kMrt
t+E3jE7UAtXZvc3Ag5XnO61n4zBnyIR33IedVSoOuWU0m/QTwzZPCClcXNpHerhs
eEUeYteNrFo2DvEP7YVDGC/pzVo90h1DSYfkuxoOoJVWUhvaKx4TDrXuR85wq7OM
PVlmBU/2XJtkVpy5AWXgJYcssHl9Mff6ZTaxBh7CUICxVafm4K1aqbs6gN1ynhv9
r1xDB96T1L4kvD9APLwiSPlkbFMArZCRKrCFFWKbN75s+vUwYr204X6qLR9LYuvc
tBxd+A29y+F7lawbHRJbd3IuTOUwe7F0U4gdgfbw078piDX88AfQICz76TaS1iHj
aCMp5KAZ4p9iQN8oa/E/cQH5jFgYcZWfkA6J2Y0kbhDxVGFiiICe4x5BaVn/1UfG
Jn9Gu2Ej86dFRU47xzH+6RYBVe0JUt0mymcczxBTSE3+V/+/CaCxKJ8d1aI+BTlV
tM86b9yg2orxu9qVZyijcors43ALunNraiVfsCrn0U7mrScu3NUp9VF1BSPoDDyZ
3fYP3rW1FSICSbb5KmLwHSaXYRWNiefc/ndqGVwo1VEKgcICqEzWR09WV2eTuYLB
yqF1FfJaRfiLntwFuYvciQ0Ju1Tl2vp/HfBE5Ik4TzTjngv6t89q4Jjzg3bTr2C8
n2enCh1BzYVpGtohmWdS1cWJVk9lyuM3BQFllmMiFuS4KeSSUuY9jfblnUD/AavU
d0/50bPoExt9gYQtJuwzP0VNreGum8QnUZD6TqIHx8YWYZADEUZLu0Uvhllvh2/9
Viw/vEzwKGm+9u62AwIobc0LPp7N85IN8cUIrWNIRR25MghfbvODC7WgBZY5n1eg
Bo/v6j0oTFWiwOML+wsZLPH6/eSdofDVLYvPs1jmwHf9MbC4BDSS4ILF3cTnhA4t
3DZ1wiu45qc9ntRrOzVJfuRd2tUfmXeddEyjxat0+9nOgrOhv/Yfl7iVgbsXOsAR
9xsya3RC4TO+E5W0Af9awemj2BEVAwvjei6j18IoMEw1Yl0EwYYxreZGs5qhfng2
REaNTKgqb/l0vaJJkhzS9uAKE19Q7p5/mwc+XCkerVjgmPFpuuzw/tEC4Qx8iOKj
r57G1dYOejhXCnmI7DUUSoY0U+zqL00IT9diXNpyxpXc2ImR4Ni/zPfza4IHWN4Q
Dl2vTdc1nJR0oPN57xD79XJlVBlKMXnQx746mMBgulgRyXJZ+6S05nm3RhG3LPs9
WSo5Gui8xxD7J5cstH8+ajhwwzVjF5uqwuZM78NqLT4jqbmonNl8MLpz2o8XPUwi
ZNqnKazVyYG016CPSESyRczLaXLjh+RPBiUUWJcI510XopE/l58svBPwt62n+1ti
MSIABuqnrcmOGMxCVh+uEDxVW1kFyt9w+sEodnesL+OSdnMn5Sf4Q6jozL51kXap
l7aPFqJmU8p+iVwi9szYX+KCitN7WOwm1WNdVn6M26yuT4kyaTLnFYoAzPaACns5
GCtHWSlu3nHvDet44R3CFi1q3rj6JccbrHhPUlfjXvufKcmJ1PgMdJEBRyuKZ4fT
PEoh/F7Nk67ZfGZ1O2/zTRGXgx3oHWs7m/kPcJNCpaD46JRdFkv5MJ11uVmkojWv
n3SoIrww0wlqY/hs63Q/X93K+/J6gAwszvXcedWwUEAk4IInPNSPX7bkavlZ5AS0
51lLr6ZuE8HXJOlvpx6PlHM85AkrX7ii/3UVI/+LjAusFTUAjVHtkEialtozNzje
Jtrcp0dnOtmNK3rij9BwLhUXQIwfrXsWOZ88vMlgkbxnzjJ6FXGUM6lXdGVwu3KI
1dlnUPp9Ld32X/CIUrT3xUn14292JLX+546NajhraUo0riZHiHbA6cRN+vuknJ/W
VANrXuy4ivYul2X9WRdauQZd4VZuXTAm9QdNCM9DuH7n4GYzl59EiaY2G9nRvQSt
aiYw3wx8iMoIC8pttWoTQ9IChQhVTk22fHQUFSuvEQkSAZi+EXMLAAVUa50hOyjR
vJoYglf/9KGAunzke2WMwUPE890iRJBBhqE8p/a/7ZhJn0gYbsZd8vLzqCcAUm49
VGwP+SdP18vTjK2PevfLNZd/7I5vfwDSzpM6ijvJSAbKCeOVQ1NN0K/Hax4aTC7D
wEnJnOYk/R1SH1U5cJQOFKrNWeWkeNjlK7z+1o1brajs8VrdbIcywVvRLnxG1nc3
SothT9YtXFWHlRsggOc2vSz+fgz5Z7Dmr4laUWXmBGJyiSR+vDhM609yGi3L68Dh
X7kjHxVK3DxmQMFe/Knb43Pkrg43CO25aHmpqBCMOFs0zHu8yq92fIzfoKCdSkP1
NZhTJnzy3x9dF/Gx0V7HaCCjS1q03t7a4kTQClPB/JVGa+5v6rmYtHhkFEmiWFM/
TPHTHyWfWfCobhdRQz9ByOPbPFGlYaUKpOXPQBXzi/aPtsWwWtq9TrmvGfaCDfpv
OTVICyc3tPP1/vWwGAgZ0bgRHD9Yc9GvmzvyydQ6uNLcqyzP/1wyJxEMMwlWyHl6
LV3PrOYN3VPZn65k12Twv659F+GIW1v/mBdtD9ooH78AaB98CMz08b4PFFh5eTTx
gPicZp2xV5tKl2v4n1qmFll6zJW7Q7yw6kmog7IbJUPQRfNyM/MwmGKNwNxZ9rzz
iZ7+GSt9z8hoE9ujuoGrmN/KIOWb97eGe/uFpO5OT6d2nIgPdNiF8Nm+yzHZI9pJ
Z/jkEkzFXR2f4bANeBM26wG9NEc1fVRlO8Zuu3qk/bvSBBFn4i7r47Fk42MtRBmY
Q4FxF0yK2chIasOYw/a+W5FBhNl3kzH0BlkIM+4N1eO5XwH8LRzJxoJEcvgiCf5E
o0JSm9FEni+oUBmoPn8US9OCkM9onQmV0VnER3On/uWoRzzBfFzp4GE8BkR1+bOH
nDLqqCPC8djQNIGziMm9GzHBjeGansqnXk+HSLdDGe3IHtgvRuthxAnEGJuIhVjT
/yGPaMJeLA2UHUN/BXsBKV0Dsq9ZecO627NZn47kG8KPvqzBQmsKaqdNMP5hXhG8
P5mqcu4IiBAUFIqlNPKSjgWzen+mrSYzC8FnAhCTX6cR8sXnbFw9AEBrIQ7aEI1J
zIbSTZjZkb/p9XcllA4djqZm8EszGVKwR7dglvsezGBIjafddhKEcNfrtZvV6VMj
slcVsHn5DUH9rweAucBjNJbSQdf2+4aDr7CjPuj+EgIAjIN+iSX6dpEW2QntoVZI
qC5tsTSvfa/nTWVc37qyWAlgVb7jdeLKRxeKfSGCInQG39P0/mLzAY9UG95LfAzW
evCivbLEm2AD3hekbw1Kj/FSfAjbOG1uBhmiSJ7yusdyXnVfjf1uNUxfdyo6DId/
UguVeEc43EOIIal4qA+VposKdhMIHkXUIRXk93IYAPYZaYakIPMH8sWKzDaaBlV2
f3hyNWYUw0nyDk5wE0xSMbNwPG6dk6Pq/qWVptmWNWLuQQu4vsu6+v9y86BIeHkF
u+nna1HX+Nf1KSC+65l8Baq5oN1NEex0c/7rwIhu73Vo0XZq3ruPnUuQUptI/Ljt
P2JcuaaCwnMcqUYzDJ59wH1BmJQEyPZZJj8XK5tmzX3RC/A9BbgUowCLEwl1ad5Y
6eCjMLiGjQwrV0iQ6q5GvRR6BSl6xNFOb6Oi+DheMIVCwU38GE+SV1NfxtDEmsiL
XnEsK6pzY6DEZiuMFA24nqmV6fBjPWNjwuERa/lhaBzi9mqULK6xuy54Pd5K8//0
oAnegrjqnrbPytADwV2uws5aU4NH5fnrg5NpBxsWHOPSii11PuNdemWzj/bseeSM
m8z3fNrEh8otcHulJMVvZTIe33u840fY9pdweHZpxL3hs+k3wGGcTsxYVemoe/7W
rUSovIgbNv6ai6axW3CU/e6qd8Ynwy7DaArVucnj/LPfZ5XFSepNb3WOdTxDitN+
1Et7naIm5Op/eC9Sh+rdDIZzHGtl+AZ6TWtZnHp+WMqTD+cnDDJWUCG8rfHkVl7d
cRj/Zimgiudiy+4/QjSPDxEs3sBrJU0TOcVPZZYeL51fFTtK/swnqFE0JgkBMB1j
a8gUnTVyk+xURz+NdbZSL7Ilkuf16nGTMxoDxef+nvHppM9HO/A7DAU5aAlELMNL
+HjJ9vO8xI3ZoN/kviaK8w2nnfr9fGS1yZRac5EBIKzjVlygPSLepECoUPB1B7/O
MuizTFei+W3xIvacQMfSDSemXs5ujAMrpaiX2YtM9+dpQhPoPEG5hvK22y9aOBxZ
oeKa+jBzu/B1OWqYD1UxoYF0b5r9r/bwqAuPJBjeA+jqpWtCvf5bA8IKcJsZH34O
4nvTguRgby/1d3tVl7byZcXVw5vANemKErlzYfN2/BfbIUqKquj4pil7lTZdgVm6
PovfzV2P93F5/DccV3J1vtMEWtO8HgH0RbTEXv4UR8EOBzYaXj583r1m6TU8rW41
MKcC0bFVPU/qBa5eMLPzXBjlQBlyLt0dHSUMZCBTq+fT7DsDVQY+Q4C0ebnNXV1Q
ql+vsi82BGUrOsLPGWnnfMdHovUwX2CkScQmb7Cb8ojtpnHrFoxqq1OP1jfKtFFo
W7ddBgdcmuvlaxFJqb2bhVqJOd2ggSiy9ARtJjTD3wHXrL9nRU6cKxdL/0jQxNhI
9Vdr7QMmw88Fnc5eemRiWPh+JDJct2Nn95egxU+gqxlUPwJlfCUvHYlnrhVh9/N7
o7Ydoa2CubM77Pqa6R6CSXZMWzJZSQd4P4f0HxxM8pWCsL6yIgRRJfp9A//ZfTAE
TE4rzy5ICIqrswnmwslWuZpRuaW5a1qNR8TFMFT4+EZbGjfmDh0XNFP5mYflAp/r
9zzBgnr9Av9Sv3ormSVyMTVs2hOZwffzevK8YYNCTqwFFHZqn7Yts1CXCb5j7O/N
ruwhH7y1hi2TjTcIfipeXOqdHO+zSAQAqTfaVbTEnw9e7GO4XbOtvoqG6c7fIS55
vccpyI/qjtcX70XUaE7odG1e4jVyb26GrZadOQ+11Xj81P66VnQRWFOf0471FKxR
Bb04AOfnc5D+L/r8TlYmCTD2Bj/ZwAhnenizuBJZzf9Nb6trlA6xif1CJY1VNVGN
BohVKa5yghuZ6Ai3GV1p2XaX+z7hA0RojFJFUAbWgyhWKUm2r367S5dDlXrUgyLw
euCBgYBqf+vDOzVZnaOPRA5MbuOVGUZrQ2Vi6x0pCtBxLjkTfbOtMuDnBCODBYmb
43FwqHLg5RmM/miWjck6lCFg0TGyW1EPSgo0BDGiu9bdCZ4Xv6vs3zoQJrEgW6PY
eg0Otw79vh+Xn9Kf65BjE/vO1wXNJ8bE358TQPqmINWyRiNZ/f1rmHHcqOcLU1bN
WxQ4G7rHxye3h/GUxvWFlW982KT4FIFF8cjFraVG4/MqWxB3IUKeTFQ8C391tEyW
tz4NZZjEiGS5f8QDldp9z8OR/wyNZ6yOHetcsWlPMBltDT1Q54nPzaRffAVqwbiH
JJg2Dzmyl77R11iZAKNxfnh63cad30Y/KA7nVspOunONWhY0c/7zcoowW1A6o9sw
AFvVYlMX+xLpNB0ulQ3N7jqvui2gL0MP+lJw7WuLeFsL7M879Jd0TcWd92T+7wIr
dRIJ/a2XLodqye5+3ukafDs08s3qApmdykbDkPGstJz5obTWMosrX7NI10royhsh
IMTQgx7Z2JtHP8Pt9I02Gq6umFt9qnOsvDDGoStXeaeqzeu0ZzJCHUe+svDU10nL
ilzthfZfBiPOSYrsrUpAGWUY8jZf+3kBINlykDxAn1bYirQWSVWrE41sLtA7u3mM
Roiq6AcxAggkfKbdzeK8zJNTOiF+Os79yyJ6cUTD5v0FU/JvD/tf251mNo+leCJG
0UF2ZKE6hWY1cwkZoFlKcvxbpTGJniZ9hLHN6L2VhV/hBi9EgdFh4u2ksLoY7UwA
cL0krZtSE+/spuxIJjcIAfWxkJuP2ASM/qPW/hozMQxooYj9Dm7JQHxAC5lTpELq
Y4qLC/cyU9Tlm1HxqBP17BVYbhKiUCOsflp7zfRusI64/fcg2qRmnjlmLqq/s6aw
qZBo+NSTuPu455Cg3XraQJc7SG1cuZbREZNo7q3kkl1KE8EJTFsaaE5rgnuh8ABJ
2/hcUi0qsuZjNVEY5M7pHBaje7YjXqFtt/B/eX81HA52SAdSaqw14UFNCK5JR/52
vaHr7vCAympPXMRw5oupB08yeAuDAR140X7tc2G1WhxwY0ZRrKeKkBUGaitc6vFK
d/Ulqlg3AKJRe5P/h33E0+PlITMSWmOva9hcXLNHIZqt8ig2cGcs9xdtT6B0sgNP
4TCHiSpBCeS52N3Jvd1XCPRnONleSzL54oob5FuxSAWrsFHXfrg4X5eLW9Y21YDF
7pXeQXPfaRsVDPhLi7kLdAkRW3zVKhQ/og/np6YvLZcZWFLRwigBP/J/62VV5MgS
81xL/TW/MXtyDv6OkR+6qu1gDGyJBxExK38Z1DnbK3ytn6SvAn2KbG8x1m1smMDk
7hNzHEGTuYX1wpCYBcW21DAUNA9IucIhi8rVDkpKYNqDsmbaLviIvYMq3PcgTaMC
0RTqoQk8fjU/onH08uasdDuDhOQgj0JEqv5vq3IJnL42cnizEbQLg0/3xBj8fEo9
eLgJmhu2StJ1VrUZgkb0p72X7wfh5u+G5RJL6vo1RiU5wcJJj9azPodK0RquWE7y
twXOfRwW5BH1y4rN9ofmZTcorjnuJ5qMx3Ksw/PPe0SiL7UgvcOxMVnEmfGDaGhV
u3GuiAW3LL1nw2Gb592s/s/GXbcTcWzp+MBoiaqy8BKZeFRB6x6742jesIEHfmBU
brAhfkA6VpWsJRbvgXVBchcarNgrppbITQSPiDO2pCAo3fqG6BuKJ31mvT/TTfGd
qpDUKz5vDqdz9+9AmftMAR2kh+QylHwe5PGwTIhx50Q5Fycqy9UX+9EDPgDtDCB5
8/eAKCplOdDTp5J/diFej5eMM41jChtEl3wLSWlY7w3Z2sWKLzY54I2/0jj/2B2a
TIJ7wQqLzui/JpCYh+F3tvv9hQQJ2H7Fuxbb2v0G9b3mOPE8456FIRCMeOiPq/uB
fKPY+q+MZU79PoEW9+0cRySPkZbr9SvBufLalhtQxL6TBmKbYxBuklL/yL5TPSPg
Oqg7rwkYd8wSCes36YAwml3wwNKGHy+B3H7MaazH1YAvMt9zbX7sWxGVVbBIjf43
GC4qahrl+d2W0srd2VCYSBcrcS+otsuoxDzxFEeh5oH0BUVXHuAKEz5IKN/8GRCq
wwhfDDLCiqSAxyQ9dGI3VRrJGGm1Mxns7A7Uf2yOgc2aDKBGOLd235Se/xCYFd2V
USRqwV4OTpIXVtx34xPm/1PX/blMROAN2S3/ZOUwUp5z4Plrv3PCUs5OrDIP0pzw
DgPyUBP7KrRc3PaIFw3/xcg6/hteFlku3ap8XqTlhLcyEmA37DCzPEmDdXXlm/aX
5dX/IIqeE/+cLgtYk9q+3ZYKZ5oM/LGpy2KgxmiGFPwfzSXRc8xN+b77JC6P5WL7
zLH33vP7emURGdSDnSACWsjojzq4FFc41UkBh91UmJuScicHWGCLshnZjbU0OTSD
SlDxvMdf4ksx6obIQgBc3aRRL66Ep7EZa1413NtAKRpLHjrVROPNTLO2wR1s0h0e
TdggpErdaiaP1oaurC+Lw1BoGV5DddQMBt7Z1VS9BrvnqRmuwEn7VUD0Kd78U7oq
mM+vyE4uLub55FonseXG3Vs+PPbb+vfXxDUXyVvNZNIz+LjTlAqiKpXl0OL3hwIP
rkK36/QjT6rzA74TSvxQIh5bso6K61g3m3b1SH7TUpnAoSQ1pKPz3u7lozxTn9yH
QAOCvwqFArR9P98HeyG6g+/eghDb+Bw4gfuYcPz1/o798D70+WXfBHJrRktwdn41
/ZCibXrpvkpUC3Y6C6lMjCzM5u4k8FGf38NoxkWNcVBbCr8Z7lkes15AjL0s15kC
w/sEbsGEt8eZZs6DdPyFT7l19+HlEH6gPHhqSmdfzXgvA+GJP3YP+y7Wn1gIW7La
T+ukm6h1OdDOJTJG81e7gzcQySO8aIhUGPWuWuSAsnPl/gOAgqaXso11sfj7LmqK
g8dDshVv5sOs+9e9CsSwKWuk2yqLOtipRL45c52zG8X7/f02AJv0cRuVTYJ9zKtq
1qeuYVYmLsOSSGe/7utbsJqDcYtV0aiEbtYZ5dUGP3V6WtpV99ylfuuCOzVxR4IC
72SsVq4bm+y7bSSxWH664g6sUSgNYxYqgjJBc467uTVdogp4u6nZY/95lWfDyth1
7ft+lmAZZUwgXC3QXjDEUrTwgjS226Vp8F5h1LDzLVBKRCi1nMP27tEo51TsgXIh
wqe+zsbI/JCSSzPhFZZimilVaEDe33rXIRjr3HPt4/vlxrbQjGKKElZ3KBi4MPIk
uUPYJBwc6eHkHcFRxyLri78UFxLKqNFeDUiDmM35+UXmWO6eDI/GWeorwvs+hQc8
Z+0pS87I3eeBz7le1fsEXZ/JB6AK46cZIOuOGl3Q17UiCOpU5XepN3X61QEJ+x5P
eJ0HxbAKLjKV+Nt4opAe7F9TRemWnwiSXG57BI2oNLB729XRXx+SRWd4rghyjwoE
TicVzGDXTjwh/OFfOJxicsLWqOffYF1HcRatJ1hWZycYJkCplKzRHtec1j4uLiON
SnLsgVzvUy5Jvzu96+wogtR+31QIh5htl4rK2/X4Ry/DaLnJLfFKuY63IZdgG9lK
0JrOjPHuzl2+WW1cNipRdg6MahGJXuuJF35GauWuATCVtk1qwcaNsqsL8Kdbfaie
5ESFq49EKbW2QyI8YgB/woCfx+p2ehQmWQdE5bz0O5/SYpF1rg4T6LxBBP2i70IU
1RljBKSkW87h6crENvNqwWp/ej3g6Sec/sMH5XuoJ+cV9FLl08qBcFGCcqE1RrIr
ms7V1CqyP1yLLPKT9XLT7dkEke/EeRPeumvvaqV87bZi0SdK608SwBVIu2Lqf6kL
pINuqBgoe3x5Cc9rBk4h5Gir1iIayCTlP/k/US9zO+3EF5+/sEKSBdZC9MZII/fW
k79AAOTTzlgCswiZCi5Whae/q+/c9+nB5dyqt7bZIqa3wj9PcTcUUeNzC9Ocd9eg
ZR/OOUkOmUTe/o38InvNmKHgQMnrtqv6E9HbJeXRfTp4XNspbTDc4uCSaWsliiDM
HweM/5RY84XrTAW5juskQCNmSXVUdlY2A+Ad7CAbB6Biap/da+XmBMdchvc5NQGb
MevygfqBT03G4K2W+uOfQvpUIMwd7imAxDhR+lO+S/QbVtwe3MjnhCN/xufZCTKf
W6ML9x3Qq96kXDSR5JFbW3OfomN/ZmMCiIzqAt2eT+B/xDxQLelRMCek1dQX9XuW
zxN3Paq74aEp3Zex2ItdMydeK791EAd7OEhRbQFzixDeFEXBZOUDr0h/luLHwUrN
3jbq5hXcKob9xQR4y1AEEZcN4kGCtrQey8NvNXb5jdAlz2Ca2qspoyazpuXQrPSv
Vs6yZDvoIg4+qNvQr8gxUSw2yiljqpe3gNtOeXNu8strfz0QCtP+Y/97CiNNw/LC
ociUoKoNT4KDH1OUdfDwsTk9tqvNELClaoh/AoxiJ4MSrSQMhJXE8jaCrJCoJcmW
ufHF5G1lK6GCXHb3fJhWx9M0kvMs8KL5vz0qN0UnSPmCTWmgisAJGDQHBDNKt8lj
EYTuwkwqMLMME5cIANiR1HbVr6IXuN2gvgyDFuXRr/LwJSdVotQ4D0yS9HsKSwHy
jNFI8D5MXsIW/iFl1h7SnnXS9WP4zbyvMCeTvSk2rDUyZIViukocShrqaR/+fUcl
N4V3+GJqTpyFqaV1M4qFDOZ6OZA0T6WsJG7rjE4CZsaugXVOcuaP1DP8gxXXoo+O
Q07xtYU8ZhOl26OqsfrMkXuRE8B8WgMpeBIAkkd43SQYWk8pIS74OLHgGIDHq+fZ
Ykv6Qe3azeZvbku+Lh2LBwoJsY6vEsv0XORorWuNxI6bHN8dUFNsZ1ujshvoQ7iF
xteJVoUppeXqpNyl7LVEbDzSboNBQo83a25LYP1zG0KO26JYEpz980gyn2M/ArG5
NIuzdzquFlTyEZiQB9DQAoxeqr1EzJD8+9+klK10KSE5//oHL/PgmDGjXBGHO3nt
fDVuyzI8hVZ1ob0CUnWegYN+4VTpnSPbS4vEzlPtfFrUg4Ei9qqgcv4HTK9UH+mb
OHcb0DAyEHInoURCrDHF9+XkNqyNJNWhUqYLr0iAe/2Fl9TSWnT6goVsS9V8owL9
/P8oXx583h+ccdH+/xIb5ENWK3/4cx8jvmny9NAwGa7nCpW64h8RrYWZw3rHStv0
NveECOve33Hm2tfhqk8nQNA5nmfPEYuiclHbc9luWUWzqIAf7lNP9M2+go4BLTDL
3TKsX9l8JnatEPTtYK5KrLD9HhmJlf1cdboZGrMQcXGzy4qbtGenTo0+SDhgqntR
XU0uVuZoNkFKRZhlnInHKUjbsS6femV16CLdt5GPvwkYMLn3kHgBr/IXHm6GYs6o
+gExW5ybQ6MBtlvvCaIdaIV8eo/LC502zJ2gpuf1kSUUd5iT92QSeGOD7nX4kBwr
Wy6L6TGqo/Bv23sn+L7mduLJFYpBSX5kdXchrExOwnFz61R9wHP8XnFifzsmJ9ta
6oyXcmI4dcqZRumCob6AVqEBVcevVvw3kYebeuYNx9VQ5YTod9ziyOHIql87bO1g
YL7BOg03+aG+txa9hYboQufNi4YQPO7SM2srKivaMlb2F5A2cehApQEZwrFofGw0
pD3cFEFkw4GUt4Ud9ckOptLpBVPT2TZqx1DNux6dwD22/sAXiQRPnVItQ62FXc6c
EL3sjrQdAGxmHWrlSbLAL/pSRMaTQsRrcVGBMPwwkWJmc/sKB7bcF+eOTuSt8qXP
fdEsHaekMWVQ1kNgTMF03Th2cpUJfW6SYMkDy090p49TA+ZBL0KUj277VUneIV4M
8wVP7OgYksIt66IZ0EZvUTxp+ApcFhRUegFPnz8xhknrBdJwm/Wevhqf5JQEjZ5T
DXIZnZOII5Wc/zQ453NAOgqFMxVbRIsmF0fyqt4D9GImpUU6WNIwkeb+4mz7LEJX
yX+JGKJ6aO1Xg1Xxtl0iS+kmUWo265QLNskWwL8WoxxDSbLQscqj6MP/3s/k0zYs
XIor3JoGvxRGuA0/JR6P3ZKv4OSip/hWVp51RTJy6Kae74V/8iE9pzKIEk9Bcb0S
1HTw+V+ta1lkB+dgV7BMHLOpUOTrVBsvDatYz7XkGXl83XX1R6LS4fy8bZgKdPdv
F6pU4nyHkwQvymhUgspuMZHcfGauDUWgI1klASUknHNNdE7eNe+xFABX3HJ4dXps
Ys9sBj+pWugPkFHX0ZVvCyg/DIAMpzHS+86odqQme6DjNslVuS7zSVhKjjvRDgdl
85WlYzdQdmHiYYXOw9fWFiN6gg+ka7jWwL8/4q+LkUPidpLMllqeN69GlLaqazhi
O/VIkC7kAm6DAGN2ZueAJqfaLxlnj5DE833uREWCA4kYwIFsTrS/FOp3NEMwGuHz
Kjq9XFv3ikZcbVGhMNSyy8jUfKpl21USr/2MxT3eHUxx6WmaPlE0dtAOzFS3q9uP
/sVAj4hCgRGdKvd/7VqtgLghdyd9rf1Eq4m2KTC05+T+0zZl68ZsxiJ2VvkKdMOI
5Vn8lC1I1X0KOUPhYE7bIZY8ugxj5u2zZ6HbmqM2xCFSBeyMpfUw1InmXZ7KjCdU
Vs+hG0IpGOqxXWaIyKMfQmlC1JCJixuf6RMc6/Ct2wZ39O7s0WkxqNzMKslKb4ep
kknPfWZzyHB6yik/90FDQcbqINeaIXCg2/6A9xLOeVgPEhn6j3UuhidvuER7uC6x
CY7azFLe4hFSdgMld3Hi2rkz+S1ubnqOK7oVMhY7hA86amTF12sziyTSDhRxNj+5
POWr6QvVHBPEV4+ecb+LC8MkZMEb717sQCwbnYPXNhXv0Xmh/iv+ddIplLJ5Im3u
j+OscILcKpgsixguT7NWJcTtLTcQbbhSdn7moEOP7ia78o3PX8pqyj8T7Zdf4qlC
i+FhzcDlVFUlCYuacKkqsqAz2Qs5VbV6Jh9KXmpqKpZCzKcL7MYTLEPf8cardhkF
hOP04R6yKcebX0QrEX76BFH5DNGLIdmhcbn8xL0Vw2Ivzb50UW4SqHY2T2hHvn+D
GTEjSz9k541vWq54CVlQ1FOLFO/VuNuvKOTFN829RQm6OGyQdjMZe5vVwu9UEdz6
vm2jzzK1YfNd+Hjxf1ANAhHbm/EQ4/2g4E3nPmp+ftZNEj2EO7WQ1v5w14VdAqDk
iGeJlWWAdh0wv5iTUtpcybfhwKLLSvy0aO1ZI7l13umlVGf0caMzQqH9PlEGMN5v
SfSr8PxarF68VRcN+Wi9qCcbUMmvfN/CeeejoZUGjr7MKTc7Xn5Nc61qRxXd0DgX
sG8BJ3aS49cDEZF3gZHNQEA1Zri3BwYKNvdUFZcg1/CMBQkGkfsnn89DFTIzzYsT
O6Sv5yIWg5Ahn+1ZYoUQoWuzFdcyW9h37giBMP7P0vTlC5XPCbDzPHUZwCMdePN9
aBHmJ2taS2hTe8rwo2OHuZ6q+SeS04PlmzuuRufwesroelnyJfI+8ebEi9NVG5QG
F0fOT4l9oZIXWDJYCgOgQIMEJ5skuya78bPheFdvRIIcnde52c15QM4Zi4spAeT7
Ss59rzrYagvTawp5lUXoRSSnlNc/nIzqF2HyPq9n7ZgyNvMShQBybSeDRwI3IQ4t
q4GrrZZD/X2+oySjP9Ib9zjgAW90WynFzzj0zRdGgOgT+zArio6J0gXT7ERcPK3k
duTcAGSyh/oNJEj0L95+kvZT6AoeqqHKlPDsvmvKKPqn362AspfKPNTZbAbCVxWw
aJ4rbXglI1CvIo8FljTLDDbuAQlF5c24W0Oz4FSyR1KJ2vEQWUyd1Lqwmmwo8cAw
nHvq+JHZKwT53J/P+DekB0ManqCa+W++55cmEa18HRh/wkhsN3THV8i765oq31eR
XHhquLbaVtFzFaO+MCodD3wRnBViWWculYmEkl/XUajJVc0VgkCN53CbxSGNKrEw
9yADVegCmGQ4vR9v5XWV9umu7EW9+CJ+kWEDoKT3VecABkZHJpTWxRNpEWozef75
Vxg/JMYY4GWXN8+emzJgfp0dsJH8HjetWEJE587aw5KDktM+ZdYUgZ7hA0J1mmye
v/+0tsrukCFu3IrdylggJWwWZjLtRtVnAje57ZOj+ZP3JAsGnKZ4VR8ysPpqobUG
m3AmOKpNMx5vGwQ8CDjCDgYUdaddZgTH8Zr9ahLxIyHVcT/V4V+4wNxQGhQJAZIt
TPCpsahPVGuuBT8ZJZc5C/UUO4fuHEjDcMSe2t2TxWNgKuaYEOjiaT1ed5LMetow
YGqqPfBTBoFurMB4wiVAp51KMABe5SYQrmxJ9Meu4zPz7CgV+LOVAavYw4Ks56iQ
ZXs8AcZYcKDUTNdx3x5ypJGhkvW7Wf9VjpaHtY756b8Vsbc6PgtcB09tj27mlSUM
uD9hQI4iatuh9ENUCNvBn3LcxKg7T/fDzVsqCrQpit7AWz009einoUNjudH6A9LF
cR+J4YUGUUVLmMy3JW0T26GIh1A1EzUcPFwO0NbPzeryLEHq3ijytWUZnS/Tqsoh
ui2XmV5eHG7h6ZpFb+2nb9WSjztNB/gFm6OLuKtjf0eidhOVZjYNAB+G1QHhXfnC
fBc8MzIYa+vsBZ0ldz0JFOXH0ZD5w+hhTZo+uSdgjf/GZnCKpC8ZPjiQlzOm4H7N
umYHV1YFzkZGrFAmjKHlhITvhibPK4bWV2j2ruLR284nD6DSSXMspKuTQhYOFQ1C
qVV4uxFzg5hr9+tpzbVrogrtm0AjYgvQ8WtzhRYJ+39YbG9XPxEOFN/vjFPVMVeE
goNNZy/nNb97RRa20JQmOu1Em/SQmXHp3J5S7lHRxbHKGJ30dcNdTER8EN1rPMtl
d0BSyvsPMusbE8ZCfkRG1uow3sTXtBgZwv31cjkr28HLI/7v86ylRn2NTVz4Omzv
HkpBzSYdwlFP+k/ALp/4eCOEYfWXJkWsXG8KGfNoyMmSfUD0gHmR+n/nsaHS85nI
BmnDIKKjER+iXBeUl8J6Os2Adx7qizHM9s10iKQjxGFdrjrDLcnnlPnAa+9GmrZh
GQypbLkcHPPGqIUUA3y1igD7UNe6aMceVizBRFO6ELDbDjxtZLTFHHliFHV0zeH0
fwX+fwc0NliMBAHb0qtMzunGzyZZWQhEAG69EIPom+QB2v20Y5eYntCBdeRVUAdK
XK5TU1x2nSqT0NVKJKUF9jBITmFJS/mP4lPj87l24Fst8sJq/Xiy2ODl3aoYz/N9
ckh8txmVspHfXNK8At7O4s9pSMByvh2ssI85izfyWOZkLSN42G0zCNHMoihIuGiO
eLYxeySdT3OrsV33l5/m7708hoyOgCgHd3Bo0wXU7trIN7rK1J/D3Abi81YaLx6F
TYbgdS5sRI/F7DdnmTJlexKRXcrewUK7lJ2B9ZWWaLQkwyHO6BP0O8k7e0oPqv5c
i6zpJm2ZJvrNV8igYp91B8nuXvD75vtchfRLd8h5C19XNAB6E7q8oZgGGvNSmgUK
3i28NIpvxRh8wpbgdTl1Vc8956nxNx2FIfw9iLikBvKQD8QEQdEdAPCxEjKhd/YS
o2k853xwPHnnivTFM9Hlf8XWfrp5d1nrZq3nBN0NHiaETTAnl1kjBf2tKOSM9E3c
3Hadi+QyvqwErf6LDNX/ZFI+5zcI6XjzUTMLRINwuXXazDsbIDL9Ll5vXqBy4IbN
hI6G5wmGxjMkLESYQM6rTpQBdMAbD8BC/JiKFW7SBPhuheiAmz6CjMlsE+843AjF
MKU8+yzsLj+sFzrDDJ3a5KuXtIKYqNZ9kr9Npw6DO8Hw0sP0uL6piLN/qnZcFaJ4
yreE2zKF1gktu4CvMUv+fE0K3Ux5P8irVpNWjtDbqa7Hv9KKyM7+tZAVI1HWKaA4
9+pegihGi8+pxy5yUtSmbAapC9FmXb8/Z1dXQ8Anm88EbjQh/2/9rU8V1fEyqxXh
9GAhHR7LwsvK0bTcLTsZTVr+JYdz+Gk4OpsmZ3wfVhTHjsYIIJCjXIl5W54sP4pA
VWBKgc3mOey1PBWDeiiusXljcdSDQTr4DD6Qr0No0pxnDzvwbWF4txRR4VIBWYKv
yP7pCuudDHvYlwqZpAdO8DpFwmwxfyQL7LTArQGofUQKlodyTokThaE7090E0tn1
aEaXiyGlojef2aTP+N6r6nTMVn6sCKe2tRb6kAro+AkogwCAxNQMRrGhligPbTiS
aABW09zxGQOjwWJ4IxuFBGSc5h5dFiJ8QgNTVw6HlPnWdplIWX+VtQstP8WNjyUw
+8+Fang0w/TOufJD+s+AW2S0eWu3QiKHeFWI0yEjDVbFR5zrlnxRnwOSGo7OkOmG
jzf/iAJhwuxteH7p8O8AjD6OlZnpIU5NkFlNBNAU1x4ROpvKXhj/DOPxetjM24T3
VPyi/Z0GtyOUXPwFD2PuW/Z5etwxE60e3Hn2erF3AU2DhciWIXie8rLW8cDzOD9m
EakrdRpgXmuYfJeHqqyA0OkBoprcfwKVZEaknMepQN0KBsBUX18gI9XpHvcynmbk
r/KsjjQsPoA/ZcNhEmTR25Vwqd3a5aWex56hUxu+goTztLdJEGC0DH94+6umhRYd
Dd4WRbIFvoVU4MHh8dwH9nQ0FnYs2Q7hlhkvVlFiweur6WajW6e9+3zWqUsnSvts
wT5+WZa+6B6Z5rpVsjEYUxETHGbgDrAcjC/ZnyHfKZyi4befhGzznaM4L+nJMnYt
6kBm8oklNJs2wotZgETS51NvCySUhFWO5ePxyEScWDXDBourS1cglVm2z1XzSGNJ
bhF45iegzcyXId01ZUn8M55hdYXERYzAadtHTMsTg4WETI+CSFnHsIvvI/32nO8h
ROj80iEnL7KuOCk1vaAUjy3W+WAcGXWOEbzm9gIGjOSud4VVexBDiS0UP5jT10qZ
W0IggbvJ8BNakGRhHqquQg4Mb+Olo9+0VeKeKnshp30UWr6zkTOlHEEm0gM9c7fk
H9H1jkZb1dbI0fN0sGVdFd8DZLJne9WI3LQsMb4+XFGQq8E5aaQIAy+dnu98OWl+
K8nr4rffX6R6mLyvIygp1ouGOq2+TpQUZlrbP7/n61OLGTDiCvjZ0Xd/Os8gDShS
ELoAtK6r7z/dT7MPlPsGBMW2q6fAPV5xvLQxGexehzA1z/2DRRhXxMfeb8d+sub1
HAY80rtYqTS2ZEp1P30FrgJCXNX3Kc9uJTdg/MI2o0SSGY7+sAeE7LaWJVYkJYdV
muXtLtnKd1hzrzeGw8FXneVi2VG2OtTirvsxoq5OtNIq0s89/Q+67JcgIFxe+Qik
r92iGfK0XIJf3WgHS7V2MBJ9aOoEWs9w3wIHIgnXMK3WfZbQzchZj4TiH38wdEaA
isnnrFP2Ebz+TMFddqH/LPhWMzcn2AAc97wEbgvnKlwfXjnPcudm+VC/ue8+fWEg
b2nfJWUn5uQHXsaf76UgHkNo2zuAZZKf+d0VMqPmw40VfB6S9QxE+bD8hHFyEqqx
L0jfANhYCs8lJjRf9NjTEcs0/pIhtuVu3KV+7baD7HN9jFK8mEjxNqQ7oTZsVNd2
3h05qr3n3cEaySjyT+UnQ7lYqc1VR4G699SAhMjhkqGsyzKeVUXKvs1gswLmUrzp
ml9ilJI3lre2rejykcHvberKCXi8ny0GxulNn1uZQa6Q3gubC5CICxCnP3IbgxFU
qejZHukMUqtkIGFzljJG7pwwLgNxFX5KxotHrWpkzoxm/37z0+ay8MDpudQuZRcC
nyeqEeXaCMhLyFXDyJE+OTjsUlKT2rXh0V8Q9vkR0F/YQPmrlBAopde5RctIiuuP
i5uf1xdU8edqFNP0/SV0qOiH//6rwDu2L8QNvNgE057c3FGV/JBX1tUBF6HWNPrd
Bxo86f1nXRzLv06uhEIIMZ/nbX1Tn+LY5D85E1Zrleh0sd91aoqQ+igxNh+7t0Oj
8GfAIqvWVz8wulcXMQvxYLUv+xgnYv09UrqTZl3fe/B0L5br0+1AhkJn59WH5eNG
JLMHGsmrgmWlO65qLpHSszCu7TJHzkwabcV7JWp0mtdqeMF04RAO+Y6S6KG59Gtg
Ef4dLLTakxRb+ljo64ZLTfdG7iS747N4zSPv6asd8x5BUeDevkjNBLBRewEKAOli
URx+oOYAQuNvtyWs1JpM2HrKcbc4qksQ0kgrUrclk35mc7U9sbwynytBrhjjsV5o
exzeqacKR4Z/MXx8qIV9V+ZYTzztOrU+kr3fS+NNzvH66e965rP4mAoOZQw883+R
hEVk5XZEu0nC+YLUbQFHyHP2+j7INnEhKKXSHXsRQ3LmO8fR0WUBSxmUBKdBQtnj
6egvFfhxFGaoxxfxcuE6BlIgyYSWnlCkx4Xon++WHFO2aMm/queKBG0GFit8mXrL
Tjw95m4NY7igRApqj3+C8V/6jyuhY8dWHmvJ9KDgjkeM7G0oQZpS4TlTCK7mcN87
q+LKZlN9ReuLBLjvOj9bPvM5NTzgjM1Oc7uZgo59uMdM8I343JIjTx6SSrJ+JDat
4z4zukpZakWXW6Pf10VRdGknzgVsM/3Nqwm/7+hv8Gq8z9oYQbAUSe3EcdiDBqCm
1uhMWxOZdPFrN6Cd5oyWz/uPMmNeobCsVv0mVYF/pGM3CS8s6NhkGNK+S4GtdZL9
3jANlt83GDHPo/haQ4eq/u+l0pL0ZZjGuqhY4hXGU5ty/HoiVxD53wNLtAU9egp5
HzqxCWvjG7gvn0FE/RRLkloLLczid5t0tlUZCTfY13j2bHcSsuSdGI4oSRa+JcBN
dQXV1A0h9oeZFz687uJnlY3AUONy3eMwKpa179+NNUH3sHk6CRHg2V6brOE1XWL9
VDRtEzFA45LB04oQNbubp5WZMq0TBRReqirGu07o2fQt3gjapja6bsciJNOMHOTH
/ygFz4AwpQ0I/XKEJc+n86F0Fw8Pq9HccoFJ20Lo8BQp9s4JFofqxKKhbQImVKX/
APAd/a4N7v7vwDKdbwNxfI9TreT4wdNpDwv7SAgJOPfstveOZWCUB9sXomCHjjCT
GVI6R1P5UyPRNLsJdLO+r84V2D+yWYA5Hx9PcQlkyjnfeIZ54ZcYUx/bT7OX6BAe
7+HFTSWUWHp2JG0sp8SQjTo24CMSJ9mPLeMiDq+Pr5XY3Ty3YDuWlfmzAQz1bjVJ
EYH9ECQlgnZyFiElcQHabZ6pqry/sjGXEj+MoGNBv79R9I2hUkQx9Tcs0pqvrsha
NYa+g9Q0HdtaQvqhlOKW+ozopjMgQrAAbQ7EnpTlP1hAMHcmW2L9E/8D84tIraHj
tX5bJYYfivUv/2qwZRCPnBiFkVj/TW23wFHyARRBVpehFTzySol/0ehapaqKp5Gz
a9AtdRp51Y+0C/WOWeZlVbNq+zZNjMTT/KMwqE5XApcu6xhxavkuiVN3jY7MlKkY
64eYT2BDmHMQuICsZF09HUQsnDd2pR4jTK5vUVmiNBOEJsMEMhpj+tU4yqzOVTg8
qaoTtDrz7zbY0uN31UsylRN4bjCZvGofEJgdho8nf0gJ3zW/nalzO9SskJIXfBXq
52QgGhv4VBDIZQphNUluMUWMmPqa8S7o6jrm07vY8vcBc95z37Ch1dpHsLB85Om+
ZFIYz98teyWcP8fpjpDSheHPuhoevFtLgjX7F3gurKptFxxWQsUc/Ord2+HGVu4f
thZUHZRb/my992Jrvyql+SBkUZdbsAiBpqXbZS8P2/6v5fNjasBlon3H0SGt4knc
kU2f7uHwqc/9/ft6E40bJuPt+4+t7IEkXINFqsE0Yfov86q2gwjg6kZLx8LXWh6B
y23yTjLtYbaOeyvGUu1c72hJMncdRyXzWzSqoLM/Rpo30vefGBBsXQxpRHFU3vy2
VQ/Cfv1QJmg7tXIfC5mOpiRwlyxPJyPvxpnBRT6KLmpIWk7BXQ9kCTy0MYOgXZlv
CtOKQ8Q/Jp/m7AHvVXfqgwQMyl5pT1wPGNg8lTtu1n/5OP7513opoiqx+DwJZqE0
8oY75/sPvBesrXAsn0KEd4uagxYXWK8Jy1prwFh0G4MZcr4G00BBltCZ1x5XqaYk
y6Fw4wg0jXiH8rsVhVJULTMFdRn7Etr/28atnIiSQN3dknWf9C5ylIkGmIawctEQ
EFcUZ08Ahy47I/sjGK2yIn1c4B3DnUvYNqXKr3TDvLfNoPEv0xvRXJ76wxEqhCXi
heAdrrdCPb/wyvextnX/7QiVpXuKzTFizKjrGZ4aO2SZ0fDkzo9ARpAHp29sbdMz
eCW3M+5OyYFulY94AhUYtXMzX4t4CBXpYzMu6riaz7QhxtAOIa4UGb8IuiJ0+H2z
wSrY8+E2X05x/xl3Aam6/iNEHU8T42VhUnc1dr1JODWrKt7Qbt/DJF4UIye70Qc6
jqgbQkiHp54MoSIps4iI45dTzLhNnBq4HhgJNxmeQ3Tbgljr6EN6g42Kwl3vMiQq
XthbbT+1+XWMZIb4Ll20hhRCXM0sg+qDt1VQ0PsGYSbPsp1vrjyxDpeySMtm6U8L
lYBnoeTzGVoxTWtVEwOxqlaykAt//pX+3hmA4eph1xc6a/xyNKiZYdsyixZJD7+E
7LHawPpl63imDj/m1mYxJgBMo2Dki0A0jax7oHCLb6mtw0sJAY737zaUmXk987et
wnA6V5oZeUjaP/M6paWWv11+PxYnwI+qiOfvzG2eZpjCyvZdPflK4HQHZxh3OShL
OZOPpH5Nhc6cnkIgdWPhElTXxPuukJR8lYbMjSEOnAmzkT7JCDny7C1TlJYl9c4R
EgylTY5BmGLiZBZHubkJOJMfLTN5vIdALGlmIICoT/EogkKmbxwj/Bxf/YmWDInS
xY28y2SE0Aw7N6DnLnk0R8WNUag2MuSudQTvKgu+/VJa83nH0Bn1LwI0zhswdiUT
a7Ky6nEZXl6NDf/keJUIsPVIXLonrqmDszwPujVSFpcT3PdsEleMXJ3paEL02A6e
ZbbZ6oUOO8N9uP3ayob8rZjCXGK/BCv4bo4bU3LCycKuLESjUPxxXab0dwnL/JMq
vmfy4qtlbyn6XhJWAXQBGP1KwzQCs1CRLkHOb+9oVtW5xFhB0UKUM7jafcyFR0Ed
dguEK/I9Ce732Z6HioEqgHhKNqd0xkx3r1x5FPqHnHZV9S9Jw2hqsUOsV0WAYOG4
ku9pzSWYKuoxDXx/zB8lPsm/y2C4/KSr+7Y175aL8GqYZ7Kj3ZXPKxLyZqM99iRo
yhMCOXgO1HS3Sw6LukaPC5dY2XJS2AgWFZ/ZKZTMVNmAuq/t1jfbNEIzu9UlNdkm
+H+aO3qw1+GzuPIhs3OKPmkB4totWWejpmDztfyohV8+Xb2WhLivAnRL2svirptb
vwNlPLVTMgAL6rivaFxBVxL7Kfn/wkaQ3Dhx1J+64wzpfHiAGeV9F4l+e4XfTTe+
iID9dDIr+SFW3Y6M8J2KN9RL5K1wICDaAbnZW0EgyAx16Ae0Xht+epbGoIVCjP60
65pCwKApCdbXTBQ6YTw130CvlYTZ2nLQ/mJXuAtptMNjeW8bjmTNnaFiFDhJXotD
eyykuXr7EcWp9EOqxBhLHItf0oGPXYRbujij0RApeguvVOyokyghZevyzmtoP21M
zkSMbZbBTsIXCNiLC7aLIGSIeKG1E7BZStqq6XjovC33JaWVHGqIfvjImw+AK8n6
dt1NP39sIw1QY1ViPY/mB7q74Qov2EHVod4TOkW8GBxcYxAjp9EFUvCXYE9voZLk
vr+bGBU8g+S0tjhtTJRusraknb4ThuvPQzNIkImuJUz7SZqlEt2cBCHU505M6N7h
SqtXD/NBXW+cG1eLCGDSKwMo0I3Q9tSA9qFGjScxNajlnBRzZfo8aGC+9BmeEDFp
khyLZ5/ya9gPWDhQWeyLNr7jbhcbOijqAQ5S+UGsjSg0m+4USGWNSPAMydTgIUhp
DLLDIjr2R3qKBtLWsta7kE27f3MAPocxaX/vsCO37sKZb7VIi6SQC5CPHFEZhMrs
S97LO3+xF2j6kDTOXWKDTTYDjHCPlSpL4Pf2bFa+PqqxPzww6hPYPW6suPwpy1NL
OvI32ig+fHB9L82xqRGaByvyNkztKRSvlHzVWX/TKHO9RXRCIlNzRymOoay+wnBw
/vYkhu06jOSGlGQZ79JHndc4MvzA2cInwAwqf5JSp+SxDHH47xgvzOAnkQ8d5RFg
f3ysEjsPywZvhS6hceZj1iMCpax2j+eOhY+JYTI95G7yg24jRSYk9pFN7MfAu85m
Gfkj+ApOSrBaWHJXJSF3c24y5ydeNf8GuqcbeIi2KYRYOtajBCQ1GEL7LKP/yAv2
jacGJvcEMp5Jgmtbwivqad5wFgIk5YPb+K2K9rB8mVxte7knDLTPX11hxsQzPlXa
1zQKaNZl4Woepop5UQIteSbJW1Fh2MKtOkUh9h+WlMO0ieZr5tc5AOC/FV5q0R4r
YAvB5O6x4Pu8dBBH+6PjHT6Qf5AMdVncUGVCSrg0Zc4eGBO6Z7m8LlGBtsuAwTQt
+ftKR7S1FjMmA532hLEK3ZhVgyVD/fGIUwSXnkcJ5FbBA0q/xTktkivNurA1J6Nz
AombEgOsFXMHXzsle9meZgpESeqtUbQKplGyAYOntJ95Q0N61w/zlf1tcMhKJsBa
N0nGkI3DMz6Nz37KP0Ne6kHo4ovmhbtIKxeQ46GVI+4Udd2yKFPE8j3PJ5OnRySs
ParnJUuIAY+kqEeOkYv9PynJ+v4IXUjKwjCyxCD0TDPuRg6MEL+RoFu7hmB+LbUH
NytGC6641AHk+EmaV6QtBb6ZqN7DDUO5YUUi5GLvzZNz7/zugHhXXAaFVtbOmqKi
JU8Tfj7JwJPeJg9vKfmq6DydG66daVf3lRo9aYhtrj3fQHqPXg3E005Yhk5A9tkT
+li664WvNYVi5vrs22gWCHm7zie1tdztRi3JiHBRva+N2AENA+DsYhuBI92ouBgg
pQI+Tcu3Uko0ZqshavBPiukqTtuwmaRvXQ8t7CL+zls6CKUCcoKJr/JAHkVCqA/0
Qqb7Eh8GW6X6umfuZLJY/7BuaBaolcIleEPnCDBYPl13diKtvtWAelzuMAV3q79e
nE7oGcy/zQXdpeqW/OGPmoqFJc8etb4eOxC09jMicPH9fBdKRMZOESUl+GxKyvV9
BqgnviayARCgfbU8pRQ33POgOD8RcXOOpBxaev85sgCSIfFO+mapkunaP5FC+6ul
gbhOEEL4Ed8yF87MfiKVPSLnjKLIcitu6Yqa9ipHi7+l/avrr7aKZ5IrS1fTsK8M
GzPJEoG02FCIL8zI4zXbiAun2OChhb87dtrbd2sgzK0qwMtYaeZfZwSREu2JKxKi
rHiPiHdALvaNcNNArfoYxBHnTnH4DjgIPd4AEASeLEUteItpDD6drdawHZ0gUdqC
4nEbGieGZenpm8VrGtUk7QQu0dKr2Hzc+dPT0U5DspjOIofHwGkBwzHJ4GaFbgV5
JPeo9a5oR0wTLuZ7S/cCfCWOdpMSEvjWkzIorHsdFXAeSIwhprAcduPjBEWKc/n9
EhQUJQY3umR2WsR3MarvjYP8cj1eZVSbkv4Y9VVwyE5+BP13O/L4rj6LonSgaibJ
ksnouYItAOp6u5kzBVunasEMAJfotJYYq2CCYENPqRl5f15tpx9hC57jSJmxSJrr
5cTX/iMkxN0W2FquYhYwxbOJu6BE91Ca5kTqjpD9lpTtVuxBiHbL6DiwZxmxNBWf
sQ2OzekHzR1bG0dus9WjUV9Yk70NSdRhGw+BIwVsU+aZ5qNbTxHLSYJJWqkhwH/3
juXXQuCHevnqEHbm1/H0pzfA30GHB7TPWAx4dlJ6hnvMyXNyn9OxIV3BBaNzBau4
GAH+NshL69UhEyt+mxCXP78CwV7X6ScjUC8lKcD7lN49jzxXjky3dGEaOfZkIwp5
ZXZ5NciGTyyy114D4b90gzaOVwMqoToQvcBWwkY+hdXL71A9By+Evc5KFJkzwTnj
R3QREt5cdWUaXR7pHiOoFs9CLYyzIg2Bp3HPQQ52f+LOfYoKi+8D2w9U3NAvWj7c
Ug9HbG0QqwBq/KEsnEJhwEuqhWMdaRmNr6siFZx1HmBSAm4FESv7W6og72oRca98
3GANeX17bT4lxAYxdvc8KGSYRoDzNLkl/CoapcoP9FHCG4b29YHDIPwb7Apl7cct
nx7G65EaMaVNfbU2wfSthwtmGxfxWVPwO7eEOK21r6igLF+gxnCEGfPIKsDcMfc6
twDLW/qqlczOExsmFW22WQZ01Z93SnaxHbI1XjWkJV3alryxl/mZI0+snWRcyQtt
hoBgrUd6Aayzr2U3s79izqSxoTQUDtYMeKyloWLGv5Yn9egbXuZwj++7VeFk2YSv
VXtoc74nHASbESO9EOtVC4Qcw/B2bNUFbEHD98Qel2HijirbC5kERY8shYmCawXg
s0clrJPS1VMRkDLiPAepDCR8AyzKX6d1WueD3+ldHTwtrpjH95Ihzz7AvRdZmAT3
uy7Uie33Hjw5SJTrBZdMlBGlbldZUdnr4FzLzw5kYkbulSQ2snBL1vrrAmkSfqMO
5Z0ApzSfZs+ZY+bEBNBXPUVlJLpULDW2ocsS9CtH0Ugn/ZxO/YO0g777B4o7PyYz
HKHj2Kp1rvJqmSJSQ1J5HhD6ZuK+5Y5e399BYhoy9Z+6ZpzaaRtUt4IkfVCrJgU8
M+RAKDkmC6srT707lhWfABgJxTTuUMv7sDAAwowa/EXUKOeBJ/y6BbEYRaWxFMTt
6pqjGKmnNTKRAx7WUaoT0fXDkTixLOLjWQYGzQf9yAEuapUStwQTDAqTcwcVEOLl
eRgYX/wMu6/o/wm190/Vu+tN5Rq5bmtoOMQNRyY31SK2iu9pt+lVvSGuMYgJSAqq
pgTlhHYA2Gp4JViApMK75caKUJin2xyziOdFquIWkpuazXqWXlV1kZNBORiGDvVj
5rGhr58fVwwPGKgY3LkFPd9ViPOMxEx4TQraJT/MSHn5cBLQXQ5zZ25TS0WRlrim
hMPZ2lj7vIr5uDVbjAbPa3WRiIP5Kfqp2l098Oe9souLTG3BJu/LQRtwuuxRkbMf
WkkCJqdw5kdEKSIuFM+vy/a/ylajFr4EM2FL67nmPcTPl621OdGYQ8zNqmF9v0Dp
FCxjVPcxL0brthUFRCU/H4Q5D59Bz70ceYc9ZzZK+ctNlMMcXeSl6SjVTJ4VStTZ
hcgXNHkiLZhYM8wcRuhFZVddkXIx0LANH3z3IDYgEIOkI8X/PzuWY9FCnlqGP93c
nn5LzAnf+IOm+ep/nELxIci+zrfRH1l7OnFdBhD+qUpCNqL/1BITtEP/XmaPCGXu
iqDz9X/1R67Omdj7Rrlc1FDglGGLK0qrkOYJBkG449p0Si2ct3uR1A4mBqJVdvQk
YVzJEzC+w5gN8gU51BzWXYWmBQL3DjmfggwRooMx/0PY1HmPPcFAklixrJTvo8go
9Sw11QBXbNVrGsrSJ2+CdQ0vBoY3ptlIiqSxmSyYgVKsvzLr99SU2QZnSSdoEECO
/mHJu3yPCEKIBM3S4nL+IevybR3KZLOoCLmoPlVUoGyaf8YyJU/zY9K+NOMRUJqc
gSCqQYUrfFoAu8h6/jG4Rbvu8gNWSypB+iNTYpkGhyRzJC8Cl9eEZFn7ni0WiAvC
OF38LhmcOgQvIOWIb16aRKdAtpRLLk9TrvVBjgqMpklAI/O8WxCLZ+8p6FV0+TNA
l6Gfmh0i+klKlwJyX3L5xSgW7MvIdMNJcb5an1lX/ra1Dszawrv7AjIBx/r/n015
C8aMyk/MI0w/oDevCwts0RG1jgYUtsHuLJgwtKPlGm38Tb3+fyBwsdFgAKyb/A3F
0XER0Hspdl6qfO8BHSIiBJOAxQGAmOo/UKyifc9drl00eu26atrs0ZhlReoDtla7
ZyiftljBbpuvWoryevvXa1ZDJVwi0SDDThAmuiqc+2c8ZWrj8j72AjMHY6EahDGH
NwgcTCrL1f384Hv5OaydO0C30gA5Z+9RUgBvS3WsPAjTNLxVx/Zww57MdJ2Zsx9+
RR0ffjj20ZgGQrNySo1iwikTktr/WfsJF/b/JL6X2oXb/JT1ffPByhR3KdZdYJk7
qCGLekEsASIZVnfNh/FBSMgrzdBzOGWaw2wS05ALkqtGn3+3FF+EruoqnPnNlhJT
NkCAc+JWvV9NeQX7mOf7h0B2jxFFbAMDV0WzySaW7seCon3lPDnsnFeDUw18Airf
AEeQf3veQChxzrYGtekvBaCacvfDT0RNCOKwaWfylsWraXaNFQGz/ySdF198Y/j5
NSU9YHHE4fTCwha6hAwbQbEDWckXVp46PobHtNkm3X13uJaDFr/ArwBztr5v2QQW
r0qKsHjFw9gmbhVjyiebP7mZpkdLJzjiGQQUgR8MGiC01W9tgfT9XIpywHXLSeDe
L1bYhwHrKeC/mXxghFjupLPEk/zbXcuhmFZs0MAacNZ2v8xPcSYFFwxrz6sYjdUq
QV0sROGJZdWWEYc0BfUgDI22rKqqa7ndDP8hXGIezQ3t/WET/ax3nkxU3eI46eqD
AEWCSRSWpOtKQy3om4dXFQB+/43Nyu5t0PPQamWIHo4wMe5+3yUJJXzIex/aFgSi
HOpi/cEN2RrKGa7mEzBiZjW2FxEHZRLZYHHcanlAi7TxfD9orh62COZahqSRpBj9
UZ0SWt9c0C+KftvmhCs6lzvJn3eTQBBpZUn7LKHI7pCzhQ9HNvIVYhbQl1GF3F23
+qEKd6nUZaGvICJKhB/+TpI2AM3rodcR8avptMlKDCZ/uv5ZORSr4xTiPxHsmAQW
ZLMeLkPK+tmtiZATEFR46KzlfJVnJYOYaoScDpZETRcEJRWTvwmWR33KvgoLU16W
CHE9jx4f75sNZA9j1xN00pG+0Molincw78aaGR4MfD2hmrWcCLzCWspe0dFMVG5d
4LEt8Tryc+Eht9Y3ffvNYwWAwBVGmtywO5p0XRjvrcGgaJ83EJ9n8HtT+yXEdSvD
n/EifNk6jfUT7FCVOLg/7Ke/ilJT32pqGycQONczDOtZZPVYJnXLaYp0SVPHk5qv
LTm9plx6hNkeswig3ufbfqK0V20zrRinRohpEWLYxZ2M+QOSFXZ1E471EQN+J4Fh
YjEbDEkuLtLsNJ2b5zqpzg0BXoEvRz/yvyl0UA9RlDTr57/vE1V5uU+zUKvemiyq
wH8UFRvfAnP+zqjMEIammiNAzpsD6Dwx/+ujVcelmuQW2feDdb7doyo3S3TAzIVX
fQ5X4tbw+ZrWqsW3d8yjKw+1bT/54TYDG6Aq2vol2L+77598sC5gvdH8B73TAIFY
yMk+jm4dPp/6MAKkipH4KaMUJ7Vry8We/8NB5oXTkmZdGZU8xqyY7hmV+3g5ym8M
zeaMqkIITh5Mgz9CJ7EBbKfU/uRNn3qGeanNsJ0I6PlTQP/YJqPhv3ASFElt7ziQ
E8eqgCjtcpHTzI9XONZzKmdFXFPJsffMpoYZw2IggUryTSsL8cuJNCUaZMO39ehe
np6LjpWjo4njB9//R/zcUSktfb3oxT1VOSWe3I4fSB+wZJwrCa+vHOpF/BbT/uEh
mIgOG2s5q0B6h7Y3UxTS5eyEgKpleuX6O6/yiITvY1aQfIjFkX37Y2JUlLh77sY0
uTEaL/YrE0PDKkg5rRKzC7ju/o0zNx+6cGnGuWhTtA0Rz4zZ6ZXv0cFCLIb3Pndr
ZzNaUolt0/lc4rmaNCFLzWv/aY6rIyHdGIn4XOtJ74paQ1WPy3qSn9FG943wsBnY
r7l9xp/yrhi9F0oMtxhDGIasMp9rB+CuJluM2+7rMPLIqve68AbKnnmvfyK4nBt8
4NIQ9Te88UG8z1Q5c+PxIWK9/wq6zEfx3QXVnRv/9v+zk14/Rd4kmCq80e5GcfP5
jEhhF6tzdmFJGzPIUKbVmGQXcUpDl/JGrCf8Y96LPnmX7L0xmu/Jsv/MwJcsTxA0
oCCG0zc09qNFo/i6RgAZ4ERpTcTl64dDvxe7rSNbSnxiCYycwWotreYDQTNknu9v
TFyDjZfYxhJDMoX6161iH4ZoR7K674cbW1kSqN26j1w8ymgmjUC5AczH4gcvdm4D
lHbLnUbiJWB/A0g7ca2HqO8Zm4durzoeVI3H02E5HyYFutwy7Nv7MVYHO/08hmu+
q7cFhWvYzIlMMYvzPRypbuxhzdkXQF59paX2YW5zUSzUf5mD4q20PjzLB5fITtg1
qv0pG+zyAaQpxR07k67VgUyADSjCqnCeg8C+U3WPUBV4pXJAmkRjMRawt5A8PW+b
bpUOztNkG1OrqBUFx9tFaG5S58otYmEMJgs9Si40AWn/mQj1RBs7n39pgABHUTDT
O3vvEfKk6NzMjVGXkIMsxP2OXf5ehPelEjZE0VvG4H61/xYjDTBG8gmUDQE7zjZm
Dm84sGQ5kTKkbvaEtIVjHEjyk5c0RPZX9qmgh5iX2Sl+Z1pIBGkqKO0ZM5MM0nuP
11xhGHdptnhPLu6Dk83/ftoiIhLNX/FRsoFUB/rchyYPFpMfmTfqTbxWEN+u+1DZ
Xsrnpf4+uPoIlQVbMHTVJfVLxqLyX3endH30sSvhNDoFmdbUcmjkJ4LOGHucf/jm
sa78WQq8j1e4pK/PVkyBrEBFn+AMTj5oVFxfEaResf5jzWxCzyB3HzwlxUG0r72Y
0kjIJmRBw460PkD/VCaziUiv6zFezQYv6wCjktWvgkoQMBgeeEYNhsfXw/303zCN
VT4uMy7zDHIy2L1u0TM+yn2Irpl7cbtzDsyv6ejBjxEEuqV5x1yx2HjT/NtwWGU1
jq24Apf8mRsBadhvOTq9fQMF8pZzaHHai0tIZ5REhyy2Rj7oZXnP9wTG11CWCyvv
jRHkO2bP/Wy2EJsFEJE26i+WEAvYDNL0dCR7v1JNcD+VgGmfG+YJYkGZD+1zdPwc
Iz9sMQmnzo1MQhiv9s9rnJOOKnvOOqM5YngNiPCOV3yTnG6TTMTHyT4q8hjk6n0W
MfYrBwWJMRrf+DRcn+cmqL60UO4LcVrXq7aH+t9OG+mlrS8ZRBBQnAWdt6ElDHdt
hYxEBHg8PFDAxC33PeiaEDzNUMDjOtXLE8fyF3kcERxX0i9jppxsXXyaPAn4LdvO
iayFfGuZfEztFlmGZhNc6A37Wu2DbwIBV67ygENWDGbgFxg7DQ+nf0XYasm2D4/g
AJ32OJvp28uyBP1W9x21gEF5oVPDzN7dlNRPhIn5YcYlngv9JaJiv+ZiJ9oQo4MW
V4VOEWfGsaBAIM+dRWEk0sIsuNstzm3EkcPG0lntfMq3f12k/YV7e3ZzBUm2/ePe
yA05JenFz53a84JnVomCT7vCjN4Z327se/2Ph2yd2QoFzE4aAebsvOAFBJ67UK1p
ZXBS+HVkJyNZlpoOFuIb2zCmCwPbnxUamnT4MnOG8gaWDrQXwhusRk15hfhinNXt
8lJua6fmr07CLDGV1bpqWntH9LDRbRIRCJlK6jkd7FCMk9WEynEGThr1rF9RY8kb
+fP5Ejazba9Ygl4vlw1fmF4sb0agM8JzUvjwaxx0Ke3watpzwyO/YlpXGKgbFDGA
vPxYhC+FJC2tRRrxRvX1/iiXKyW5rhWEIDZ/V3ifr5HC6gHSJFrsMfMReSmlcZ99
ezlWj+a00XDPfsJKqqBZxDO/iZaF1+NKUeWePNyO2gTfjofr27codB5tgPUK9B95
6YpdRrCgDdVDh0VGxc+1CJb6myyGW9emKHw3qFI0jlbPOM4QD6dp6MYMqq6qx0ve
k7XZeRGFYZ0kdLyhPsttDf2JRS3yRjWXHY/YC4cDfX79E1i8mq9CdVcoWrA4kv83
wgH+FLRfKYfEMLJGqIhNqEFfv6eIGBJ13BWgUoo8NuWtrJ2yWwsEfy90onfQpJs7
HAp0PC2An9+8hSBe0HopYanIXbsJQklxjPggXN8IVtfr0wewFcYiWtG0iYSPubm2
OZnVKeI48BizlKOu+tGotH6GyQhKkLv+zT58Fyuzd5EJWSTw4RsiiXCru1h4Jpst
rZXiVTLMKgqkVg/QOig71/hy7tqGd7u3/wEyFTGhVykuI5zXT8x5G3U1YpAREJ29
T+PsbdQ9qTcHATwhKBt3UQb+gL8Sa3NYNS9w8D50QD6mjX1ITsYHQO6HYp3A1QYj
DQ8JY9s4XH0t9HuUKuQBmI7MgIk5y6dsvyTXBC9BWMgMrycVi4y9XUGa6kv2Bu9e
hnaKs3lj4TMJVKu5MWrM6mb0pMYwd3sFfuXcB367735nnaM9KCnYRi6op25pM2UY
S5uNZkZ4JZ7cHkA0rFGf5VyimL5FCyO7JnnRLFS6KSEMmKLrRj84p9vYvGl93NSE
3sr87IFuGMk2AfQNoqhmdgyveQNyWXfF1edruFWzomvxpARdVh33Ea19P4l0GKJN
iR0DENUVRA/LXXhNheLftovETVzme+e+TI62NZdWbIXsRt+xMV7zLpiMT0DHXqOA
uzAnoOP7X4+0Z8vlHl61PsQU9QnMmw/ARzzpl/8iIP1HqvOqxK1ucLke2goPCeZd
+NPUP+3YEaq/POHN08I1dGpHbDVkLU+H1FqLpMK0ZjRO+PncyJGfc+OME6x8grDx
/ZjTe/yDbMKCq+UrOdS71QLG38b8htQEKcJhFBlk3+/0ZEnX61u7ViAC9RZQSOSe
0D6w1h2GMjkHm/FBagvggXBfm5OgwhUihUBvrtjjR2lmcJcjxafqum1978jXJzkA
flIr9Sb8V5rAA/4d6zl1weZpy66UkpGKygGZ6uHPDIlTdR1ZQu9bj+9TgtxHDypS
NNPB1Fq3EEyLCl6d+KLAAPPZ3VoOqtzEJT92UJ3PngUolPwKfLjqWsgRp2peA0R5
JjhE6zxWat+g8gyjRkGTnzGx1m8JoA1Yc3PiQ1omGba5DnH6ivsuo4azZkpH0ZiG
Rf+H/CaNhC2BF3ahm8V0zUBZoTgRm/rJ1oAn6qH1kNcyW+Lmyg9/noPZ64xtn+Ze
pc3LGD2m+70CJSiwFFAo9PslBXcaukw7hyRQF4BhPgKKk5HAQoQr5VIY7K++cBeu
FBU8CSm6rYsCOke3oiuwDCvSUy2fsNJECLj6vk5GAAuo/OCHV0dXfR7wrfZyFkIG
LIrPHHvjuZnwlE9s5AFvZeAuRm5AyacUk/voZ+0Izvki2WQhx04ghgBY+O840a28
ZwC5l05UeircEarlV5ofD9Z1m5BWbDmspAeapV0xvRLv19AVdPjq0ET0Tsdwm5EC
os4wf+wHwhTuoO9ggYtjgQKowpTp5kLI4WMLsekDf9xFlgKBG8qAdna1vQZUYGsd
wdjNWhquIuStJJZTssMMvjcc+4Ppbg9tvTm0mocPz1C5eSwl9HsuGWn7nsFAbv0W
rNNFcprHOiLxCpK9pBeh2D93vqFknmii1doODYjyXBFX6YTjT4oXBHNAcTiV+Zkl
qc5TsWmtGBMSG9XxadMY+mkYL3vBSYsbcOAmxGS4T/Aaurc3eBFhEculApDVn2rD
nWR0x87BAX2RiXxVGChL33zDmsRV57GtDa0EigmPIpMam/Tc/mXMYHbK4lUeScb1
mVYr+OJRF37DeuyPe/o/aQKDpeVl7zCiF8h9kLPo4W697kvFW4/IdUzFIIkAr7Vq
MAKrjhDB9I4rxMBELOR8wMBTHedNR0z1Y/U6pr+GWOOU2ymK/CeuAs+TeO1Q51qv
Y8cyPNAGFxf3sGwVDGn/sDzk4Lh2J9wgId+spO1T1zTi8eu+rByP2QIxzogZhs66
6tNWJhwKESsRFeNJp1i5DnKHouFp/vwg6bO2POkN+h9Q37lP3AW2XI7rpg1dRTPv
ihVZiesRWmygG0TJhIT4HmxeSq/YlvPU3WmMCRgVisU1WcReRzsCrH0SlevMOrib
eNzdpXGqYSHmFIcIhlsQcgK3e40NHqKl9ChcB5EYX2nsbgAXRM24djYz8uNxekub
/Qhq5NaoQhPOQjfUNINsZDdL/9QE3QzGFVE2TCrEvCPPBi5QHtvTwfx4ZfxBPBPV
jkb3+6V05eU3jsigkCRgXq6Rb2opglogCMBmBy7XRUgEG/56Go3ktyUqfcgSZCeZ
5raqLdAiU1UZG9E3pko81TWlpZPszm0i6hZCzMYj9L5nH10pKHKLvDeRgvRiA5SD
acpZ+nlkyRUtPfLOlP3W5L0jMI9vxyvLYPeZ3RmExA1i97sZ9/Q9gOBaKuioNrO3
VzpswFb61Wq/BJoXOcIflg1Y/pdx/RCEzxXSvbj8ldfC6thihg/K0SL1nyleFNrh
0DuI/FQ/Zj4gJK9SMbylf5OqpLqOM1kCo1J+l0sol6JsTO+g7MNdtR8ZZpGz1FQY
BZuA3YrkacRvW2sk330HqpRc1DCdSIaBDYVy3jDvQsoNpNXl6/O/Jeq4hQUuODbs
nGhy1YmqZ9rATDCjkvGqCHCuE4SHNaoCvUysFX0ENDV1EX03ZDKvedIcElvLAw2B
bFr++C05vrtQvEu71hVILYf75ZNb91PUnglxnqeHzoZgXEYFy83ArLo0Xkf417Hz
taxXJ4Z/STSi9fv6PqibIy/UziNSQKF86EHNHkii+cYX5WhpoCPs2Nvsj5FykrwD
nh2V2kVumDCx2NuKpN90qv3KZKCAVYkx+n6a0+v5ir/PVldv8pQJkz0yunJbGX7l
SwwC1u9cJzThwcZURhJUNTJFHgx8oIjZXfJee78Z2NH3wVO+y3/hd1GffeM4OttM
pQOoXk9ROyBlA+vGCnFYckC9pE9QMbaAm6qjpMGNgpiUHaeIfANg/H5Dn0vEs0c7
eWbOkEEbTwWkDmem7lqv8YS96kFr84dsPrjZgTm9KRAVFPGMx8SWbWe+TtRPED8Z
dht3cMrLCsJbEHnEkac8Q1dayX05EZBss+HSxbLJsTQ0kqRVW8qDdXqqhCIQhlWD
H5y6Sb3azF8jehukfdoPY6oqXKdgSwLKoRD1l1VPOrHFHgGCy3RoyEfYL6VcwW/c
ypV9ZGUZ9vrx3MjnUlJGdMD6k90y3pFWo4e9GYclmBO6nNZJnzkQDHV/g4pCJo2D
v89AkfZ5UNOpfcjRBimORPWv9hcw92A82COkzg2qBmSzIMEDGyCk1JIenkL65W5p
kz0DfUeNFb7Yn5+djjEgpEPUclk/mKQbW6T3Y0cvcAJje4BM9Koaxg+QuC1JuAvx
ptmOrNxHEeelA/zdVT5HoAR9ThUA/33TMQD2/ZZYcgrztMnN8VqxIOMdgB8WKRvV
+xTVWZt6SoSXhqtDKvk5GUSwqWMkXHQphhRG2a8fOo06HAhgBuXGrk3dmfoujxJ5
XW0e7ljCuDamEoCgzzwuKCnWPVXufgMrgPWJzi8cm2+i4adqAcugeUChGURH+lbN
syth4vpjq55BTRaFC+cg2xfqsGg6Kd0WVB8p8wJingNZNLoBKCmPTFpnQyzZUa2c
Gkvt1DZOJbHQQQ08k2CCNggitWWReW2lYwO+6msbkxObG7wva59OJZ2XWGQ8ANIZ
VRY2JBgcIQQEZU67+hCC9YRCxOJex9IDRlk/wzorVVygPoIQVZAjY4odCvjWV8Yw
RBI3sVOcb/qzmP9IK0sy+KOKxyqOlwAfGkENL//zWGpzJAO1oR0EH7eDJbKyQlQW
zUMj7ftIHif+nnVlA674RWPez3mQAoO1XwFi3AtAr3sIJFrV8atDxeMPu9tm6tOM
6gjC8iEBODGdSVIzK2HRh4QgedciC1wt1uOZ9llZql9mQJsPKHWTjTJF24A8HAwV
sDZTShPrfj0KYFFohAowMOtpce6+MEjRSdb71yYtChJ7Wq3srjPF1Pdc8vyi5oI9
ZUbg1LCv38No87tiScB2khbgIA9Wfy/E0g69llQ47x5J/PnsrQL+Gq1oug9+T68P
AV0tOEJ9JnUY+mN4ZlGXDNEMgbMXSPyWff/LGlZYB9jpzy18/QAcuyvsgtdPS3Dl
h3s11KMsJLHhJu9+b4CbMgjsAlkYE75CtzQnCjMx63MiMB3UwY3b1GpyJE8mYbdD
JVwlhpJpHVMVqDS48u8ViXkA6xngRQrp/B5CIkSvIEgYlHurkpyjGtDdGwCmIOZt
u4vQEVwyJ2Vx5SP4XwTI6mGSokwzdIujouPp0b6zVMoJltEgx+EYeiNi1EWr25Nf
GsG7Wuwlui9NF0X7y2PCAYilQBxwaZ51g+QUfYfXYnQCSECukVRiwdi9iS0benhT
1E0rnwSUgXjEK7R8LblUtBrY25mPbVTdlL13HCbuSYeFitoUL5yHiZI9Mg/JsQvG
Hsbcu9VfVaJRT5bkRvv3KHA95JIFFtK2kArSRgNZLQxkpkrEudhTND38t83FpuEd
wbfizqGRi1aqxIoQB7PJN3GhS6ODoB6szspH7Jfuj3WpvDA8DFT6GZULsKxPwN9N
EYG1xLTNuFqDx5MaAC+6fcYkrLC4x1DPuTvE1gycecIw9xgDj4VADjr8l2Bou1q5
PaYdu1lALRxNmAV8vn7fdJWStaGTPvS1bSudTDXGODLEI9n1ouCHGz5EPRgaB1kj
BSFc/cpRD3/JLH0xqWOUj+r00Kt3Bcs8gA+GANCYowioRvrdBKPAj+O+6tBTy2Pd
ea5FI933I6PDOcyZW2AqIv6f4UNdWmZ5pIZW4vJ14nfdysCM73tXa1cnmZX8aH8a
sLlatzfavl4s4d7CFMiALTQPE3u10g8Vgdy3bcIlZcqjajbT2sa/k+91fgbzjd0+
x3lGWStuWIIG7g2jPGwS6v7kzfjBoDgZTqBbnFNvVInDcQh5weqlPWJu5pcsPHF4
s6KJlVqAKcgoH9nm7r7wy77arpvyyTpxxMUsFhhQtk7nsnx72JQavOoblUywJjc0
1STPk1Rk2Wv2QsQSpHlPCpk3cGyaxwdYDVM1xQWNqAmZ3vXe8DaAe7W8L7sPM5j6
km6JBrbuUDwBINwHGiOYc5QPj862IpBAdbeRiWvplblhIe30rDxI7M7bLITrCZvk
CHCz1dnettUCrQKX7vSQ8tCku19zGimr2kpXKLnprpN0FOQASPio3OaBF+++wKDh
s0tqNgvK10wd7LTZ0x2OsXwazCJIe8iSqy6ypfeGcJRflSG92+UmKj6df6g49DC4
gdtayXDBENoFlNGnKul9oXW/kTTaR3a/yWpZ0zRwot6eMzzi5phlPNJ6KTIqcRgF
WhUuWWmyP/7EhFSE02F8DuH5d4rUiaxuTCUcYjYJFRFpC1r6d/es90JeYkNajpjS
66M2QJtIyKxdNvFAGZENjZ2El+x0B7jNsVeF4DFKJXxzQf1v/IqQOdH5zjIBx+Sp
vKrhHW9gjyoAFgFGewaUemwEY7y2E8wDFTpy8PXZ1MznqtxWOKR7jNVLVYN1fOKe
OXy0AismsUU0+cJZBNC+UAWZWCbCSt88JsiLLw6TwFaOnGgAz+VOuLnvLHUqFQAR
PlTASMiXKvxbi1oeahwmBm7hOp+DVX/YN9iloZlbh6mzBfVTb1oiheBrqheq6f1W
x5H8l1s28EViI/FefAgT1IqG6FfQ1TWL17qNoS0Ny2k1WLC2YtExWC60T/M5qmRx
98sQouLaedL4nrr/G0s3Vdg9sUhTcDx1KeMRsA/C/pGQAfByjf04mBMkhMDc/sst
yg7f0i5T+++yFFvUKQZGb0cXzNkmXnY3h9bxeZVW9StPhBozmZ1GQIbMe/FVJkea
WyH0u7p7I8id8X3fkDs+U8c0Uxwdr8LLeuINIWPZOoPMiQRzLBeJrgGIuj4/D8n7
vmmt8EHMyzraQQsM2Lk/h0Hk/tkx0nnYw8TzC1KgZN69xk2tnk953nPQNguesFAU
k/Zbr9JcCmCrTWjtlQd5LTRHAJUzxfft+bWhkQ0C1qhNRsXhnEe7/mThL7LzEDrE
a9qYiukq37tH3cNHRKGoJbD1sSQbIUm/eusM6LcIDBQCWtNmSPFEW8ky0O8Cfigv
C5gfE271HQiEaZjhm+k/UgKBdjfZOdH/mNXg7IANtMf5P4s/WyLq06KJWTErpqlB
AK93hrAMyPh+ATf8fqxnYfhFsy1SmbNc+ZOrb/COXwKSXvvRRDBE/wZPI9O062ij
m32EIsy5DCI7K/5+xS7zIuSId9S8xzrcCc5v3nXlhIxWSDk+XkH7/1k85dgE/b4q
+MwAgs16hebu0cgyxj7jwi6BBd5Ky4DbQxL3XcaQ5CAbl4VSU4sWYUpc0ow1tQHz
RSt7L9rgf4w/fSMZKq/MXd0npgzsOYkIoUZKp9xC1e5CJr8Ae7R2AvLz9yUECscT
44cJRFirpf8L8xeONgkwg9CUDYfujK9pxyqHeUYh8VOxpoyF2Y5PRDGJM++z+zv/
GMGQO/5g2dDuv0rf2IZIe5aSPb9sUNOws7wm2PxDutEfzpxh4xVFRW61T8a2SO6K
qMDKy7XDCj1KFxGQ+qV+kgMNzKm2vRJbjDbxfIUnio2WSyqhFKFvhAtW4GUoA6YK
PtmMfsf6fGxKFdWn3PxtNEyiLu5QhEgfAbSvWlTMHOppxboTaQND4bD3urBjwf2K
m0kqr+bd18smq6oWsTek5854Ht7tmhZNWu2CvbL0KpgL/p8SiUEUDI+ogUBl2djQ
APiPPujhVBEupwsoqxYwsXcAfvocqDt3tNqBquuMrxCUNLTQR4ckxBlzeQ6W3VrD
zZ3dce9MmNJYNzzcic2bCafBsAg+rpak7mDFhOIOw0U3AZsW0Y441VScvAwcc5QB
l8FYyKDcTxZn+IQFjPOducpU5D14Wy1lr/v09WGx1lOM/DS/vmhm/i+KCV6VCfh4
ogCmU5L3l9mdIH2BrbhFApqjutZk9OkC7Zb9o3sDZb0PA2FunJyxXClNxxggaeB3
Bnfuveyf9MCxtiQZBnynUMhkaiJI1psOAni0Qex2X23dcUclzSvCmtVoyAGDFY5R
Nw/gTgfrd2y7UxMZVx6CZB8YbEgDtqK0J9hM8oz3OcUKEp0Hxx5mnZ9Y7akon4Kr
4qcunHUFF0TQ6ygowttztW0J61WEXhLQCJAIJavipSjjCiBA62nU1Xm2FjcDfWXD
3C0C5l/MCEFQOqUDkr5E60e0C1ZVPQxvIJvB8NVBiccsRQxsYunfTVT4UQ0JRsoO
eWSROwfBS/R4CiaIZkd6+AhD4yg98TPAB9ikdR1TuAKue4Zo4LYTkx9pirfPv4iX
3oDYAKo4f5GVfD+JGZY28caHThD+BUYS4Uv22ZqWZh0BcEHtcBdi6OE1kBDAcJj/
AmUYrFqDIY8KFFKsdvx/cBwGB5ncDuTjQIqzNsVbZu/9S41/9aRgybJCbLOAAM9B
5hXleKBmx2fJA2K8z6sXVzjNA24jmcHT5ey1IKLOjEZYjLDoJ6aAsIojN0RWxm/W
0DtjV4xfRQF7sRs+QGRlSfwMWohVOvEO333jZfaWlsT7gQB8wA8tHSC4fvTHP0Fr
V+4UFzXVw6OvfrtKjHVvxN9UksuDaFLgkrXHIGE0QPMGjmq/7IV9azFw6CJ21hy6
VERRI1vohFKyYp40gReZyjjWUhtYINvIT3whMPTkv0y37+RBxCvJa4I51swNCn2O
vmTuMR/a5dmGcXwj7ajduwWmC3xHaOFGXMVztwQ6ZXjNHu2Jz9n2/w9E2qsLwfK8
X7dgBF3nmrDIw8uB82EX7spUb9RLPaER9xMX/0GH6YVLjeE58bOrFBfnb0EFXX5L
/rpiyff6YXhCI9ycCHNs/w/iZIJn2zG7IrWOZhCZKW6Li+X3qTuOJQ7CRUyvEgIJ
AK3dnPtHmuWMmQW7JFIXLwnw5ga8rv8mfkULU0TTSCC/7aMwsC8oMaxoVc/+SbVF
UFtrE24j3UkaxPrOgYuDSKRCBT0wbYo0/G7GfSWNKyQkXM3Ds7xTCXafG++0Iz+6
CY2z2Qb9j+gALPrrFEBldXz1+4WVMeFGZMaFGj/1Oy87lKLoi9MmDUwXoGQIueRS
n/+p7cEp40e09mWBLKzNk9xMu2+0ICzSilgsO3D8SXKF4XkD3x6UgAmGlKnSfTmd
og2ahDaT9LV6nnw5FB0WX5rlwhwCNPb3mhZnvooDw94+BUjuOJDPlKi2LRmwh0tt
KPqlOo+oQVp3CIuJNpxZxdV06iBUkdTCS55KyLQwyMlEjzlYots8NLXyugFZfNke
+djVLzQrdftGSkh87MH5FBvNMR2OxVp3yoeGRSTH0ykytVStHL/yyIHASBHmgTKz
TP+VPo+YEfnspudo/gvDOKU+1jDoWkDm+cL8A98l3clm78vVpVmXNIRUCeKP9o7g
bJLgN4ZLBExEstAwqqVpKYceFiXFRTdgplFduoKC+mlsxLB9ssRB0rU2biWDvw75
BTcf34spOD0WKJ6Kbcj5EMlEi7ePkrA9T9P/vecvZGTuVOnVfkGMCD9TySFpvvXt
ndd+exF/b71rLW5jubVeZXMBNQH19e1xX9lyoCMUZa6ZXqT//79zwZxQdH8bCGcu
7q4RNVqvX0paUs+ss3gGF9SbMtBpG7xc2aPSjWp2gLN9C5ykaO8hARdxcisc7uDW
4hyW47WNdYnKucVspfsW2R2AugEFHlTqUHAMEXvdzN39l0Nknf5aWuaYm7pZREb/
Zvg5dH1t+j4blNqxvbgGacKjnYlUjHrVF0OSbngMjMcVLcN1KRpxOgUSJ9ynqKHt
TGI5VAQhWqRPsLTdCzIZRp32XgcBXltRiDqxUlmK2/GJyWztWDHVt+eXf81v2yTl
KMbFmrOhr6OXigpZqxz6jJUH14/U+JWHyv+mYSzIyyK99DRrcr/5HYE2MYv4fY37
7LdOleApu/7Wvj9bm/ftPMY+c723qVFv8BEHEUszMWrVwgMtfshY+avdbFaZUH2T
+vKQ1LU6cxcwG6zvwywxbhDEx2LCEJoqZvVNmKlh8juTfskkoaWQD0GODXKlyqxM
NKPsGsxm6OF9fQTWGBYqDeCuOSzSYE/QUbskOIt4aw6dRtKKMS1oY3m4Qs1JP/yp
P8v9KsIg5wYDLq7EejnjQXi0auTT+zQvl/f7qpFl4fIX/PkS8VCFBJMpZHKBS170
xzlKuKnAJwoQO6sbeSN/ZCSPlNAF5cHHvQQpaWBf7Ix5EsNoJe66ikA/k4GRjPHn
R+yoS8k6YRYyABXYt+SbqhbKqkLtDQZAQ9777OCMsWZfVIW5gMBHg/DKpuS/DcnU
csJp315uZzLF/ujA/JfG12DzQZvCQzAKdApSmBALFYqzEkp/psScUTFv35L7IvCd
MY+ho1GsZLW/Rx5JJhUaltoaEtHXZ4Oh+wQiWoqYeGlTkvjTL2rvSFZCOicnRkLe
Ho4JnboeUDyrOJNoOaXloyMpoqpfCxErykcBC/BS/LtIFqPxAI0PgMbARfu2Es7Q
brJyrcCJpRRqERJ/9g/Vt6G1jCyXDl8HA+iF3aI7UwRIXM1zW41Qy9biBenuIlH0
SVtfNqyMwuHZ8XvHZuxtWqojFNom7DxLbPktjlCnYmjwe5Ywz9P4Rw9ui8oq0Yuf
hab9gWaepTVN6QHJct63idnXk8Ib9ogK5oN+HfWhIywV2ZRw7eL0fOnXOvyeNCwN
ACK5r1vItDXlGa8iaF5nSheLbf0gGZK08bRtbOqir8ezqNW5wihhYT/xAlVn6ieY
prO2ZvegdmmKoY/CTjAkA3cReeO3fQBEvDQyNFR5nzziGWdQaBoparZJ+jPABZHd
tE+tfoYYfSMmVGkUJkCCYK85B3lXeQ6ccI5sGkkF8vtt6VLgWOaa7QZCVbZIELcW
zSon2HqDQ7V01FDGfPBu/l5QbDfZHGFo9q8sHI/bK3XCnmMCgUW2bZKYSOF4W7Ou
aZTFRhPCBhyHPSNtuwKDIlY3zq5EzvuQevi2iVcDtvIdn5Onn/7lkLceJzniiUB0
ZbKbN0C5HR+X1RokpAx7v5MVanSdJW34xgWZ+9Tnq9qtWPwmCl24iDSav7arKekK
j2mvMbFumWwYW/XR2XOapzzJo6bxx2chnbnvRMJmR5PllbO5p20JCJL/UpWj2Zy2
QnCH9kPsP+nio9aV52Bg+/aNszPNN1ram7WpIVW/Hziow1uggZdTE347kGYQiTNn
tEJLJ7peW39Mc3KMq1qCWLNBCa2t1cNhBy48Fv4EfZWA7RLU4XpBiVye7upMfIPr
CNcHB2o7d/1pIF3Iq5Rb2fS9uXxCTgVxfUhowgQFVdLLA3djyF7YYc4T/eRZdvkm
Z4Y/2jXZTY0Y8+66Zewo5QdyWi7ThJ8LwAlAYuzbHAP/fYR8mCac3XmrE3DXQlbH
wtX2Q5YTjyQDOmhL5egkdZg6P3KGBqSttlcyLj0dBsGdwFz5oR3eSO6jZoUrwDlU
JeiVKwFDKNs+H/PTQb5L7bcBjmD7Jro9vkKvxhjFYhTlh6N5xL1HYQpsx5O/NE/F
5OOU/kfujiWFiWtYmwfrbiuNOLFa3reXRtXWKut5D2g+cHPYh0Hmi2ln8aVC8Jjx
MgkocO6EDObOA/gL3aJGQD+ZhNTzNwsrZN9xXdhKI/6Umm4Pp2jKencI6d6tY+aJ
+KKqwvWWL60ytCgdo3a+//ejIzD4r3KhWEpKo71oUZH/r/qY9TZSHKGqbJIjd+3h
g6QSp/Pi4t53KKkFNoYmdPLTXrod+2jKa6VnUVm+zawAnKs5r5ZztDfJEJ6FZoVk
IKiIkSHOoqbwoM4BbVi21J8kqQ6AmiX4hPPtxNd0nVlzadt00rjtcIGReNh9y0Q3
iOHq1/KdJcVfqvBSGT+DSdsKPemOREBW7CKpKp7yhOEI6XCfQzUXcxDbCF9PmFSb
krpiEZjkVbue3XlZmEzUYb+7bheQzVERqiEhlEr16Oig3aQVFh7T9pz5WDZVwtOJ
3eRIEBbx9n7fbzqfZVw4eEl1nDq1rX09jS5SgD80QnzJ16yEQdshUotb43O4AIba
1/Id0jyMdEn152OE+ZuPyo0zK4TDpmHeZBhcCJj+1t2cHSn7l2acUtQqLOKMcUqa
ovL6nSyM0JAwSuQPegRDzOzlKMw+C/09IwN8qZIMndjtNwYylChKE6f++g/U7wBE
60kqMN8blju77hA4ed/DZo3KWqDDHjddH34kqqTmXSpfPGcGc4NrYLwev6D6KU0R
/gb3zY7iG6EGgwrcc15f9Jo/lyMxCWvPSnYMQRzJmNNPn0cU8r2H4Q+31C/lzK8V
lm6dQaaF/TqJ57SadMi0zKH2ue0M5UObQIR4++I1RBbGigTrqEt5ErqoYhMkRtp+
yaKkIXrGel+DnU4o5FSvOwZq6nKJ3ei/QXJ03iAJ+JPilsQ+uUky6nz2b7lIzH6A
bglcALM5Lk2iU5brdcXvr9DeEDMfDGTe+HIaG3r/dcPo33vO45NyaDqZLaEkHs+T
kaSwwT3+ekBDZaRa8e+jRNOE2za3GvGTe0ds8+/FRhNH/2BpkLzOvK+0zOBy11U6
zcnvEBjrYRVgkSs8voRy+ujmYWWJkp16o+p2wzE5lwqRdPxCrS7139QNU3L1S5Y3
kFAXa2R/65IBOT7K4ULmympZL0RNvahTXIBPMb+xWHzBrdb4Y12YHfBQhvovrgp7
zmJ8EhPlrCUrjk7d1HTbAo2023ZZxBb1V8mMdCVbjOKFlPZvzh7/LkGSP5QvbAbW
AHw7BVuw7SEDrXCioH4UUsy+F3S0zc5l+OvEzwcBz68mf7xz/5v5idbDSVuBYtCZ
JNYrS4ps6aHJK/Gz4AH2X+krQebp2HoLqndwDXjzDTc65Z+N1LhLFkhTidbK7Wli
VJ9IUT77YchcwSQ5i0WcpnZU9nvshO3nZdM33qDBm8dn0ig6eJLM3RwbHJKiFTVz
NioEEIHEi62oI8iCU8akjwKbpCaBBTJvSUACkrNI7kMlWxB0+dTLDwGmQifLy9/p
Y/S6mIEGMsp79OO46+4wAvYYUyaIfg0TsAAmamG01uzIV5KyANujilOnsNCSOc9a
mAWOeyFHa2+FhDirhlCuwC9nUyTgH8WIUIslsBvYQHZLdcka6JsND5VYOKseXi/w
th05FNay3XBViHlRXdlxGWyknF2OUPPxXbpQ4/1eTrGu2VmsRvrQLeyHekbIX6UQ
3wXPIvAKnxfVBYmlFuFhztXBIDdOMc/lj7QMB+ZSQv1rs8fVK6UqusfzKYntPIvd
isDnhzejBIARMtGfsdH4x4H2mQqtmf9hz+48wX+NCfMgZAiIgX+YbKzvAvby1fpo
/q5AEPPPZJoDmB34F8/dytQPkslpxidveOiMspnYvfL9hxQqprE0e3z1GR8+aM/A
7MX+ST+3vbCv1BU5BETHnNmQ1AdcTJcCb/idcjWrEty9NEhhdo/c6+nRx4EbsBhe
QsV337ReI32MjxXkZ3P1yaNBxeSoVdbQOID3ufw/vcbvm6IZ6mewAzKC2LMPbQnl
MGTXlUb9r9N+V3HrPUevAMCL9TlF/hvh8M+En5FQq/BA5u4GojkOgiqjLVAZWClA
+fvykI9iadis1TOj6FIrly6BJVVGVUkp8hcM+48D98wrO/0T13rfPk9IHHnsyTap
k82qPG0dOC7Km2xYWpid+pchhGfS91dx96edXRhsIAhYqpUfB91s7Ws3H+wNOTW+
kermV5jemMJanvXU5u5Vi1gYfC21yVQhyFrmG0KCU+gmgUlKyqjIE7+pVHZhKkfM
HYLTQFSbryNKR22UYXFa2R5HoJDAVWnn6fXS1X2KEUwTMamj5e7/IZvWXHBZLLQo
3CRemwbvH/cEFXEU1a8ISYP5VCbP4Dthzgr06UXBPmT3A3lDqmkwBVyr/Efk6p3C
uCAHyfkYQxQixJcVn2CCS13c8/c9vYp+ARG71VsT/PNS6nMpWhrN92JIivh8H/vD
xjBFJcBc+VuoaWjveI67h/QY4QS5TJJc7pMQZf1/JwQB3tW1JNx+HrWXdJTmyj7p
Y1BIBOuyl5HXKuLIWn9C2jeNmRgkgjgn+YEo/s2BgyPmwQKabsMwc4sjc3+C5Iuf
d80qwdRueh6MA1lJhS0PVe1suU3UwREvWM5ZyZ9+fv+TPTgnxyNuB1iBTX2fByVQ
+xeE339HmeX/AsIdWNpSu0zfO9eWAwDsJMQmRtjtTE0JR1wxYUm5hJe5SXvxSpsI
JXeaOA0QzzENlXxdOEVX2RqPkb0wQEtF76psL3KHE3Y2v62YMYy2PJ+Q4Q7+dq4u
x/xETFYulWBLUtvo5bDACSpp7Fm419F1UmjubotWXKuWx18gT8JPCgw28iNhxMKj
onOzMPb/TjH+Jf25enB4usPwM1YqdyJYPC75yBWDE5s3s1d62B60VkbW9Sga5hq7
Rh832ycwCCP4lzvOpJ9KSoWHVIC/DnDABuSRkuB3sjpfa7g5f5hCfQn9RnYMsVmz
7Jm+4B4Sdu/AOp2sVZ7wSD5gtICInIrXm13BCAbZm2axVA6XvvBdfqC20rgfZ4fF
v+duB/WNpQ6iagfj4mdogfu7RuBekWt/5JKeHwiX93YGcBxGg7y8Az5fhCU2RJyu
1DOOjXzvxt+Xt23BtsHQnp19ar5wDWLUYsFc/b8wqukjKHN+bwEu/TbQEj3op/ja
e06GJ3m6v06G+91HgYRnyy1N0F47gSz42SwcQlKeteF1Xzjz194kd5M3yA/SH2kC
s6CVa+kqtKEuUMOeZrUZmUjxNA6NAq3Nf419HRXhQud8Uh+/MfKlVbrJY5/QpZjn
GB7NfBHjCdQylR5yFBMc0VyZekkF4Qtvy0EZA9A2UDJWVE/qXLgRTV84hlurIcIt
yvTqa50rX0Y4PbT+Q/raJAupzFc8O1WSfr+v0qZm/cEnnTRDDfKI+fuGG9H4xnuH
u5o/1Zz7T0oDqhel8/rhxeF+Kt198aROPMwm8o/u94VSjsc3fBbkLkCFwPkqM4Vy
C5s+atAJs1axanQR9M1zjLR4/1X7eUuvLO7H0yqVQtuy0epVSMo8jT6TQi40SQX0
2ei3+avy0WxOFzqDdMeIdnSw4q2kZ0rpxeiPCIuX7tcdlwkOxOIlXryyUZ/yMN91
GD0kiJpfeYH+3AgWOz3wZji/1c+tZNmUFtiryKwKR0zySMMOmk7H81dVD0pCAfKZ
OKRxqaqP01Gq869zSCSKoAg99VonzdA2uQeqWSrWduzm3IQors5Ul5Dbdu3j05EE
KMcOag4tmLz5ZKcBiYKJhbbaQ4kvc1o+VRj2vRpmlBy5/EKNIVH5KKcIiUBWrfYi
abKfxggxzaKDHqNUvkpnIqQAJDQYpFrNTrfFdz22OR+obzYJ5U3pLSZnDOv4NxKO
1VnSPxQBoZJYeIKkW75IlRM1hBtNGOx2/oFTppSWSJ0wf6JjbbYyv+FgV0oH9wFG
G6AN5IG6tNUTst0Bm47s+UaZxuj996FngD3NiX0yk9sKljdTsqsJW4L7FA9uvScf
qPxpUuKO0Ayz70DcJ3YFcNRnNPmmo9WEiqXq53/Myb+wX1lrrXfMViqLlMaX/Nl2
rLeDR66BOHys+YTF9fA+yMNSVzKALljGLRZ2oHl5MOgc+/DiIIFlq4qnMNcwiJ1b
UiuoCWtNoTaHfaYGjF+fhNN08DsOzxqnFtMZXbapxX2jH818cYf07xFkBClHYQZ5
ooVpTGExDnafV0Od/qA10Td7y4aNI1SV6yhLx1A3YlmkRJtdfutdU40Ngzu3RMBH
RPJAqRTi0/Lpo79JPwKRs1nEL0nhABV2bZpIXI346EuKIPRrnCkR+QVtEVafv9Bd
tSX9DyDnmbcphQqiBKOWlJrzyKYHsXP9b5DbGUd1vFFd8gHOhbzIJM9Oenm94Koj
pBu+SMHktrNZO1DkB8BEbxHRJEJdFdSzm6c9moIiXl/grIL1o95EePh00hQL9v96
EuGXjLYUVCGRXbrWLXxOTvk7kTXzpwXhIY/gjqlOZbLR4VWLDwa20g2oLierbx2V
UQu1SC3M4UKfCaf2LeQyic3+aQu3alnvJpdH3r92WdFGqyfkQd86rgCapAh+/cZF
ABB3QfHcN/bNjd2aouAFZVC3l9gOp0Y6GDvQTi4Tsp1AyuUhtZiOp6F0sMY4Qe0y
HARG/tcS0ZfmUOEviJ6eD5M4HkBZ/QrwDBK32B3cRU17QFZtiHmr4+j0zJalbRWN
mA9cNIRksE3SSOjVuXTBuNm7/36MS61GNeBAgXLWMWWtqybSvCd5St0bRHJZqTxN
UqhYS2a2rGb/N9NYzK3fHk4LsVHS0mZgSc7Xf4NwmiXsT2joTRQEIE450H6ve8ME
YcR8saEdNeP/IO5/ap1y9g8lVN8WtDbbXqEz1O+NX1jgpCcbvRYwab6wnYRILqsK
efCAQTlfGoQvSAX0mh0UYtLfLpbYkmo73HDb8L47vUnmufSDhsX1zVSip2x6pdBC
ZsKzqBbfOExd8UKerjFvvo0yG4Ry/TLPApTkaa4UaHqdi556VeJbzHBRAlOPlfQR
ioOevmrKwLqwdE9Koli9g4x4dDVrRfcZTT1cgDjarNn6kUcMXw/i+7b+3X6skzl6
P5X/lWHIqMPdxu8Ssy6sCgULR8XmBC4CdNgnpGY0sYmzseK2E1swX79Z+ScUPmq1
xIabakjEKxKZ3/K0VxLak+Z2BG68Z/fXLWDx58c8tgYSHpOoVvRCfXQbU2C8AW/0
i3cZkBWhLq6GDZXdtiV8C0XOhsHBiGLBeX79TF51aiimBjN72v35t+BLu04SyMzV
RX2H3D8zR6wIShSmyuNCaiuFbZPJzSd1SfT1RUQMPRJsMcD/osxnadND56XcKiO2
7fsb4HcfcNMVS5eFcwDwsI3ayu/w+IsK8k9H55LTC33uX12xdFJRRXRuScwstpfk
gPk0Vav1lvkdLW/BszGKOaO2KOB7zcUtlHSK9tJfLdt/DekvEXqtzLs2eRonp437
9sPEqWNDJvkXSJ7cWGEX/7bgwW0OnCXCCjwIvyOegUQCls02lMOgh8uWx2sD93jj
S9hPVhmx5ThdovE+M4fyHxafOhccj/bFxyDwkLP7DvGVwNPAME996xLwEpFVNLE8
5lexj2Y4C/BJjqI7dnGWupOcjMedw0GgyejyF+eXKKT4JccGMa6gCSYHt2bRRQNv
yXFwEUSzswvq4/CE7g4GdubB4R3iBNWstS7ska8FwIoEnvGM0ioYBXFTX2Ufrosz
MzkgA5Q7iUPB4iknk3VcXRGXYUyJMij+3P6EPqMUYOLKdPWihwGYgwNVN0i4osp9
tp2eAyv6ixkQrzkrb/ovTokR/v6tfN1OEAUAJQUJsPiykx5MY9ZxBwpblDBZvQ4s
jfD42hamJxzIvfuXBxHp1J6hfQ73Sd4mUzMRcdRi4gQQWGPfIKLiHSP8UUJGnmoS
+t8cYdk67hQbq1XoopVWlpEDThULiFi1nBeVjE7e8twAUwnLluEvY2KkyFoylDFu
JdhEyhHfTx/4nD6miK3JMcfLD9gdX1EW21cWQAIyxWhjDOnHay5o5knXJGeifC6I
WrWnuuzc0SJZcZTqGkg16+vuP2iOdnnXjREWInwJSkYOpwUR36IvtJEE7yb3npdh
OddoZiCjppiBkDs6CJU1+raPDHH50JXJhVqj5s9XGOSCXmVgdfonI7gjD5gmw0UJ
TCpxAFA4HLZ4+z60MuLK4rN19qkx49tj0s/0f6PL+S10Ii/YJpX81dfkl2cjLyYn
7GPPBkiB36RcjZ4BnAYn0pCuVw70TURq/QmZsIXlqhnhtcU6Jt2ZSzG9c9rH7rZ4
AkygPJYuM3qluJDVxCKb2IAEdDU3H1R2FGBfcxx/oogHc9LKnTO78DF4REyL2l8r
4vR0+pd0Wwiv4w5swLrGVoIzcHKc6XSBhgohIf50K5yMmQ5BE5JTKnf6VsEPvhG1
dXbAc90bOEQF5h6FsCaqAppb33IyhQ2qu3nLLbl2dSZO5nLsMs8Ny+WjpPD4kDnq
W+qLofBoIOWAfrz6uhcY7KfgwbUrDoDmC5Rnvwgh4lsK2DbTfKiCT2xh/dqXmBu4
3gaWaYro4SaSp2fBWVJ0Sn5UgJyL6TMMCBZqBnNTG5kuNldmg4VvZ3QLpHqpCy6P
8OIuByO2sbxd7hiznJK6Tr1G7wd4t69g31jt70UWlIZ3gPIjtDIpGAND1v0h9zdv
nK2fV4UdeppL9I/96w/aQka2+Z+iNDNqVoCDUSlfoi5Yj9a2/Ffstr5Nbq+j2b8c
/sv0AYqyrtt397Bb04Dj88cRhNmwexr/wMGtocruWMpgY74/z1Q6ByQAdmcRkJVb
zdjCt304rrp9SozuEVThLho8nLcbKPuukqugzFr5wUiG+fwEhfY3Dy/gfi9TbwXf
nfM3ayGJ9E/PS7CAgCN86EEaDSzqUrLK+FDugmlMiccvbF/qkwgv/1OXO9IFV+ki
E6AvdE6sgiHcXv4Zp5v1wSxGIHRNG6fwXEoexxBa+NmjONBFxtHPlc0cl3QgaFoW
+lFfU9k6c5BgDxHypN/pbsirUXK7ze1dTAE09qZOv7EW+WV5vCAE2fPcwYEplG4c
FWxyZqWFLIkvfc2zwi4azYtwCGGS5oYbHzwfvPeACpHwQcRpb/JzZTGDSzpA1AFr
NhcH2DDOpV0ybDt95Msf2tQXtLKGfQlQeUmRsaqDjZPEU5AK/xN72d0KeNjRHJGo
im5N1uKktGyMWmzddrtDUcwB4Bd3tnrvKq9xfiyJQxd6dcDq9wDRIF3WOWt9vNA2
231WuVKU+kbjTxth8OSCBWLbAQwNcBVpy/A1tgrp8Tq6D4AV9Ighd/2v37OjX7V1
xYC/3MiYSFQwMnPBguAemzN2GdkUIrUMnGgBU44XsEe0Xrdx1ptTMRnpMh/HYgSp
zEOMSNJXf0Pp4qKE65mIXUx+N88NqRTjzgfBxkllanA9r6XBVFLasFD5V+5qy+s6
XTuwaU+Zy7KjLAcDZaBwc/2Aq6jHdTb+e7ksFIl//yQ=
`pragma protect end_protected
