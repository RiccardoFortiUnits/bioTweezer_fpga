`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dg2o3hEQV8p3IEpgzlr6R192K0/sGEKN18NbMDaUcHnRFg+AycoG2FshZKwy9ZGo
z5FvXEsiFeaKEwRFWmpEip/gDLN+E2eeHt8PMzbxDWpPIrm31M8nDCZtmZytdeBp
4zzrtERQ+4EFn7Zekrg8R/nREyaNLctqTqPqm8eaOr0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
IYjIZhlcNTnDz0gFydA/1kei8oRRXu3GnTRYxG4ohsAQdDB/H47UB+EEJopEPMEx
TJohR2vyNnYE5LskG1KzuFjx+rjtQYsVZfVrpKWsNLFYqBc50sV/YzF85HhoVuNh
v7S7vRgaqjKKAP531cwXUN/9yXepMCbrIiKVqiHoU2VKNVZFiXY6NqvKLKhn2elq
I3WUs/BHWHNI8VW0OYnGuJlxMcta7VUi6D9W5YRQR9Y14/SEYFL6tWcarqa98Qfj
GqmR8xvOKb07allhamuseAOefE7MUpENuWmQRzAL551+1yC2cITCcY5rxsYJoa9P
jtKiGlPh8sm4xXbKXGzDV1h6upzZG0AS6+oybspsJ6MnFpTl+MlZC0ZvOMviyz3C
sndMr5sPpQhg+0+feQuIeEmTrkZfFC9AfGNdm+54rBDtUQAtO7EF/XfyTCCozk0L
8owYowG+1kaWftEGw05fhlgw1V874SpDwi+fixtNlh9ATcFVdCTR8fsftSRc4qkZ
dRROgvG8T3TNyILsU6DvQUqwoLSdr33gdo3pw+qtyHmLYQar52osxfb1TfVJLxD8
m6FPvdTFZUKb9TYpxVJQwhuxEbiMsZn+/vYpCRZKklAEu/PIBUNZRYhuaBZ69rV4
yfe4WhysvjvgEZMtaQ1Ss02YilGVvEV2JeL1HRGGUznLbQpfdxGyNL6P/EX9qPMA
2OBIhZa0tKy9y7wAMtHLPNnpp2S9IhulAFp/O1CeEp0oAhhzQkzHRFx7WaFFR40O
SUZICUqf5m+2ueDh/fQwQytuuyKP58zy4dWGKb5uZ2VKa83pKuMtA7KuCUMdzDnr
QZqzexAJBS5FbnssnEIKD6th1MDsv6NQoasa6Grm7Ii6y7w76HfgHx+D/rzopTzf
TVUodcNJ19oYtPj7Q1zep0WPGSQn2q/DlPz2VojHcGrhF7iPR8EDO2Wgy7SACGFU
EXlouYy+qT2GC3uxRC75Sy81iXPpUoc+dXlRHAJK97gW2QxZlDG6xoq6wpSEGcV1
I8q+KYnY6d/kIZE/6ZNy9pGtAYlPh9h/jnQ6fPiYANF55JoWqgSGlnrJwu69M1Oo
8QkaVjeqSUKus331qxr19D93v3UD6MHo4tixs34zh5jmcljvxSHCF0Isuoots/KS
FlMLelTMrGvVVM2g5tfYFLmbzsTE4lJJYIN11uf9kFjcLVAD+ZicEnyQwubA/Keu
UG5Pdz7B3Li5CTiGbuPdTBbf9pSFCB6juWdQU4/+VtsrCzQj7s0nyTTmQufQ9iTS
Zmt5x10Bsy553XsGGaHT73bcRpf9HugKLe8H/FmaMZCvk4fkcsGx4H93fyYdkr1o
MegfzjtGZmI+EvN+I6oteeV7NlJHwcRrkEqSSxmVcVEwuTa2+w35pzvVk44xnzqv
KmaGkcZrza9HsMq8CmxDpkZJZh7utR7lsq0TI64mdhKXqqA1J14c9FPQN57w/02y
HdQefZw2pgXVBqtGpvfVJ5N5OmPUNSeJ4Z1k3Lk5Lbww+NAjnx8cnUbcxqCrX7FM
EkrGVElaW6wGcCSf2Xh5b1kFueYGsmGMPaifdGbCxf0KEs6iu7YAidmmty8Hu6Zi
mbCBYCkcXPfOZWh7w+vi0MOP17C1CcTA8kv1H4evpCO6UT+AwLg0RVV5E9h+MVUL
J2XMiYOX8auxoQBArGHLqFYWAYPkBTHmjEokTkz2up98Onx09RvVFUtgKoWGjcGt
YwdOALtU48rqKmovwm1k5gXc4j/k7alWMP9KrEmIFH5Md/H8HuN3d+uZC082Rp5E
oqROvn+qis9pEHvsXd+QoJVXPSciuGfbOXfFvYzCKbGqD4jArKl/kj8RLVI6NqH9
uJi8SrV/DccT8bMQ35F6FAbTgofMD+r2VltSm8xyVEdOncnpD3QZFeXKl4qb94P8
O19oWXMcmm7JUbzR78sKQOwV0gPBxlpjnJ9dhtRW+LSWzSGIZvDZkPhheqW9AUef
RXv3b/SWtUJjHftNr6p5YOd22ryKuO7R6HaAicHBZJIHCxxKRWRpGaCHoOtQGp2f
W/KfO3Vka3GjTOgo5oHeJYuCBa3HfKv1SJ7tAUG9prJeKeIrJHPxA/kLWHj/LRom
7ItQwGLTZJu4qRYSwMV5xPJkutSg54ULZpqKoiwJdKNZwuYLvnlcFxSgg6uXIbs4
9R6j499/JYRj1+QH0BAOVyWtYnBjyVR6UiKlf+N2K+hlNoYlU89bOU/wnChvUM60
pXgMHokw2YaPEsVAB6LC0IaKksJUlvWsjhm+PvPfaWjIMF4B2kDSdfYSsj0f7i8m
9F94QT+0Fv1Fc4F2HMeBtFho4jDVbIyJHseL1TkPSXXkyn4oTwEfviNp4NUQDe27
mTi1tll1TCvVG8R81tqQnBKNYNisf7SVeRwnf87xXUACo0do0RogzXW0vd+cYpMF
DWrEMZ2fay3G72jJBpTEIHFR9CrmwCZoRuU6jg6vxZEkYofMx7SeGEZFKguHMkCr
Sq6Vg2EsDau2Yv8sCtDjP0GiGVCJwNjj8SOiVY1HpNz5eF4Koa0nYh6oBKclCV15
+Ls3/YelCX6/cULrCE/cJFnkVca3OtOMZ1pccEiBXjZTrHbmC0cVTeDz1Sx1JrUH
MOwIS/FZwNDkJXBrjJ5P6QExWKp6gDtXKV6/NxNvqrvH9lHIP0zzvmvFFCgU2+B8
AbyKcLBUpScTZUXjcO+rVz+gSMLM8wOumVdmX5ndNQFm809Q9FNlsGqUbbkC6CIq
m579lVzJmeAjeyI4J1tTfYlII8rjaoLXqsXW1ATPc515uNALCK1Ql5Ks2OdyIy8r
ET/U1LY2rvAoukDk/AIc1hqh4GgDo30m+rswj5lc7pgLLIPx9z6d8V07oKaTXQfc
UyJy6C22lfdxuoRg2f0ER7JmuQYyBirPNPwnRd0ZNHqF49zytX813Xz+VmGe2YEU
wTxphbdkUTdMa7/g4op4CohExBhN6tFZIqQmP4XZsNlw0sCpjc1qVFOb9qVOBI2q
Nvi/4lukbs6bM2lsQ9rSsZ5GBuAYk8HHqpbsRY0jd4RzOA1Qe/SYTMbo03BWkEzn
/o34FRrRizN2gDRjLplPM/OiV9dHEOZqre+bE8oH1NtnBSJ0h4QtCM4rIaVa9xLu
1dhEKIOemTNM3M1pWsGv4bzn8fXfw7UE346ISINPDusvloSVVRfd4KDrS33Avi+4
0vlQyvmYJb0XoaB8UOWE18DWYxGIRF6qUq2tPYZyv53/00oM2F4KgN3HeKRYVwl8
KASNY8B6BXoaPG69EldwheDCvSVwOaE/eDzAvPUoWgiQF/UoFXF6uKl2yPLFlLjC
YnETvoVZT6czI8swPBBhCLLmrHBeWw/5o4Egiq6H+401X7Mfh1dHr5kk0/XGTneU
X8Rg8uEk2e2M5JrmHWz9CK90b/Znlx7lM0oMj1vAMOHwwebuOAhGrK8V6s085i7R
g8TpBO9X8Y/Bh4SPOib+AZhTKZMBSVhK7yQutPMBNWhXT9LfOlkHrYx/zy7AtRHc
/72q0OPZl53id54kzAGLY46VzjFkoxR17/DUab8SwBprSFPYAlJ4B55q/RAr7vft
XQqcGKTkYoC1LYfu5YTpc3qP4Wvs78IFuU+029AbAfYOPEGqVQEHflNm/NeeCrrD
NXGhVx6J4PIGCQdToTEEK0jDAKD6tPlGcIRK58QOARaW0/+hNQphyD9wQoDNT8bS
sVxRIidXNSDmyAZtK5W1yTBueyD4K9f72tL36bTelVI+yNpnxUHDnlqrI4WxzNhO
xmItCQXmy9Hz3O/hURPjUellCzUZsTljaQVkpakk8L2p8FC3WEWyramdFRtMpCuy
BTdKWPanua2jlyXUvzDYPTlK/zirBM0jTFJtKncpvfScape1kw1W6N6EpXcLe26x
94QnWGWGTJ5hgKx3h/PpvEE/EIkn83IueT7abL+KnolKZy+UbquSm6gIZgd0mbHe
3tRbhV+BrvS++CDhV266vw754dOWKNgjX8QLodWa38rl9TYqIPFfYkVEJyEDeY1+
R/2JPvb3WIrY8uZadOifdA==
`pragma protect end_protected
