`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
thHzM6uo8aF8pUcqYej5RBw8kcL8af/vyLCZkW8yba5WB2MIkM4rRQmw20nkNN/C
lqjHSjy2KPQYSdesmIP2GIJBgcV9cntq4HvdW9kX6qvsbC6M0j3+ydvoj6+mFge8
EMpEjV0z12B1K//nBEfpA098r6gQUsqzK7IM4JD1WZc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
E2KtU/PIv7jIe+Ep6/k4jRnLXMPW+WmRB7+ZSx59iuq4qb20uJpENU77iw+B4lep
KV6JdaPfcDXn0UMYVbn5HI8onj16V2fX7AlkQ8ytXbufSHAnV4bQKqoob7Sdr7lH
aajEPIUXvBW/GIk6RQq08YknFnbt5kEIKY6U9g3cLkmlIa6/EtD8eUwfTMyDXgdr
BW6X6noILxgPGXw4qsUJ9+W4MeLQtYPmzzBbTZKST4y+solQx3U/1+V1lJ8rmoYx
YwREK9G0Y1eC9zOrwKEZfEjTTwJhJ9wMttPXKgwBDEzkXinD6sjFB1FTMrqGxHek
EEdLIjKj353NjRFdTLYXrMFs+s7qsGhW+dN8jxd9Io7GPJiAcXDxglegLhyshVx6
B6ffX15mDbkSwVe8nDYU1tWZ0Ng4mAlNakBxfF2OysOF3eA/paECi8GNCqoBHOqt
fg7swNouX+KP6FGd6iFfy9TyGDtY24Mlqq1+VWXXbu1ilQze09fwFVeN2LJ0RJV1
9JbvmpsRvB2MGSrmOLXa1Wl3Ud9DrhzQXfCRuzPKSiZp4GGMTFStcC5jlP3UPLc9
hBhk8q+D5FCVq0ciUyc0dkhG3EMx7aYmIupjkG2dDwRaw1sJ9fOZ75iTXlGv/f2v
VIka+qgsN6FTCqH12c1wa0niQmmF1xz/FrYqeBo1rBl67RkwhsRalg6AjkpMJz7A
EnErCcheTEa4WislegJW5d6oJi58hmLhy3UycRSZUibFvh62yo8hldMu3SZNiuoZ
kBID1p3xhMARgDKyeH7iEvrrVQlUeBi6qnvPn4LwYJn53Br1U1r9YRiqTU2yvpoz
Sywd/NQZxp2wG0or3ka/DQcW0nYJsvF1yoW4g5p0IDGYpnLAfT0FEwY9otQAlFSZ
HjDZTa7uRpgvBSY+or8UF+7KyQZo9fU5QXBH6fxtgwAaaWcNuHbPU7lmIU2+22d6
wf0dCWSHXVWoyicBjLg/pSVL3MXyI6XGU/gCPgpB8kPFyHbHTVWrBBkFfCCmjYhC
oeqILVwrDu8P1rwSeUcT/utANp8ki2aQyU9esMCvacxfiQd8OgNaXPR91994gFZx
SEMR1rUm4dkU6sfwCS9ikgqOVPdhE//ILI4cgq6UcG96n7Eckw2pifVOexbcVsRl
cT7h2diTijP0ogaH8Fg5grxfyVuTYWgBVFJKuAun0EJNS0l4r8r8CA+ZPZZJ2eOu
7XtfIAMxNCblfhQh4/afcPff5qzmxxw7jUiDLRSWKUcjiDUn4VIJ9pDICLYEAVea
JnLS9aC+TUq4joormA3hGAGmSWYVNjqXjFL47M3tJdWg4HOHvKqawthQxYnfBTyk
CCmqBTyLNlG0sYgXUyKlRfwnYwD9AKMVAl9FXSq/b0d+PkSuuQxIonHfB9Iybgb3
RRPPsp1PmjZGRaPO1thjhpOTAxhlSpnb9IWdOhNt24rBYy9jAUsmkfP8cQLVxZN8
skVOmIn191Vu1ufsdFDZXJ4JI4PWCrE3gtsVVTZucIr+IsIeZau7Mb1AmY4r4lKQ
eqxOZnBX5C90dgao4ABxA01UURQnt4cvcAWaEy1YHKofAoGSJGSRR1C5MbZ9/t5Z
7GFJAqea1mDOgACfUdcAqJYNJbib5KDrX8+kcgThL6NR/LSvctJytih/Lgu3D24+
IMwdE5L5XbINGgvlI0jTkZTd5YEBYJkG32Qe3akpVx4LvT81r6odJIdDzgoPDWDw
eGKtL2WDl7XXL5Y857/aOseAOeaZflDk9mGvHkj4sDunJkZgPiVEVB7RQVaxRTbM
xbU6ZuD9ZElokExs18BFdqRO8nnlnWa8Ypxh7MFM+s3QwHDHRPzQUw5UoZMwbwyV
ANLP46mHKjSf8y53/b4ecOl0sQZtcGTX7C18wxVXqvg4Lkgi4jhoPH0t7EQOFKs0
1aVcNBDFLkovqm+4HQkhfbYOatRZs1jr375r8qv0Fto86/vUmXVup97pMeRshDAp
KR/SIjlzsKM99yv50S3XAcMQeHGcAdGjVLMXpUMJiwtebOuGjxOWD67iDyWyW3Nk
rj1SO7HWb4ujN5JDuyF9EFU1x/vvWy2H1qnE3m2mvGOm7UmPrXCs9ax6Gzy4o89n
OZZh1pxGX1nti8yJ/sLC371Y57AXHGPR6TdKsw+hHf6zXCiddXlUEWf1Cpf6rFpl
GF6aFA5HYH11/V/2XFsjvfS1U0z77SOPVt9qjIdk1xgEl78D+j965f5oPcB8fd+y
jwNozIbh0o6qnHr4mpLgiLj/5whTebBe7LfZYJ6SNyDs4GoK3pQo1BEnnWAiX2qb
kVz1dGPdQJNrksGQiUEUvmBZL+4M/bkD8zf8F85hbAOvb2x9aVfV4qX/irlwTGoC
I9oyqBZlLfK+aRSLV3Q1qJrREsBstKLqz06rdQUZgy4ZxvX1pW2dWBU3rEScHStd
NZw3i1kQqvAfCOhmab6LIZ4G56GOjna/wZFshr2sG6x0O5VPCxYN5YQNfHNECBxC
hDELzYzRBZLm8Bp+EjmvpgnBcQHpN4hJZky1LC5lTx8ZhNnJZG0+7yVEPZMrdmdN
KOkFNTPLe2bMZg8PpGHckZLYC4isSncWifYEG+kyhPG9vmXcklo3Xv20v/G+rVXT
vOO5JPSCpmNbiTvTRvxsporM5VQUDrjVMqrFPHyluvfJQ9cl6Q96C+ZaiGdIJDP7
1yTEajCeBfF413fm8S5ZV6QPWWFUg+wsV+SqZot7GV1bONpdnuZvdEGQvurN3nW4
opbzwG9CGgkk2NcLS6cO1E1DKMEJHxffO/8gjhmMa9iqItqIfzE3guSWhaX8MlMh
7SZ6wgabSFCcO1G2Knu2GJxkPsYED4lv8rn5JU2TsS8zxCCGByIF9gnodhTw6YwC
yC/5qo3ZYdmb1aDdzYwDDDu3XAmu6Y1VbxsLIKaoce0oWdieiJ9O5oqhz7Ww72mK
ZBgh3K8uovpEYyn8C4lNvCQxeBxW+jg7VPcwbx3XdWPa9+C6PpJyv/vlTzpVcXuq
kLusWA7oKEbBFNDAlG7ZloQo129C/EtkXl349uUD8wdu+yyYqmIYNCUpZpx0kM2g
+JytP0avv2EgInOO9oNMpQPi5hap2pf0/mVVvOYdjtvGxAAL4cizu+iGHHY6xyHz
CI6hTsuuaSqK73S21WeS1mzb22WIbftRdLjcVjv7cvpJY4PWoEMRZIPxjnWuMumx
DsgPbzBc9T0IZRS9+PToQoreDqVKuHbRW51uELRHho/lvCHjtCdLIVx7wqJf2DmB
wCi30nyZ4bQpDA10WAiF5bz6uQTJ6cOET7Ox3d0x6hPskVfvsdGT8TtKTEe7TPog
f91vFL5qIR3ZqzJ4/kBTXLTcbVQxp8rt1RFaV4rZQL7TpEOh+dSNrXQzLTBlCPAc
SHmgKIDK3mBU/MYTitXlCbVmRFQM444iorJxX0zF05SdCDoPteTbvwFTrkfRtlx9
QzqizgFE1NyZsbHg4yyHCDVT+GVgXSj+gXeM4dt6UOzYMvnuuygAd2m2ho9hZKR6
cEmW8diyqI3N4yr5nEFolFmOVBY+X1V9GJMbSDFxY6FnmqF8f8raBmgrZWHnDXwD
L4sCIy96U99FOJfUAHzuaWreCzCibfKtqqBSvS6/+sGwWEcGua/xdMigmsnDhsr0
KtA5TNIU1K10axP30naofixsXtJxti5NuTec6qh2JON4VcMBabiSM4+rcNdkNASe
Tvt1GxVWWpqPhNTqxyG3878gVzHl2gTrgbU5pnJduHWPRq0bRmPaSWP8BNIpgkNV
nbIs0ZxMUpz8upOyM8emQWaAY6DCPKwJ1yRVaXJsszVXhybKF6fTTKdCNKxOH46C
JIIJUJi71w6LE4RUPjO+/1Jwcpxwwv0TCY0EhBtHzlE9Cn4RUtfSDEAcBQna+ymW
kXNWA6g8RQJOPLUyYLdNi7Z32L7Ma/8vXIOZG15XVUuZCtTAF1HWoj8KEg2oLiMo
xVKqBzj8ofuCSf2+yZVoIixwdXcvuUIUkfS+mgH5NFFeOVOy9x6iiwqm39357JY7
KAOAqFs4860m9v/2JZBQEHRpv9Qn7/bU53DuYsCrJ24XtGvNCf7ft9uvaMFbp2kb
77Qfe888GgvEqAItqBgxhDUc57ohObK2mTJejV3KrtZvsOV/EGy8sqKL2ErTD+wq
aL+IiWNZ4CI1UUz98sOHG0K3T+KglpPMovBWd99Wy1e1RlbLZmOR9qEpcLyo3ytz
yTwSHlQGVq18dr+26tLUsOkWLN1CQwFsFqyMToKQQmBN0rYmHPLdjdex129e09We
rIpM2uTKjU9SwBWKeK9KOL7TduDAGk+p0KywUVeZLrPto0UqqsVBofQh6iM6iLuY
mKUbpo0kUw83cCVWvyzFvbdFMm4LHHtQ7kb+DS5jbUeZMEK5hKQJcrn95TvNx1Bo
9Z9WJrUVe4awacAw6ZNJJhR762WZ7/nZmLw7Ysy594PLUzwIYQeQSM85PrMTjI7+
kM0QhLkxYYbHwQzrYr8WejyfFozZAiG98jVOqU+uFRe2IczlutspCXrA3e8jyRvy
09cFrHuQLVd2NOhuz9jgCEsnY9I90MIfVlSxJ6naQvCTUeHalF/H9BqUYCp4rYbN
VriTC1PA9VRlbsHoo5UPxPqlQcYpyCoC5qIHRknXssttV0Wp9196c7qx59J0J9nw
R0cYVLsMQGjQ0eB8nZMJH879Sn7/BUDMEI2dRjePex8ovz02R4l+dxK+V9qaYmI3
BeqGKvRz6i0Wy5xt81YOLOW4VJX3+/LeD18e/tBPLUpL1sAKsjnOq/jrb5fcRFgI
rCyJgKOw5QxfIru7/Cape3JD0PnEN79VqqqNlXTHtEw4aZN1/ns/MGSZuvAaq88x
8R0Q4Bxkyj6t4RJrpCihfs24oneHcfNlJgQICaPajQz2QAVlpoeVDaPfqAwz1hKX
tt/+3z5ONruZVaHgHoImpKKVk3eK1H/X9rTNPbTY4rDnUF9HvmeANEET0YbX9N2j
AmpnvUCih6VEIhVO+UURrvQyU1xtsXm9kX5KvetCUScAfCFaScYyxsthH+G8A+ue
m/IYpFdIsiis7kHGIksjuu0cgooNT9/QIMIKEw167ndsXE+bQW3Naj1rpuC0UGjU
MEWKNP89M5W8GWvaVsfw/LORrvBfqTywbIHasfp67UPeU2pgdaIKBNSAOo7eZy4V
5mUZQs7a4EKtODzqD2w0VKSiFJz4T8bMCOLbe8bp+sgxLDVXKHJszgj5bFIQ4NUd
wRpO0+6+97Wml/xMEqVoD3vz1Zy5W6P7zHnRJ6aOP1mNqqf4GiwBW4tOTOXs7NOn
M82aL8ZSkefpyHEjVTohLvcDqkuNpRpLaIJU7CuRGU2s1Is8RDPDsTgCaAYdByTY
zDEOqRXJOvXPcJdkMoSnvmXjuep8FnFptEFbbHKomYe2hrTtfVkXNfgJFeQTqfyH
B8yDwPK962em2fHQBsnmMz8jmCyP7NYqbK02cWQsJB+JzbPp1frFjk4nco0B2h1T
Y2s86y/46cQ8fQmBAC4uEwWAN+iuurQgSUwDGC4IJgJjXyD1Cj/fKdWz99J7imLb
Q85BoAgtHylSNW2puWhQ87yqdIRseQilrj15OxAbSciQjX/lor8WPx4XDxD3V/w2
n1kx7sYfnyg3HGHSiuq9lfY8WJ6bNY2v4S2BhkMXjUJVvS7Vjw68vUV0AKA8eAEE
59YvsLIm8UlNCxjpUtyuRl/rShgbdYmbbzqBdaTAhDX4/OY4F7gwB5U0t2r2CKC/
hOUghXDhmFYT7ZeqL55yo3jlMtmfsQgPewO/DELJG9WbldaexGWgc9DjdXk7t4Hr
lGEd4nVCeCzOwuCzvcLKHOvlMwKoLc8dMgcllIgM55EswPaQWqHaNIZe+TVqbtTr
Tm0G4EmKGXz7dHriR5/FXClBG0dvrNt0jKYpuc5DhV6TL7bgoI4CeNGPhxHfcP19
3l31fa9bFQ5cPU4h1RTNCZd3cw9dg5MuXWvhiGJu5akTkBJmbhxA1uDRcd6pgmHQ
nrShr7Hjhk0JX7ZS25AVMk9DygfwZrg5a6HIS+2x5SQ1sA9Y9wWAUdVUV6LXQLm/
5hU/qzYZVUhKhA1PBhzWyYgeAIBsqa692du4GaWbmVQpRlmVRt+dKCz1TYqqL8ZS
qd/tRsaNcsjni6BTDzL01ewYQmPLIueG3PMf+kH9ViLSTp4kLzKRrpfpESjQpGLR
Vur/dUaS2nZYyZZTVu9H0XNpEo0Fzlg/dq8CrzLQpjYIs0DaF744OJr7i/KZiLHZ
SDyCS22KjYNL9nxajizQCHLkyn/ME572QXOcVO01kNGpnT0UunKbv11Xod/uWZ9q
qCtg33BmYAIqltSZME6Cik1cCxbyxnicnSq5GzGD8JnqFpUxF8mFOOTy4TTJKpz5
ipdvuQshcSmg1JanfKmezWpcR1/1qD5UaLMsFLXKy8vBVgfN7LlW4uEOkph4BTeL
5ytBrnUHnbguOyZalU463tJeFvSYdBUprgu8OgsyYtfgpYFNypGjwOvwz98c1Lw+
j3WJ0RcgaAD+Xg/JHYO8VkGpaQnH2gOGAb56DHQ3UNgXp2/5WHObN3jyi/S9cxOf
AtNp9eVnNbyJQAcx9AC+AXT53DXb0Pg+rKkfEDai5UmzTrIKCtuU1TZH8gxkCuj7
oQd1Raa0ymwmqgflxHTQzV7yg2Nl4AnBdCtxnt9q4JoEub8PzTmwSGO8lTNFp0S4
hIFEtniIduqnqN8sxvuIUBqe4lt2i8lPcBCFe0IyjwpFhnalh7rqMPpuds5sjZLm
aluubTHTe5dsOhGHPstXAmplNAZY2dmblSz8EEQp6GNfp1/1T3AnHaJ7Ujg4B4qd
iccIx2tWx6ucR4RjdOFUDUlk2I2fWkE9Zurst+IqRK9Q3yrpR6uDEsiGm8mCQKFY
rhQHYJ1Bzd0/BIyvGJzJ9ZnAUFc82jr39k7ryeN2/SMuV2HjWN2ZtyK6mT01eJ2Y
l/WiOxB6t11IdW+ZjHxEEd3ohtx1WtC99NVrpU3UMbMgaH3hOm+heXRoQcNKNi0N
uiXUwU9CbyiuVSooY5oxxUJgaw4iy3qvay0vz3T7iQCNjZVIUkQvqm/86EGbbILH
/NQo5Z49ivtgNKpD4Uaz1WsHsG+kNvuhPxFgBP/asM3oqubP3Z2yW8JIM9Yr1LtU
bWlsc7bFGH/sEHAJFMWmgz3I9w9OYOjR9aHGyq4DWUHTDCK15K0R2fR3HjSM3/aB
HqQ6gsdYnsEfPdFOENRCYpKH6L3elSO93jDd2fOu7muiVG0wcm8IEO1G87/icJRZ
0VMjzymdATRkAlQDrBz6Xgc5Y/Vt5TeF2UX1UZoeJrJwY8mKFy2yFt9IjN3gk244
OVRR+sXjJ2Vc1LsDadORta3dz79wPBHN+vMsCvaQArfuZWM1KcHFdQbsubAbzkGx
FczXdtB8su6Mb+ReCWVg3EWdMK5Ewg/c4Ost78abfn8=
`pragma protect end_protected
