`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MB0Tx9LGisrZkv9g4Lffcn3Lv4mve9QSiHvK0eVHtfB6wTGPTwh68DkIA34WPnsn
xV4tH3z90DZlQL1l3YQqBkWqC/ewKwlhAqVFetFegA9P4yHHoAun0NcV46hY9TWJ
lt2HfeqS4levlldnkPCENQgmJOYyh/LSQAhKbmufOM8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15680)
U9Tm/5FPK53A6bmZCRplbs0EqX4COzTS1GvKLT4yW3B7QSntOPL/l5qZ1GpPMb04
7cnA/+WtC7IyhTr7tZmizfeqXXk/mSGrBjQfJ8MK0CBwizTTiPJeZ+qRFpIxjtI5
GdZNjRDAylJNjmJGtt1A5MhHPnnhleUHf47uXIdRuJUeZjiptf2cbGDO4u3PwT+j
BqId38cI4x6Ke2eUiMayXipJoP+Uv0b4n8GXVzjomMJ0QqkWReIIOha+oXVsyhum
gEJ++UhssvTIRVBQaeCpwOWcMY5G51y6hDm+jRLB8GXOAzvnLF+croe8bFAu9TlD
GeAihjDGlQYcjz5+nDy1Rlgv9r0LjPQVsPWtLRbUopWckB/SpOAHIE8FLxBOtuM4
/eVFfi39hpno85w98r16kllzrMli/2JWkD//c0uOppNHTj1mX5mfXG51w8w/qU8H
TH+Od6sDd7R6T1PSj/Yn51a99lZO8ek62BsszRV0fcHvYSFILZZ2KsccmlpwNGPO
kQqH4YYMI04jaYHMMQ22iuHGgKsrDqgPDYIMPBgv/5sAK5anCbwLCZB+tT9Idsed
a6g/0hI632AntCcXNxtf8bvBZuKodkQqhowWTrIn7A5DX0LbzB6dpOyUciI0OBuU
BAprfN1TaFEykVpgwvbe5s1rIkeYQ6b/BzlUKHrkBcIOZfyDF8MFkXZgY0g/iouw
AWXfo+/wi6xehfnTX14DqQMrRFDqSzU/snzDoAhUJ1sxYEplMOnI+8b8yzV3iIqO
+on6fPPpbNvuj9Uc049fECHGa3cbKykTPak5pCmJ8yaCO27adhss4e1AKexccTii
jJ5XPN2roB/HiGD8a0lh5iRH9OztFFISZClpV9xze0A0fLk8NafNfSBpI3bonbOq
5jAaLN3TxTSuuWniytuq46bWor63tJoHII1BjzVhw0cCvKh0wYX3OnaPQLLDG3Y4
hsqQyr2TW7Rw2R44tNGpGbhikF+23DkWCQW4Xr1EcvwzMQElACKvwBMrJIoZyaqo
C67cZNDcJKFfiA8jo9CP7lTVQg7a3jNgJjuMSVjyLUCm/SqwefZB6cUdqFEcnAUZ
SoQKizbPXs6GyJfPCWVEJsBkD9cDfyWK0ezHnumRa4D0r2NcM88Q6UeGSrF0TcXD
10K+C+Syg7DgS+CwvtH4wBhAWo3Wg2yXcL4+k3XbQSzyWRVYxlR+RDGvH8fTR7Th
l9/S24iZaWxBZNKL+DcfHUyH1X1uirOF/f5Nw/mSZn6TcelBG8s38drQJSb+ZVFr
cmJvscqctLykE9HFfP1dVXaU8YTzG/vdRFi7ahxnTi4Ucl1XfL1a1YDzpJpkJuJt
J2S9RpbeOl9CjgjWyoQcYjb3GKJunhQrI07HkUOwhuws49C+XX2E4wAx1hpZsOg7
UgwNyj/2OFqqyXEVhXrAA8bOylG2o+T3pgDYiqxe4xnWQPzOXUPrRsg6p8dKPE8c
invU83IJROClG0OZa/fE1p7zhwfCqhFE7xah9INDuv/eexfAOlL8YogwI7/250LY
/VfHeq8aO8uOYVQrVLUfbxIzJCzgwRldhsh0mCuK+2sYyN2dEGxqEPAODrzYDFDT
zWcVkn/Q+scyEUnuhXJbsuxQza+1z20T2A6ekqStlODLdbahrAbH7fWO1/RYoudg
ffsYuM/hQ8IqZpH5V44TG2/So5gJDVn0Ba/D/HdRzgDJjKxW93OVQooRtrVUdv9h
QP8uDJIq4qU9Dv6k8R8z8TOpIPjdpj22D3Y1rToz3p7RkmHi3IIeDyThsY905Ccq
BFRIkhzCWToB5PVWH2RuTZcdgZn2Pc3UnFM56gVcurJ1sKfzUPUeARgrlCNQFUxZ
EwPKYHDyh0KVE05G9gpjCRyggHA9F2zQKUhvyyO2grur2Arui7cCNTzg3UlwKC8M
BPhpUx/4JjfCH+675MPAVKpird7rY04pvGmMQKtshWDdVgW3kE2XCsfPbSsZuZcg
rHXxl8dZQa6mfEQAHpWXh2lXoW83mQCXrwSuFOjC0a2TdTzEt1cRcSN7j1J6s6nG
uPIwdlko90cWm5gE7l8EoYQWcVLyTfJXeeunVSORP9G85/oCh6Y9hVGbe1WvoUIH
N4e8vGn7n9zmZXS4MmZaS+wv23gbwsLLGxCvg0U3hgmJmwh1QIz6hrbP6V2nkEkn
/gPTaQw6vDx08F/g0foXu2cLBAD1NQ9FpOSQKMvsVaTWKwc7ny9uOKa7Q78e8SiS
DPOCL0hlu+DxwEXjJWnFj9fffzmiqofR1NTAAUtJk5QcDVvJsN53QigK99Ngdyc7
sNj+rtZDq0TUCcXy4O1CJ7bx/2G7l7snp4ekyLVd3wCkE4xMT1jnbM48YAGCRqAU
Qo58WOasf2jgDK3HPzDb6oM+LkpVtRCO/Md9zD0yV23fMbrUBAswLApF8UA5cm6+
wWU5kiBhqurLk+Lhvk7772DXwdWGpePLP3Z0lGLohUTooYqzQFXtEWkoji+K8cKt
YCBimx7+/sMFB/HPuktFcyF5C9gMsa36VXaSB49J1emuEGP8coolzymHGawX7lNs
yvsjRODoZjjnsETxKT5jByGHQlRt8b0vGm9F/c/W/Erp30sUQvRDDphT1lmtUAd1
LTjMp/CkEJ8UdPjiant7A7B3Ydi1DmGaMNzqsApcEQMt1h+9LfmFI6QdJFCCV2Y4
PsaKkgbQNC9kfDwSgIn5d5reSJMg/QeSs3pMGSIo7J6oaUCml85X/WCpuI0UqRft
gL9YWU9a99r1LhzyWJq7MxQFl4aDuWuMfNUvCijdvIQ4Fi4XsUsm7Bqt33HZR1kn
9CtnVxcR2rVQcuze2dvCesWahp+lANOV6W886iMdDL1JDl3X/2OGQlpQGLPw7toM
KQChHHscmknE029k7F5PV+jICdPzOkDnk4CMdsa0jKTBVipCwVwPX/wvdQW8W/YF
JhxdCr/IT1jnq1qTWDS/Vjir0f8CVnsUFUkvLXlbX16ib/HCM0VIvGk7LTCmHxPV
NK+c8mGyxR7HYkXevTQrHz/k7WmqDqvEGfNBVF8+cdW1T6Z5v0kRTuP36L65Mve2
703SnmEFFoIwKT1OYOvwbFZ00gc5f+6xbkLdzrxyD+ZL3YXeUJakR4X0vLQmPMD0
tua8qhquEpiLhh8rwUC1YZ3Wxu5++iW+4pABooEKjl/6zgHeizn3qLc7aGQ0nPrY
OfQXB16tc0RxF6XoxlAxnob6n41xWh6DcD4i8VlSJmtV6aPYx2FBwqqSIljLWDN8
ZB8TklvPX+th7PMgrxwDq10fd8bTVLqIThyZM3p5JOYHCZQfIIzJlWXyetQEU2Ug
ZkwUR25cjsaKlTU7mNmUGwsztvFek7ano7ykMi1mfcVtjsFV4ILgXbAi17zdkKuq
KqQ1Ts9R4XOgjN2n7wC2trpt28EjR2uh8NgKVHYb3Vf2npvLpv54+Gs/I8Ammy4F
GSysuyZdeACSg0ZhBzTDF1nl3AthZe941WX2UMiLxE4w+w6I682cca012L44NA6q
ZHD2+DlROuy8Br/7eiUQUkUq2DMYia141HytjypdeBjikjS+dms+oORbbsdFjjxr
JXtAdxcdDpi1FlkjFwPOZEQDY8wRkBmxtYQhCajRSqPlv+gNgsulVh3BcMK0yAaz
vTdAjS7LL6Ew7ahNenRhhKVbSX0O392j6NgOS4rwZFcUyLoZzy/bh4Jta2jgsmwe
umc4szOKLiscf5a/IYejNAE3sPoXw0scy9JC6EokQaA5VfbTHuXozePF+zT0vF/Z
DzZk/nDM9Cn4czslh5joVgGhx5frn+PSs6tyf+nzJmnIZ9ll7CVW4gHjEY/oH7wU
Pbq/QcgDF23NC6Ob3HWI9zNpfxIDJD0tSBL5Xfx2ZUK3KHHdh4VykLfSnZevKRLQ
PETXCCTwVWUh7GnOqk2pl8VJkaq2oZnHfdBzugPqlJPxAzX8TxLgkKkO/qgjKjmM
JKfwJ/Q6KwyxZsGfLWhtVtWt0nAJC1opj0Itp+GiK1OlfOZqpvbHgDFzIqMFsqO7
q9YD8Jo/ur0x1MvLo8X6fT+kKxK7RKN5vvDnhX7GnNKQCZAertdKr/1iWP/54Jjg
+Tmr4uWZ4FODFehOoK1gLhLHZc2UYuuofFdkMlK1Dcu/f3h9rXkr5KBD7y8E2Qoz
U1QSOWA0V/78kbTX19ka5uWMRvLvkdm2cenFOup13/9Vf2eMhJYzL/6SZyyFO2c8
n8vd5O7af3Xg2p4uAbBsv3ae8KV8nGeJAOcQiMNI3+ghTSHEgQohisCtmGu4QPuX
AGO/OOiaCSkE2pT5x63iypMT1WBCptoPy8eJ6j+uCKj09b0s81M0wEF1mxgaG/N4
t7LuSSOCpmUF0KX5rv4ngS+qRTQt5LE1oK4Dye2J0LbHdk5YM/HEUPVh6Jyoy5KA
Z65dfFKq4XsxcTJjIQYPQ2CtG8gmo7twVNjatz1VDZIi97OZxHdPcwkqZ/11jdeI
+JzhDVNNWf7r/w3kLoNseLi7RdCHTdhe1EDRtwEmqU1ldtoH4cqNZLp3GxHEmZqF
N9f/xaBgwZ3jQ42pk7cTx80SVOB7qu7Zw1oCgBYMaq+HUbr8gXrJHeysfZsvd9Hd
uXNTDehScPYUF/T+XwM38GPw2yRW+EAeCshxc5Z6T44D8tuZv820+/ozQMAQG8Aq
IVm0K0XZ/kMb7sg+RZsEZTjNrJfcnN6/c8PZWyJ+/cjVSygweTea8kLfQrifyV8P
G+G6eQJ/z9R0ZKXeFKZjs/NUitvedlPL+RYPKS3VcGfy8wM1mO9Tq5r8bUD4Jd9S
nrvx0xZKLl8Uv9c1g33UQSL/T2n9b4Q18mda6JTWP40XaIMPpXWibaGPl4BbtM3v
UCFcU/TingRsaaC2u/f+uUqUQPmoZxxtq9A9IZuPUqF7PaqQOBkdJa37DeN2sdyN
1oRJ1TvRG/VarGamqym65Q1qWHyHOctkduaODj1fEeZ9HZ/NggCOFry7BEM8ROzL
AfilV+v9PT0A/2VDio+AdpjcTztsOQqg0yWjetJWmrgGbtzVPF7ZrYHZsq8jalAl
Vgw8hCyiM9JFN7sXMtsYw7Waaz8rKdt7BByKjKBlnYQgEnD7+wFsllBZHNqso/iu
VByH5gNmO6IaXFZ2CWSdUFEHLCQEAvDWjxLpBHoGRrbTLqMuq2iAfGSfjLdiA+e3
KRNmxOEv+DHolI4gV3Ck0eB3pZmkUlUa0kXHsnJQ9I1k8ma7E4RIOAADYkfD1w54
TR8WKiu9X7OzN9LxvP3AT/jXmsA47l0QnBamlqUQYE8COnxWCYz0mbyfCkhSvbnN
O/MqNfv4XYB6+J0pngdipMudj3zSdBQLZis+YkynmH8NOldl/K9oTQsGpYlpXKt1
mi5q045svr9bXVqA1fDgpF5lzES7tyNzpBwS6yuuz/Ge9PYCo9Rr0s2VzAZoZr+V
fv03lSUX/+vTkS2+6QG4zOu/USFG8rXIqJ2Ca1Sd9w7O/N+N2pIhmLbruCXtzPKT
rusiU9GjVuI9DsEuwUTrY4Wehuj7MS84GarxEoSvIfC2CYm+WE+f5wAleJJKy99h
Y69koT2WxEwfxMF43SZB1qFrcg+neFoqaWDGv3yJ2b+0oxPwJqwEjTtSvMok7Hij
UMb/b7haC/gFaZ/He2AH/2x7OQoq33GxGCw3TcM4KfCrosGDwZo3ebQjOXWtU9EA
ptXXDaerJ8fS2EqQ+4PXFNa0/ZhULCwMHcK+BYl+RoZBbnD5URLm6TpA/caSA6WV
s9Sz9YGKEu4DP4aH5oZrnH3KYKQNGSB/bfVIRqO3o7oaBNkGI6ffQnMtXdaLdyof
lRDLXINrt64V651h6r0gjEf1bZYCut/I5Wrvoq637i0eDjh9K9gCrQV/qdThxpsD
RD4GrtLcX64mbkuSXjU5v5VxYe26UVUXrCAvYX/O86yAQaoD/swel86wuaSzNiWY
CDnJTh7FYGhWi4nZyQCJQI50wNmpvs3G0Mlnp+26LYzwHM3fKqGOHWsqZrsdqpg1
IHd0C0BSWHIB9jx4At0Y6uGj2416ZpWxUy2I9VE8J0w5DFzkAlkPFjiToYkwfq+6
FXiIXUrZFzhOsyNmpdi2imo8yRuNmoTsk4G/ObQuxHchSHJ4yBxnu5ncgkCZkS5P
u6AxG/REsG4A1XtpjvM+mcjjQ2QOadWI83wtTBXqNfiN1MqDLtBnV3hDwWXhftEW
iKdi8lzJu3czTad55BqFflBNhT40m7uSYXRKftVxvuPngk8teN3Fg5kqwYCBzVm9
2teE+B9REKTCwE1e/zRMdnQwuJHwI8KHM0YBoAa7XkE2f1g2JBh7oNXb/nrlkb+U
0quyechgGo+zI+m3oSHe/b1SB4H5i4UgdErVfsBZrFUQ1I1zmZxppuZKExd0//da
sCE/xPvYoXttUXSugYdS2I6x9HI4lF1/hVMqP0/nn4kKHiIEw6DJjUT7HEsQKPAE
H31rZ3f6bIuuSN8sdfdo+FLUpsHCKEeqC9pXhDoUslrzR+RMDFirREavv+sOKZoR
AEEr3SV/6rLbeX22IU+UKMximpjBARI2jsLHaQJB/rACktvsRoNgymLICJ39tUAA
d98fSWS58w2y2K5kbtjQ0V6m7vgzpxo4K3KFu9QZVhKq/SLXTKq2Owm1UmGqVKEe
ZIfVlU/8F9QxzPcm5P4CYPN+c4vNxAj48e3G7wp2YYlECyIPiqmemYyCLneyVJyW
Wmc0Z/jGCmDFc/4h1qrgjCvECltz1BqMXph5a2piTzfe1wCvRZdh7x8zmm6Jb9Fs
arIUrC+uFLphl3axtzYY+ZK6eRBUeBTkmAj3N0936xgT2MFw3TJvZK2VQZfAmFeY
D8REOrOp0t9edvwh7+8W7cGZOQXMHYmMXHyNnSW5RsdBAP+GRul+vxfWX3vXjGbE
5n5arrBYjAd0dIpATQVtr/jnVbTfPD1Ql0yigXveRHQbP21aB6qS+4c2erfEH7XN
GUoC6NfJfYcEsvG7hndwKcBSYkjZ2MowOx4oLtIXk9JBKDBjcxOe6NKzM4NutJAm
Yact7ovt+2W2Ivhqr2bRWikEVlx5ZbGP4Q+RwXu2n/MIGXCH2b0yAGsa/8D8TjB0
dZzIBqY9X8UxRWChtLjJGMyVwAivycaPRDbZRCobfarTMcEf0i6ttU780UxnVS83
YswbGFP13i4Vi7eE+GTtuP5wPV0JONntQW8vPqWLdkHcPRt0zJXMesyJkLDPi897
ir5WzziBbCDZr6Ceu25JLjwnDLZ3GUey4p+ppyZSGWt7jdY7XQ4ZIXLJW6jyYcJd
U7JE2k5g8a3BKjLXdP5GFfPcQegkzfe1dhu4b53ghtOzyIZmQIls+TDrCANIylmL
Z4HYJDetztr38GL0xHaruhD3knJRKRsaPNPufDFRy8ne+p81LbnxywYk6Q71gEhX
7zM9xjotdeDeydr13kfLhkmiCHAVT3R5LUY0NHqleE+6CnKO/5e3exLah1Awrxmr
glezjVM9oVSAhxm3/FrFdDfvxb1xPWwMdMfAC69upgdu8XTlszWb7oAhDJNcX1Vj
lC/NaA5x0xXMCxprtzBpYzpdLUTcr12LeQXbJW9c4JpnJMoqXASiT1nM8fN/yz9F
INC0BSlizM8maSaTmYv/zWAni3knPF4iRcFM6YdV0UR2qt+l0pTrV918dfCvGgfk
50iME0w60kAiqF03jfCkMKLoMI8R4a+JF2DKBePm9CGFHHOlsUukyq13R9p/muKS
M3JVn33QyUfSQZWAJiyRvVxjZuCr0b4wIsQFVFbzjwkTCEaI9AV7cE5TQofaC9QW
2jWPcYydDaHZD1X+JOXmsm649N8nNlUfN9+yPFRDrzVnnEEYvMvL/QdjpErdv4tf
cvpJrVJO9Ta8B3ZCnRjFEJY1Fwabl9SLXGiaL6NIqXK0Z5A6JM9sbEA9aVg2CDPk
D7TxEIPKX9CIaAzbrVWx6opD6vKhs1JAzFnVfEJyhdniTFNjMNKgEw5WUNnRjoDR
fE4YJEPnd8wz2bHzUbGX6BDpeP3wtwdrgIsf41pkIhtgeGvuWcDo1UvS4TuZefUr
TI9RyokgP80K2VjxbPS2qfOB0l3D7i7wEoerispRAVWSMZrNAgL9BkmHOqx2HJEO
/oU4Izwg0eO4JYFFDGeox9UVRGrox0x25qhukhrrmgtkVnpwsv6eA4RINvf0PvMa
89jzq8WbZeD794jipKvlWeIAouvXLnUGq7mqL7Pbz3cGYEOP877yoDYBucmRROtZ
QZOkrdhV8JmzwZTeq72SGirmqih/Swj//rxTZpDKNADWojLK+72BVxrpCID21+gF
w8aGBUwcc8yhqew1Y+oPZsYqe/7ri2pY5BjI0/ceCE4jcB/n+VmMy4T7n+ukWFwk
XN2ZZGsZwadpHD1sRHO/ObZeG1JrpUNNYa5UL/3lB7rbxcDskgkR/JTNePm3Uzuk
g3E4cDdNjtT/GzAny0aJwPu1hz7OoY7I7PcW7YqsFOUWbJo0jh5yA4MqS00Yq/C0
KsgGw40oMiraeN99qv8AdV4E3x3mSlAifzOheXbYiYHtzAvBFXD9HUsfSzW/5Sfg
aBYVLLFuorN27tIZNEH5SH7nvjxAgP1w9ulTWSmChsaHBQ1EfKrlaL4bMfESbqOq
tKkDawCNvx6/78e2pn/7543ZD2txpzVT+i7Onzh7J23us78qI1SejdtRrJyKu44c
cEzgA7138q0x0x/v6uYJP9XlCsPjhmcVf5H2WRrXhudrw6OvpoAaiz9xgosOQXU6
KUPBmmOxElv9ohjUyISoqxZvxK+gnrah61+a+SycKKgzfnPrieZqNP0cju+cE7R9
wcd/KXSPmHE1mDF2rjYWJJV7qUR2EFfQLb1nHMo3KMw6ouJEtHNxsdg1IzlzRazY
zLV4rRDmBwTV+Vpg1lZZw218zqGFPhDSuenqAzs15N2e/jVZ4VMnj7dUCgcdoU/x
pQ3ww8qTcz2PZoiFht8zanRzAiV7iYZSP++maotlo9bThQbkR7xtEpON/2WGVjag
dZ2TRUrKxJihtXJ9MJR8esQYdnJqz6FdFq5DlYSSsohE1j3nCYqSEMP+/WAmPKKm
ga0q5wBgQUZydoErLRNskm81NgIwzwkeavGG1PSw2ISkMT7U487WY6OxsVMnaWmx
pdahyORBvra1gXsT1+PnuQBRoocOgi3IfFThx/sO0FUFysHZckDf7nknCHhx8pvx
Z/pvnDD0y/n6ojme15D+ChK9+egNeskiZRBFHcC4ivGotjvzVTFfZc5WrFrRINdx
z8qRoB/iU0lPCkrRGfSQ8sJa8DZh5xHzxV/nPdw+nwE2Z+k82zugwz6a7XcXiVsa
gO8app7db9iDl9MA+bcLDq9loFtk64uI37OtcxFbhAZrlYxIPumsBvFATSBe5Iwz
7RVz9Cd17ZNsC75nXr6oqiVP5mcsYBkFQ1dED0/nbjAIkxxuN64FExn5rTTLg307
zAg5RtAN+CkNcEigDRSlnNZcntlM9yYIwHSKmxcpsN1i2M7FTVJYegqETC+1+lRj
jsdJyDtCpBABHZN/znya6UfhwytZOePxAsFjuUKEi01IWEoEYCgvaMjwiobbGySK
Jt//qEVujSP3Wnayyfy1V9n3f01ORrnF+aljACqgKIvKVDchiUHYHU2TjKc1G1xB
eRBhaN3EZj/sXsr5QFYC3qTcrY8kCny8hPrD7ZdgOrOVeX8PnWr2ZBszisorCZvO
7JX6xc4F+YFZNFcLNYm7YG9d7N7XX16eQQAtP5SF11AjJgayLPTl+/iGnnnKHBtn
4TQq2AhJfIpePiMQDoIDTp6YsWlov++ckQPE1kwcxUBOms6qOYAtfq7souq94h66
uDJ5Aey5E/VHzK1JM77Akzr/5uqeNLJpQtytXwXL5gGDlfrAgJxUqYaEzLLKot0j
Aw4fglvWuJV+IOdWGlNSRvwIbIUO1YccXdYEKNm4beycs9ovuFWK5zJCP/bWkLyM
6Fjly7Xv7cnH6IjPIBQ+jJllq1oe27Hs+SwNgbog63EPdhVsZkUk3x23R+pYbcEB
g3l5ftwlt11Hoi2gMPIqWntsen6msF0R+u1HGMjpei6ydxsh1nSFQU2d5gzd7b63
OXXUdXQmsJ4klPLs2TQlAbIfYIJZBgCIW3splUw1fua9hJ8SkYjawlh7vH2jlH3x
2+RH1MTO2OIivs8JhVSwJnpbTiucO46ouXJm9HCyUz4zaDltAM2WR+tO7g6SE3qf
SLGAqgtzI+EBEZZVNuANGGx3FN+J/JuA8Vcn32Fr1W+ds6QsiTCg+eIh883Pp4cC
cf/EcwJ056tE4CHA0tHax7uM5vfJ9QFJbm80VrFOT+bklvmSdn64Sf4gwJP7Fqc9
kkKtFl1odg0ymenMO3ZGY6m83p0oTHCbfxtSD89cUwBMbtI1EMlQiqgWgNw45Sdi
cPrW0ubrYbyFzM6dRpf5WGL6LQZlZkuUewAqvUProwFdtCjOHi9dgOTs7OJLCkdw
tXUxwG8SqcgXFRm+OgiYH28vp7ngEeFXFRzNwhdofQC461QboOFHs/iCLb1toKlV
c+xVPc/60txbDFbKFR/UQ1a8vqEqYUFuMi6HXtzjfMRDTbRH56c8n10hHZSCxTQT
t/GRRnLpRJfTlafGP94IrM8anGUe/ZG2TvS0tIEu8Es3xwHJePfI+0kS8EHjxPPJ
SG/T4EPr5r4/ItLvMTCD0JsufuiZQPbMTHMgw2Q9j6qZWd+NEUY9HKtSPwBTUB+6
GDha2n4qSaeIwOTTLzQ3y26oJ1BD9qacI2nmYUHJMj8eyRIBYQ7QgoW0K4vXAtpB
zL/LHilebwN+n7fXcdU9KGeekVIuU6+dhqRKq9omIU7PSvuaYmxuAYP3SmNODG9F
PazyL9awn+q4bYbPF60xgs3w1LKNHxMSGaxUToWXWoR3o2SRbCkkkrlwoEHA4r84
eKD5Uo2F5qoKVc39WXDOfqYSp208ELDTRqCw/KY9CHGKLXS1ktzR4IMVBVPAHx3y
+GQsNKDO+9iXmib89Bij95wKqgZhTVKfgiOGhkjn0W4HPxfZRxlFgm2MKawVjszH
Zgo/BdRMQLhcwExXrm+chRD7eRkUpIzZzn+9HNeFYa85c9rUhtIN0YmqFbuZUQKI
xIqPKUcvvIeoFQpfp3iDJQiQEste3f1hXuTqrlUZuSVYkZPG8KtCQBFrFDINrH6n
EAGQNpcEmXdV4UkPcn42j2pTe6wiU5t8yhekkGV+BMiKow5uW9qBKmjqB3WUXs26
tGcI9ilwalPKhouekuJ917XC4eJ53ooZbNAJ1ZdNnFtZXKB235HrrxMOeraS89Vi
mTJWPRIGDkj+5o0W7yT289aCoN8oAuXabvGw0OSPHGr5D9XP2UPmc7i5hHCQMbEq
qrScbtlc5sHV4UIfdSeGuzTnS2fZ91G4n9ixT3IrNti2KUqBqaaLsm0f7Tqi/6vA
wp9YrXRggLR2UZ9S59RXY3AQ5GqwPzLT8eNIRPQ1rSHd5VxWkVgUjuBgDFUOfWhn
emCVUGddPT+pHkxI05KL5YvBuzkj7lnaGH7+sqqHtQPtd0mu34naGRdmNbCei/RY
S75Hs7k/A4L5nlYxlC0G9T7dk6FrZ6j7qPz0t194qkVai0PkWxg8jf3KxSjaKJ0L
p4P7j5OrRi9nnmvTTtuMjzteWoqRQubUgzFLtH3C0M+PTTPJ6TSAMaJKw1UIrsUD
gLlfciyYeiEiEKfdriIpEJh8i5umL/eIdo7PexYIphIevo6hb+4mwpHlKPRHgGen
otoBD1vYC8MIzp9XX0ozd57iDqwJ7RIPcAQ8fcC6d8Mp1dQ9PQtXWpuTarGlnK8G
+XedV3kdLp3CKiriyTiVW39o5QfI1rY/e9ZOYIum5xoxrIxKvVJbJa3Bof7Kfg6A
lPoTULfeJHt0L1HG6kQ3ymEeP4iEA/z7z9KqRsVVF82pkhkboRU4b1E8LAAlLWWf
73KlnWCQATjvREtr6mxtvPbcAhLRw8s24Kq3ka0CCEUaleA+MgUM2isMbp5T38a3
erSBjggxxaFORZiwFRf5m9KVS4feDf4is1zToQc5XulBRhybekPFY4dkaUOUFvc9
RCBWGBBuWiLFmHDzx4EI/qnZo5dltkiXsKJLPlOWl4dRYCsgfyivr3Ys3yM1zaz3
15UmNRoUtdJsPxIXnC2RWqKMVCwJlz84mntwenh1C38sOY0ikqmAVPYWJhf4tT1N
gDfbiku47jLIIXRZMDz2be1X618H5FSHwFaL0nlFTkyu4L0tpha7Sn92hq9b+3df
mTeeRAoj7gR30MAPDjXtW+zZKv0BDR4HOle8An9zLHFdqohVAvT49ee5HHWo4nM0
CcTwwkMNkWLd30CusMcydktRz+AjIrRmam2c6F/NIv13v0gfsgumRkAKHD9/N2M+
Qvycjd+GxgVB8Q1UgKZp/nyGGE9QnFDXApl3i3GGwxfW1WW83abhRovqzayxrBqW
FBxTi6/Ua9xBGluJe3w6qnd46i0ZvK1APy3dFP8LDbcPKnV2kXSAOBNyyFikMZym
0DTYvmTLMaeR3Ld1LI4eWiDVL1OUjWvhIUuSqeLCluMLaavB4AwWR1f+IJpO9i+I
o9z07M/XrPFk1dPhcp/kyxriNv31cYjmVvfAb2Fxg7vJN2JpPo6pOFaKjonCb6y9
OAZC4LO9UhYEYaSwZGevRYrI0ipHl4d7G+Lfq5FONE9ytWAAhnIFiv47twiyW+wn
aFZmeEh80kBhsX4YwahZn47rNTZrfRfh9T9hjDlL98E9sFy4s3fwQwg4gkSI1fms
H1MYKeEX6+G0C/lXuCIC2wekHG2Zjk5UUUSm07cINM2tqFxIf5a3KUVO5RBog/gu
Zyi6nLNReJJqUGqJ0SbHgj7OfSaNApuvXycfoCFhz2b+xxq614w1RR/0/OpQ3n1l
GLaQ7pCdKMRzceNl2ztxnGDsloJe3TvMtDxDUMUKbjbJbOadqRi1wfkp749dX3h7
yyaCT/lqmTNo+G6Nzeg1pnRRPbgPr1DBZZBqufaAEXnjpKjsEBjmt6sjXtxju5YT
jOziwH5CwyzosNU34F537QFuyRJZ78i/8u2ll56hE44tAoT0QXcApTMn1tiPFbh/
WBa+fJHPFYPvwfhZoOgLFgP+0YQ/VPWnOCZAIn+/6BFnLa9thx8Lx0timRu2yPAJ
trRvO/qF1J3ntKEzZc0kLqDJSx238/bI4/9RtXXSkfXDJ8OMCg5fQowGgvMarC6k
9IFPgtHFNmdzh+tCWOaAdvDycXDAoIpMixJkROiInVEiDoGmvZmKPT7ig4ka1ENu
t+GLFPX47nis/HH2whdF0djy3/aYd3x4tLNkk66T+ch6nw45kBarztg7vy4kCUkB
7TthYptxQU0cIJDw30lq/oIfOKFNIknEzcKMZrgRF1ZYDXMjxSSJKhh+EcgZIELl
WnPjGH+vg9K9NFPAxiQkAGVe+hA8PlGC9JJobV51UKB3A1RQeLQ//4tGVCpdoL2e
cY9s8KQFqxOanDTwuO+KH5jB1OB1hmtpsyngNnZiWeDBaGEy64bzA/LoIdxNQrRJ
jPu6sBiPXfiobS0eTINk5EoYqrJ5afW7yQ3/i0et8tdQNosXcteAzJ8BMEuO7bSL
o2BDxIhLosPJZL7g9GPlrjmnxC9O8hjXi169a2GZKb1X9/fY4Ty6H7XAhNI210zD
1JM0WgqDOLLctGMj2lmaXoS7WwdMGaNXzDIKHFAj+Uk+tnr0OHifWdXRYGAa3iiW
HkW031/iuBnP/SHPH78WOtHX3psOJp4BTuW6dz/oAyiXVhIUPYwf/lnHvQtTnKIE
ygtWhH/lDbDZksxghWpJLjs35NQHP212x/CTjaWqFCaTH0EeNYJpE053hYwKs9PX
8a7q9CKfOhZmeecqU2898Hbe7+KyKfHY2L6WCSSyzOMermmtjQL0SxcQIv83HLdW
UQurDXC6a1h6l0nZheC5a6hN3PIaS6woe/qiX47Zk77tYG4uOA4idh8SwtXosXi7
sY7dpS7jgwZ0VAQQAzHTZPBwQGjRUoTeIftj1sjY1sUzPuSXH32tAcLf+vE6iUpk
RiqKCS5uu+JcqnJ+bhJbekWJ/MDmRwGXMGhGJHqSBtEPS8cfpIlEy43Nx+THFhaw
k/FFgJv3zoNsL3ai3pR4Bl0m7QGG0AM3UtSKGuO0kfyZcnoIwwnX7DH9BAyxvNO8
znTg0NQJC07f+3vUGSOedD+NQD8VgFiddhY9nW2KgXJKpssUoWzlEV8T3s+cEeu5
cpQffkFyRvQOBX6L8tFd4KyOXmoi0bkdQZaFcI8E0FM2TocP5UfyCfJ689ENQW3b
VNgrO50WPk5u2rjigHqSn/heK5Db6BLo7st3lTRMHVDhpsqjgFrWnDL4eo7xSDUy
zMFN3k6/bFWCRb82WN5xnrb4FVKrM41CasNV5jOGSl+WxOei2CJZdFxzVLfqPDLf
wjZWg1aCsCB7a+B/R2SgKGbDZE9z5XzW7WocZI8Kzk8i7cnC0zhPVScsahgmT396
tqVSqnw1mj9ZZZWnhfMF72AgHs3YknS0L9zAKV8UXtS0TOZncabwwGLpu8FfmpLV
KVzPUT9FBhEk0+jpWRxH/+fSpjmMQqYo42kA+GgZFCfjwyFLZshEURX2xx7J7CTB
DJ4namyrnGJXYX+LgUVWve+KV3K6U+yHaXURp4bgNhtgH+WgTcpTwI3S0cmZ7h0C
QhTzHshVuCsf43t9BqGNTLF0ddqFKZukC/m7OX2dhFYs0DxqDJSwBeYPnOX+t/Yh
0oB5tnh+IpTnOEicsXLICrvtv1BX+KMw42o9vHbOP1qzE9rpqchQ+uJkLs/ei0T9
ROEIWrAUySFNdc5OAvYTeCWzI1zwR/g7gmdMT+8RtJRiBKu1Amx4RAk3u2Deey8D
GMA3z/CNsuJvyx8PhbmA/FQXtwbuMejMv1K4tWFwHRC0skQ5PeuatZYNA9u3xVVF
4feupMrC2W1ZK/dK93rgaSBiUx5SBanpMfVuh49+mJ+QFtyBO4ySwitehbx8Eyda
aJNnNGu6/vqCvPjwtDaPQCKC3En0drKZvEFm8q8sh5teWeZP6du9YcgBZ7fjcfI5
QpQM4omRyTFnCLgHHC3tVnZ/4AfO5Z0QwF5EDCJ+q/mKZ5tdBRTg5u5b44eD5JzF
kUsvSAxxEQkECu6ODfdxIjWaYdxQxPFjD8O00lDY9Yh6I22rhNNVqF1TyQ0fJafk
v/YmupFh5BiE17eN3x6/sKrGbFPunb5fz8qwI5awByPddbACheFc5xNA2K1As0Ay
TsqAPS89xcSr8Kq3kV7J/v7R8Mem1RrRxQoW7Ls2+u1SWKybCUmyXpbbCC1xjRfq
G6xUEW5iVfZFiLLN6a+X2TZPU9MmXn5bn/vbYCpTQ7mx1oDoqd9y9Es2OqEi/1VI
Q7f63imJJfpLb9I2QmX2UbYSF6srBG2AiHaygjpbbO/UUmps6WhaiGE92Sk2Sg6e
9fODI2If/fqSbYPPCZq/NIm38Mlar865Spcy7LFmXzoUQjbU/k7c94lBtRtnu3Hl
yGxhPCmMjVkDQ4h1bXDAi3Ur7gJ/JIQ98+JLIc6KPaqCH/Q4jecrHhIrntXhbdWA
AK1c5ZLxYv/SFJg/nfAgS4/OatQLJaZPsaOPKU0sBymZKBVmHLRCzgah2AIO5lCL
pzgSx3GfDQ901dN9CzP/n7Tlc1EWeBoxS9Q2X9tniSsKSQ2oQNnuQW1kye3wRpDv
nNSTb3LNQ0xXVELwgBlvc9Ci8r60PX1oY5wmtjtghT9cszmkTzwrNL/u8ld7LmEI
EVFNbkUNawepIxQ7H1u4XappJek/4E96RZpcMYFjkw0e006tYDn2tjmQl+aXNkaA
NkcL7/NbHwyZ9eGFGnWmOeUaYUDDMoQXDAGHmdUI+WRfpHHKfk+LvCSN/D/10FME
ySNNewjY/WV2R6n2i0wkrPdrSaEi/CEOul8Qdqq359TSqPT1vwMTH6CCWmnNQH8I
HW9HZrMgC98sdyouY7AikZ8SxlZ9aOyq5kCFemXFGY6Yjl9eHB4dJFfLaaA72ccm
0w46f6kuGFyQHDsX0xr+2qWOOkRYmgvxZJD+Ucq2MCKru9OldwMB/Z/XrrnR4ZC2
m6TBLSCwCyyaGKTunl/1IcWB30tpnGPbzRzJb2KNrSSRMCmtCLsUBQcLQEY99d2b
mHpPVYfhIjZ2o153Rgiu+5NuWpmqIAn3WipRtqA3a37TCv2756hCROA0R4DAWhX5
sjUtd6ghJgblWlj1d/IebNjftbjkz65CfxCpi8NsTlPqBiCBvdBXgYqZzxM5b9X3
66klg42f5fQi7fVegI7BeyiwU2zradeZY3d2c4K0UzJ/2D47/6bEkaBjvETVVpld
c1A5oeR+NCg3iIaiQXKepSo8P6Jy5a3MmV28vJLO3qffTzqp1dRbFi3nSadrPWs6
eQCZY7pTWRmcKxDacanPBNBKeDzIPUbLh8sNImb/baY1kDx+/pumRVPqLxbbeYU/
DqVtcnMdTZYLIZHshQcGoBfwudg//f8/SynHokfJ9JlhFXnJFcQocGpJDKugDkUe
ciuVkD9NsWgmN8bKbP0M4eD8O6LI9cd1bj+1qag+bPfn5g89o6SHe1AI8jOqVTyd
ut1n3Jy7Z76Ji+waorABiTylncsOkVv8OxtHz0bGSIb2Zu/HySvkFQMLF+GVMROz
gJPwh05NgOiReZasYrrtd9MP0OlaazhlbIEBvFRLqmEnZCUAAoHRaYhBJTKLqQaI
4JxStpu/vI6poc/FjZYoZ9n+L6pq0R5C+JPmRLw+DLsARzU5M8JFqs8bo60deXCV
v639gu0aFHAls4Kyrhk87vClU1HwnorGrQcG1CCgHxPJFFvrWDHtjwwVnk3EPPaJ
pf5L8aeXFxVlobqOPWfGwHoBb6KmDi+JcWdnhvIXYhixcAzHQN+RoU2nZt4ITnic
FQciXwvZv4MiZWdJydXraJraLEgKGW6k2PW4qqUT9PhMWBq2ihrf0NPKs45G9uDr
1vyyPfGdjRJmXNhmZdMshWQFttq/S554dgfcFBADwhrCYNgkfG63Ji0LLvnQLgpI
fqvZGBKm11FqX+yoNXjI43LJZZiu4o23/6OVUuY4n7VQTRMxsa+G8ScxQqZ83Wju
oIk+3Le8x+FcBnStaC7PSlf8JlAQSOnBaYcrorMXnLeCMfGYHvlXV5VXxGrC97oT
j1Im8ukr6IiOe4CfT2VlQENLCnRV1hsm2WIF1QJqnISHPCRXPU3ryvI6ANyMTlk4
zLaHQkV8Str373kWUw6/R1iF7TFtZF4DmIx2bzbTeRU4XMgkDRriZp9daAfPk0b0
EV+iS6QB+hH5+yqrC7tzDuZK5QfHGP7v7/GQ8O3hbH98Bcmfwv8RR5v1VbbNF3hT
Yy8CEalXplBBn3b67tV0OqEYCglVcsUVe2wrAfQWFedc2zbd5N15cePtU+q9nlY6
P8zH1XHEA/WLuuAp0ptuni4DTdH8D+AhMnGCZEVbqqQsrnQ3J0+C5kpqCsYSlAy5
bZ2FYK4X03BCuqWUhMIQ5TxXR1PwCrSikbWz3Xq3HQBUs3YS3ZfuRn97zAdmc+FX
cYXzRX8ruePeIGRoXbAnMwqeSBDUzef5gd6WKSUSLpM0WQP5pKZTKSd74wY7B5zl
832OPulFVR80nIjab7cts0YJiMcmXYJ0Ds+rwm1zi7l/U0IH8kR2GL6JhrSaLj9d
NnWkp1ebSdSRkElASXYVaLxM6/vCrtv3mF9+vHaTbgM2ZSgslSH80MIJNS+sVtYi
NQZ89z/qUvEfTX/ZJUyesApF30AfTMJo1QjN1usdDx1YB58wOkhcPb54+Im7YjNb
Vswwdn7hfknzexbRIhMvlaCr6+pkf6ksxkp8C/Di76YHpjv6W6elma1whkVsFLuW
dhCTDyVF8pOkAd94fHItZZhPyU1ymknI3+dhlyDR0t3KcgfybsjogiuTxkxi6qm6
hCpcWo0t/9ImHW9iu4+TpoWKidtxjHGHwDyaw77JX29TRGKMOiqhEMgkV/ovbHhf
D7Gf5SqBsrKM38hOb1/arytYKRyIF7cxEnuFiRBHiYXcNFunux3g0A6a59ZBJ7i8
p+lJiTbGaAw3n5+kWVuyp+OTLM6fyYEOTRM/ul4yo41vPMpikWAXTSsgp7JPVOpM
KXDEdLpVNiDhb5etLx0XhgaTIaNF95s8ycgvKbM04bm40kKyUO7ObQwD7Y3USBsr
Pa/EFfHOBIgpDMIbNDPNF1V7Qf3BEBNfn34668UsF2zHOQ0JvowlcejX/rJEB8O4
RkuRn43JQbCV0PTiFGh6l0hhbIS35xT2xOFyTbhrAhGSK647GyTofgO6jZhn0pn5
C2us1RIy7JVsp4PgqdErFnQVVToIAFF1NSN0DL0MNBopYU98qUIfoIs+W85ZHRiN
42AHVrhZXzc3WScdVsp5ubzEOb47StauykshsUoMcVenNRgsVPdNlgCncQvAHZ9z
TkZlIW3yrDrG1mcSFQvEExgz5rZGma6+ro5c17+8DDP7iNrjJDqaRtJmB/nIrVbT
6Mh/vO4cYFGI18xXgJUgVCE22Gq2iOtlgtsl162jsObhzn9DN52pk3YonxYqPfzT
HKPLM/GNjs6ICf1ej+XEPZv5ASHjDvn3k3cUdden7n+rGEl5BzQY9sXKNibUuR30
H6mA1Xkkfn550N/EteXrfRet+eycA2cQtO79XlBuWC+q4WuHKLOjeW7IUyq467zO
USFjvKwUuyvMYoPlOl2riQFzuC+lQ6qhsB8tWNMasdntG8ry4n2bnw2DQvalsa5t
KgnlgrzaFJP2fQOwmINAn+hGdW//ygyQgvoDijCPnjCsAqGB4Th/c15iRr800t0p
4fWfqv6t4uVsdSL0gFXX8FzmAPou68fwrPXm6YBSSoqH9PGUJw8a3OLJjwtIaSfW
jLcbyTcJKpYSki33nHB23g+clqTn1Oo158nRGDuOhmpj68G0zOfSlD0q2TlIYtSi
Buh0aa5VNfWGOBCv8fCBdb6p0lPW1BOplxM85aflfJW6tu1Cx9T1huPB2zitInOx
uj3j+ik9vuhUu3sjN7WrEgbMmenSeGciwxcyu9X/hzrNa4WblWd+hQjRu/MuksLU
HkkD1Q27KjYdcJhlA3CBVnUVdtWtHVK4YimqYa+xnPlLMYztCjn+c7bUbKw5cmlO
MkkWgGutDaTVJhpV7e9wk0+QqVklsmuE1fkOPpUSxIHIQcBQtCb21IOMTB9U49mu
gxGcipl0NgslpPVAZniEZccKcuEAtTGjwpZ59Ro6NJypX9drfbTuGGuZ0fdUNY20
A7WkvSPVSmTQk2xY4U3Yy2kkWeOk8OKmJ5peAVQPlQDTtaI1Ud7MtATEzPpQ0Utr
tyl036+rTh+Wm5T8Bd9JykmwEGeo2JAONTl1+5nT4V5u5lnFACdxYy9fbUl+hRaW
DkN/KFcJLCr9fx+fHGSLgv676h6g8tZCRsoEc7HfSQDDY5KphRzPaUQmf1OMpao2
fSmQu7xk748try0TfbyVe6Ra0eWkRc0+CRCw1Vaah8xiumJSUTV36ogEobVQZMZU
DQp7Yy97qwvZ4rRNLxfvCYTC6Y9VOoYuQkYQFSOpWobQYjQ0TPlJKT/Z4pWdmJlc
ohVgcJdJUtlOBZlLOUamZ3Gg5m52zk0wRiHY7lTE5uxAb0gpNLmi8jmxzJMQmKEx
tBPQTb622+Fx6gU1OWZ4smGfS8I0pxx2PKyKoOjmBAOAEiUSM7qhCj7dSWLNL3i5
rRYZMNi4G13c958gcw27yIAXePtjMd0UbNx57Q4NjSfYKIbd43bz218YUEBH1DyF
OlcdmcUZy9NtnCZrxt07DDifGIHr8s5NY2fmuBd1OmaO1Cx7pyE7kIanmCyJD9Do
WXTWxOgjWW7sqQIfuzeVzUFxW2adiP9HEu63felORUMHi8Km0TMQtLaBmjTOACHT
ZxRbih+vXtN5vIwe/ANv8RoPvrkNo9371wP+ZY/5uuXFxt+SovMtyqgz9dwfNn8G
jTyanB8+J2/Vg1xnqhcKpahMawKhAp6cHd6mpb/HMrp13PKqKGOmVh0mYts+r6yL
hbTAhDKJYTMTWFBGZ1Pjk93d0hlt8T4mRkFXxIfC8o5Fx05R4m+8tWpzm46+HhE5
0QT6UNpj/FIRNjygQoDQpeo66weuD/c70pYkAbou1H107HQcVdqECCkALGMcWPYf
AcFnHWdpnNnDEudEyfqzluO+wWo1upMa8NWWXh20cL8VjFy2buXt3+0IchtqfegU
M6dDu3cldkjDUzL3UHzpG+PBSRd5BEdevcUOpj6XhHqKIN0tzxEISm3sQwYYY6Ue
mkOcBmlZj3TzEsZEn4VqywiRBVhAvy4u+bcs0UC6mM25FXD7SKCTSLX4CuJ0cJtG
YLI0X9vhfZsrlORQQb/CRKbITp7cQ3NZRQLfd53vBsGyAJPJdOWnOs9ij+8J2Eqi
0U0TN4SMW2eUMNYT/pQ0kISu4hYnLQ+aNtrJZTKlECeY4ml9hJemzW3c9P+Xyf/Q
LVtPAASV0vIyL3Oi7ALaAFm1pbZwHRPUnBphtkyvpo2sCWw6nuHBwO8UhsoXNFRR
nyPzJ9CeukDqH05izCeePx1soEH3CKWl7R0SPq7/GJuYigBPHbYOrMJAdFwFhej0
Yx0jI+/Q9MyKkyURBLEMC9tmaynGiXxkBdniSqs5KRHceSD0hnvFroySRT+iXsK8
Z09j2AyeRV8NXx694TeBKqW6dCKDNg04rEU+H/GpAccrm8aUsDPLS8MeX6PT/JYw
o+XUUQ/jgnkmPTyNmJ5S8TsRfLqPbT4NYnBqPfZSqgILJe+pHCCIT8QwdSDX9GOF
UZVixAh1yGLRraSTKL8NLiJ6X8/dVlCByr66SryQhjw=
`pragma protect end_protected
