`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sAhLpg20C+eoRBnvnq5k9gBkdR169thI2LKfCTKQ2hK4ah6/bcC+m3lev/6B5uyr
5XYpZDg227jXmO093Wx28vkpVNpwhQRcLZ0G8zIvAw/q5q5ltc6sNcL7XMrKBkp5
gujbd8AcLOAu9nV2Gs+3WU/F7UKhZ4rH+ZBnkrU8fno=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46192)
tsgKOhXhTvQQEvxPljtK2Li5nQU9kiRk0Iy16LvNFapTs3mR48Ceo0PlD7YGnR1I
RAeJadJdgNWvBjD64B09rqfZHxonTMlQp6EKMeXRXxPq9dIp/c1RxIvpfgd7SxkK
jD88bjRXdf9/egJ5jsdVyk5RdE0139tKgrEpX2Uws3p+68Zl4GUApRySqPv1b8wC
0aZ4EScSQvAY6JA4qwUFEsQPkjNgvq5YM+Z2wjYHKUPqZrRZoACNjcP6CRPP23nW
psmeL7FkRhVLvZ/Oa2T7i1r4kLtIlWIny/whiNza4k9ctqB4XEqknNuYGAohp8Hf
9B1UhXectGIU23ZaBDdsL15F0nC4K0a5I1s8lm09U/sjsZOJsmCcgpr9XjVeYxY7
0KKYoITg6ejjpI6/2UqnHNcMA0IowkyVIBG1mHIrB6pXp2AYJcCr96HrSXWVru3U
Gad1cw9nfEMtq2zHjclfpvjWdwiUC8bpQiABxoDFYKs4jeI6Gd6EKC+Prbu0WIgZ
3WfBhnC4AeTZL4L17OKwnFhC3+ak57wDJwIh+XQabNZUmxA1D7O+LFZXu/EuVAvF
odiHNGVTzMBUYJku4eM6EzlL1dTgLHQbuVY5OV3Z3KrmHudERb0BXjC8z93ONHnh
o++fukyqtlCTwWkaPfWco3Uyd8QFzupRv3eAQYUrVYqbN4ia83HE03qd0Arxlum+
CuRgFTkFnviO9M0YUbWV0B85GLN6RsdGBClheuqbz7wzSlb+nBjfcVygr224TANc
NeCE/I9RgQqjZgoVHBizSb2TRErJhMUSi5DNlbb1KqBxubNJfjkiwyEudBqspmxF
tfwsbkmyjBHJ1UwJVQ6vmLTjNEmqeMHUtUoxlCPCvcfmblfCCFJYWLaMaxT++vxB
Y//QM3cu2RwMtB9EWIGwjMO7cXPqvil+jlNgK8h5sFVpmx4TDWcehuOlEgvp7YG6
a9Q4gvM31jsGymQxOkw1n3c/gjfZOSHWji3yYxY6UA5n90SRYIl9c/HBA+EpZ3NU
9DyO96HNmnlHchuV9WeBV626oToL29ZkXSsLU4Io8SYik4+kTUBohGrO/25hnLw8
5KuyFrzqVIKUy7tEgSRT8/mI+2qfKoLNPHXtJz0R3b8lPHTeKE0t/bM6hLMlOi1B
345V6gqA04Guq6cX6Vlpp/YIrAkyKr9q4C13LNEydYIQH8DFP7BnmiAyM6ajNjoh
osbBC/80sGgZPgmTGAidUsl4+AcMmln0cJYRBR/VM7t7xzF+EeFV0NUc2eUt7mDH
edF9XZcPkJlbKSz0jk6qI9UVx01o3Cw4iNRhL6sguz1tNv71cXKzxS8DNHlBp6Ya
Ab1FX821db3nNLBkGdefROoiZOd2BYygoh8n0l4LovgFAYIpJgZ0LiXSDBLewo97
Dd9ER8MqZKYXSzXS/MQYB6up9rd2WvxHtv+Q6dRI2Hk47Xq9KCHd9MiyfcwJfxH3
ez1madg5gn5HZz4zsPfX5CKlJ23tGGCKxcLvU7eiceDysdT5HD8SeQYZlPeTNpac
NPUSLK8lUcj/GZMEu+uK8uO6Tz+CSm3Ms0wyZFhnV5fhm7FpJV4kD2K9F/iz8wjB
v85wN4XMZUZ4ueRdiuwAQCuLzEoeCdXPsVWY76jKpbqRI/SejhwIzwLKGuQEc2zX
EPZZAXWxH9TSKKZZu1qvqrHxeO3mXvgJbxFjpRjkzzIo0gilRT6MgyurpCrO3pFy
tPNoITfWjTxbZMz+6/jgUawKHGWS+O8i3UaPievcNuBCX8MZ9lxwWLDrdxIy5tyG
b5PML20TXxR/oHiwUVHk6an9udVolFgcJWngJeVh7+Pght8/WUkDvIPmarxqwqmt
3BFDou/4s4xtozhSaOWxi5R+kjabCjXo1LqjJBdvYtmEc6Wek5SSOD3Gz6CjrM61
ra0/D2N32C8fBSP/2ytAM+7w9Ysc1o98vF8FR4pyvLlnItJSsusV2ViwZcunzoOj
Sk/yiYTPif4BeL+1clRW2TrfQoYBnp7Mu8qkl/7/IebcJnMkMAQQR0wBH+afovoa
PP+YQVdOd6AmtK4mRzw9ayXeiSXBrPcJQFa5tt9ZRnzTjtGCTcR1Id6MiboGTlXL
z2F15zEkQ3NpBMX93u2+xDt66KjyDYFZIKQ3yhEaWSgOK1fkrZmx+9GnyA/bQG/+
9dxPV/bMzNaHccbPIzHJb3US/0+OEKuo+K/rZ9G0Ls4SLT0pM7wrt5d+yRns8JQp
VsO7GmIAqssPcSBWkZvsgU8otekYhtQO0TNytm9EI3Li4jDDnxJ+O8W7KgZ8dIC7
45sj5dN7bD0x/ryDTFVHTQafdgSUuaJwEdTEj5SO4X9ku+uVDO2FoKu3FDiryFLq
HR0OAkkLMxsl5F15RmD+fFzJZ8Xez0SDq0X51a+1ir9cFg8bVqkIT9NZ34RGlSMD
caaq2xjaBq+PtDCh+YqGpRs6g+YL1OzBGSMS3ZFzqJhWUGqPvUMFcTN4UB/pwsod
5rDJFfe1z4ClrOkHJ1L8rx3gP1MBZywOr7aly7ZUSqmf3wVIXGhS2bXl8mB1WIYz
HSVq1yuBC4ZfpmY9mdssI8k6ZhMyVtZeL2pspV/KWu7Zx/e+1KDSHYcqLIcBd66/
QfHlZedHNZ4KTUDUQP0GSmdw4m707yQwp3evzd7oPiUEDUxfIu3RNVZGkQ13VwJt
QKlzxIe+hrvWlPb6EOuu6E9sEtVL5ff748m9SC0Fp+DdzOP9fQR9URxDeGAHVoyC
HA/vLW+dlrsv8ggAHa6R10G5NmMCuL4S4575BhaEIvODmlmfJBEj3hpw+YJvhlnF
40dudbgQYslXt0cBhFokd/vFLePByG78OvxYAjLac4t0z0pR58xq0//MwoiJH9A+
eXRK1PWU2kaewGnT9bNe5GUMW4aM9ff2wmx360vKxORKY690v90+WA/8a612thS6
TlDYQgb51Nq5XfoDU/zB+jc93EUW3vc3GPPP7vEN43p86F6Y9GgKJwYfZHK3R8VG
xlojJCihZCzd1jJvXxMaDKhcLse3aXq6AIxJ2BkMj4geGbOWnQD7HWlruJJOadTn
u+GOdh9pBOzIJR2jaeBWlonIdZgmMeg3L38eVW3w15lM4ju0kBS+CGEH7szbuf5T
0V6/JImRTRT/3ktgMOINfaXCWToV+FyWS0g9oh3Gq27uS58bdribcICpYxGuvOgt
M7e1nHMc2oUcYMwMPvUnts7eS/yL55r+yQHn7w7S/zlyORtA6+Qi4gnpC9KRTxz3
awcaXG8/mIT1Wt9IZRa5ihngggTbDEtsWfnYjqrFcbJ8lkawQ03BA/YDk0eq3ciI
R40Bg0+C1yOYgL6Bi0RQTdqIndYAolcF15Q0h8BT5J9JvwZSvn1XIM2Bii7eY2za
lWA4AIeCvayUU90gk0lV+hQw3CUKR/JIQbpccWyJt2+c/EjVTLw7EnmnKG21sVfu
sh+vIOeih99R/Rw+H9I0cwhMkZeHywbFOYt770RciBwmY+VDbgjpj8ST1/WF9LHb
hNdpvuQNqN1gq6/xR5alpebxA8rDopRilbnYbZK4wGQXqml8smXacYtS2KFe+KVg
I0bIddBgn10Y+tzhJklrfAuGVaMlsvwFcVxYdC7UH32n4OzTFMrVs6Z3Kgx7FCne
WRRkz9RT1G4bzNN0GZzEVEOrWL/ya9T/GF1gp97uIRlgcvKQGP6RBkX/3n/S1pCC
37ojbXunypHdQ0/Sx5qtD/uvVxG8HRdxe3oGDmJu7Z4TtX3gQrKwxDUcGlYvP2EJ
Zkcve03S6d50aesm42e8sYsBQbHAL91yHSGJWADWo+atFyZqOSeEiuvfWVySAP4u
4asT66rwk61ryDQmLPlroi82IgvpgAaWupWoZRPvQbNzOp4tbxgdtRUFToIO2iBt
qTyVBrIbDMp5ubX6UpbbqhSAH4I2EKIDA678MJ5aqSKdVwnj4WDA1I4RwyWg2gl6
Mn86mSe4OqqcAxAnsvSL1L0xm1qucoAw0Zs1o+1n8vH1p+TbQbev2bCJttWdg2T4
arPBnZmic/BUU+I6cZs8sHq8e5GYJqjyrNvc1DQzxh/Gflm14O9b/pyutyBDU+RG
cdsVO1wGLyRpbbYUls3mimCm4BHe8uwsIYZMZzYjpt5tfeN+N4MkXer9CW87jr1Q
pqWT+Ztlv0XRFnoX+qgw1RLJvX0KQp0zkm4HHN3MFkyJIa8AihWtCxI7iPP1vIHy
ebDPB3Nx8fCnXDORGr36ehRm8lnrXvmZdyeCTqWLT78W9GsAwD8sapEXiu9QlBe3
gI2hNUpImGifA2xXsSR3DJkjt57Gu/ogv25z+Obp31WGrUITW0p5TIzyNVK/y0mn
QCg4iImA4/1iByG0kd2D8TABut+kFSmf5h8kvsv9/oJvtBJaAEhQ5vFPPOB9odXe
5xmq2lsX5K6cbjkwrOScfUzB4PnCFl25V1qDoph+qUx8TGh1W6QFpMj86sirBaIy
sPrnS+iDQ5rvp7k8h9opQriWZpIN8LB8VLtOpO4vJnS3ic+Q9VLsnJ3kPx7oZvTV
wrP2rTmiIqhm2Rwzrrzz4JLUAOnYM+69KvoBPFeacSQk7lpXm465MDSpc8SLwChv
55t7kq3VNMhz5ZCVsIPUD07B/bLMzQ4DemRVPrUT5W+wB5B/OxwZ8muX+sEwY6cM
zZzd7Qo1gv1CplxdxA0/YS+0mKAxqWwZsbbI/sVsWURyhV8hfZvrHCo6gTzipk/w
TZzlTo5z6Sg838WWFE481aNJPDZNGkoUWdbhauR9ifNiSV3b6Sq+EFG7VPZjEM4W
W6wr84Ty/S7OifI7mehbw8Vin1RN5by8BYt4ZE/lmrTHqo/nW/AdQznQO3iGBZ0l
OnZNqerGUXAP7JUjuZa1rrc0NJblCA7Ua+e0KsGDEfiGbU8J6iRMcwjozRoMelEE
A4H+pJKgDZ41jnMHgeEYXPslaT1sEgynahkL/qmMkTU+Cc8P7e8qZC4V2OQ8/UXn
9HfI5A9W7Y8fWN0mp/BRUg8LJlTKJAfSemRsMcccjrbknLPgD8ZyUAXif31aIRY9
1G6m+paRDw1cnl7/x9lMTL9clvR85v7kcX+l1MKZQ43u2V/o5DWkpF0AbSCg/rWM
N7brHpAhRnLnbyuYZi+72/cAXt8vm9xANU8b9yRLp7MmJV07BHGo3uXKH1jM1J7b
KVGzUCyFWYfNj5RetHar1NpJJ9cg22SipRuezypB+iUbI7VYRe0aJun9j5CW5HJP
xQYx9MS92ouM4ElCzLdENdQKSRDdsRHxpk5uBAvyGZbwa9ukHtVC4UmnALSxUqvO
JSJfclGPcxD3AOEzFhKGOigH35HlqRjjcqCTvqj0DAVbTLDJ9RmNiJgmJ6lTuGgE
rKDVmZl17atTMobtDiAagv8nMdFnXVfj98UPJoRHu0FfLO1eSmIZ4IiRgoyyrPhh
/DTjdyYdxLovjOu0iuEaIQWImcZeh9UsNtLjLP2B+apugVtuy9REOkynQaeLuLYf
Mm3vpe7gkpmdUmJ3wJ1OJlsLmY4E6YD83vNFKP/US30BAI7oHBl2RTzCY50fgBWg
uj7qQim41QRU5nsLycXyXy9NoXg1n/EapbdetdEtZ3BS5PRjeExnvQJ9OSEmALmf
A3XpfTn2W/bGnsmHnOrFtZ0vEJwPdVUwRL0efueEdmJjaoL+xrKl4RbQ7Eb9kmVJ
gwYEKVVXjGPkNYFJm1zaHnFS8Fl+wtieqtUXRisN28wBCBDyOoEEtS+DO0i61Wth
wq/UAULvGFfu+tfCc9zzOs5qgv4R0CeqMyq+CB/OkLZGRC8PiUmu0Tr0YzOs3C6E
iRFUPzMJtuZEzqd1xZXTYkPBjTsni9JjC4pglJEPuo9W3/sjeEF6WWbStr5FGtzt
e9oTlzeHFJ/lfgrUWfOTGeCF9CvcuS4V0n3uteVK3FLz/xZeKa0jIfC4YvLU+Qia
5n9s0XjqXV+iPeV7YETYrYY86pVp0EZvfIWXYWieEntYGwUmEMdSkF7bpqVuGCK3
Z1EubzvXr1oetnw1t4avu5FhqULwDNxaWHDvw/fbARI9x7SBJyyi3YTIgNF83zMU
2O88nHoqq9hlO929cPbqOU7Rm+eIe4FE71N6hECGxQWs0VWEVuuVA6OXzmmePFRN
B8alc3E4kAnOHY7YElhurBww2TyGbSG/WZpjTtGeyWnpl0vY3wP/Yq1aer/Erfw8
26s48zBUpj/DsY8afD4ac6HSd8VaIm0wfwoqymdp9HtErZYXVANCQnX7vTf1m334
iLRLqwzuErN6OtjoLGlfnbg6MEjITgNwmlV9BLAhLyHWPLc02gBelWfIVDafyHKu
RpCTkR0roHcU2GKEvZL1YWCdzNH3XxVOSdZHQIi2FOe0xwsedukN3vwi62ZHjcno
sOAd/brj8xte0YzkHElTgQOa6RKCsUf/mIFheDJfPWlMP8ekyV3mlqUiBXpYxyVy
iJzZlG+N2wAfmkOBPtLVdxI82gPbijDKpmafa0KJuG95ulMh9NYxsz/vzuQdmMrx
/s1Rnf6uj282Ea/NybhSYUqXpHA4RBOmK8g8On3O/a2K8UOMyZ6EuOhaOl1TrRMs
EQqCe6UOt15rt6PKKhLp0KZY3S4ijgjsq5dV17E0sukp9j30V+ysijKbwUZ8R5MQ
HNCNlXn35iaFaNa/XFuPJnpX783kybXeFmar7Cra8ybSASbMqNPbPAXq4lXDaxX2
KJRSGTLZnTbdR5I3E8LtHYXHwOGHwh2O7PFUBZLNCEh8L9fnvDQaqWf92a+TrLt/
Bw5MlM/cdSikf8gWG4OqhlXy9VTDcJykT0U2FmovtC22qX2g7JI+Inm5xfx/+fyu
qFMabx3mVBWjZiXY7afjVqipQr2WEcymfBCJzGHUMWyL1BSvkn80f3FwRDNSFoPM
xdeR7bmlVXibmKUfRCkQ0OR+KesazBnUD3XIldwsoTymdZxBnw+I+eG0oct+xNtz
iABY546V5V+jynmaCDUFfYyOwTft8sjmPhLBBN71xTXOugT4UMHKE6cH+RPiFGhh
iDedQfy6vTBbQoQb2Yx/eijgMrWIXtdaXXkhbrYsLrTrSrd7Lbb9NXkrVPxGwWgz
Ee9lJRmAAh78MnDkeCPAgDq83g8A0302wOQSvq8YzdKAonNdWwebryxwFRvKUQw9
E2Lc+82IJonuYLRffCEN5lbFz/g+HhFkXIifYwm7FrUsb/rc2knSxehLCWJE5ZjB
Xuv2R0ADmXZYJJIC2hdeMc5u5lZObGwClfnseHWNIEtWfgLQR7/R8p9xonzBz7NG
Nkja4kOqs3F9ZztceQcab+qH9udA0RdlpdlWzjkhexhWKylTzxga8uqisrycPSCR
VuJFgGNmmdmP7RjgQprBsM/zo4pTCT3CFs76nDOPIamPeIqIsrsmzu6n1uTfvsqR
rLpnTk6tUOptNv/TP/sUtWBkBV3ybefAUjUkO6AP8qwgAHuCswUn9t27eIfOgQed
1H4Ei3oCRBklgJIWzt1uxMXaD+EDcOMA7f5+kCsjROo666FUxZoG5boCKczI4HkS
h7Cb0vNd/f6/ZTw+kv6RdO6s2tZfCG+2h9XRIaDIFLzpdb5XF1XAkOJq0XJU4uMb
q0XNiwaNvNYIURuCrl31vB/zKIw7dAK7xG559pH9YoNbY0i62U4axtiHzOa/Ovwj
pF0FlKv3OKDnf2lfGQvcR2JdMn0j2qw5YjJLQdKbJer8rjZN9boT6TC5ymgGESFp
4kfYSbR54895uwzhcloj+9cwNl1WedffvX68v5YOnQzliwV0qh60XyTlLtdWKWcs
f6bJ6/BrD6RpACt5IaqBYvhhQCsNs0ZdR1RFHw3nkvwHU7HwInNSRRyXMk6y6h6I
lvjrroZp6Y7RMLCblBVfO+fCNJQZPWi3SGR5cRGJ9tex8FUFkG6+3hOG4FCueWr+
C8PCTcMC2witNntFAwPU3zDh3F5HaXEvqt8NlHDJXxXLVp7ij6UcXVUC/Sxk2SEO
FgFYJfFVtS89x6x/leDaFcXtAl3Q4uGUfOiWItufqvLMJDeONQBXNr95B+Xfd2Pq
P2shseyi/EVIgdZqyRGpT/WVzQucW+TMzHjH+Le5yNQZRLZOLX+DBlVyHcFjSMoT
+ViWkpqoXWxKdGgTq6bgifdagU0sg+qu341pBmXtmARsC/clcSM8Zqzs9jPlwNrV
MSIHYK34hOn9acVx9l/h5aH/4SZW9hNyqfg9wWzE5gC8EG5It1ggNdPWigaFiATq
xlYh1smRHnVawXuRtMTKt/Ny1TTPObCUOJbQB2wbrlXSwY7eJvWaf4N1zCT0lNY4
ORJ6MIUa3QTteqoPgkD76PJ5magOPZrhlJ/T4Rkc45aH/dXUU9Y/LszxRpXjOBK2
+u+766/fkr2+gY6u346phRm0/mhfuiX5R0+ZPTU/+mVOctoa4ng0YJRQisYXHZED
/rZUfUDKGNo06L/iwsrjr21hOSpFcf5GmJaNquQy0pansecFfA5j4nmYdPhjlpzC
5LjwN7o0mvYcOKXqF5QThy1+0hqIQdW/072igb9Dygdf7zRpgsW2ClAS4dWPBVS/
3Nli35qdsV1Ox5guYe47ecdZk9+84pS/yQ7agVEbBgvkzuXQQIREegLZbRqJfEpQ
8yu86UaIKj2mNqEMoNedwkx62G6vvs3C6Q8y0jcrsS+3xiaZX2mAoz6MVnQrybg9
hf7dtfmKbO5Yw8XI0ad80VwpmkpliiIzcymFb/WZGY/+QkgomQ1vMrq3X443Vp6+
Foy3A93e0n4nlLMYHkRQZDcAg0bDUexqqQyYfk5y56j1LiIvH9VHgRqRGeEP6eom
5VtaDEmKepV4HTqfmtiHU6mzof5B6MQGRJtLJFY7LXZAioVub+A8+dw1bRh3eaiF
FFHslCtHqjJfE+dENPfw4MCyq9eO/68fU9WSPsRT5FiCPwiNmaAU6NUXxYD/LsuL
/XjDFIB/uThWWG28gkedAVQ6RtwNxc1vq+5ta5pIk8Wy3d02wki0sc0olXoyF7ug
A2MGD+Em3NPBeGlC2JPrvwmrBG5xZe0bprDKsxgitEKLTYpFUQEW9e+SRlJkMqfp
sY8/jaZ2XGFCl9hmaPosFqrSnWKdab1MnDcdzzDUVxdxx4/Qm2hnf+sQuHF9kjFq
ReP5s9TYm+DS/vQBPAPnuWaMpG312c41Wnnf4yvOgODhKv9ikgJ45w1O419ojaaa
9PZgV7JV9Z69NLwhP23/m0OREx0xzbuBk2Kaz4+VxaLZReazo0ig5aUL4GOrc8zO
zjrS/f+/xatmjOWIlydKtRByMClrbMsuwi4xYNOvYuVHPDY1atG5R1hqfF1fMws+
lY5U3lGe6ES5JZmBSW62e27F54TPI7nhRsNCBTO1TzupGor1P2kwoY1Q4QvRV2R4
KPWZvBs8iMPaJcHYJmfekyVGiaa/eRmGMGHezK7v6UJQe/LuJ/OqL2o1j5VJaFQO
uDWaJt17fM6J0/cbyfIhTpuYe763212pqqndv6PTe2Jkpwupf030uRILzKpkxU4j
bT69ELaUPQayzqGDtZU+aESyOTNC4+lrKC2am7IdPkldbTuYozKelOx+HksL4vR6
5VakyArzD0Ut15s1Jj2Xe93k0wzZ/hba5XepyrI4biDcpqRGLpZFTxCmfNPBHR4e
fvB3lJrjt9WGRA6WVQRorImBeNs1k5vyd4iOBg8wfOu3u0xdA9J0eV0A5fHEIGwk
V1kS64CzK7MJxV/NK3WK4N/zx7oPQtL70KTLqtAefoaU/EW9sNHWmx4FeTtK8GZS
UPXta1VYTkaN3EmZYpyJn08LWoE13L0ngRUr4ASkSi86caS4Dto9tmHJYzXuXmBa
Lwsd5SmI9nKP8yCmWjSCO727kX49VIsITaX5KNY1nQEXqP9kPDRsN14yIuKoQeXz
t2Lj31zC4hcwiiHs5n9seSDPdLu6b4esJEEkgcsbfM613HwD8ZhaHg31ONviiPQj
P/ZGgBfII2xY6GfjreXuhxZMjcaqd8iKA/MWQqifWUbt5hmwvSTVMN9+tEoYmNXk
CwMgjUxAqLos4QNH2RiHsY4CWQxU4dfIGaTkbuIl0pXUNjalWNTBpGR2rQoZpZb8
2PHixfklHH5522oGHmrF9KVe25vtabm1qZ8OAFFIu3lnwZTFVGRH+EeAISPmiZY0
bY1LJA8swmM7QjtQSpFRYG7G5j8Phog5tCMfkI1cVLFVoLnRTio/CRPyeFL/Ghps
Q03I2LX/Y+qttP1H6rnpIZuvjP96STV53q0DDlaDVVkhuBu5F5HbJMNpWVQHzpko
lMNWl6kLrGTo1zuJQXcEs5lfo7osyrb3XWto0fR+fBhTx0/BEdC4fEWVsbuNbb/o
XI/jFBh647TZxTkhZufnASNbQ3zzHjmILjjKlvlhz7QCyZVjNGTvCDClCQKUQg96
rKWTbJt2OIZq/RxKm2Ot+7F9+x+bftrvlpZms2hSvITwchF/V81jG24kM+DPAaF9
0S7TyEWBWLMSFQF+rWuXyonh7zo+SaDa7Sk8t4ay3kWrdwlIjThinY56hbFEMgwH
i5IlhXd559BGT+I01A3tHsiOtXgfMwXRF0XELqrcQghHf9c4CPNXt+1EYhF4iQo2
wPN82kKPlShr7mBJ+Cqz5gXDDwMsmAjeXmjv3QxBw/toaoFyGIgwJdeXSG2HBmKx
cPEyQJm69C3jpBk7NHHcLDNvqcll0LKhDsF47spZgqTCUWUnrLWi6chvQW4XrJwa
3zEpwHE2+qoVDbpUJfQvjRCY4GveCAk91JnAR9+uCuF34gDyqHUgxTvqqItUbhEO
mXTemJz+C7LPI1GxCOV/2nkCHLJM7K5Zu+DAs8dNUyW0rcsRkCwsOh6MMTS5IAYe
RTNaGTJ1q1uiY3p/iuFBRwcxnxH1Pxl1K9iFmC7akzINYzm3d/4Ma2kZkuOVwlKa
UjSHooHnOg31nt4ElQZ5xtXkq5vQPWHVhh9YHpL0C5wftjm/j0UlxNVCs/BlkoW4
nHgvd8xVtn+wWRLDd4m2ACurefvim18hzy0+tnWwtZE+IDDpIj9B2JPbqeqs70ou
UIDMQWo3xCv8bpAgiJxaunJOmljwBmC57/hRRthfNvOj5Wf+8tg9hknxlnF76vzy
0kR0jxwssXe2xkCiK6HogamRtkeGetuFq1tqNQetIAsfg+rz1wvmkV/yMXt6oA44
c4FBwfov2kBkD1jHeYGhFjR9urh1kDUugX5uaD18Fpg6AuJKYcdA0utYJ91Mrc+R
5FApr35hhtvM4O7qjTwJVNwzmLVZ79sSZOT4b7Kk63JowQcKTy/rE9pmDuNianVt
qQPYlk0mz+3lzQtrVStRvViEeZtJrejXsQ4G/EAmu05l7Xust69h5c5spmrsE5vO
8iyD/t4/sGzkLAI7xCdbfHE1saF0gx8jXyEtQYkEomsXMRMGS4P3h6YNWSj1KsLt
zsBAE19nnlu93bMPD+yfsPMPNDCo7gwyfGLJ4sv+zZBekv/6lf9AE2a/VnvhmAvm
EKv3BibY4XFZp4XnNZgbsrGUMRp/jysh4P23IE6jTCKZbcDOulpZEvd2+GpPTH9R
p5SwvfJy3y4q8CiOc4QAvYS9I55TFMrvJI9IoLMDY06O5uyfaDpbGKOBxcxVyzrK
g7Vr0VeLnmjY+m2Zhvr982Yg0R0P6Em3Lje2bYOan33oyQ5wYDTHGoH36IwQ36Z6
f5PxPUUpkIHfXBkRG1v9SjH9DO/C0WjBJzLMuShWP1WLH2W6Vdo5S1rxqPEr8hxH
pKK8/zidN8ukPzvNLf9WEUxJA5QqGi2m92qi/lGEsCescsVOlqaEzb1m5KiA1/EC
Xfsgr8vE/d2UmKJJHFdiaZD1QPWz9GORsV0o2PBPsQhznQAoul3Svd+0tqnBsjiO
RwRuQ2uFt0+1KeXy+ONDHqKRJROtvQkVTwFGcIzZDici2kFVvnZmLZHGewCeVVm4
x+H5zq0kEenreuOJM8zVWXMENaQ13eUtc68cPnt2qauqHuqynUmPUx8ui/nZdcoi
kdYscHFT4Q1TSnzF7VAxBYZ3bS64z96bRr+SEF6CdAwLLJCI6XG8yNTjfhlrrdDs
bfgNsRNBVidcy81/zVrCfg+u8fDxkuslGz39GiFy08EBDl3oBs6/s+A5IzHKt025
WEst2m20TXaROUlJe1wV0f5+mKrTZddGjDsGWyVKk8zdrGr+sF3CEcgWtCbONmaJ
EvvjXckzQfkCLJtRH5Prlg7e1k6mlLHdJ3/jVLhx01vAzlvKHE8EqiCVyQq8FI2n
DZYQ69/lQdGyHRzcCIs7ZTzGsGTeWIDOjTCqKwBKPrns0j4gR2aVGG9MBAjeDzGa
6UFGyrOQ4R3cLtpOfbN3HoUGZrFq3I/deutpNg7dH9L0MjAiGhFcaQRTpZxyn8jh
Z/I8xrRxq5fHYCEHqzNkisTEcPc0UXiNMZETP1JKLoXLDRGXu8lXxrToCq6JaTRX
7CwQxIHm01IUMCHAbqxF41Z6QJWdzbWxdaKaAGSYytVkyP+0aSC/BVGS2okA8F/b
SVWZlWE5paaOLULz08imma6JVwXTFgSlrNHuCjPiMNKe8698ypdIRml3qF0dtW/j
YCJVdWViKmxcpjeDNKk0Y8GgkYxxD2Wb5kHGCh9AtFMzOLH1yGC043lrb80SOHda
KPWja9K8BOcZrozX7SLapb++jmiT1+zTOWOhHuqhX0NxDcoLQkKKlZRstmJH3hKk
hsWTmOGa4i3ub9uPydp7t9/HuI42FfQ4n4dRO+S9NTWk0R9zN38LQS9mIOkx0tHC
zAMiI2CtIixH2yLMepqFR64EisA0uDL3/gEGjkM5es7COxwQSEJCjJNYz8Y3txGL
fIVzVP44Zfw2LzGGE9+Y9O8XSJfrcsq/DH3306cm4Dd5q6wxRDVpuQ0U84gkxgVi
kxrSs83FZBFmNES+eNmXaLXL6zeFE4gSc3dVwNHi52Jrd8DDx8ZB9CgbdtR31Eqc
/JBfU1F7yLKrsanzuXKB2pQJcuTEVrcq6rsQkmUVBJT7e2llHr1rZJdKrtAGVrh+
T8dr4EycjTlrmOXjzh60Z5YDFM/OmeLCRne/snF6+2SZOiv+Z4w+okDUwp7MuR8F
f4yRSFiVteIm1A98S2BVDL6izd3yDpoU43NyiPzQoxRVinyQs8QfbxP9rK6mGJ+9
kN6yiXtRGDtGd1awEuqKjyI7qbtOtLD4qS5aKFkfVdBsnWjDUNBMP8F1EFK92rx5
sIq+kx+Re+ouuWE2pGmNFoYRlFDwV8Xx8cOeDWHzpqyD/PLJUnJ04cAHNAzCx1d1
fYBJu8BVT8LrGKrrs6PgYBMRHUNNMo23aHAYcWnL6pj/yQlZMXpoZOBz1cmyiBMK
bSqDg2pvREbGM9wZEdfQnE+QnYbqZG6IkYjSQkfRpqmRe5egreayAJnT0Hv7IZib
3p0JZIA9HLSUP3k+eKaxTiHMLf8bSjjbTgZX20pOJWzoLSiFFXOkh1f9rtFe7pK8
TV7ZfqJkU+Oz/xMvyQhcnixnMKh6Eb+I7AVxn31gjEEUS1ULKQ67WbQ2a2OXvn12
n136fY/6lHAB/ueZm3LOcgMo7JtvUYUsW2k9NyiEyTySExVAiEg3KJZYWgU8b6f9
GHyQRk9TzE03gHJibklXoRzScizS2YYbkvbaFSMqRh1cpCZC/FqmLNCqy1hDM4Ky
GEVZ86IfJxIkXMhPcNRvVikZivb05d7LHazp5oWEBYOJwSdmnuZY3r/Zzdhk7aeO
/8DCgr8aXlrnJo7ZhVtrAYlVq7F0GGWRbSjXMFx9nchQuwzJfVxoTcrqA1beKrTo
RhaNbbB7tSAmIDn5LoNGdAgDiuM8nLU7+S/kKl0ZqzlwKcDEfs1IaGWvh+alM/nx
gFVidEYwaHlRq4pI6/wwChzu34zvAH4Gaj1t/q0xr7k2L4gRp8+9Cl7TMhgXtw5a
/80GgxzRyLeOFDd2qQ+fNOooVa0d89QyhhahkgBfncN0Z9b/nFvveoFKVPJ/KN2/
WkP5/wvWjMCEcTWdiZMvTnKx7ko9u7o8roWVha5NWI7lx5i/liImReL0Vk+U8Sfa
OKg2IA7OeB0WV0SOy56d8FF/2/q/wSj4wo1pGCzaunLRJuC7DvI5gR+T1o/5D0vT
oL6yiQokDLmScUUEfkmK8Y8/8lP54cmaWVrylRvRsdgzWn8i1zEQ5w9/RQfjRj4u
9NfsmKQbfr+4ADb/xge11RZv5egHdje2cuHVX0O9m9J9sTz9ZdNWHEgBVkJomwg6
cNhgyEc+jUbz2Cy6mF+SBT518rQqusuJLqL5/N2YXsFnfa2RAKFpfKtoCz5oIKNh
NR2nfwQ0A95D73sOEMSkJTQJ2FpWPxkv9pCotVcWgoHaDdzG2r0HvEojLpIaLXEX
x9XDlrzln6PXql+OxWM+mmffeAse+QbD9XozS5+rRgA6d271w+muIaKmLLtlzEaR
Rsqxow9/kc6qT6//pWEq0/NwqWmjmtt8Je96NMkVFT6zcY/8aqhPG5tsZAUH9fAp
ji/Ic4fZVhoCg++BEstyHdMafcNgj3CtzWb6zK7Nul5AhySsNMnQt8K0IRhVn18H
nC/XXcspQ73YpsHBXgd0AkTjYRIPrvRTKPi6WISDn76CG12Voh1OLbinn9y+y2Pm
OaZC6JQxKaczWIhHfANVW4bZa1NH1TFawtI0k/gaNcC0X2T/CzQ5IJfkXhrWpDqK
Wls8vHS1kHSZNRW3ZWTNLSY9ggcG+psCPpMMH6b21qc83lD7PqnHeVqVNhB1M5vo
h0+pn//KWNLsDV8I6v/XMZHBKb4yvrZEu8VpOQL9OFHIQ1KgN71X3cMwa0fy3tHm
cD74FgGv6B2vzGv9fq4iyPrI4PGBY8rBaaYYxpmqAsberFjEUfjpwOqeIPhpSToR
CX/pvecxy6/Yhw2oPOTJVBzQfaHphkGKwGEwwMGRq07pZ4eiDeNbFBFfyJjt6IcW
NkHpQNxC6PUSvBW1eQyp3Gg/T0AlCW833LKkPOUrkXz9s7c7nGF3PToqrBubUA/f
5BWtE7HpiOPfbmMVU6wwuiDPEP5HmYDbjGsYaquJB3wdR9eeKtwS3b9QXkAHvv3Q
SrgTBBHR7n3xNMv+mbyNiDNgo45J2YcFDBmOIgo3g5PtXuDDIxfWxxP8uaWCGCpY
/K3mqjOyMI3BP6hqcifiKY8k5hvKPVGeLP7q3B8JsDmBcPGyzJZPs/597VbuT9ud
xJ+p4vFmpM+sl7Fv56QKoqjgzm1l3DahCDq0QVkoPQ/hYGMrcX/ELq0xsnOIZCPA
u4CrKYqLp4hp2Kcm1RmCutE6kFRIoH0DJG6MV+If47I/XClCRzOIXutBns06b+kC
mooepF6d9tUMcaygwG/cUiE/bOZ7KLRGaZvzKWSGrv/X5yWCHky4oyvTwbj4UIoU
wtH7YwCn27GTJSdeGRFJXoZ34s6qBUTfUMm9t6c38U+e4Jk0bMJgIr3iJoKC/PL8
6aheijjtl50Q92rSg4aztRAqec4P6AJgxxmVvKPxvpkmmZQZuyMCVcG5NMvbSE/j
mYPgtlYic0XsxjTcU4NNMVROq59aDmxyc0RMj43e5yBhD4Sc//ZsssfjSCkzlYNw
AG0RfjzDGW1DebxZdMnZSzfE5HkNpSMEVobq+scrZWMrGaUFUznGQteLcmZbTn7w
1H/fjrSrmUDvE3V8J22DgVsBkvo1W5qr+V9mAxI6HyhdroOwV4aZ57bycWWaYCwn
3nC2cT5Bz4x4crwFV4l0az81b7LULGiVmEkqUaA/1fsRXkNiB04FcI62d+rOm3Hr
1D40MDYhmCc353Bc91CT4zNU+EckGoDKbdOGFIWe9w3Evj073eEiA7litj7U6yzp
H49dmV4EyNbUjtx0aoK5Xu2mRByBpYXye2T/CS1vkTOs6p1sbw/Z42GU2JRgCpOQ
0y6A2+Ez8uEFnFIJkSzN+W56rWMbiNJYd5XU/pOdEfCYNfqQitiQNwndLtNyNXal
qfrR3FhQjNnldjwlfZ5JtyepA9yquy52i/Jnlm9KkAfwgtxSnUBNfuF0FoTk2Vh+
OP07gn50OYTiUlFcAIOL6jLZfSmnftKSZRIfvEF5Qbdh6ZoAl13laoLXmyUm2O+X
IzqM3uDgCwto4XX/hHwvNGzvpbPsglNZ7YMTnkXTJ/r9/6WKEbWnfKyDfieg72K+
w2vcGlL4D9VaSWdR43bzYIfjVpXczNVanMtb02s14/OjH9pSAonSXIUgn3M3Iar5
BO/1PnCdTpJhFrhoHEaODZK/LI3oukOQy13IXoMP3keO7QcSyqFqonVnQ0wxi9nS
kt5Ak/brjMikxxZmfMXHNYjnmm3KrXrhoOfrE4Se5P9/prGSUbRDgAUV7ufb6fzx
I82M6rI3prQOo4fFB3Xt+gyRX8rlVzBGvW8TeFSLzlzN0Eb94naNRkaJM/UXkxys
6vWcYUEzJ77GjLeJXIwiR+N0UMWmWNktnAJVrRqds6Bgia/YyuFLhPkZY+AIF3jb
vc6imxh6ezhPKrgA4HeTLsmich1jPirIT88NiSVjSmDhZlp3OqTWrFkS2dOYPFxn
0qFCcakGn4Ktwv4m6N1CmgKA0RhLk8FWQLw4vHRFiHOKhY2CwVjD0f2X8xwNuyaZ
R2PtQ57SHb7OAzlEqK/M8l0RCDBQLbW0+6mJxZ5izF9QQX565xA83W5CkojeF0Fg
O/rUrkvN5q4GBIET1Htn9z0LvKqrvDMWoxpMLiigZ0L6HoPHUeLP3emhfMNjSdCv
KQB3bksgBbSUkEBVk8bNPqMn3s4XmMu+QfvGZwOgd9bn5Ppv5UpMppqjcqdeY/PE
9fTaBma4i6PLzoP85yrXW6VKYsgUQhRT/ZY39t5PQlqqSwZ9slPSd20aFPKb1pJc
CDVVdf3opnRxo/ai6BeffkFAdtKzU/0p7M0odP8pt/ViVr8Vruj537S5yEjNZUBQ
NjL13FVq3gxtg08D0KRPIMFGuu8yTL6Y47IY9S8LGPWRt84zihSp2Xxo5FUjL8si
jBq1kCGe73dFhS4BZf1n/Xafk/Zv9iYu1dQTTVUPs+qbQUwRySJccBuECRDwXyJX
YiWKc3xLEnWpECGUsHf+IUGZNARhcYgPYGJGdUhEsA99Rr3O1jhwWqAcfva32PjG
p7q8PgEaRh6j9nugR5GDGWnqkaoNTfNCC14a0V6XbOEwlzvp98UTpoZsWkx9PRQx
AQ6uAYowW9oWw7mOPUaZpn3ty9/RAaVQ0sBtNz9A8bKSwPhUKveAGOCsiSKdSuMH
SdKoVBcwbK7k8Vx/yYjTV/aGhj9WCYBjxV4fmH8urBaiap7CTAWYmjMt1NCTJndQ
Fi3yz7gnXtGf7ggUwqz5xlZ2haAKSUgF5v9Wosk1JRFA11eR1iVLpP5Bmd+Ftwue
dFh4EAlBj01FRrD56nbpiK9Q5pJAc97AGbQHbdEkj2c7UGWuR5NUl/U75IKABY5R
40Q86+cXlAQv9mLBolvD7Jly0NX8MCgS6LmbgJAi9C2RIFnGMXfp1CJdZiAsIbAJ
/sQLX1Hr0j3g/Z/IWyGUgi/E2yNw5jCsM2VYOsuVNqRA/Ygkc5uM2OKopIvKJGD1
V8856qlMDPkeDjHGiN1Sis/3usj1J3ClU7EfS0MRl0dXG1vLm480fZXAbQJihtcS
GThDgvKVsCXqN9lE/I1oL4omlePRAGkzXp2KtUu0Zp00E7H6UJpetyvBndHIvt/h
BjCWfH1JJ6xrpTfrL2idAKB/ZrMEaJl4xEhdU2ZwZc12OT1HNn5IIlSLN2vzZsld
SsV7quo31ugrkWwPHlL37dNq4XhwVT/55nKQdfyDfNgeh5YCvRug+bZW8NN41zdi
+QSx13X0pQJ+GmpgA2T3i99yFUEE1+6VeVuYU2WtEfIaWDwxoBEwuhruc5qfdwTw
gcSGbTTr9aAgJ6jSUqTMZ2ajJD76Gb+3rh2zI45I2VMmzBvt1qeFHcJpmhHcunzN
oveFlLKLc72fMcDum7p1tV051Gw+2dzWh9DXL0VX7y32nHk0TrElY12hqQEbVF+6
uOe5LDHTd4OvVFMrYSlfAe9cCP3vMn5/kvBQSj8U+ZTmTjXolYVjE05sNVxpW+5m
nCnIoqV1KlmLYGnWlE58EbU3asfLyFUFiYn+GFNdtRxY3nCycppQgGWclUfanDmU
Lb9/LAbOxJWcZ/te4+VSGAN0Kb/sH6fEa5HkhWr8dCnke5nrK4Ws4PXAHkDksurw
SCwneeSh/EBDbecHiEl4846sl4/qNBKdgNdGi7hxa/d0g5aJXtiJsFTlhZgPEyq1
AiRyLezL6GmM02hBfWVjogZZGjGL2KjUhVPaKGnc5+vvMJLTQhYbUwQk3SpUdAHo
EK/6D4riYsb6ytC1s02MF6UMe+GEeODss7pN2DyOjfIyOrNX+634E+eA9gYIz3Mz
g764kmj6z+DNODsb7fC1LXE1pqWhmr9H6y8EPEQPkpO7d9I1/qXZgB30mNCQ7zY/
2nEonX98P8x8aMWEBL8hvYuL6sOqNRwFCay06g/YxwFhoIWY3xZd16b+91cDINMy
F8MKgAREELJ/0WlYhMLXJWON3GYmYTe6nR6yamaqFrP+YWHtrqIb5sfOykkvnjpj
Un0Kgn7R91MtevZwcsHFWMjibWEbmTpcQRptsDI+eicKEUEEEMBoBQWv7Pep9Vmf
WX+sqtICV/TM8srv8Rg3Mu0SWKdnyhkk49ieL8GdVdQ2hbGXr3DS2kTVKKIix6hB
UUHK30e+l+A2zKqZLtHfXDO2cZLsVAdLuPHTdTj9e9Td9v9cNTMPRuNP2bqiGe4E
jZdDxSYWfmdlwe8DXG1+xRLarARvu+WAkJKyEVSOPhVANL+BKzk8fFgN9nfcI37V
VEfwctcKl0kBu8lkwh+7NtVFFmHFJkjLRKJBf5ZeeHQTSfIVXR45M7mozNumehz9
ojOe8nXmu+uRHaSFMEXaYZ4hR9SsWkc4iFoFJxT7yBY4TdvN8+6NM2Ca9bIi0rYx
20w6GomoYFffnXAYdtcFyp4qdx35umD0p2I2WLwKXenINaa1ncax7buGD4t24oML
JjEnhpb/ADfUyvpqNsEHkaI2a1tlcY0VM/aH2+g2fk2J5imawah4nQTiGUkOsV33
DyISePW2EwKDnOymUZjefsiJV/2pGRPNYr1zCqzL67J2fjtVDMr+EflrVF8YRTSW
sGqjUoVrF6v09gJ7C/o7TZsKGIqOIjD24VtH8iejO0UErbs/NtpPlLcIsMW2PWt8
epBlB+8RTf90safI+5Qlmi0o7Ih/vIWVpKIaYQMvgH2/XLWnMaRDkckz1dt88GpN
j/h92SKXdZyfu1KHhOkLKIZZF9Ch6H7CtC/lXTWgHsQfQDWfbcTvohQoIwLP5G65
gKzLaME5JNZD+oXnXxPnQ2DxGMKkGjIaEYxDhK/5r5wr0i2MVuimBas84QYrhsTC
2wB/x9j+Iy6qxZZvuK/56QnDRdggp7+57HN0SdfpaO3IIfLPjvHzeVET/4YOGa/P
AhFb0XX7Q5YMHAcbc/kWU/h4gy/gLxzf3obsEEGkO3d2uuNxHVZ0N433r2zivmID
9MhowQABCmw9/M0jqS7IBKD4YRVuKQX0elMZgbV0gWJ5t81mjGnSPniUzbF9Y8zC
jSi/4BKSHEyuhUXIFs58HW5phfCayFSGwrzcdElT3yxny9EiJqdeYbDCll6U1pGh
PX/oPY/XI/XOWYT6dqGlK1qJNqpRsakYDax+llA+Ow4zlFwVJtXwTrVG3wpoYxey
DI854a6q89xCguuFKiS0vrlWybDffwmQndaSztF0RD+bJskixioRxsKmJ3c/bXYv
2W7o/yK/0/U8ghatmNMdmkdxmq3BuSgGWBFi3J3GwUXP3FVl0sn55NRiSOnw5our
PBeCh48RVcZ7Ud2J5ocXpAyBY9CPDlw7TA+gHtlUrbFjWl7O4dok81goVqMzP8Qq
Dgv2w+VQSQdEJ6VrweyzhZk2QS5jbx7Sb/hZ8DXgadrUu/uKl6iHqGCuhAjWnQ6O
LtajRRyi6m8ZK5phzLe3LCKModocKf1EOmm5oz0s/18Kd6oQgCzKE7htIgq99d8r
ZwoCp0HwdmZpzhbJklsO10AbSm8ea2JsXTTraosDsDe+uyQQl2D15QVLqlryqp/K
9IuoyDyI/jsnt+lKaOfMwiBad8XMJjq08WV1rr2O3bidkM3vAMz9pUGlZNsXfRAH
Td4WRUB5vmGMLJSH7jKVutK4mhyUkPMfdd8smzp0NxrPvQszbSq0n4+ne+kps8PZ
K5K6d+4wRPvaXMCdOL7v2MbjWX5oa4Zx9uOZFOG3zkGM78Vr5WGLMr1fgqfWYDwr
IPeLdOzs/4N0cga8c2H0PDySw8uTgCNT09Ljo87aKBbKU5fDBFZCnzSG8duUMMW0
4FT0cAj2n9g0H72JayDpB9NjznnFfqra8QBj4ATmTV3BmN84B5iqG8c3RF8hz+tG
8MykepQAN1W7AOSB6moXwwfNeJthi4B2IFDKJ9UxOqkkQfxMs9qLkmsxrVET2L9G
y1CtKRH6QJi8WGuwnY6yVEe1hrjPvx3bD2+J1sPRQKw97ROG8utFDbN/E9HNfIys
59PITbubqSloSDDjoIDwjSYv2U9lIxrk5aOw4l789MiFAn2S8qPFkV36xJpKSoN+
+ZbeSVwlbb4HtuV9QLTzyIUYodIiYqAZOecxBjyKk+SK2/nsbbAxtLDTFuedzs3G
I5EqGLx2IoW6qfIxNeqxwc3e7fPWhKX3D1i7rXD8W1EYIn33YgFzjAmzIFHf+XeC
z/StyQfbWjXorKNvwGtCf61YMSVPOHUkWHcirOvOWNFZInVhpaaG4Uap2b4pgSs4
83SXICHIfS0xK4vgfFOlK0ECCRZD3WA9eITsHV2KKemld4SpA9LYmvF0tFUR+k6l
khmH3cY8WbXegj66RQ4lCAth1DhsClI6UPdgdjTHvtvwz08bOSLSspoDroL9b1aP
TotxCaIEn29bmsGTtpBsMZcivykCKlJPbavt5o480CkQSjxsD6KqbOQTcQdQXM2p
ap02B+02IluHpENHCYPU2k7Gt1utNzphyWkgNnRY1YYjdrdqdUhmCQxrLhEY28Ia
5QpPylh8JSVZro+ryICHzSAnVrSFtjHuYnbeuv8G384nWE6D+NUz+qVzbxKXwQgX
icxdZzHdgBBZaIgL0S8WP2xgDCfrilQzZ2SOBDwyZmxboQaP0TOKt/b8yfyRR/gM
gbYZ7fTQQ2XI4ySfWo2UqAGSrhlGL2L8Oa4fA0CIqu7hPJjGbFy0OWQ7vzW29nZP
b2TXHhCsejviwjN+iXSWXFZcHJz1hiGtgp+qVA9BQXP2MYNauH8qcpxkR/oUWC3v
skLoyN7WLVP1CBW49R3ygBKOb5xU7VZqCmk5UTupIiQBs7fs9l2xCVtG9FXwDGmf
pUCP8VDBPeaX0VMeEDZiJ/JHUgWjmIAr0Zmbbndsu5sx1h3f1F5jatClbX9cD7GB
8z4ZhOri1G51Jy/Vbb3llpAT5twOMUsz8x3ygbUKZIPaDfSYnKmMx78TEKYNi+Kw
5AFwA3uUauJaErvPnjbUl2Ecd/GF4zk31d8xDuwz1LGezgkhHm2AfE5ynIP4Odn/
isRPSd0yO6P0MToqOfwuXVY/8QwWS8GoUtXQpjT+3lyvVaNbTRCx+/y18RrY1N08
R7I5evMydCqvtx/Zj1lLKPV+1S1cymjdQYbdvNh4P6lPfKY4BA4afKw5LuDb/k2J
IptQKUUruvQXeGRwhg9mTdlGeYEb8W6fKDvVZkn1UsLQBNuKLNjcchiuGJUAdWeR
IBKps2i2DgEg4ZIyl/GJbEp1JtqXVkPtvlA9dNGU1OogHJpRAxT/zVAt6Y7WS4di
izn5eb4RwYxQe+TqE++uiZvAbecKB3Z70WMdqfy6CQ087M4JMPTkws+N4FduBIIM
ube88ddMmM6yVuLhQ30VKG25gKccCakm9CtyL8/mUVuUewE96rtvgMpMVtY0+ErG
qgleFgzwTJTLnjqbzXVByIIqRi8DDs72rrBHJQtJeP9QSGfSvoJGlcnReBAwu4iD
WHLTBhboudFtKwmqzOH21Bkl5tCaC/hrSYGYwwSsGI625CBxxcltYbXI2rtcE38f
udfzbEVqeFb/WLcDT3UjoZp7iMuErdSAAj0SoVtIfXnSfgRV8IqfuoegjAMh+GKJ
k9N/tcerozY7+WmBuedvzrk/vyjfjNQCSpCZI++Es2jwzLZqzVdqq3LhHgu0/Lv5
10Cnccm/dsOeOxf5CgEdhHQh3ivd7uX34K+oycwlsbASo5MWA4+mQTZHvR2znP0r
QNo5ejpS9DzpHFcRPL1qiqwFQwdBFWlewF64bltd+h/POZ9t21v2aNMOeDxDqF5Y
8jUzg4a/AsG0iGXdRiiLK6kfHFczGWs76mObJP6Umtx1lkxuGCd/0m1eybeEzMns
/fxYKq1LSLgvGB7xuYllBSOWk/jkwCnDr0xoLGDkupLp3byO/sckX4AzzSYVB8et
Ip8qFUfLjD3ZwkJ/ulRpeEg60vUnpBZS+bB/o9EOYzmTgYJPG04Vs1FZfa2G9Biq
j+3pzCEY4NmWWRcqZh6lptVeDV02tQNtr9QHdxKEOrEek9iVYkspYnSDGxYGgXEo
EscPtinGRi5B5+U2vtM4j4Oig30zwl1oh+DWcgwXxL9cqiTeifpqA4fNtR/HcRf8
9dx1jtBHHNhJFRmaCWqg4K45yacBzMJp+3YNVG1I5qAM6I9gK6sXVHLa4qpgxLMr
VveM9JJTCaL3nDho3ULEsnY4y31vMdETNRaU3CtvRR3x12D7Hg+BJ0gPGsQTncOO
iMEzlp59Z8UfCGRp2zrtkagyEk2uecrlTnOGvwmAs/OjqJgol+Pc9dZHd7PlTn+C
2RAhHLOjuo8E6NZ50IDl4i5lHzBFWahKKWPsu+Us+teW8N+bAwlOA+WfQK1gQr7t
UHZq8FqkyOA2QpWMx8htNAS78orZyQ5DQ1BLcA2ZaLFwS1tqyBMacD+pMrGasgV1
0VA221dswAcTKEVbMoHPUgHCTefQ2P+vig2meHRyd15k76hiZ0lHCQdAWw7W3roN
W065fka5VQW8QaxXii7XzN/lZ/jh9zTleWqXceV7BmAp2znhUfy0K/CDaf9Zotgd
1cnO3hKwIXR9k2idQeQ9OqUBVEI+C63zg/WKs39/jFtd/Cct62KlqmTo/kHrZwVa
3keUe1qh2YP0KUErwPLGdf/3UwMl8g1ZuJuY4aZ7LgKXB2AmmR9MRGV/+A2U6eNw
hmNwpFbYJ2HlvXXd+tjev4BjN7VYM2eNRgAhnOa4KDTeZDUr7Nb9lfvqpA/KHrzN
qTvgwGteklEQtpA2LHIQ0xscVOvhP56k7A4ElcOs4CYu9sf5nBgyd8M3Azz9i1/y
b7IuJ3uA6tO5DdWMS9WdnCP8K9IQFiXM2KB6yM5HW2CcNl+9sZvXH5jzVLULZOqn
Lb93yMCnj9sifU1L/Nztado4x5wjUnCmIdHf74OI68GKKaECTjIqbBAqPVXVUTr8
lKkfNeEx4Jg0ZbAZgHg2lXQexgFE4jQXLL5TV8DIdgKL/EorSoVo20iI1wFmg792
s+1cfPZayNRST8Q456tqX1Xxh6kBgGtb2vgqLeRc5BwPNAkckTG7FpTZ6Ly8QE4E
IYuMgbzeuu1Rfw2i3hzme4kxYZpIWfYiLt0gW081Nez+TjtjPlijrmPVeNe4U5Oa
HZLk5P284qNrCZ+/c3umvBKHbjEJRCNV8kgsPEU0GcUKOaBvHPuYqz3i0Yjvpoqt
LDPuYBuX7QURP+QXC6kHYWc7dfol2uZ2sZqRLl9fbL63eseXxzIGE/lhn2SEf7sY
NtB17nFp+YewdMvXGX/17/IYjS8d/4MOIaVkOBYPh26tI3empgevDJntG7Nss6o1
xiEv+Av06/rc9pATEiK/Xi1MiSC1PU0P/Bs4hPn3pK2Db1k1AniqkAjtI/rP28F9
QwgtdjnNJzHKK+2E/t87M9cjaG0CWC21p29hY9jDfUlaZDMg6q7OEdicRjLN1oqN
lNrNGv3a49/nOWKjv1MoNXpVK2Vg7TznRrPMHXNHQ0wJxaPwTMZQyZZ5xCbsthvR
60fWLaV+gUT1gOZfiW10yDgxLww3WtEYJNycvT6A4dbYQsXio95oC6amOSVWUjoe
zakT0DsmA4EcTia9THt+yFPAzvuAbi3DpYYyOYC84wxTez67NYmspXwV9hBjYZhT
XMf2dxh9cJKhZy/L70JRYLjEen2E47uR+WcLWa2Ete0oAxTDBMDuM8dGkmCL42DH
X+27uzBWkqZHony87VVcB8TfDDQL19fukqXDSICx057IM8sZSv4ulMeO4aLx61/M
Zk9p6LOpv+YPtfBfQ2l5xm29h/0s086p1uTRulL6VP56U1M4PPUxZ/nQgiwQWhsK
aAkAllOU/cejqaBXtWvWdeCgIUIoIeBPEnLwJGiEMcGWJ4nFTAok5xmrnUtLNPpj
lzriDvy6monVOZs+GNHArE393h+D34fY1ibDFrMcQeTagE/8ZFi3e5DVln6lYEzB
Sym2zEtsp3vu5pDgbJz1o4ls5ccNfHYsH3OZaMDojAOS9Yv+iaQsl9zQIuEUWCzg
3OWpNdUAC5vdt771McV6aJzU18764YdP0gUMdICUqhqEJZsiLN0CvUi6Dn+bjNrG
m6gPifOSwibLe4/+Mi2AFKpcKakSN/eP6RAWcjUQzmK6frr7tehRDKcespCuO9pV
090kCqRfcIzh8saZ2g7cXlLD9i1w3S3VkUdkVTw6SbMjcOOY7tq6vhlVETtCH76P
eNY5qo7yistlLdeQ4G7a9ghluFofI4CqghB+s5xb2VUDQuv02gK3WwhUeFPfujFB
i+uw7acLUx7AC7HdeG+6Zh50lpDmpEFX8j0Av1Q76MmUde+WGkt1o3Bkr/aodXAX
37fmGDFAyG0g3Y4e59Ea1al7pjT3RFEtr3b0Dxk/FkH8vxKMMhXidzuvjhsuq1yU
A2vuxdGR32t4GKbRwdwt9CrnTaY2t6OnqAKOCNBEi3w6fqI5GQ7ROvzpwUEZNevl
xCCYsNf8X/yGMf45f2UalyABLNHEVUqeWu+cGGIQbB2xQoZMLP/uloLEi4R0LdLZ
3tOin9L4z3DapnV4CZPHTYa+r6N87jpZ2eIAH7Y4Iuk527YsxxtpNCPmWxfmufr/
raUX4AccuaNl94X/YabMDCpj/MbfWFySYy+S6vWSGWCKLkc0wnWdsp9efY65Dz9I
o3SsaB4GVe7sepFZw3DlvObz5tv/aqbmH1tw3Ylvb1lSkrOKkIj+mpBJPbiKs5pF
KkykeZnQyN5E0zYSc2281MlApGOJyOsixt28Rcci9PibrVqVLaAnPWH+XQe42jGy
JmJp4dkdfETwKtP+ege9EZLkpO9EU09BZZjtr1Nnz8/cIKZBd9zXJUFteXwX1Y+7
7LVbr0SO2nCV6MC3YordayBo7QKAJ1cohu5/AZBkprvNmr9NJO4PG/cCn3wmF5wy
3c+IhqbQ2nBCvvjqdu9Xtu4Z+u7TGUqVLRXQnzDbqK6M+Ui3Ku2Z4GXPyAMesOP2
sJLcGRwYoophh42HyqQqIGPk9qZ3TAMGuXD4VcEnT/xFE1TpFM7Vgja1tdb8CuZ2
BXrlI29QKaYAWCgeXLBGyyigpur05ZE3zgA/WuHzaarL0N00Ny6cGBIWXYZ7doJG
tZg4DWpuFdwiyv5+/wHzVRLLW/ulDPJ81b22Q8teYiLvsWMQyRHxe864mUqBF7uA
SfUeXfY0M9aWYO4T0SC5RfZ+i2EpChmhoxqE0OTEwleI2yOb/EGhZqlBwPFHyyVm
yXZoHJjWp1u9xvswd/aVBo2fayrkZG5Hbhcr+PEYNVB8R9RBn35mFbwOj6NKgHIm
FOQMtXf4O6VXfzYFCaShPaj+xs35dbWd/CyyIVxUzX1wuvsh3LAnnTdPxn2auNoK
xzoeIIR4bBes+cbtkZHpW5Rl6FBH9W+Hri/IHlx9AE9jOIlgpjouPrmTdsK3Gr3b
tm8PvzjKETdR588x8uch5UGZmnA+W2HZSb34ozwgBo3abKStmnFeDsf5Ci1TGPQw
yLfJ8/9NG6rb9kNCO4xQA5zfddB+CU/C+itiY5xtsEiQs7/syVsPcF4+amUrZi77
jrbg99k1VG3JJO5U2pFVEXbCpuKqkOZY8qMbs2J47GBVzAhJynCRGuyBF8OdA5xp
YIFR3ovl8t6h3rPWloBMQs7RXQzTAFya62KJYZ0Sp6ykPO5CSGzW4rQPd3RU/D73
waHzFNxmhZDBeJoEUeggctnDDDfRfacMca3TYKcLf/eJrHVWI22jZy3RsMYGDLTy
CDqwb2SY8B2rqolZYdVriRbA/L5Oz3UpjdOkaLedA8FwJJAM7ep5RFjJxO5rn2rz
4ktjAGt7Yp8qjfbR22K3Ge3IRRC6qPi1zx1UPxjnzrOUkGy+9NEn1JrheieuKJjH
RSabDZoEbTvo+5mev2GAter08CQXG6h7nu6ONAaqQzK+3Fu7RTlaQrY5XSHBx1RS
mkBI51eg0pt5k1Eydd5T86W/mZG0dp9cs15ymv2KyshlRbIqjlDzZQ2e+TGjG0wL
xCcTox56qsL29wPRSFUUF0bexbAP2lE/0JQ8aqTcu5jeqJBuhTe//ttJIdPjXG4m
jvd1xSqdqkNX83tNQam44PDicZVsADFQYikmnWg+e/4yiAlkrYgyJ4J1Y7hHZRpl
f3ASO3DzUhE9rS3fAzn/czF7rvs40ujbeXJ3aLvFyUgsWrl2d4zALrXkTWFYG0x3
arBxqZvrqA9z8ztpOvYPh+MDcwlA8aX7N8f9IPf4o4VT77sRkHbe6EetJsBfCLtb
99sHqKiQBquZZGv8OnJY+nStTJS5lO8z6+2HW12E3f9tlkEqffV2kdQ7EsoheWQm
YaRpRz97pKRO7lcAQMMZjqF13+3e76YIdIl4bwTiGbwso7hzAdak+A2erQE/O0j4
UCWJwzuKh1ob4KfQOio5DpOByd7X9Km6DCUBEEn0U3sGppMJjO/j4sbYJwcVeZGS
JOQX/Mo+8RIZLsO5ocMUZZaBFqkwz3W4jpB+airbuX4FTMthbZ5dQ3st410jFNdj
g03jC7qYTkOjT7X5xZnIBmzk4ZoVlTVYUZjkTooL+mYf7Khph7hTU1s/S9TJpxH+
302jjMmLibBRHClOT/aY8KxR5POGGGok1i7UMDIUQplq8wWa+cIartId81eYrfnE
OTF9zeqBWUdU7p+gaKu1BtCo0fFRRmZDnQR/T7Di7JOXPXeBFgb2Xx7oHxt2C+4Y
91Bbm1EEcP7ZoSWEWSxBJR6YeL0eiBDn/dyU+ibqmEWKL+pQSpG/4XmJ/w+q1OOD
8fT4kXeDEc8/eB2j5pwOzUesN9L7sOy3f0jraeGBZjCgZuc2Q+QTgTw30Fwok4ac
t72ORpX4O6JQiYfZXAomzwhmNlNpIamTGlFCyi0iY1YyRhQBH678EG/Y1ImPOzz3
g+9fsz9heOQSKC7FF8nJQBvzEttuIzPeKQFThMJfv6MobsBVpIj66oc61z8/1SrM
spr69sn9m0dNCT0gvK7jwNxbOClJIu0aqyMPgpwuYacG3uy/K0OAvKvuI55CWIXD
yU03BQMwL5RM0+41kxh4TriLwwDzoxoKo0F5PsAtM5qk1c4ouFs20NxdXpMmGwPa
5YJUOSJpfpqWW4O+YiqWqqY0OepkGBAkGmqgeaw+JqqbozqJPshdru3oXJ+vq7/5
g4y72/gtHtJSuW+/a9kAAzWsGiEa7+rweznTaeHgrBYz0Xqc6dgF+A0xfAhvbFbQ
83HB7KRpWKpaU1vWzD28VxCzwaLGrTD58djg/bKLQSorXrOy6RiCJFgdetWJxd7L
LJ9ZPyhmCX9HM0RKdZYYf2dyQsJK1P0jO//rbU1+bSYf1rIuNvyVZgTRGV5BcEjT
Ip/cgwODjSOw6zw8seZGAQWrFnwReNLI8vPrnqWjeGafur9wkfYY7cb0FUNYOBCq
Qzcnco7goB+VmztUhvdC0XxssBAxSj4jAKgZvJ6LZhiD9Ogpx1FdzW+jHx/VluuN
UxCK9IfhvIxLxwSvyiuUe/QLgqPQPfEiySdh2zitk35EBpySlmAVTrvWMb3Fqv+e
/sXy9y+egy+4LkbKrkeBL8f8QdZ9fqGp6S0WplOuNqYtq78bGDLpedCWyfrF8ioY
coennuRAaVHcX4dveRbXe/sk0FqyI7OQM7eMr7rqzNAlefE/eMBWXQY33iVgPev3
iNiCp3rSmd9/BYrJ5nYyJKrtB06V/DHTRfRbClk6usQrS8fjD6K9WxVy2G6DMNrp
SiTFcADkuK8kMmHPyc8up3pTjtRawvwsygjgG9hnXHctvnLZO6A77FGLBeKXIxHQ
TBtaKvKKi4S7W8V+O9sqMKBZRqQ1zXbQj6Um95AgDql1VkYxcPkjglkxp5rszrzn
AISapDPnBQTW3zgx1CfjA60hcn17KIQppQJASw+SQiKlHFCXBp4a4HsTmngyVPNM
/62BAt04YiCaTAFlEPLSq2jOlc0JnXoKaDj/e+/NbL1co0T1kTGg6uJBabCVtksB
etcxtW7PiZGn/iRv1bJFz/UEkY9LJXqe0d/VzRdgdjwsBD76R8yWU9PEUS2BTV+s
E29DX1vzpwlUcKqaEHuznVfehDe3GN5yeWFUl+a00ibOLulxWHRzKVNK65QuPZR9
gPFj3DwocYt3N5/x63bMRsV7/n3mZopgEbo76uqM+OnNI3D9WOz8ItCW3pmlX+Sv
6ycxNumktO4qvsmqRUWrPQ/lNnwtWC/5Zjfmg46KtUu4NX8/3RYlQtuE8XFicQE+
REU9/CQEJ0cwKQFMT9Ss0w1Ax9FEFa8AGWz/vdIDMAbR9olPMs4Gz5g07eSanG4e
ng1LP6oJ0Vm+uokRRYKvgu/i0GOc150gfjB3R85Hs6wULlioC/B14B67gm+J30s2
tgBCoDCMxowGNHgV4eHxsSo21L+doE4cD2KkTKg3VqXYikbkV46wqrJSuAbnbdP4
krhleT0HQwyq6HHA72bQdYT2rgrYJn3AYZKG7z4ml7CahlZjjzmdSddI/QfuV3N+
FJOvflUzJAaWz9NRMVx7CvUZ/TM89+E7JBNoxBk5wvH46I82lby9hWTQ2fQCA7pq
iyh7Ptm7YnQxQ5MAGrXhW0//hkm4kOlpM4sREsPyjCIt3DeYyb8q8TxRzxMTv+pZ
VEP/JtiK1vvz+uEzaPnvzH8ev53dZl+YmsYj87qZ0apWW69bIIhVGEcZkbeP10o7
XVphY95/C++qxgJIZsI1QFZwLghYD6LRUeSgtjO8UbORNKxaCn14zjowQYCw4wgO
ULoVsRpwwaYpQ84j8HshMHEzObKktmJEVH+bBvwXlBkC0xFY3yTGjHsMypKoR6mF
28dgJKhQ+Z5j9wZdPSf7nnfAB6JvrdlyF/2VNoogYKV1ctZUpB8CiPdiK6oX0Hxy
0kUCBiHZST8HI3tOI/LPZcgQa9rjFJh2YCBES8RysTRxIOVOIRmBeArpg/a+TF28
WQ3JlEBOaOKMAVfaQFqXdypxiTdp+XYc1xVRq+SRCQ7HNQJVu0iz1wfZGa7GkpOB
5RcQrY53F33K9MLJweQpcArSbe0OrfbK+mAyJ3Ifp5jaR3BHKEvItjCoqXQ8NoGi
R8VeMF6NKN2zN+zGR/Ug452BmAvRsta6rAB8C88/AklaqlN+Vfxc2SE+O2+gt6Rz
UvLY7adFkKrD/yqs3q5FA6KOS0ZlT/OWEE85AKUdTPCj3Qc4WrJpF7E/IEpO7Kpk
9dhpKIxpFFOUiil1aeAqiVjZaSU6oZpbuqCja+/Ya/9mb5wfl4cs43ecBK8wKgXw
v6Y6w61PcCLBQ8tYyPRTSNvJUW9YsUDVP4QF4l1UjzNFOTuNfRu55kcfAJfnJPXl
GTIipPOxGYKrZC/UedelZtBefsGX42Z3vmDMPqHJpKvR3JnCzYwHDP43tuJtQ6Qj
IJFe778oFlhlZmJ+Vrx19oVUe6Hu1OxJ4897VhwpCJeIX5JZQHN05wpnL4x1Q2eJ
Xa2XyFdEV4GKz9UJ5Ozgiu+n+VfDswiDMgIe7moF8DPm3z0YnIhP36g+1W9Nrstw
xBGhcHhru0eNaFxYcSYmyipdjtRN0+f3Q46a25ry3mbzRto5M1qiD7E0p7Isj8NE
9F3Gs872IWiEHRccK2T9L8+8var/c9SipHkgy1C4cRAhYE3Hl0spREdYfuDhJekK
jtJl3hDTJ45kDV2z64PXOx7LrCJ+CoYuXJEtsN04yoa6Bv3fu8CLKDAYt+x9VMed
zt9Cqu8Ypj74bU1sYJ6jr4XlGiinuNjtA5UzqozNIoNQKy2JV/hN0uj7PvmL5O9b
qBHHu1fHc+X+aefHCL7KMfDEIaNfGINZdXLqdIDyJ1yzCtpbRVvWA9zs0q1qxIkc
yCADo1I+HKa82pKbfBCRuhyfqew8ZDj7JzTC/vKU+ZEbZO+6IXzOFR0YjdKPDdgi
RVr2fPaqa8KIm3L46aDkZCKd2iKJqlOZh3xER/24pA5D7Spfs2VMjAR/u51VvuY/
JkFYvqfB+7TQiJkbV7t5PUGyMZwyj8Vvpt0WLIP5PtZbLNWbEvt0JmWe1gLfeOiy
LNZ/vnWOEmPT7J5mNoNoQMFWC2LIhU32EfPbso7V1Q4H1uKwR/LAyRXaREtIGXcE
Hi+C79zvy4mnV07Z+wQssw/2stuwMpq9c6FslO4GLzmCVRE98n409pmlSFWkHzVs
MICRuuWLDNqtjvx98LzooS0pZjYjXF7qXoyZboGItcdjgydB6wYdbHzQckCVcsAP
sW0OL0IkNIHhejQtQCpBWuFOLy4dRfC9l1/1C2s5wHK9fcMwUcUoI4L6uKABIBbM
hjVzyhaaN+ElqwMo8UFp6h2R02nQHFIwS6OVIHeE0DJ0DzUMhgjJPKXPzRYM9oj2
70I+uhDr/O85mCgjKFLPwVRPfpo+w6NfGzvZbpGEhZVZwMAvVTGohKxzQMriTz/X
B4yW3auLQniKeDvcHaaoDtQcZjAx0U0mm3uwTAp92Tnn4NnEMJwQ+dVTCuNEAErB
qgSLBVIYGLro/sJpFebfW5FnB3Wt2Nlkrdq5ciHjWSB76A/mWZN56F7nmd+cy3ZF
XOU2yGg9v8hjM1+hsIIwrgpBUKxMxti1pKb/DJV/xuxSsqF8xF4vAznGlAvNW6iT
7QX/0yJpbvTAoKvTzb83nmSwm3VFJJwxL0wBF1vVYPF2MZuVJ5r8xHb69jV+BHsg
8l+PIMhia2MTizYMUsvRYNSgCLgLZHOyn7IndkO4mSrL/1aLOWe3RfLlhiIG0t/d
7md0VN1GXgIWnp21RKpHxDbUyn6Y/P30z42Ca7rUA5Cn69mTOnuccTzJYnswrMgN
XnLJZHFGH5F6S/nz3Z4EPOO2ODCiGKwvDrDS+qcjP1/c4gdTO9hr0YrOALM6HkPd
luiqfTDwYZGKU+jlqNvYD/5pQIN0Ga64IDZWAYA0qVp+9Af1ieyXwkHK+e4m7MZv
7Van9h6X9znGHStRHg583lkuZwRwg3ok5z3xdt+W0ovR/uvLn3D67ZBPzEBeQat6
kbyKgrDY83GrUTE41PHYGjAMbaL7iwu8IGt8d1Hgx25JP2GL0Jp55RD5f/lSRY42
Eh0WzgFvnYbyISFizxsODFWnuRXgUhb+GyARw3RjSXE+cSLvJ9kzVNYp4irGZieA
7LLfH4ICY13QcchPAHoaVr+w+K6/jcf1ueskJE1URLTkRtpt4AdWLVoSTmZbMMfm
ADwOQEBl4h7Pax2aU7bUVsIf2dvlgnNC/mB/eTDp1IXOzWTToPGrzllglIm/kpMq
6U6idJmrVS8va/o1qu8rjJICmCgRTAhSAv2ehGzzMi+5XDqGRUDLQVlBAPF6IFxZ
ymAPxarewXfpI3oY92EdNLyGth4+VxUVRMzA/63SP1IxVKci6+yizNlOb5AYJort
mztv8Y3gboMPalCcgoz4NCGIWNWgOCdS0Cg9Mn0aQSCc6KExAzwhB2Y36TwjszFb
AhzXN1l5zJ0JC5dlNfOU6/Z9Kyybi+QJrbNi6mHx9Ln/5x6QtHTM2iwWvWZO15yL
Nn8I4z9edWsBdEXQm4uv+Bt6Geai68ymDylCgr8VPxZu/qai6I+Cyi6H//14oPwO
bcRUUAx/hvbWtG6ehWEm8Mgs6699M/g65nJBNvDxN5Io7IzxJJrP7vLb9hL/6tOz
amkqn3gzVynlfswg79XlcdPckRygY7LXb+WjTi6IWwNzIxPm8H5fwYvinTlsBM/g
Nb4tvirQ2SrQ61SICDmjILn7sxEAefaDcI537YTDmOJoznZSSXG6bWiiRggXJlL+
VV8N+UlpxtVa5Y9HKQAC+tDdUC7SgirmTRg8uWmA5yr1pfGpBJURKlRV4acp7IBc
aBbuKuW7l5YAZs4MzbybY/U2h8oslsyjNA73r7fC4e9iFDwYgLhzy12iQbaMVNeK
kZHyMNDFu94Zq1zisMtbdehrncmamTmJiIhgeCc0wEwlY7DjOhxNs0iksHkJVojO
gV3BHOAs/Q4uwnk3+mGKUPDpMsKWeGYPQIgk4SJ6D1iTgUegxeH4PHWVgt9SMKua
cOl9HOGdLlXINjmD/nNIogEm02L+SKcmmGJtgwP8GEtg/kGOfdU8DggCHNFUXcQ/
8t3dos2yWltznHFvw+YUrfmqlyuDXjowzO9rmhrY+jMoeyLpnThEcKcdfVJlQKJC
z32rdMJ7kYVvKuO6dk/O6kY+F41Q5mqaBTqmfV0VzOG0A4FMdvfDO7EzP2Ea4+9D
/9/b/lYEQQxeYPjrv61d8VJKvzW8bNYlyQ3SM7UQT1QFEhIf40gwwnaWoxUwI/M/
iiz0dGwBt8X0ADzhj6bNLKtGSrpc2keMnbnFk2SI+9oqK3LEbHGKEuErSPE9vu1i
zFjVuoENoq9klkkb89RmKOLxjF2rnodgmeT3yjqGaWtgsZibsVCe2zQJpQmkwnPs
R3xTKzIe0f1hS/RkyH9ULCBYkBQiiz08VL/KWIstV7TXYzO99dzD/xE8I23fK6YT
jn0Zj4CouO+66P2OBQjqaqWfKQW/WjipEqBQq3RxrQnxY+xifRJFS0YeNg964poY
MAhxX3G1CizvUuu/DVo0KrKjkE/6iunEQ7Ko8pVR1lhAgD5nzt20i0waWjI1ddj1
j2dd3vqxgVN/nu6Q+/NKBTqy5MtGuOIbkE/oCWppi0r5Ooe1DUON5wtLcmefmVsZ
O9DE4AMUeZYv1CAyjS6zcOZnZ1sgJllNhrTe5PUyx8fHDh3Q3y/erV4GBGpHl4Nz
qd+HcDAh2xFUeVJFtWG874DNcB3EGxDfyEbl7mfe6FeHi1vNZAsBMuyBHbiC7dkY
waczS3jmJMsaW8TcSFH9QR2DPTB9UxrUIDduu7CvAuR2XfWHZbFCjQj9ZXgL8oyJ
PzqzoFeY1f5lBwmZ8UoOLS/WRhi3hceLyUMVsWsoR7ClTdahrPHYsusm3dJsrBRR
+8S6BbPBsLcGo4pOZmsmiHqMGAoMJdUi+Xc/SnlpBN/sgiix7lVQ0g4rhlvOqxoA
kwYooDxlCtV21TpyT7Diox7XBz+Z4inWytEanBrfuaQ2nVperM4A9QudtUg2r/9/
S2/7EpaDPWc2xahTdl/DX46d5/7Y5SdsAkYdFA5Yw8yM2YD/y1GT0sQZ1Kt5SzOa
01gR/6Uo/dttG3pl8OiQynpHR5XFlv+oKZNFWZxBMf7A/xpyLtpB7Nn4veSHaZXH
dNGwVAVTEBxAFbb1j+NTj79NV5TAhH+rPmx/TnqQxj4//vXS6iQ0V85ZIGKTd8Ox
J1a+GAzDti4ka3i6xIhs2fvrjulP3vitQb3DX1230USAW6eWmx10Z9VVd9E6EN9Y
wDSKoYezNFWyLPbKn+9awBaRR8Y8QtrD3M8hTqK9GYe2n/MmggAxBgx/vwGHxGoz
b4HCE2HbQOCq3Tv06jHC8y1YAhJEuN5Q3d9Gb67VyeiFa/dxRabZ8DUKwnZ5stNz
jV8M1ypOf7XdFxYY+3ei8rBnynlz4TAK6p0fHypD8mgvGVHCOkdAu2AiKtpnI1Mp
t4ag2shJXKVxr517uE2cXvADyyybs5mUUauMJmoRDaDWsnpXN8C3axokadro+czW
XcH9lv1IEU0ecZqChtJYGCQV9gc7NoYFFsy4t9zCDh42E8lvv/Yv0JFgqlogowFg
OGqdhCMAE3eGDP7+VOq3QCF1TdrtY/HN9+tb6GBEG9aEIpzTzdovTKgSwEancVkq
6PjUA+83dpCxuPZseU2xwKqGe0nhAeP8TRp4kk8ESLkpXBuSoZRXh9mVGZdr8Iq9
0nk2BW+sUTpS7HYR8AhnVekJNkTjowDQQzpBzaTwY4UOoT2aHI8R51JU97jEfEDi
TW22Wdojov+nf00lQLH4ew0QJkskpqLOeU7+krZcyyKx9oeV99nAZS5lMDkp3XAV
iQFdSD0kUUjFZDjFFiH/+MYYaZmBzPemHaLJfEidwgHyx0asmhO/eSzAzHqXdKdT
ZA2/3EIWY6FaRGag/R06djx+pHH7Rd9+OeixpzqoNlmgyCxin6ZBtLXVguLdHuWk
PrPFEFw+hbVS1v3gIwdX9+6t244muh6MuEbHeHeFu77JSgfigfe2bz5abPa7yw6c
C2FAqc6VWd+UmJj6layCAfh19+CjSVT1E9Wu9cbNbKeA4TJLWtfEyWNOa0/sMIRf
sgPBr9s1H5Oz0pypBzZ5xsV3ZsuZoJDA40XOgKV+0JnlZwF4a7deUxMH35OaBFFa
qMFS4Z4G8wod7Zoa9zd5UFJVs7gy9amjf4zSYLurTK67/Pw7fgyUw052l3vgUn6O
5P1VzDzjz4uzVFkcUX+2oubAgOggKgkJpC9m3RHmme5YVWQ89dPkpjXrU4FhuF/t
vZnAeJRHf4w+F44J++XAiTm5XckkPaVFKApj432qsTxsUf8tbfyhqe3d2W2S+dbg
aDvUy05aoJJ/Lw91jSas+tmRB2qZBX9sZGkvqvtMzVNznNYH+eZQhvVmxeiQz4YJ
dGFNwKZNBRsYskx3iy5ZjJdG4Iis5BvBlWhqak0uyZkRlxlpT086z4rzmTrV74cJ
JSEkdMZT1GNVfacBrk1+jEj39OZN8ZjPpJCJllVw354GpR1XvfzyK7CIn7+SKgEX
q0EK87Hx4J3mmlZJtDQj6XJfzvi7WuoRWYHTSHrDetjXQOCkhOFfTg/V1s8r7sHt
fuJSsXez2e1QZnpuiBlO7HvPO2fNlYhutZGOqPvUC4Vvsx6XL6h+W9KLF669wHOp
dCa2jmVSHwPJqZ2qfU/uG85gXqJphDl5WW17obX7vpnt3UCN7YXr6NV0fq75Hz8d
ZkyUU67tv0mkwKa9LyGvS+MS8Tq6uuJLTWTJEmGMRqbFnISIPO/0JF48DKjizXzA
WGvGkt5TrlCuYkonespIFNh32+onpbi8tMsph+/cc7XigLwV6UHLpYY5ylmUixoE
h/RH8oiRbGUw9BGwah3Xw2ewx5kwht/Iz4WFasH7J0HWLj++rkPFu8iX1m5ntHY+
yOEfvX688Db9rU6ThUhVafW7gIpWZq1v+ESg2M7z4oj3ZjsLV11OO+hyewZDEtnQ
MpeByN8TYHHRgTm1QMlSn+AugxbutyGwKB2NShot+A0mpceR9gXCga9+PcQX5eNS
wuY7a12KK88DwzlLdoq4QIgUybdcX6EL+7CGW1JEckm279qYO63mK9dhsSWCndYK
nB601KDJOHIfG/ixluwCImZ52g9L5nm71uZDi9Tx6gYjORt3uGMSsj9ym7fX7lza
pL/ncf/lOwxG7KiVs3W1zknhYdsxnSHQcLhce336yp9NQUJ8xZmio2aDZch3F5/p
MFE2HWvjHd3JGHs2nPkDPG691oaRh/GKrd7mGhlM2Tq0BNODxSnpUYsMjSvNk3Tr
DO0tFULsAjreD9a8+KPB3tmzS5AGGAgbwahXhWBZbtUA1Dq27fEgbRdAywMRBaVt
ogzifgoIrzr+9kBQDq9pGe8mmIUSvHk4U9NRSnCmN8MnD2KD3IvOwV4o7ykEb3kU
hY4SG9OmBsAt+BYan9JhP+0WvAHaJdeDHQGTb7v/vS+i7fRAhzZ7u3AvROfx9Ugl
no4YWhfNSSgscO80HtWyP9CCieFH2iC3fd5g7rgxTrB4gwEcV5BcGveF4dIVeEVQ
/rOlst2Ovgx4EvLSndxSEbY0CEnvVYU5ouc+h7Z2jTjgoyJiA3jnXObp8IDn1I6O
6Pax039RbHJmS28jVtENZqXQvRz+TCW3ESXHG0HI6jOZyPhRtRZGsXtAAfECdo73
UCJjyFQo6jLXcR1XBTw+HKU5JnYUgV7QdpNP6KP4gB13l0pHxBiUzkmMab3WoD5P
n9ZpaIfpMofuyA7b1ibIZWI5v/CnqxNQqOsoOXq5lG72ExdEA+4B10aHjSseeL1F
xth0qY3GDF0Z/0mxMw+ojz2Z6bgYX++p7SYd7asijwBO57QhRbdHgPdr4diJQkrM
4caotkEa2r+wvM2D7WynAFySQ+jAO0EnG8XLNFTOz08j5JIgQjo8YZbqKAxsqdGs
zYmsDjMnnSLTRYweygzOWTt1NqH8ZHTpyWQc89HqfFUMp7OSfoy0BAd1499IzaLD
vuu0DGEpCYICMLmZolWmEU2nZZITnUr59/aX0l1X8yUvPuQRSnZk12v/H0aGJEYt
VSEOcVPzHHc3y9HZbcbZMGYzZ4QT9Wltqfq2YUsnHrBKZaNRJDjrNtXXFX+SqARD
f+LTqytdjSGWC+xUoEXT2/7kDNXu/xg6Lp8wErH1vjnEdisSHEbs8c2YsREba/NU
8rhIeAalK2ynPzyhf1JdeoDXbhBJyUyfS0UM3qOSd/SJwUOcNE0trEEfQXfiTdOz
YRrOCZdva1jZO5V2xTvesqkPkFuGxqYIi9y0rEEqT4i+mcdQ/gvHxTT06ubu1VCo
ILyYWAkCFkuNdPatOZvfe6nQHkAOUQypW1cejHJ+QnNAQg4OnAN8CsiPsFjM0y12
ggBrVYFFLNNaK6zuZGmAWZ7t47A1UQ+LQE8VAP42qXVXqfxIXkHfQmsA03wzNuso
fU7tuW5lqvnwgofiGhYARVZ6QFzSRh80j1nLce5f6PwQiqK9QpZWKEfb1BuQNMv7
BVGKcp4arGEhkMlRAGYiWoYTdOnZH2EWB4icZuB6Oh8YLcc0UxOt370w84/QZnR/
FkqmejS6MNkkrRg2RFaV30g5+TGZhZwZJNeyCEo+oj8AW09cJQ2KNnPHFGDY5EV5
pmht267RTEZbBpRS7To4vrD97dBX+PbZa/g3325KAVEPJej3fOMjNr57bk49U2UD
a+l0yWO6n9V6rl4D4ZWf3iIWxCnrsafcx0JDrrjpo4bg/S1WXgnm/npQRINB0MJN
MbQbVNTgpQsq+E2q3b5biGzn8v/Bl1lyDJuUdMaynYFQDWRwA8SAIj9jJ5uMx7fs
IjL1PBozW0ncqCNZCiapsA0zmCG5c9wRTQa8Cz9sIeBVYWuUADd93eIlqQBowQKg
2WfONs5XAA9qj/pNJh9I40bkYgTB1fbdiqc6ZisVeJsClH1ELBRPfQVJBwOrBFOC
jhpNBXcrqmi4ajwnM02vRjWkVVIwvZLsh9UC2WXsyMaJQBNvTkerpz5XHB5nCieT
CKvPFBoh6vOsNMlIA0xKyXNcdkOCOpFVpFMU0i+MaghhS8oCtlzRrYPETURxdeHs
+foQxaIpGQoDMnslGHqSwo/1E2NJ2Y70+RA0ZqFtA9KFAV9xXO8e93QvP4Z/rW67
oe9JATFToUe/vvP6GlTJvko/ny6xdry0pLCgJEP8BavnKSXeE1ZwQ70NauRC+/28
unZBDdAyqsriVnUy5jYTQDa8W/nYuj2AV6o9e0+LTI041hKVOfQVGngsTr79RgZJ
sl+/5kGIooQM75J+DrXNXaLU3BaOasXhc8WBIYAA4GhI0j+w2roTIzLJ/UYHQBOh
MGSRMt4tE/ehpOudSeYfchcAwZvdMeJWcAIuVJO4ycB2lX8hDT9gB+7ElXfMX7/G
KjtqcyvDgHMQLtAH8j5I3hjiSb9ivnARDEPTesJOC02sTrjmbi0D7ArTSikqlfAZ
CNp2Swa74x0gg2DBF0iN0U2YN427PCPiawPaKOZLVb2G04i8PULXIP66esD76Biu
8HjtVZah1cbxW2Ebh4uGlHzc3qpMEUCBXh5JDHs/iAK3bfVpxQU6yP2ZEAHtlNoL
xNg/reLbXiGQSFqqjuoQCOQxoyb1IrW5oX1ie7ZSKdJl930bkm8U0JjVOWF5QL1W
l0jUzwaJLjWBjQVr4x3+G+PMN9d5WkgZV06siwmBNh94huNqvqgQcDCxt4GNTQoP
6p3KQPAA44cvb3opJItLGQeYywYlfDisu011u8XOt8LLMsWVADqbTpYoepDysZRg
q5oAPRYLdVCApCM2Zyai0iDcnYuS2kxg1FiEL4o9ujvK6lyuzNRSZKzViPqz6kFf
8WBJivdHsue9reJ+yLXB5x5pMSAShg8bHOB1lbcGdi+qn1ZUKtSv2kFAGb0Zvwhz
iMsZDNFSRgXsbDhHMCc4QLhZFJXNo1MO2NYtepXwqgSSxbXKu+hhAAqvnPVYknU8
H6Se4bDKN0IAd+6TYvISC8HPAqVa5HkCGizGNhNaF7kU4mSw9DvLlC2xATv263Sb
8AiDSk4MgLQQgcjWqtojW11VFZHJrYymX3Li30mfqUsZDMUIFjka7GZnD4OFibOL
haDwo43QLdMUjvh1mlCTWrjP2Vr4fHljD8+BLKsHsQSPlZ1soO0lNR/9lY+DH6Bh
zhjK6ComOd767oyk33RiXVTwTVme/TIiqOrWAYmYrB6+82Q7mfsYTzwPMWoP/zkq
HUpz0/GHTiKqmAktLDiC4/VBbmV0lxWes+9WdaEYghfv4oqOfsZnDVCbJAc9z4mW
Mb+uodPB5OiUjAfVt5bp2Il3KwHYNB3Vp9F5ZD28VPljgOrqMbidlWqANuVOgZvT
kBBWcD9zb9mqNbbPvN/97js+BK2SpymOISyGapTT8M6HueNXcz4xOtIdFAX8kZsZ
DR4VvDo+b7O0ltHSWbcYjbiZO80KxddUYoXDb5fKAxY3wKRsZ7lko+p1LWJrZA9p
KVB54Dp9ri+KUk7FSeHAM8N18Sqw/ZAsPxufxiA4PQWkqcH5BROKCEYR/DBQC3CU
87WmfT4A/27Pomtc+pekoHb0bF6WxrYoR48M+kQsAxzMov2jIs8pEZFukPl51Nb6
ydsWmOD0m0Aplr/VBSrAAPMo4hOg/JQTo/4YF7HSPuYDZ0X71tVSElSU1E76JA61
As9AXdzfdvaHyKNmWcW+fMveH7yGQ/SkwhyqrIWCQfvMVSVPi0rvpFkI/QiHS2Ne
Aigv/vGblT7j0Suy0KyhpHknrIy6eyd2rmIskrAjfWf3wbzJgC8iZZ6o+4IUU7pT
47N6ybOzgYGmgoiWKIx3fL0br4RxaNhGNJ5Ut3s0/RTaZkRwwRMdBtwT2hSQJ/lX
VqNtN6ky9K6gBCiEQADVacQ1yDS5HCKwVRiAAfEEtN97e5tB0QKd8nwlqR+OlqJ4
SQVnkG3ZThdkWNdnxFyhErx7QFC8CwAjV1v0D7HnQT3gwl6NeqZxt5m6psdLu4Jx
zVTBGEeoaEb9kbm2BjhIUShi3jdUcFekjJH44a57aeAOE4waBsEzkaLwk1f/BP12
sIRHM7DUty7/xfkBq40j1UMwJCXZyRHEUrblc2P65mraugJDOmgzQCdcaVq67g3A
1SlR5EGoRYYvhSMthb5aGBLcf3ItMkvJK6qrrRWdao7bD7r8A0mTi7PbaVAZq23t
yhSpQnOJrH4J7FnucGXrV1azSIZj8fE1lSxWw13M3zgkG0WRKgoD1WT+6s4Z/K0C
GuDSXU4aeu6U6P8UyhbttfQGsFbFTv3/zUIa1OL62Dc3myJP02FvR4B6cLZzvIbi
6tDr0Z2pvMkDFyxaWJ6eC/6OPUFL2BJtaqasF5+30NCoGtWsgL+EnwJOzEJGb2NH
sHhAkPZserKJE1XxRFp8jBOBi1v1BgT4HcIfxXUYr46v1Wj3CZwRQe0wOU9U3GmW
+peAMy6/Wh/eFFVUbXTef+azYif/42xV4ejUeTWGDCdMXPhURwcsXuL9yna7aoRp
d32/w3jkw35bpN0ILXDr9YFoKp3IfeoIpOH+31/FeVlUCgMFw1voKPtRbbQLc1cp
MPwa57CZ74YNXOS8Isg3biDdLSGyXHOw+rVDOOZ2niOUC+75eEW3hSGo5kjcK4w2
SUElk63EqUPOsb4l5QrNXroQxWpfAjaaUH32xo7A3wZ2091qFBkkTOOtYj5BukfY
rc4Y9iukws9a3yFuaSeer4+ln+p0GkYJdxCitLQcAfZE8h7uNr63+woTeIIvz9gZ
nwOkBYT4Z2ahsWwAvCl9i6O8Udnqhwb6iqGxv7su7mGiBUxr/RvQ08+nkJzsS39f
nIAjPr+75jeKsoyy5/z4P5ZpEeFWMrtfs9L0Z8Dnv5ZYjV8jdwl78xcdV2fYQc/V
svLdCnOKPIiGn0O5/m74luHGW1dzFIHNDwG3BHEYpoYmB8OAc0cNM9OUXh9k8taj
3Da/FwX2mpP1xLDOnoWCuWEfG9TbmW3dV9NJkmyQOIxp9Hz25D8FmR/W2nGGh7Sz
k7lzUmoq/Tkfk/1k6y9gXku3sA1+xQZ0T7mPa1q5NBm6HmVa5y1V5BP9/5yHL28n
jDDK8nXf7vFxPcXnjS/oUDelRl8kVTEq1yCuv2V/Jn5aX8FG9eP/5WL8bmtQI2sp
i/5tjy3A9d3MSfmj6B18gv2NHfpNf0tH7U/N+aiNLyJ2aoX2pluewcz0kCIs9qMH
I9DW0CX/atIFGQ5SLCxfvsqQV1uRDj6nW3ByxP0qdnwhv5uukABQ+iHsxOViW0Dr
Fz749dRhfrp6fhd2/r6hZvs5J/HORAdxQRRUECE5Loza0S+VzXyKfKlPG7S961xP
MjSthzRDupEVcjHpjL4VeyMFs911T6GEAUPnL81Uf44wh8/qKnhhKn94+aSVsZri
Vcsg9NdNoUbzb0liMclZ9P+qIw+ZMTLEWXqJyxOSZjHeZujb0Zsd9U+LI2k40px2
rBsG0eX7xQew5+cruVAe2RtmA0PaV7URdR6iVRFfxRuV9f87Ska6gNBzwKcTjEz+
4fpBJXOAGn2mxPTu0o1NnRi/nZWaTpu9osTHMhuIP91RWJeA4L3EQYgXVi+2b8eb
f9QWLS+6U86Rq1r4wf7Hvo5a6y9uG03+KcckKF3WiARBaUeNx5+9ZV59J3snqOjz
xhCVDoQPhSX6HX1KKScU47xC8MOB+UTnw7mlQ6kMzDFVwSDo8z4mVLlGF8PkAf3t
AiH39K8idQtFtj8WonGVxNyNqmZaxpTQXO3akThckP5ZWB+y49aYBtf6mBVahKEw
UGgiAwWgdps15zJBePux/JyYcDeJDL5K4naa1UNAkhno+YeKOxKzI7EMrhWqmXYU
oOCzNp5PVnm7N7ajD3gJFmuCRxe0IeB5TZMLlYyDzmBwsFp/FUFe55lu3CwN12Pf
4MtzFo0z0ltDKknY708HWwi8r2vPbeCnEemmNZVjlj8EkWUDB6Slj2NG7d1aYeXn
60MarXU+gagbSGSmioF4MXq4MCSkQ1foDqESLqCVEQfNyScTPp1vw6AqA/r4I5cH
TrPh0io6gMMw/iPErhrL0qnR2QBw3Uis23AbQHuE+xnhF9kzn5tt5cuvqmTIjl16
GWWpQedVu9s9ZpD840PQLIwkRYpRksUaHaWVHqf/Y8wnm4eMDmXkRwNHb69j+Tn4
JGmI8+zq3X496ws0AHALnM7lGVgsJX5X0wEoKNtbir+U2ebRtzKoDF+5FRmsblK+
A3CSWwYB9edxvhoGig4EKiLoBMCp8N2u4a5/kaviDBPaNGair0qj+s6kiXnR4p5m
sd/VMKnhEd/nv1EdsOUwneQfZI01Ea3BLZ3fyemotJAHQLcSRrwnNZ3YyrygyDa9
it/Evpil7NHA4YAHCcIlMUoXFk58bLO/PBCUeIEm3bWn+5f0XUxcCQANcyW47LO0
b9Cnfxd7toqmYG8YrWD9UxGtLDIhtwT5WaNaWMgLgOC9nt6GkxwsZrMrxiTlFZHR
krbFVbOECxx0FzXbcMcq583adBrqQVvFjfzC0m8iYRLrPW0ivB97x049VfRKOHU6
5JDYyH6KaZbu9tUxYgrCg/P9NUp8ba34R3NFytcmnde2tpSPdOO6BDlrisLIKR0w
HymISzS0xg/O195SnRMVZthLM2wJjqVqRsrfBq5dxEuu6LaQT6WIOyD9ElzFofEh
rdLFsaKJsocp9Is1avaKQzYpHzTM7DSZETkqh/kbJcRUQiM1lsWUa6vgb2C4elzx
yvbWeEo4MXDiRticRDyXn+BwQ6QOWH2KKELII/S4u18G/osVvIrqsmMiFdetm+Z+
n23jHj9u0vJtfXOobvl8VTiZsMXOJkyYue7+4hgkqF/C7+kLBeFtoM7EviRqFsch
RDvqmwyKpv3aEwtYsV/zS39rPjwm+6vzY4PNP7iGqs6TYLg1YY+OS3vrofRzaec7
jQrFf7/Fo5dyjEgqghr1cnG9W40J7f0klhEYmlafzOEgILW3Zk4lpr++DQ5ISyp+
GXr3Phj7ffa3ri0oGi0xjZinPS9S3JX16EM5hBdTO0wOssIgrETlDBgzQvV+yOMX
npcTfnxas7fiumaZFGqUObWB7rXtQ/fS7FGKRTBATu/kYqamC92BW0O9J/iM4Df0
zSNWkZ4cn+RnbAokwSc/zmgUj2XpUVhHYk/8f2SdZb03nHon2wFMlHMN68LiQb9G
tp180U4uyQlpMlE/IuKKepWjsHFNKNnVy2QYa8m/4NZ4aF3IWpxly9k1LcxXo2Rq
u5xxs84CxItoch5MNqnPBz3aeUvlmFOm4J9OKeCAbV4eIX4LuHoIqDDSa9fr7njk
prfq+t9ZEdPHDaLK8akVAu+/eJ6Wjmrnj0SeRzw73/BeHZnZLbmtJhyXw2L0Mrlz
SMm48x62ZYQ2dMfNF0Dcd82zuX82B+nFIzfKfn7iGk5mEOupHzUVcZN3bJMXCCE/
6GtPk6asZAdF5LiGUiI4g6IgX4dqKbUZ/5BiC4/Lv+le0MFGZFzQPxJmXzLCHsEe
P4IUqMAz2zLEC6l1nyhmnv6azmI0xy0qZnHbAsI2nTnE2WP586I3+L2+uoeX8+Km
GEuUeyzesJamS46T/ngKmQ7x+gy0TQWkvxn9/n+2H2wmZ+b1T7kyLEKxUCzBP/UA
knD5NT/NgYmzQmMCzxNdg3Ym2FkKphbKaCJmcJVOY0OUWA9E9/APP0BYMruHwuhW
H98GVd44RJ7K8oliqI9lO4en7WkltBfvdH6/JxofZoqn/uyUf0LLeBNBmq0HHwsL
RaH6tNCyqPdbOV0Gd38EkeIADjyE7ckmydJCvpCNoUXOr8WrNaP4vcLqUe9g3LFR
Vy1FL7D5/re5+rJN65TbKWcPg78DrzVxMActrbhD7Ya8wJgDenkzoixqAeTwmoFY
BJRmbZ2cAuLGf6Gpe7F7oTa2jwKkq7ph701RPiHNSMP6VW3vQkGOPsNdYXSCxMEz
TqtOYL/HmA0p8TV3XKUI+EmTOR8XH+5w3bg/OSl0sacor8k24ZNUjvegaFVNtRBI
Q/cqidx020NcSDP4bui8w3q0F3TCxRK1nUevNGKPXmUtM5igtFKl7z3HYBQRjlFf
FNm5gOjOnRJ/PT9mQhwrbQya37kWC0IffvwJunFeY9GcwAo5uOFscbaCfPr+ElHj
DMJB5YIuZ4bE2+uW4pXpYgdt8DRnz6DHCriYFOqtNjTMi9LxXg5R52Wfd85DxHfH
7mQEqEP131/pOnzGUCdC2YJYfwnOLAK6CO5jWXjJWBr/iQUPTOpI/TQvzL+XNXfw
YBEDKd/lqI9/CAJuUOB1ALEhrq2fAQ3gxaCl/9rwsI1WzcbSYGMv+TGdRBxQvj//
BZwuQ+X5hkejHfn6dY/2xWlk2DIpSRAopIz+ENz5guxoC1g+A5VC7ksoS+7nwS8j
C98UY9Uy1TpBL6Nb506bOTs45/KHXDmBws63xQU8/VFyaFNuP9CSqV155SFmeuLy
sf1ivl6K0q1cTeW871aOXUPpFyVWIdgUpvFWFHOzVrIIQJIZVt4+iiYzmzI+utac
S2TC9mIPCASq7NYp7v7RmaZGL8jVUpr6ZsLx/t1ftPKyoc5INeYoDuvFmiYFoTOW
RRdy08gy0WVBLx1AoNQf1Y18sspqy74hqZHKfa1RWoj+Vs6cS+bypmtDmmoSfshz
Rq18GHgb1U7oF8wzRldPuViRZX9fv1XsJjjKDEh3xMkTeZ6jrG0Ap73jL0NUzYK3
uJTEs/XAXv0L0i/uMGd15bokdh+8rH2uQteiKvkSwePBHUG8q880bx+Yo4WoAYQ0
lY7U8xOrjIq4GCEHe6ZByG8tpGK8/Q9Uu2YC23QkZIY8mYh3Oss5bLRaAyEzE0uU
/Q90fspBDebeQUCuyOO+H2zAdzu4ijbWucNAqGiOr6apzNHW3MoCZ1KhEVO40p4T
Aj0bZ2wBPmePKdTKt8gosiwBXxsXiwROQhszFc5vQTWUbrG0/aj/Dv8uPRoJGIkF
71cydvUk/RCI6/VDeQZPR8fuDIfsamX+TEBAIePFu7yDpmjYiQ1DKsZ4gaRaIzi5
xx61FAR+pidFubop2zo0VcQUVMgAa+EQt8PFZdrOI1xnI8WJZL7bm2jAd+QzbtrN
QiWhRjE6fEWALlLZzmpWdb6BLEllglv8/miVveKffXRfm5jkzD/+QWyYX9/mc3Yu
ptiuRB6m0BtHuS8rbHvouYIP0RYpcyDuN4jdT4p/3udZsw/uuKQdSzdIoJ01nQvF
tZSwJ2VBrx/sTAguxWfHqza2QQ2BF+QRmxMWbbb3uGZb+a0/pqdPf+3xHXxg2ylD
0j0YripDnK/dXHdCyglcKOivhrUC7CsP/BUMeLvdNvabtyeRVqlLRckI8dSBK3O4
VhYSI47+s1JmmMVPVk5lTC+H0/00OhszCD2gCc32gA53QK2qy8SX8a+lBPBAcdHA
lTfBQBGvp7aJ18cMg8FeEj/URpbUY45oYD6HUPj0banlyJap+0cGOz1RJZAaQOkR
RgH9TdMDdSail9YYW13cB59hac+j/TIKW7t6hndlko4cihb7ZeqY4FasgChxQM1P
iYmrvHdoUWwZo7R+wwp2qvZvFWZoZgm5kHrmYGqfRQyEX1Fq2trjJK0jSHOW5YRF
isiv2k1+7VFryrCTqSXD3dUWjnXOYfQXnhnvodM31ETyUw4Zy7KOk6Pb+4nX/0/K
EXB8+ewgEwBMgF7jin2y2uyG78A2HOn27FvlCQRH0AkJ1ZeBQnT9t9GKLNfmcCTY
6C5OTNcCvKSl2vcYVB7ViBi1zUZkrpye7CqbPRmz+wAZlNi79Hf3p77Vdc2NUTiU
7+tsnxXIQQEZFHGhPO7D4igeEnZYn0pBx2fwpj7UEjqkrhB15b9S/ccHtmP/meGd
DuYBeIRe8kRZsuDhTDCO+jzkI4e8EeAiVrXwGde9ofAfAi844fmR4FxkhSzxEQpr
dV9VDbPxZHpB9s50PwR3K1EDGdKN0EwZu3Wu7TGhABblABn6YGvLk4tBwSifakl5
v+A+jG9xRpzYAzWJq0qJHkYHzPGrhgMQmuhGsINqKaa0F7SI9S6o5DhJR22AIadE
3GFtFRSOhNL9Cncebh0ZdLCB7l+49LgnAJkJ1eBVPTH7QjBaw3DQj3eoTb0gtCA6
qwLLejY4t4cS+5nGz/RbgOluNCroF4e4OntuYgjIvrEaY5adrcygt0Vg45I2jhLp
MCSlNRo131x+umly/rvxQ7XMQGmz4JR+Ej+5H69ElXHjk8LRwq4XJfNf5b2XEk4/
ldRUUdm2oamgsC+6OcPNnZtwu8oGeBoGNfxCYkz+wFa1EPah/RJFrNI1e1EIfanM
7+AgvaO0sy0beBhT4KfPC0QfpJ8qaNNOYzjyBj9GSLG4K43iivy0twfutd4zuLSB
cQTCTUq2qjAbYP7M5b2AbSSR8vTzPs5CkAD/R8V5dvbJxEl544Y5BmQSdI+6T5YS
oOqO/I/4atsc7Kzq4l3iYea8mTtLfZkBWAl1SQnNxrJLcPzQLWipvY1dglQRPx4p
mE7OuTxzT5IwxKQjsoANi4zNAQ+q+94tv4gGjCFG9yTgEyOunO5EaOV8bmIuPhHj
k0TMm8tVzsiqEZkhAfUpiyCNoNVs7lbHKNZcpOFdVdl/128oFrPZomQDAK7NyoVP
lt0CMkewyvQ+2sA+3KfzMZS/RDxpsA0hH3EYptK3RBDtUTW25Lbd1dw08zv6gWjJ
DzM0s2aZQmXHoxDzwXG+bNOkE6sj9u+3i59i5Tw3wuSJzFzJVa42mJ1iX07/ARni
jQ5nf+U8dg4ABt3C6yNPSBXlEUsWc5ucVVZhv1WqUHPUAstds0XF+SyVSsJA20Q0
CAq3oNGdB/9/MulC3caAvBdb6PcYrDA7byPQSE/U8KyPL+V0jUPeyvm1gL5uUnPL
4ccnDtI1D19vD4fbMvyemTb6BZ0h9qUS4dpI/rTsc39Qgdi+ERLNk8GGQoqyvCkN
Ki3dyqeukqnSI9A3unt17O3DitucF9ht2+DkXSWEXveXSlQ2nBARH140sZbJdygF
qAzYxamH8MShPAbVyWAdpFEMD+xEEN5XQEqyMV6ZCn+cD0wCCwWIPEZitKz9MN6E
zHe6cmAW2PWsxA0rZsFZeabwzNQN88vF8HuJ0/YlpPF6GlFaLA8XsgAWx1MexzTc
WNeoLkLufWmHRLZEudXB/9stS5fvvyxi0vw0nlsz8dx0YkPBlnTvaDXntB9XQSpA
NHqqXpQXQ5QDmKpuC4ZZGej9eAe18c7cE4rsmLoJU0zX9KNueHMzmbrWavga1d8e
9UKvqy7BLXvJw7t1hmg5LRJLd4CyzGF5apOAdPenRo+HL5uG6k+zK0mGIiU4ZeBN
7GMjOX3wSjgNJn3RFvdFrKg618W11mcydn/qycQVxF2eZrYQv7x6uXjyAVHhByx6
oOJmrRdlNJqbNS0RFCrHQuO21OBRZFIr37JJjjGxYzO4eM0vzEFNOOgp2SCSBq+R
27908YIoGZXuquoTDay00MXbxVqrcUKpU6S6tGBd3zchclJVFszxERX+r1JM0MQZ
cxjSbVFLvD16C8IkC2aK6SeFMWgy9ygZxbd3wzif71PINBuJ+KpLlnynK1zxh5ro
MKIW8DuTnkUwqw3YcLugWEZk4rbV8VZmaxXrG9w1PQyblJf3yIYe3icTTWwk778V
Ed1yAUPnuD9VCXJYm80H388S02swriv56jBtzdm/H/XbHWJYQZwzTKqnslnl5/Cl
72lLIdyPpYlJjw8Sjv7IjSq9u2lWh/HuWVP9vWM2VbCsz7o2+IR1y7wfV+cDYiE5
JJOnUTAqU7WdEZWOQ1pBPAf1NHOi6Dx8RvGdJm67RHMo1ljxIiSifoRKH6PLtdPA
p2CD2qlCymsY/z75yuOiYki1TwGGOINyLrxR38qCyI0WG03R9/I/K2QhT28YWg6P
8BHCQYx6mb/D9KxAP9TO4vrZsvV/wtZwQ0G3SEVLIS2DDlry8bodBk+l9CLCFjnA
w9mt0BHfjX2BWoR8kU/uzjKD5x05ZoUNLFgfsV8GN+oRepRqSxUAyImChOglE2nO
pSR5jDAAm2E0iVxQbJu40mcHxSH6S+gAOhrCveOtJggVKsnPVMSWJy1tUX3XoGF6
E7cCDL/kkWF0DVn5Bb3st6jN08y5DgDjIvW46YNgKYBWavaHti8qsO4P5DDwR7E9
nktAWmJ5QZQrFD06rsMg1IFxfhSuo4roB3axeqnZkmjuWqR7avSGS8lw4rLK+0G3
R4UAjsowFyw5FcV0ccz6N+sEYPSnNMedfxuE2G+o7Ya2IZd9Js1O/AT6EjlEDQYj
VYei6+x3Z+dJjTMNK6DZgHSfFMYsODq4ecE78fJOh9ZT3+T9BEXgTSqYaS+0V0FI
7rK22J5RTf+cuKNb1mwPWe1UKaqT+7KSks+AxIf8HyCtz1KdXxu66KyqAnP2XlAi
qAgsa+Ige1lMGOy7CkEwbbUJACXZ/vatb6gzNwLHS2krOlRz1LQHK0bDlrefzu2h
ngJEXI7m/WhXB6lSlWyAjmQODng/aFFXNkZPOnqvygJKg0IGpDG0BibaU0XJcPX9
w5IsXV+aCpbj08VjhBASztIaXsfP3dC8HSD8rEMoJAkvCyquHlpd8dPF9mmwbIbJ
iakIeQb/FDzosm+NiIIjXhE2ob5SvvjQGsTKzggClbMMS12KWtLSR4pI06qAbmU4
nP3LvXqfUoG02up2UDrHh3OuMN4/WH3pmMbXo6MXDnc8UoLXaRrqKMX6gjVXVrey
nBz5mJ9aU/FyRIZyJ5tQebP5AZFLgcETQdHTNI3PWVuxxjE4OWybY7Tu2htQn+so
ABe0i6rOVFS6fRHq0VwNYfblfeYCpOHmnIhMllGq84FyMl4S5QVXYQfhBbldq1NK
nFPAZyRomp5B4ZNh60hyda6WCiDGzZBp3HWAhjFShdovMeE6uUyx5cvfL9Vmwbn0
ogEtWeSQTZa1ikWP46ScG1524zAdwnbxhsBK/8mbrYs8YYTMZ7ptEBnkd0YhvAcl
GUYpRAssSHZT2y/YTapoPjBFvRzsrzp5U0jyAs9YMPcIMtcsPOh2n6rzMQNAtyG1
tgDpFLAvOgamFTO/xZZs+S3B4Tzze0+Oqn9BrOs/5feRowthfhrjd81rer7ry3D7
vcpCrMcHK8mrSgUKymgbWrTAKx76MLGdZVXb7QxuLh01GAI3+zrl2HSbgkB2llsn
IGnK8Tmf0fiCiMkBtX5L/LXTH8h3bQNkq4rBj+IlPve77cgjEGuxPsW3pWszPn0o
FjWFR8D7GDtaynJXq0R2pOVm3SRnNNE3gfQ6aIAXnC3d2lLZ73jEoq3jFY8wiIyW
7K/MBi8LyS9SEi9cLR3BnBm3UafhLlcCHC1BP5ZT7t+HYx0IGLIa7fi7ep2Jmy62
Clr0Xm2lRDKsOA1FFRbr/g/T0x5TJfuTu6JJuW6JWmk8OWT2IHq5tfyfXi8AYa7A
j81QmZ8gHcgGRv4Gu0q9SAlDt9wmTjD/mLml6d197bvhPH7Mavt4p1zsZJyC2uvb
0vlqaAjxO6gSZp2UsjgsUJt+I9KbJGf1h/BFIEHOS4It86HPZPTfDiNTLNyJeoCI
MYEQiqmjEKAHSF8t/Zf8p9JCEt6igxaATDb7kTn98UGDKxr5yeccfR3vlhzSP2Qv
x8zXAXc50bLA4cGL8ECJklYT5GUR3PUYSjbeRkBRyMO/BNfEcJOKjZcV6g50dnQt
BV5Fm+u5FQm61DTz0i9juUBmOkrwR9J9vNyOzoz83hhpxGnmXQ9y7JSppZuKw8jS
IR7YwJZy8x0q6PSX+Yf8alUgDNCiOsUj1B2gLExuLar+vADXghTIGnJMf70vMdrc
xgAfzOqqena8lGaWLn7gzffYpqx9S5rn/LQNt8+6GVwXXCAV35gG/Cuf8UwCDVkT
DmDkUtYiyhTb+fhWQ/sJu5LY6LqQeovs4lmC3gEnG1Un2NamYTdC/IHvxPjZ6BKT
ICoCMfbdt60Y924Hfv/hONxMZqdSm/kVL2alh/JwsyFA9N73b9oQd3SMoalKFqRY
vhanpkYOky2QiJEG8xM5YsborjDrSVmd/e5lHc9kSewSYtpod5+Q1itX/9LiWA6V
qYSAD5BP/bOJiays+Th3iDcY9GF4FSRHgOEj2rzFiqs8fK5+oUMI+eP8iOBcePRN
Ktn1NCt+6ig8F2yKjGVVyhySb5n7m0CcB/Mo1tukYsdsBo+mu7X5QBigM/YPbi2h
U73oiaoA3MGIppvliGZtvTwUuGfnYEy94ltV4yRnQeHu9tFx8/gM7wtvzPXWtQNx
OjCb8mZPMsql/fYHpmjvRJrRhSRazFsUWcn6HnmWg9hf+qyhiXkxxgIlEAfdnF1o
5bSuNbDA9dA1UBo3ViFQJm7E3zdZgoV79b+IZ3DBeTOMhndG2U3a0R9ByPS6KYWX
gKIrSpPmCpx/3+Efu94oiqw9o44vOi7JQhSw4xgS9sAOkU6ZyEVNmup+oJ4eKzYm
M4Kj7E2WIJz0w2XN4X62qDOggDedoTaZDV+IlcQGfq9IrPOmI59hWx+0EYqls77O
62iYqLN0sx00Dvlpg4LggPRfRLCSdubpQcDgCqBc0h1qhMW66c/52S0lSqrxrCno
xPQX4LVbMkkKSeUP+le6JKII/aG/Nn4Mrj7mJFyJkLZePrVWoWGdbuh3Mj3KAfEW
3U5pPHyGHRsc7UyGF33kXAvaa2KAhXyf1wa270sriYtEfW0zA4QFlO0duFS+J6ml
MEdllivR3+aMrQy/JoEV3pJJ0f0qdVK1IlxpP2zBHXjUhMQ7YAwNyxHCu8UHzcXQ
JLeIrxo5NFoSBlmIWnYWb+6Cs+gcxRP2jfYmgoddAfY7ROUzj4uj5kkWc+CtjiAl
bYvB4abZbB3S65OjLRzewv6xSfzA8Ik4fcTbCHdGeEiHEniLg+06x3YCw+rde0fF
RQd3eVnZhVqNWDFwjmmEzVkCKxFISozXdCUKij0Fm2+wE1pFRfnCVjsYKQAFhhim
H/HdMzy1A+1yTf663/5f4Pe1OSJLirs2gJHiGmg99tfR7iDgL563EMLifwtJRQIv
Idy+4FilfFe/aAZph3Np7HVRE7ld+KqXcQb9raQ7YT931Mr8CU7GFnP/qQWgoMzm
NA8r2Jkl+9DG83WjoDLnI5EXAYL5Qep2PwsZ/Cg5mnZ5RideLWKlKR2uYTOdoxc6
gxfXviUCRdjmY4xJLIPZIlTvcUOtsBYKgnG0pFl+gkjJNQN4x9gs7+tKt8zb/ltU
BSeZ21k1SKlOj3LaVtgnK17Nfuyig/Rune5J9iJioiTThsNqw7RyRwjMbxps2kcc
fFmVvpyiSDYxzmKtlxxmoJof0im2qxBrV0y3/fCpuCJbwKVTbOWtWcvVDe1qvknD
0/gcZ5k58h7IPpyvkjhzP6Y96QakspZD1bhVY+eV3/NRZgA89kBR0WgwyNEZC5dq
vHS8Nox70/4mIDzPct6AhnOcraVSlAVC4leescJlPRgxkWphleD2Y9lOuZVG0kF9
HQEMJ0x3VYszQ/zYK9Jh8mgZZMvczmTfclr1yCsDvgqrvQyOfArw+4t0JF1nKJTH
kzbwJUxU0xr/nHfFKCfZ031ecGEFAdQF/kN13VIzMXgeJtH/v2jIXM1hzP3huwkU
fJirPMDqNFZ3W0qddDpZYhChg5V+OhGrcoU2WevhgwKw/sju8HUZkXpTRFoOIFSb
bw1YoiTohHpozGy5jbYOHpFKu1fPVVr4JXkYO4opTFF3xPBdc6drIKYGDHdnARXI
ac5KNVB1xjE7OuMXcrzAEWZm7LETBBOd1yjk9+fqDpo5tlglHuzj7+Rc5bPAsRgP
l+pVGtADBjTVIX6koWqVnupYoGSbHcoVMSVmIsUnluEagvZ0OqEsxgtavF7MVlyZ
vaklnIwUrkWoIfVONU//JLyRQiTLJf99hcy20tEXh/JYj+izAf3g6Byb9xOvJnf5
Pd+2Hie3l98ugxVvX3QYXQJTXpSbOl7zFqpcUmzGDQg5C0eTcqr+5bgenIEXR6XV
zqffepxik56e/mzn1hHPMyd3Gpzmh4wGHWvXSbVdkddkIP3BCy3T2N4dUWF+Bk43
FwNzUsFIn9sg0fkW3+bZiH+AkBxY6S19ljrFrZacax3bAkXrOjq4KDhL/cTgc0Gm
MMe1oqkY7h/N5smrogIEY3BJFLaQc1jrjS1NsUwlhMlRHJQUbtjcI0B0FMHShw/b
1VP1TuqKXdZefFFL3e82ekLuwynl+gXI+I7xDYkY+aWlzweuUxpnVwBWlDhhKCXm
jnGdda9pRqP06M4VO5RZQTwhf49pF4HVkt/kd+xTJZE7R/11tPDA4FPXAYJrb5C9
pDOp6YtTepqSzowJmaDzBLvM/6SXXSPxdPQ12kDtaRlSPH6dQZjcU5pWix/EX5wU
/q1KlR6QjyfBmf5+95DogXyr24WIsuP+b28XoNiJfhE1mWmaowpRB6YaYC+pR+Ae
VZaXXH7mwRGusoyD1Qeojwmf2b0AhCODTtspMUaTrGQkrdysAAVUPFdiCneLVJLk
hNsngNh2E9Sk+55X9fpL5kt1wljwltd7XSJAkPDp2djODwqXOn3VkVnELc/MDxDw
e851S/9APhiX54fsMa/r5YrA1cUPScz4l5gn19xM1d5AxbstqrPuQyk946+xoSJb
q8KrCGMu6FuT+H8u3Yv6D2cO2/QHOsksOM25sdZb+kYk10Io2m75URkGiMDDQ+T8
RdUcT/HZwKFAs7s2AlZNwbS1oFXN6kbZcul1GJxy6rXXbqWZKPXSITB6DeXc88iw
t2/zAKD7BlAWrsYevARwZ0IfVLeYikmzkGaXiYyVLhSfPEmTvmujTu9usTWlNo2G
9NkK/xM/rBcXU80OInOsDYo+hSlxkxB/tkNDJEf6rHWAcnEsNDTs3sgnX9sSdymw
/32P7B6YRNo5tRag/IJB6xrXV0PEf/72M5vD3BCwfCme/pQ/sVF+4dsA3d8H9vhr
lad+VHRlrZdnPRzMUWUgp9zQ3PsbWYl1mVjn0uSpURbWfY8kWWrpbbecZXL9AijR
9Lu5zwrj1QDKV6+Q9zww1LT7Zcr3T5PaYtE35wH+w4M/RH6Sv2TJeSrDDlpgFrLN
Qpw+qB3rv8GdUishF3oRF/ui0P0+ReQ4cHl0Pz+N/mbpBHAp2PYLbHFbmjxXHlDq
7rT3adoUTbXiTJO1j8VAffCOuwvjTSQyZcb9fkAPB/be7P0d1rjUISCKA01oAZ1w
0Co+h1hpnBl+gad9cd9v13a8r7aJVMoakMUm7z1Zp9UCun/t07PMY5JU9gPFPbnG
BmBU8USaeg/se3gJaBxHKYzCPtYb/nhgBW/kBAvfn47K2u1tq/zGm+V00BDd4Uz9
hfYj9o7mOVHc1K6CINhO+o+5PVF2Y3LCCAbL6XslKAw37NNEsrru9PpKXRUA7JlQ
KG60/xtlkAyXh2CTobi7fBpFhobWxh4Go6iwvNJahkvYIWXDA1Q8oq3XJ47P1mxg
OJRcOtQN/9kZOagR8qBvHVBALaSMDQ1GmoHjUVpHELGcU4L6iE9CaZPwOmyB4Uc0
VAvciKxNeh5gf6+yTKVMjx5ZD2Rbb666TSjMpY/TAcUAvaDC2z3OTPsVn+4DLNA8
+rVL9OIffJ0DiZWGnW9AO42vSLd/ThtoT04DoHs5CczIV2xvh8skZIt4Bah9228C
JOtPY9OPX+XtnRP+PM8utW1JfgnMiIY4c4Hcq/stBrffJNIfYT3hhOI8wGQloF1j
/H2sgxf81arW5TcZcWSDtUJ+aW4bhCRu9S/UMvDOBVf3BgsUAiNsuNwGsfJ5q17W
MfZE74+plXBKWagxupgckd7yhnF+kYFBLppo2Ddxe/MWNh+mL+pzCp0WGdzvjJ9f
11M4ZeaeE3AwqEW9a4fgLMJLFqOsxBDU6ssmvhsq2Gg5EmyplNbEWbZYL0PJya09
9fYjrhXOCi9wgH7cFHpXZ640S50LYFJvA5SRrt8rGBWCXczLn8tQvmlt/vb8xQtN
uiMtkYkty/2XgKACwpCpRpFZ+GWDj7wKQ4Zam8U9tfysPvxn3myfM+KNK3AT3NTa
NLZhEZGRGaDM5Y7qYJ2xNxsQsRgECgL8ZibF6+OrQM0swUybnthz3ni68uzieOiY
hyT56FnGRAXGP6LO44WkJZn01ZDTPHXelOdVdNfN+LhmmivNspc58iZb8eVPWvyc
boFii2jy6/MWxYNNrv/c1HEKVR3YG+O50E4oZXZGEltjnMfuat+OrmtpuCgbr67r
vWfqrSaCcIIpB23vUl234HBCGChYOueaUQ7C2ZqAWRM2Y9ip+TRh6ZnmROSmwxXT
T8HmfFO28OjKRKeXWs8kxNy11HBxaX1Mu8X81FOWmNm6CKDnB1sSdxPaExASJY5e
9GMA5SGT4aZiCLzLN3KfITWsecun6rUQVCoQuqGXoVfYbCvNXXcUQmDVw9SuxrgV
uquBTDOjeUktS0wz5/YGtPITeTLf0f0FON78XdFXDW11SJQpPcD5j5sNlumB1z8n
w6zk/wG7lAQXc2q4vC+CLS+xoDSn7kEbSNw9sno30ZE9B05V3KCrCyZxcgw6i8kN
kx7+m2D0nz1dT5EU3KeKt89zlFPc1pAHmWEIgtwSfuFYGT9px3OORiEueXQOaXus
MhflVJPyZmKgTJfgraj/YVBdABVsVRzW0iEYqAA/JbZgGzC/NyPxTrgq8U3Fj8j2
aulx/S3O2Hykfp3cTxVZIy0IuaAemyPLdWXh1zzhqS1Q8+BcWKhElsYv/TASnTz9
sXxj0OUrzEyUbE5n9Mq+eqPyCBq49xsKOo0GCGoSQJf4tcDVviAIfBwkaJsSWs6+
T3nYO2JIpuxx3gLeeBCNAUfA0Gilov00iFpLaWxFR2lrp83tSFfxw9WeZ+QsxaDq
v3up9jONe6Lj8qwywqpcDRuyWirpHy+FuA/fABTPhzf3auS3FTrVXTJeSBbt5A83
WhFiQLkLJ240U7Vqv8L6TXsakCp8CRi12uztETJefcXnZBs9P+D2uvpfYBq953zV
tEYioMXFazoApzIuxcLlcW8pbLE0PgCJ9BkOBwjpXuX8L+vdzXOs9paRZCvApG0I
y+8jmkul0VC5uGH7zBJkhdP9WjrIo0MFL3U58f1suovVPVYRY8LSaUYcYnPHLOiz
xPb6rDT/cbvV374uma3jdLSfAz4p2bQkgcf5fOI9qxMHxA2+CzSH3Ojqf0nwvBCS
1isz0Z5hySW16mzmXud/SHPJPOBIMwwDj3a2OpNabamZH1nC+knqZFHOTQPSommZ
jxghQUBQDpx5o7QfwekpKp+0CtsWXxo1MBGBwVFx8h4GdS7BoOXr9KIOHnImtHHH
v1x57alTRryaPkJCjLngIebUqUyAFbZ+rlJTkS5cB0H1toYKgSd6drfrsz1XyTqx
nphvmNBdWPWkxHc+eoVqPklBMk9hTwCc/rB5hBj2y0ZtyYpRh396xCqDamIuvJA2
TxlPjbIx0IR2K8c7JDA6pZW4jc9lPLAVehmOHU0v5v2/hxT1IYWmb45Jr0gh7AdZ
lGLKb2KQflcT+eZ0sW9hfExVR67EvRNUdgzdoO8gRxppbLxqnfSxz7JUJVOK4cxu
bNtXjrNeVHefambltI3/dcGjjg6V6aVRucTkKaiNTI4sCqdEMw17QhfWvE9YCDiJ
kr7gPBnGABrpOCLLA4+f+wqpEC1B3NIFTbg+j027ftxQoO4Qy+cIt+pi6/BP9Env
oolh0096NNdUNCp5x+7ZciLB8BxJQWNDZhJGRBnIJjmdIdQQ2jgy4WXgoAgmx+Xk
lZ7g4T6/aS8x6ja4GsWv+0xoq96T9UQGp+AIdXrY2mqGa2rcCuxu9BDsZlWntoNc
3T4KQyhyUvR65zV/B551CHVqS7Ew042+USUYtuBt6FQx/GZiAvnR9r2mB3KZf/qc
kFs1/iKjJvOkE73wPlYcgu5mlSzhe6yEUdDHhEKFLK678HQ9yWEuOVhTb4FLb91n
IsBr/m1/MHrhwYbQ5BHciRadHWnHikCEPCnnho4SGQzcebX99kvUWoawN/tKXXhj
Q3q02OBCGrXkMl9576j0HF6t5EsxX3GBHy6r/FfeYlyiURjYDmDR2RzxNI+5Z366
6CQC/giVtS0EmRtafHVMaRYfbajKH6vjOCtMOxKGrSmEvhM37p4ibBkyLY/sqwJ/
dbUCGcPuJgnXGWUnOwn4ie/TlYBBWhZukSoumdZN2oqqzdsvkrHQoLTIYP7zcBQL
ijQR3Xe/zpjwEcsi1r/aDxR8M1gfzXw+/fGcB3hCqGLazUPFXoY5+f1E6qYfReeg
OW5YHnXh767zU59XuHi1sIu/Lk8aDLgi0RRtfGJ8HeuQiad1kTp5AY7Zml7oxNYz
uawRjQUn4QleWc3FCzdB0ikeeIwSVp79Fbje3lfvf2yEtir598BSxyEQ30O1BiYc
D2c227FoI8eJC95nhrwVSMcQbr1/OH+Q3Oa56ZXFfO0ghnZEVpz2UTGP8vzWmwO5
tEdKWdogvo1gTMjvFb5OFF7LpYY2OYSpKk0jpkiEXJLf3X0c/GzgrRDMZodXx39u
TD5J+m6ZNR9lW0UGpL4e6W/l5sBYygz+3e3Ttj37lclSuTEPTEkh3U+YssGtr7Xh
yRlRR0U7qnL7KzPHtn5fzUjeXIVikT+wzRLuurFUTBfZARe4l9eyXtfuV8ToGnSM
VTGc9MwKihUKzY6YcjcgNDC3Hz/s3OYEr1YBVvV0tPAeeG1o8KRB8EyzRPhOMbpR
Gb67DIC7t5nFww1NV8Wa1x3HYGA7DRAYuCpXmNBnqSU6zLmKekjHtRHMS1Gz8CO+
2L8NxK8JQLJI4pYqy4cSyt1UFFugiSffehSIiZizlhG8ofKqjgCcKwG8T5KOmX9f
BvldmZG2V91u6z0m7X1vOXlRRER7MIoC3cXr+KkwoQeFsQ3P+flDpgQ0PwKqqcFP
CrLOV5Hb0P7bPkDw+PjcSKpAtvz//hVgGonmc9zHMYyU5NV3rmnIEbB62mBoMyfF
M1oYp29PMdS48EKD1V0pwOMq17dYhfGtnzlkfvg6oetR3hfyuTRh6Pnk+LpkJGKR
7ghyZlOHpeu2P2CKRM8TxTjPyp69Hmw+a9kURZSAVlNLyGg7EHzcLlfbWcsnNqS9
WHApDl+Ggk45YtZbhdaK+q7WW3JAcmW2Y+DHEPFGPcPtY9r6Gx6cv4jjZWeDsZpy
n3leEDvg8xuHNnXNAwdz+8cZwE8MJKY1PO9YlWhivaq6fSkxGgq/AiQUkZz06FKY
j/IYWPgvMyc3G02bIS+vtlf41nLbOLJijpDmBlRiybq5LNorp6B932j4LKOLDl8Y
FYV6rCr9f6e6QvXiJbfoTC/2LYyUFdTam89qIfBiy6vemq+hsyrYdBPQQd9m3PYn
EpUCh2tCMbmYVKgdr8Rp6RRJZdRnxoT3ir9xwIT87ft/b0RBK1jQpdw+YAUMWT82
MHAeNGMRziVqgZV5ii1pIDTnWBJefoXJEGQ2r8BOccLNXecJUzWMrMVvUqUVJEuy
YKEYKNJ3X8SjfkJ4Q4ZoU1ciECw0YR88Ieb5Ex9OSb2qpczOE7+/ZRAvKymNOi6R
QZt7mHsrMeEC2o6hYBlA24XRqCyTHDkIe3xWBO1cAl4aU0VaQuUNaxCgEsVUtLvO
t1PphVaOSH5uQJgENgIu2tpZyqbZu4G+CcPxBnSXFzO/za5oA2HfUk/qK0iBNxAv
+vHftIoguR9wr3HP8vokuY89JmtmX+13m0npLnArEf2/UY2cFiduR6DlDhZ+LwVV
GYGG8Qwvjw0NC7eOIddA5H1pYxqYvtG2kSMRMvfKveBf7UnFebQ4bK2NskiMED4+
B1gMxRj4HvJfuXluVYwR1cc4TcFcjjR4jQ6GMpSiSBHkyE32O3u62odKBjF4RZ2W
/H/qJ4+94wozgck60PZC+zwbcHANzL1Ur7C8h2mttQi+Y0cJVc6K+y9/2GbMYWV/
JGeaujQ6ew0/zDZtXtjqaJ5HFU3I1qxz6fkPFzDXvRgnsboHzQQWmVzR79/Zjy5E
BnMNlw6LmS/+AYcgJKeVGSSiSNUqob7sZ9IESQSjlDCxKNHaKHADV8bfgaJyNIzi
6mK0+PLtDv22B6wTQmLe9cXrZoTXzq8SsaS4WFVzpOrSRXc9TQLI2WADHKEpsrhW
Sz+iBtZBq7VxuF3zRfD3bz+MAvnV8x3NXyPqr1qI6ozmOdKl1WOOJNp6aoKQcgPJ
wefHCqc+cdSOlHLvvqL3YGmZo6txTlaJuLFcP/UKQqXOlU5pRYZlp+QrZcQ9gIue
vIOaS4SgEhsuFbbWSdULUPjNsiTJX8TqzSnxPMrqbOFJHFYjyFM5J/c7Jz5XblwT
Iz7kJOMgHGVxzsQn8EEuco5/u4rHESzr3eaTustYmZRO16b6/nsd2X3dwVeWkqw9
JDM6OefiuuLlT+3byITDLEw0Yi1JLoayRC3sq9JMPLYWnN8dgT4M2OE6lF0rLWc6
CziitgW7cCVV8OFoy4auks+UGm08RRBiXNcAwoRLaQcudP1kd+w4CHtOaYQHY8Ur
ax6Vv0zxEqBJDdF2Dfwtds53/C+knAp9pbhnu6eyB241wxIEvmAKqwqrw/hFV7Zo
hnVw1x/TB4vmBskrfAtBUXJ2L0ZMlX01Ey4F/ZOMp/95MX0Tm0j/mTaOrD5V2x7N
unyggfBoiqDb6o33YPcpYRiu7bsl+9WIhkfDRwexX1CZoFBJPpChG/qegWWQK7bo
ZFWRh9MJkMDZSbZ8jDtepEtqF+Avapdzbxc3IvaIwJHBV0wG8Gnn9FIz3iQbghxO
r45WsohI2UimLhXsbbHIzgKS+v3GTIsl5OlYX/f2jgd40OAnZyv+6gX9szuUIbrA
3cJC5L2WPjulFHjOetRhqFhaMOaBqmYIadT/9khjV9T+pGfvJh9GTlxY2/1/mxOe
m0RB6DtIjJvCsOHR/cUe3RWsrSUWH9CHl4eSnZc/rTGVqA6oBlbxsDX5xsicT9Vq
bJud5Ci+nD6OYE8Br9hGCXUm+Ux8xbAR4sWEwPIODfHqbUr+hWm7i8feukLasTwj
gJ7A0qqsgqVie+YnWqtuudM9MiS1+gO39VLq86096BXA8wCyPJP3hrvQ+MmfFSPv
pMhIvxufEc45yNAXAlp7QN4IXflevC+mG/qXw7Mca8YSCA1wcEsy1tXsZ0ri75J4
AU8mkdZYTuT69wq7CdEzseF+ls+g/PIaLfR1v6GFX9p9D02V0Au0leh30C7zc3NO
aB5eftxlA0KY1pKrPwJJ5oyK+iaLWl24Ay6aMuSE2R0IqlRMC87mI9sB3fb/qjoy
ls21MtHYgWCiqz1abEHkCPAjUERa22CnivaBj/0YYnqlhsEQavPLO6+MOj4grKrR
YZOWcNBCKJSY3vZ0jF8Q68ZB9cksknVgWzR2nS9sy7J8A1SUZWgwwKl9S3dn4zTU
WMqNVe0TGtleUWiQQlozNRm3QdwwVv1WfOsZsNfKp/wrdHWB6ryvT+/iM561j0gE
OLrvwlcVNOwyBvfjnJgb6ipK/8+PKU6F2jxt6WXMqTO6DT3fAr3Leiofqib2Z6/g
/CCQuWjoaAQnIF2knoiyGNXFogqV8I2EumWcOpNN5akthobVnF0rJu6bOwEcbenb
yOUxww/qhXBcmuBiXfO+zzgtddSI7cQtRjUSl/j1GTzcOcsKhGrYAKCHKnyWU2R+
I1ipN2lT/gbLtBKxeP0UtP/MMhoWrW87vpi+B4Pm69kPD+zdTLuihUvW0bE7+Ily
46C4ON7FIZ9DXkMLyMvSyM5Lrh8umTevboUPFkHQA6JhEFk3bSRRQptbHz8AeITM
xDLUOvfZw8UFl8y8IQYIPMKCSMcsKLjm4twb6Xu84XTInT5FMPB5Ue+AULTi+7YW
oLdmtCg2EZDERVjeFop9cU1SsqXsHPyJlSmgnCw6fd2Zgop+6FAoFLJTA0nfjWUt
2mRE0pBLfr0modhXB/9qmOtbyFO1aHOALfTyv3dcwo0qZZfIiRHeTmyS/Q0n728c
abYO7ZywSfLONnuskY4o3xoL0GLb/Ns5oxRZ3OEi0aMRbzvVg/FNo1l4umcjgHaT
PJjQ/uGhBqLMudynTuC9PUJ9jJtsnQN82UR5iljoPQonNZpGNKvdVMuGyN+lmd34
2KEKX9Vif2Skgg+goGXfDoNOk4DuhVFNHOhYdwzM0s2cOasWYM8fUSvuseFGIx6R
LVl08JEnOZMjOYTkiDQd+5TYwlUr5G9+rT8XyXLx/xBlgcDROsUP8/D+tJi1ElEq
qdGgCRTaAVicxvjgEhbTwlTtIEwOJbtyw1bAy3HA0RzTSPZ01PnK9cygEaKY6X3P
azJ5Ce4ZgJgja8eZpKe2ZeUzylzwuhTPP0MLIP8v6SdSm6P4EtkuuSm87fNOAj7s
CjNGwT613eTxJLo0C2+xY9USrr46eZjjqpAd+VM4oPKPV+ofdzD/WSPMrLvYW8vI
lurXiUDa4ive2xSHFb1+iDdr5YG+Fc3ukXDWwsGdx5cMtUBbB+QiUY09wb58pGZG
oKHh4wPIw8MmVhJajrZlpR/XWbhQyrNBavK+w5hNKO8uVChpDPZUfDbJl5o5mCLW
3YiTSMYDUjSacZyJq/Vu+guqVIGRSCaBFgZ4QHGJNEZMFyO0PYd0Vn2zWYkHRJ0s
0ywaw6xPLK+CKOka+KKuge1iuIDOhVD9UK2SCn4lZ0AyUgZzOC+hRiMvHDFG/shH
uemDJ175z6RAY5G7NJdWqRcxGef6yvdubwUasxywwsYwEl36sh7CAMANf1lBfm2e
CG4MR9Hh48h0ULBM8mKwoGeCx2RZmmgAt5egUc0QJhVtyeBAP/tjGPwd0pDOd7Ua
ZQdEs1Aa83spoA4PBa705c5D2cV/rkeGS1PdkpfvEVshp2HjuxmYNGwLhZR3mCbp
+F7mAj06aelH4jJtlB4wtjuL1TR8dPqDXhtlJB2y2DTKv1D3GoxQxMCY6miopZQm
rMq6iIQNBVBKYxE0giXbgHYz9qp9ghu5GEEp1LYXioaO0YVZei2XEVKiU4tDgkqK
ofoKzOMHZfFPSDToRJYs6MIQWupvFqotLOgwgG3QY1XEtbG4zn4jsAkakXG/3ZRD
j3TycB3uIEe1rO/ZFM5m22AMOqoTcbkLmt/yDlgY7HGZn6d5QQKmSXuPFKzbUrJH
LQm+FG4UvVCpCfLzsR/7rEHZlfGJt6B2oxy/JLFBFMS7XaMYjmPtmdB5Ol238KSM
LuOW9rJYAbfIZ5YoqA7bagvZuttN35yQ8H20Pz7Ha0fN6gX2WdvM3yXKBd/etZZD
dD3Fb5xmaIFvoZJLTURqah+y8tnl455CpxlNoZ5p0zgWZdgI2+3cz5TDCY80wLs8
Y5TCewiOMCE+l0sjgy4C2ww8x1xS7cL/O9LOq+5yYdbiN+K0N/A35OQxSuUW4TaH
yk6m2DQTUXpy1IuveDu4izZh4ucTy5q3nSvlBcA+9qkOOv86C327z2T2/H0RETq4
VjcPRM2BKNZIrYLWriUw0CcnjJvCVxZA/jiHWEY54Mdqbqq7utxU6fT+mMwcvMpO
iBRsUD9ZBsvgf7opaTd83VVuD8xS2QqG0BnB/eBGaenxuK2I1XpOn+iT2DKXyZ5B
6hntPEDdf9ZFNMt13Cp8952+6f8TxixVWC7CkMxqNP13OelyisX4NwOIaKTrcfyQ
/EUqgGclI45mLKgOCjT9VR5aV8/qeTmUTwr4eqkczHjOa+fbxpQi0LXZG01Ole1h
bQzcVlRGVVBeu9SzpxBOZJ2fgqrqo6dYghk3H12V60JBWEei7cOSEyG7bAMHthBc
otYziowfPtFfRqXWIj/M1ee8oX6nprQJMlJNcMOteBCfCteZgpi9i/ei6l/T/8vH
SMKyOfBoesYY8gW4ljDP5A==
`pragma protect end_protected
