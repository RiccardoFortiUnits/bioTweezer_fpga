`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c7zcI3gfMTuudRESnB90gimkwLEWqFwg95D5FC83/kD6lUi+a+/PMu6enxQVg0Wg
JEQOKZGzNsuNYtp5oT/VidpM5iopSoeKx8J71ppei8gefyqMHCtz7NbjRiMlgpol
+eoa6Zf4mkJr0ANwlGgP3n0mdqAC3OLdCtaKtfqMiiE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4416)
D8B+Qb4SvCEFAna46tyrCKJjYfAInWGzsldBmCCHcPF8AKzFldpWRhHgWZZPZ31S
sbRZd2i9wBqX9eyCnGm3yVHqy8K85JkkvK122tjcus/2iX77FPrBAiHo+1H4paCI
2suqmyc4CSEee/gq2LTKoofXZ3t9P/TYvWLvA88GQ6TIoXZAT421Su8JFzTPJxak
3IdfFuqKBUHx3+szqLe7DkjnXQfcGmPJDAgxKkiYMIRx/ohYodm8yHwibZqtzt2M
6Bl87dEHG70wiRF2T+Iml9fijGxPLB+ULrOp4mKncffQVZyRI2cbXycUCZHOrnjV
hVdKH0rnWLpVy4vDXCbCNolBAB7mY1Ud6BCx+BDfL59fCHecaF7UK/f7d1mfEb+S
jpaVBh1kPMn9bMT1rVZRpe23GZfsPfXAYTwzvLb5y4Byi//9J8nG2bx/9+EmZ/Uf
/DT8UfhmxySmw7Zr53tfyLXQ6P9WLtd2MZuqdsDSnEFSqJ3b/fk2sCzuXDPTRVhv
uxooGU3I2GPv1P0Oawq3vHEXeBuCab3DBZlCWROg0vs5lzWSxolS+AtKZABmuRi1
AuywgpeIZ/YTNhQE8mZFN62i0J2Y7RQHhSgn2/opH30X4ShkSJJSUiKISpFWQ5s5
7d+rjNjpwJR6y1tubHrzKDTQEo/BPX0UyJFhbSfIAkRumlDqaXK+Ag+qQxZ8jic5
v6Lo7kYU/jjchgiaOsqcPs9tTOKMelJkD2TnRnMd47PhPIrR0hmjj6Y60KNBy8kR
p39dNRajWDmGqP7E6gl+FJfnyi+ToSu84NwVr1cJPR9N9X6Ird0lsb6r8nsz7KcQ
A+dDuDr1ux7ScFwNIVVM8xVB6+6hX+qBD1bxeX0cDYezHpdnYfv025q7L9n98mzv
mkZOvhPmegXuvFKF059CIFUKRbmi5ntmiuagw/NUithQpy4npwBNMBTz6T8/z8Lc
gHFs7hxrZMqE5nKnID7Q6pHGTpdxgqAcn5WZCnNQT9zKncYKFJCLivzwhd/sRr8K
JGKYqAZdeEKUhk2vvufYyDR/KzhdgXUETK1SHzDPEClau4DvhiJI+z8uPfIQ4kqD
g/K8rYVU2jBK61fv64X4JdWiM0jiMugNnQullUMkhcKvydZplwV9XdL82G2rqweW
aHd947qY/LIVcY5kEtfBjKVPBMXH3N80BDa9fJi4nmAcuLE7NXKGWxfAS18wwlM5
pQjQiZY2OP/y9D6PgIn0rrtX0ZQK6Iey+Yz4hVf8qqDXaztuEry3snDxuNOvaFRP
XmP3o1P39vqclqpna3VSHfXe/sCP+zKttcZxScMMjuk+28AV0R4nLHFE9dj7Sixm
Ofa2F9g/zPgmXkKorlSuG+Y3kJkKNxQMyMMc0X+mB7HONbq6HBXLVpB1fJVJU5UG
kT/QzrPZAyJpORDwv2Bdc3zXZtz9P8O8Fx6LOhCZa89EdnBl7SorH5JxXns3FjHz
VDsj+G4Oro7MLlKPz+M0jC77pDVfzCW7RPjxycCe8ol074V2wViFJ0r4M/CW1ybI
cT/Vn0KqGXVi+VsiVSz4RsgPoGpfWkex0UHMrfMw+sTMQN0mVcK7CUlclGPpc+NU
DuRJBdy1xih+3GJ+1QLDoEJYfXFWeuLtFCZIZmz+k3qhonXjSHUKiPFb5V0jNn8U
8cbivS5z6CCA/xijOno0FedOJVEJPZyxocOzELx+YULoJ02ULG0cFjr0GXbhYNED
Qfnahh7DIKZ1qBjL8t+hLA0EV1SatHtupg19i+hU11B5zp7P9TXz14P1MHxHinkw
sA4uV5E6E4hjSzfvN3JsBi0JO28N5swTweuPTM30kGT7/89bpAJWZDIOiGgp422t
9CQQ+sY+5uP5ivAIQJNgkDeEh6twreJo9BxDJRw9fkSeROcX6ytYPZFrNNTBwQ/N
A32gRVDm9e7y9RUYadtUvdHVLP7FvTvtjn0tF2n/hlmFhMv7js1n52alb5nmSAFr
tEjZffo70Z0GyztHgStDYBLwGmk5uc2US1bGUJdxNriRIb57mgxOi93Gh3NK3lGn
s73d/YBNwJVJSrry3qxTPfEQZs0H8dC5vfoBGX/NPWJojqhTiuFRGX+aPgSDEYHd
u0tunZuKD/nuJUF+kgWISVg8SxKgafSxSgrZwqs/HJc4KVLJF/wd4WA6gRfq4d5b
jxq5jxej2wJoMadzAnl2WKRPV+Avp4yGjafAzguHzWLNGyC/9Mh9FK0P+mooi4H7
KrytvuqeaOUwn1eZP8dhMLrJmdwOWr92mX9w1+TqejBm0Q0CF7/sUXh4G+jevc/3
gppBURSlLN7vWpxY9y0a0lAcOF16X4CHOU6+kFCSBwmD5xuz96+Ts/Xupfchrp9m
p0hGBZgnudpboEJnaenMSFUPbpfB0nFtG0ftdL1Tj9i32j/BcMOSqs4kxOXgcYsq
27ZKQAAJsm7najILBezSkTHn5UPY+9zY/gctjVvVEP/5kdhP66B2yn2en7UGoslF
ir0XK1K7BVgb6jmcciTYDLP0B6f0dWIi2UnHG/HvG72vR5aqwwke9L2Pg5T7HFs7
2PHfiLlrMe+7qyXj2Jtk7hE+veYHSNAWPX54EysUUpYlz8YwpkKzN2PC1jZ+oM8v
VvGhXjfxQABt3jMvTvkJUiveHxazdCcj7SPlvJz+ve6UWefLRze3pgHNgSyodzis
JBKcelE8hzLSzv3gwgAFx7O1lCushzWk+9jZM0nHB0m0y1FiNN2VTndU7AMkCbjb
NvBco2QcG9lBK/o/5uOK1YRYxwwAlLOE1TNUWnF6GQEQNGZNpyGHfejUintnNKky
uA02Em1sZkJ+o3cep1Ztxz4PY3rlIz49OoeovAA+4ORKlrjIxw6uDtNbydj02Xfg
K7y8iL9a6XBvMvwyys+FotCoiAvOd0SfKyO3vQMi430j8UZJ/kPVTff3KulbqtsP
Gr+bXqXWwwtf6RydN9lUWOPPs23uWD41qj11TEKWmtjkl5NtQChRFLQXNugfSJ2b
Zt8IG8qpteIMlRSKzYxXQy0fp3MG/m0miRO5V+GgeUfRtoMfafCIImM81yIAkX5g
6sqpiEPe1yHznSkp6rVG3NXehY1bfzxCQDqxYkEBuq1qoyaVxfCcgXB2gcro5h/E
gYe+6RdLEx6OiO1EfYFvu+vGzHhU8y/rNHdrTejNHNIxZnebFB6w42G+bloL+jcJ
9rFm7nxoNAsJYTnsCNq1KbhV/yplvfk9C7duHZ6YuptgtFhvCqreRx83yEJUK52K
2TzVLT0+wcWFnHrnV3PWKn/uaVkTWkqjgX7LgxcN6owBcN9CB4aoFW2gts2T273/
mNddyKDvAC7Klu7/sFrMKzWcB9NnmaBAdhK8kNoKOIo6+VGoZ6vNA4L7dWFM/fVo
2Tf5daXsMhBR8X9CtFow1d412JRqD0gJAW6j1TZj9Dx0X+QKcQFaSAdjnS0vRtFb
62UUmlxb997MvraKGJi5IWy3z2c9ERQf727XCf8Qz+/wdqKKEoHezEPgb0ZMxvmZ
OeOQwKpKjZdcP0HUOwzNW/fMx7DsWz1U7V4dv1d+rOc0Pm1wSEdcd98TeZsKB+vs
PTJNv2uDyDa2mS4yKlIbfahYzYw6OPxpG/8/C5CWrnYAtrR1nhFwUcdxD8LFS6q2
itC/Daza1WpspA5TIvkcZ0Hdse8migwPi12SxCVNQ8XOJ3LoLRhpTu1DLBBm+Af9
iEjeSXpVHA+WNhESAuMpXDWlGyd2fLhuqdwGelV2IuvV+Mm0GmzBYRhGR7fLIN71
5dMFFgYXIIUM5xoyVM7uHoMWjTsu5euJ8EKKBpNMDqxVk6pena6bsLorV5LBUrLS
GZzsMpNlnfFdY58BGlspGosjlhJg3ruJJXqk3+3uBOus697EmUlc9etLKOLLaguz
+VZs6UC3Mtue4+88hwXOZGGx6RR5YDuVuxQMrE6hY5ZzFVOiNcfR2Wn1ebMWweFl
vpm2854w2T50nVP4C58PIjCHXNbFhAdrvNTkDJ1xODdMoIoiFphol9oGcxeLmg7O
M5gQLfyK5cJPU0VT+mmZzG/418INF5vJe/3JOjZMGQIy29ecAhmulV+wihTQrQLC
7G+RLXGE9GH7KDQW1GF3HpIwmW5Q920otWvMCUw1Wg7RGSUhy3GnBT/tVFygvskI
IciCPuOHBFKMbN+tjFuBgjPc1uL+0xuH4vBmno1riqVSbKWUvQUUS8yXtFvpgnyg
72zywjEFv5hXkLKe8Scp6ncsLCXZFH9I4WgHkrj8s2pg0ErYPBHzo9WhbPGLMXR0
/6pmYDlWlVZ+aORXvh6ySNWlZqqYa8e/wyLdi/BHQXxUpybY7Lk3EIMEtDh7xJVU
wtvPwFzj/CQcZAgcGcM+ONihfThszMbBCF9qFi8/qROTHWGrJkrU6eWKB/15hVI/
RDK73g4/fTL8AXq88NnHz5L4XVZmYWdor55csrymkJzjQDUz8DI3uMnvXmp/RCWj
G6p5iAVAyK64xNg++AsTivWSP6CimbBWiJ/XankqV2YmgPTA+jTsvRJs8kvFtIHr
fnFlyij5e1QkA55eWxWfCOTeTjwuPyVLydkdnpPcW9vz80KcUpDbOa7ML4iqlgtq
uedjCNh2+9RauL4MbK2ozWfbhu44Fx8ReM6eCj5mggiOoU8NYRzCMgiNu982AjGq
At8Sx8DAZ1lt0s+UrAoKmvWf2TS1YAsedI5lTTWacslAYoW/6e4JN3AlIZ/Ebcyr
cbyJqfoEPE0732Hxb/L6UUrA0jks7C8Pij+K/Afp7v7FL5aApLoyWKeqysmrgpJd
RccXanMn05YFD6+Zo7dfJ5C3JtUVkiYLx06hULp0zOrJ+1WNmz6kI3bryVzZ/4hR
I+I5YENnHiXdYuUW8TX88Z071pFZCOGhBMTuZI3znx5AcQXp93f1CgiulPBzgjb+
MRHH/WZmuQ2oPF91XmmZxXhpIX0avtVc6rYqDYIybSa4wy9upDbW3Jp0mlEIb0vR
9tZPCiCeWL0OQecKKtJEwZN0CNRtrymAe+BNem7Y/Nqi9tcKoI1UhHdys4i92B4I
0HjZZU5fQ3YkdUwO7UYrXENEfF33i4RnlQABbjEkngTqT1wKJbCRTenlkfZ9fEvv
bTRQCi9FNWBRl07vTrHhP/jxW0OEBkPT8dHx9aQRNNST4lXezK/mh2a/grZqculb
I0jR4flDfu+JK5aveCMrRTTZkpkuGwjM+OSbPv+Eu13DK7rB8J6GDZZjcneBqwxj
rLcOU/GbAGsp7lqAmjnXgl0aRdq2ahUvOHywnjkoCRh6Iha8pu8XcS70ainKK7+u
D16qoJXPKcevMzMRyanYDW+S0k6y3/DrAq7aJjFlv2SQLApY5riax3zS0STnmidi
3QZc/Va1hvSLRHpzJ6vZxcoyvzjp3Jd7YhZP4tWQQvFnrlnzlAzmsRVJ0PDE8EtZ
N/pQXlAsM7630KQDgHSQfm70685ZCz9s4g2zUwboO5I8BSV+wkoFCLSHpHa80xT4
Tnb98DSlUnjPteVPE091IAzD7prarABfQF4C9tCfNG13ZdJxzKMoBh47qlyIC6K/
bQwNY1BS/cECOowfiGzVrElaSTXx7u/eHAK0KlL7Gh3b3C22TBjLjL6HJnVM/G1d
dFtdhd0pWZlo9bqdknFnE6G8b8/rWMZ2ZlE6PjCS9NFBKVxpE+O7fU2j9kqi9FEp
U0Kc3JjKTKWreDi6Oo8COl3fIINPbxDkL2n5cjo0LKi7SZJel/vGQNQ+oXLY7uNL
3bpdv8RKwvOyTz0N8IQvJsTjq4dwaadBFeW+jTDjDt06xn10Ecn6/Uk0T2dhoHcm
CunuBvrHCrfLYxO64Wh5LV98rwFl5yfYwzHD6CdGhCGaFEgOYHCKuNHVRo0IvWIl
`pragma protect end_protected
