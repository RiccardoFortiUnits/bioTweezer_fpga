`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XjwcQ0COaNil/xzoJRg9JA8Rsx128SCneI3ID7O45KtRZb2d9CtZyXNhHOMOvSVQ
rie8T2le5Gj9rs1yB3kdwT6QpcVqkCQO2kPasgJmmNtUos8UsJAzitjMgsPrleCW
upflDI/ylZJSkN1cUDEcXck8loB//Dupb91nshaeXw0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
CWGfk20iH+vV5X3bv8wtUrhbK4kM0kRfGiig4F+7yCvV/JMW4c/cGSyZQ+4f3913
ephi8ClqTC58eExMn/G7NHb2MymBi16clF8zv+5q4eqAQPPjma6sb8xQ4gFEsaW1
L+IuBv/rljMIR8TsEE2K17HqifsMkqwPcMbc0w1SY5jB6rqO6mQuvcDice0hcw9n
lfYB3EkFgg5qYVQFtuReErmBTzYjTcm22Yi9XNXu5gLPSNyzvSgzlBCEEaayyNog
GzzKR2lsxQisU6qxPuLgJRxVshJkA5251Ow4ezFGdK3ldKYJa2oyvm0v9gUrRPwB
mevUza1ug90NOCOcb4a39j0EJUyAAkqIyGCaWeHyloj8ZzUCgPHoCAwoMl5xappZ
bWhf2gGmhzqExHqwHBpWS7uohCXFC3u9+7CKCkKCXgw9eIaZFkzoJBGk6URrxbqG
VKBE8J38dbrOma6aS2gZxuqZbkWeNzvyvT75oXwDWCwvbs5al6afQjJdAaX5ewOX
9a/LlwT6eCzCVzChrZus7WzCyaSP/uUZnoJ8pRvljVvpVsouWbpoXgixeV3lF555
IXq8YcmZn6hqg8W/9RsiINFC7pvBSxDCpKEZeoBKzGPYIiyJtscIZy0AuIdgBZTW
HUwHAfCHV8Aq0DtTiroEwOKgKd5U9RJwmcjcFoq6+HNAmI3D5bnkHLpCK+kQsYHz
guYzv0mN6fVJEQMq40aKo/9mWTv/KFbsn4BrynZGzUqWqhUYWDsxFk/Z/T5CtQr4
QSun02wSUI1/3Gew+U+17/mSS+nU3VvnuQVJCuucDoQf5sMUOIP6dJ089Z+TLzEk
HYOnJz6ePE3pSCM1xHu1TKw4FKbKwtsQNtZGnHI0WoF5zHR/cMsJ3JcqgQNcdMP6
hOUYS4D4fuADEwH148MEA73cFtpmB5UFJinyHanc2jCjsNhVUtBNRG4a247mrl2L
m4SaJOqzlNygRIj5jClA1aPDpiYDMwSjREhX7HzJN5fLvkQBM4ffn3nd3fDHRqBO
UOL66Msaa8EBuy2MCnfyhbkyLB3udDRZBb8mbylxBX6Hec/s8O9VY10/TdYCBX92
etNHdRYZc8ZK5TyMVMu4oPXx8wg9+W13ipMYnXRWnccOeUNFiPCtgULuzcoo+J3M
4zTj8Skz18WfusuZVz7XuV/X+n2x7dhqx3MOajb4wjTRYekiQTN5ER1B0WF/RG53
ghbKIoBG5rjVBtLEYhHUU5rLaqm8OyhAwBVVY5Y6Lr37xdsO+6MiGMFf9HV/vBjf
jLP6NXb7UhtyRNo0j5ZnySGt+MvMFg8Wn1M2hCSj8bvZyNaCC8qO0404wsFUpaGx
EAXIcrpPRw0ilMm8ea7pmPQEn5g+4CDA9uUVosV+hYskENrxQ7zOFurtJ+vDe2Y1
/Aupv+6Oxi7q6LIZjhR7+wpRZuwOpKCqpQMWyxS1dmGcvnOuNTTXzg4UKrsc2Z4Q
WzyzA3rLAFCZteNfywlOHrRuIs78i8ZX/sUIa7W7bQ5scnfW8QyYfrEqbzXyWwJD
ZspGLE4hauNPXm8lC4GYDrZSXONYpWEEHe4mVJa/iBkX4f2vBk0+6/cdLu6m+s4l
zOLIlop/+t4yy0/pYuRcNOSqezlz3JRj5cefBNuSVpkMOVGZ19PcS4zhS7mOLol0
4O5V+mpMr63cESl4UYuBe7pqlMFNQN5BgaWZUv+yNPtD+2ORI7s82bHKkSc7OBfF
ZBNbBG3YfD2eILMdjZs+HrNJjMcFpenZ3YCZo0Ovw801Fl/NIIt45XJ+9EGfIe2N
MNv13pVJPknb6JzEIU2roBr39wTfGAN6XKxSDGkTjqp2NghNdL6dYDAzjsGQuZOr
Jc9Qa/9uUzwlt079CTfrWvVRNxMXAovIugFsQV2lmZ9UcvRoBV1jWeonF2ECJvWQ
9++wl7rZvcvCgILclvoCy6l111Q1DsgiUvApDrWLZK6/KwwzOJLS9tIzKwjALYkD
iILg4MHfpa+jYI6MMNMvKemsckQrlcOyvhYgMjw2AFc5Q8MjOHkj0G2QyFns9LKN
7l5h7N2XumKZjsVZWPkyOZcIEj6elFUmakZhW+9GwZjGl9hRA6+otPu3yo0w/XTy
AabCm65rTEWWcFeRIqK0uSgbCkDlmbEcfJ+u5NqxbKlyQkcxmcLpl8avv6cEOLma
qi1oyNWuqHtBD/OYeeC+YxNJ3V/vybjs2hcIOLNLfoBgy0gsKRhu3/A/CgddKNl9
ElAzGCC181s8IPkJ2N+qRU4eXVE4K0d1cvq0rN9OnQ1tYu7fVrlnvGNMtVGJbmQg
nGLq/vpmoBRIiMHiWAXSjdEa3mgjDpznkCE/HgrVGipLbfat3r0X/VU4BIE9/kML
AavaVIvh1ANy3zDJUxbBT+lLnt0WRA8/uWG0v2LXobHKCCfzqELt/PWxk5XyGqQu
69pBUVcT6k/K4RrlNzthTWYHMB5H5dZaxILtPLNgelZn+gHteX4ciorx3fXEdjJz
pqdNjwzD1jYWS5Ur2UEshII6WBdGUVCJfMeK9GIXJWDKzC4RUkO2iJK7LGxQTb21
0F6fwks+sC+sLBE3KZVi6eJDVWR48wHO4NYVoMK3hpzWFMjtYfPS+tNinw7mdGV1
RuArF9nIBVRZz9CMko+E4AlN3aCD80HoA3ZAcowZolp9ExOqPgIuOsvFxwZ+i72J
QbgcLMXitZZguSbgfuG+bDEzXYd1ZJ+fmXlJVy8kKowYydM2MYqqV12hthr97gZs
rfmRBYqD6lGcQRB36UrAX+MBWcw3RO57GWCpU9FEZtnplBAd23psY4OJar0VS+su
0nil0z6YfC1zMwCda3V/eHbipec47ugz5IhqtZhukb/opFKOCkAXP8UtvfZvp7Np
ZcFlWRd6HYw2hoaHI0GGrh0tI6JGpO/GKbxyoSsYrxfTwHABE3tJk0gU9FFl6n2m
1NwkSUWv4f6hB+FZ6xrQLt978sHMST+3hrmjIsSe74wSHApjXy+kxKVZCJjAPhie
c3hGAkt0gqHR/HE/uX6KX7fegMz0G8odtKwvWvNN8V6oCUiA8aG+gHcXEE6/2ihR
IbXm7aJvWulKro0wHuQGL6vcBsQmXez7qKji5IA3eGaxED8jEk6pX2utyTvuIdh8
HHmU0iof8q1PQbxWnlEKfo+5T1+tRc93OAK0Eo2ubZG5NzJlg3wrwW+jsBXQmsqb
Wb2Jm9Nlezqux3ALFYixO+ox7G25G7j2xPBTYBtdfbkID7ldwYidQrwKQMWm7CCe
is7v1tTBsycSbhkNETqXJD/Da7Jps/gE0Fly7ZwCaq2QyFs0etPPxDbur8M+Gd1O
jvs8ocRwz0V3d8bYV7tC4Yo7RuX7O6Ot8oMBnQOk9JqhygNNmNmkljxydpCohdGZ
Fmvj7QWtugWtnOWq9gpOaLy86HmkOiIoB1WpOsg3N8qtvoBi1bXv7zFvk/lG23Mm
9DMJfqDBF6RGEJx0uVAtBOfM9NzQk15lJX/ff0f1jpdIIW078Dg6xHt0PldqKUGj
4bQgaNkrIzNpJcI47hXokhcNklytDJ6gl9xkWOzKXSd1MRwW50vrZZpuNdqoi3H5
susXoqo5QNlUWQyYYLyjpmrtXp4umMLRVqQ6FJE2BTn8VsTrLNZDIaRhRoF9eo/O
075clT6Qz116E4tE1Fs/IBCE1zaNgvl3+GHvTkClY4L8UiuXZDyeS5i2w/FfSa9Q
1vhjyNRp1NUKk0usAtPudNYfNQCyVrt/ZReOGJBdbHA1e3waH24Ek2OxQs/zIngK
h+MePQG8i0ESf9OZJDYbIGYZz9s08Rb6QNW5UaJi+T2JUPtnkuyD5tB4xj2tFKxS
gn2xTrIL/2eQNAn9q97CRisMfmtkElWw6IbWVcnsyBd3yE+4Obxemjh9xtZPBDH7
mbyRnq/105N4i1wwodlBt17WogbbmltnvZHqs6Tj9ufs5Le9P3QY8M2l+4hle0aK
6BNwMnzpNMnq7JzrQJJWkFneZIn2xkFnJY+bWM1NSa8qkGfkv5NWqxA0rpO3LAyD
He72FnoBdno+osLuUh+Q4e1FDao/7fKmrBwCUTvGQOM6/682ZAiXgqic2hlgNUIs
Go4LfceDGEAWKzrvtYDp7yrIwWrQHYtlHzmrBjrb7F4XxaZjBQdywNKIdnGWHgw+
4CWlGr0rRyc4plOl4Et4T7zmwfVx0w8165x9aPyJUQp3EYc5BvK1syyEL1cLoz4l
XBCn/NfjSGhhobaRc7lwzY9+KMNNuaiY8x52f4txlxEofwyeWBAft60NoLgGTHl4
kRH6fZlNM7e5q3Cd9DAWtNm/FZJoeh0yByHcwIjAphUPdrmnejkF5rtktZtWddH0
iwCoafFDaikXmID8k2W6OVN04TbYT2s9tejd7+o3XAT5tK9dQjzSYzVOjVDnGtbn
C0iDkwuGRv7NYjea4nRbhYs5SqqncyIYFXGVTiSTx+SnRSqIh665q4lQIJ5EEdSm
AWH1qJAVYptykQLXJr0Dc3UMfye3NQs9HoEZIz5DnGXx2ptrHywPDBvKHC9MVuB2
UdP0FXA62YiCduOg3EtcN3NdaWPJQwoXfkzZZI02HUmgLFnwURF69NsxlaJzYryo
dWY5aUwC1Tdfuysc2F3asTQ6hgvuY3G2gfPsyqkkYQpHRNDYziUMUVMViuTlzls6
FCXqxSyhYgtFE9BRHMwrum3izBBg58j8ByNUBngRU8AQx2TXD/z/P8Nt+r7Zluyq
Qqs32Jvm7wufO39ifYJB/0sDGfP3+Mx/3oTQqAFRiblCcP09HMvAHitoDDG/GHFP
oFaUHwj6XF2vo2ZblBRmwI75Tz/2BKl0XscKbresawGvD1eSJPsA4LeQlTnNPDJM
Cu1kLV9lAt7JRd1vh3JbkKehvZg73w2Zodsb/LrbO0UfywQiA5Iy4vHFLALtUDrD
+Yx4Fr12Nr/f9gPpd6S91XYvplt6sV50kYPd3bq70tu4ydDwvRz2UcRsgQoWU7LU
5t8vHy2ICtZz11G0hhbFhprMhw2zBLFqchwpeOl1CdU7kZFJBUIfn67jw3YyMppM
Frm7Hl0n+EEm/jyRsefJhRx+ziW/JqDo4epOHIYjC51eFnOUTI4H0SIPQZPbqScK
8MKgUvNn5I/wow38FAvKlnvn2DHtRXrlClyktfBv/KSeGxOwaSQHb4KscoPgxd3W
pQ/wEjCdmwe6RGbhkvVpi0BKCGLzRZRy1++anDw7nXPOA2IsPJNKzqx5WJ/MTpfd
635q1xTbQBJ4rtIsxkL9LxxuC6JlzL7T0c1pXEPjdtRAsuH8taWUaIg9eazTbNwm
mqBecer8MypNhx9BLYcxdXpDJpfRtlmb8g/AW9KuIPmlsAnyZQhmUZ7OSc9taJ7/
/LPH/cJ9hr7XAtbqGe1Lp5zQoZ9Hfc6yQdLQ18E7VNrlD/PDC+z1SSMyFnToJbtm
tf7h8QIY/uQpBep0h9rK31c4zNg18Ra/38em1LsPmm09NtVdNw4zHr1/Yx8QdNBF
LsWKmIeVIb4UEyWB2laFEgpdsGmdwGZu+aMpM//rl9oq+cqZZCd2L+tDt2YLM3ty
aTqRkWvM61F8VxRx+lg1LE6tqzQDAFgu2R4OB5AtjSaEtN5HZ3cT9AtuFGR8zMwW
aDXLSyLJGIxBHQ2v6Fxy/6N+JZI75C74oNZ5L/KvjvzJxOXvPTKFCnVJPkqYiLqP
5udtvt2EyvuiyYKpDXAw4Kjd0/g2TjxCrADIIo0WAmKmBBEOX5O8ohSpGP3HYU7j
rC78B8dzeezaJs+jiujCaSaXcw/zzb7/KxOX3Y7vy78ztllSc1SCtZx1UGMXQK4I
kE9cJOQjUHbkwR7G+Ki0H08CveOYrt3UcF04dx7OIuCl7ZEI0kp22ciczsxnk7lF
OsK83yDPzmPeK4BEUhxf9gxkWyHvzjGFIN5lGWK6WNuGGHGdYqStagf08mnv7dt3
0TcM1r/pre/lft2PIzMrJ8vX+PbMLLW+6B4DA1aNdoXwgCmjZX4qovg4OBvVkJi4
CWbcchL9XoaGSylANu9oPSsH2Cx7sijGhbuz1EAUp+v0T+tZ/edG2GM+N/R7zyEU
8/0TNEQPDwq1rMDnlOeq5KYX2YkDDFifSo3l0YRRgVms54puTsA9WuuqTBKKN+fQ
0ZeQEns4wV8VZLIoqOHtijfzdpBGYWG8u5r347OYT93y8MJqB8OD7cbGUt9EudgD
1B6/QONhIb2Nr3fseAAN46vZyFikONgqEjpXapsLvUKqzOjFJxB47wm+vk1qiSpU
kaHvSVkQABR/nQ9QLlYA0CbQzJrQHThztYv4XAmFNZWKWO5qG3qh4y6xJVKWca1Z
C+G41zPD9jsfrvhNe1z+zeIma5arsYJYneGx9Op8nQIv9HI01EI5yuU3wmcU2Buz
zAve0T1gZTV+YOWQSqN2eB8x2EbwGzvhLL/gHdvC2+wbcpahOahVpCy1tPukSfOd
JnGAzkeqHV9JdIvDEUgrhOtPfebZvg1OYSVjGHssHwp+otGO9qWrbToEKzvLOeA9
iLc+0vUf3Lje6uAwWxywG4HcJ2nb7ZCkZRiWjWNBzkBpVaPIW1sa4L2UCpvejOvw
VDHp/RlDGuKoxSR3gKGwigXpXJSi1D0/yNh+idhiRGH+uEmJWoN4hWU6g8gI1a/D
phF+8lp/answPcmoyGvukY/jxaFpz1VW83xjFGB70Sc51AMDmJ2sDRw7JdfZyNa+
RJwDx1V3nHVI1+Bck27UAv+OiX3pD0/zN64BZ8qN8Rovhs5U3NGG/E9RZCyJNDVU
PwQ16PDb57X7KdFig/upCDXz+fryI0ioUqIM3U3nfTiM/TpRwNrZxl11venczOkH
RFxLUUpdBCVoxOOXTz+Hb9wL/Z2htYz7Ov1pXUR2p5+nmnH29WQ+aAIPVBJ/IFrI
bxQ2G2KWdwEXpmpm8XfDsMo6xto9uluGwvVYsk7eNnjcdMc1vrZLHQ/aTbYDHK7N
0v7khKKenRA/BIkDXtfJjwkQnv3ERJzA1NpDUDjuLSuCbtHOcJlK8XONsg/acpXT
fapxadUPSdSrK585lD2OjV0A1vbFYxjybRv/HQoIy7nYV+Oo+DOt0jxqaQpJvwtv
kc1C6XMTlfkRrfCQJweEZjTUA+qqu3YqRPOTGFBOOFA0GNE2NENwLuDac8sSLdBt
FhFmvp5loSFgK9oIwh+HnoCscPV7GCJrna17CWEL8Hg=
`pragma protect end_protected
