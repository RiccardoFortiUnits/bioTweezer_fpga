`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
E6v2djzMiEFAzT9rlg2Fs5b7UZu53Xl9rOdjPhF0KqrW2sDnTEPd2ddrFyONr/O8
ajaVT/uKD6RfWiUpOrid6wkHNAqgER8Wvnqm4m4VQps4VZs85jmpY7/pjHHdptoh
zeCPZHbuji6mmj8w7r1rgU0kXqbwPZFN12IOxOoWMVk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26016)
az2xVu3vv+qTEGZMjf6t8nKcOEV442yU3mPpVqdYD9bpmeB/Y1K7d66I4O/8JXWC
hHRE9L37hnCm+hxEo6mlpHa6WkjNKqV6seug1o65xd/CVWu1jAFRrcvroODpxwgb
5OL0DuU2bBBEAu1BsHi8hksm9nrF+mP6sXtxCGtxuz45j/e75FMLiohUpASxqTRq
GrgV9QbwWTvxda/G8ImxnIPnKq3SwxVyHSaFmgzpr4RQwNPOxGIbDRCsiLAkmqNa
Ml9qA78F8ymHaSfSOVjpH9icQqcpUoc+A0QdKLh3/TJgzMYT3rtOGt5fGMR9GDcm
vWtjbf6qsGxJ/og8ev4UfvTH3Og+eskOp97j9sGviggHeLaSbf2unOCycHkLT+UR
FIL/GypP4dLiROI2RByCH8MI8frTwiwBYBQP7Mm76cf+UDDNYb/G2izQDOq79IBz
v8jgRqy8C2e/02zB6Yr7L0HvknSGyuj5AAI+YdRMttnQc99Zrkw518on7bXflkqY
3v/Roq2OO7TcH2KvHXswfqMteydsuQTs0i01zNBZVX5Y/nPM8naMouiBptikd0Ta
SehnYreSGbLS38LUpEvgZ3Lc4r/TQYbEPJ9wFDHJ5dXHusXNPPQvWSARaezfE588
V456kK41kVNQdKZQnJaXpWbgWheF+tu4Zr1hUg+OvtZ34Pm4OU9Mr0zn9OiV0e9k
hpL571WLBOW6hp74RRmGFPs01Ooca+8PgYQ5xeZG90fd8q+m6a5/S9v8nRFRJrnQ
X91vgb09Ecy4/sfVM2XasNUzPMzeRvr6gf4k+KtUXVTaGZex/uXWZmuweaL9wP2Z
iZWGbgXmdXhliSha2zZxWbcalRwmU7LDP0a1V/q69UwtZbBQFzILVNRrbYkzsUSA
pfKfMB7QIczZHbTXhLnIjCTWgE4UO/25XE375aooXa3M9V30DTT2iJsxKqKt+ul2
gOhaZbvKmR40UaH8502DE33OswHOsV81byEIPHL1nvLYsQ+C+fk0vRbcOHoSXUvm
+OYI0u9ncRrTwjrkWCc76bXJFA2EZ89w/A6QS/qSN1+SvzykpI82ZBJsAm4ZRuzK
FIgREOFISdB1EpE5QXIS2E/J1kHDqc7UwKe6AU1k/LfRZByLz87w6g+QZTejO1Lk
uO3TrdDvM+5+NHeVn/hNDz4QXneQ82bKun70bcA6hGFwq7amyBKYFT64fkfo+38C
05QYwTtAvivi1vo+8D2as61fwmLPO0FiyP/qcRobPJ6sf1lHY7jN4BU09RTOEpuL
LdiOwVUW0TcM/qZebKnFZADZhc98/XlATtE4aIRCHWe00B0osrpzV50Bri61+dPm
+NG7yoxDhQskzpEnlFsA7p6uRGgZb39HSqaP0X2jhAaNcovxdUw+42OzK7ANV4zT
xmfr0p17nMMDuHa4dgPtnGo3nPmUwH/SwQK4vFIm7XxstNK1RoU9MNmx1KbXHmIC
ntCHaHZ58P4oRm103x/ciNmnTB+Y9zKUSj4ng/I52nxn3IvbqUXxZgr/wNvrHz+6
LBWVZOP7UVFUY52neav3CxC9w5SA0EgupqHZUwSDPkIb2niBTU/0Em5rGyPwzQJ/
XzKMr1FZD8VxeuPKCnSHnfOZuxD2AqbrihX2vW832GlDrTKurkBqegIxzyS/ZNuq
jkI/RARj1kI8FT09R0QlQPX38xWQ+e1LbB0TLEnSuLmCfkQ2JFoVCTbYVZWWDhqf
+Mwdr5AWrU2Q9bHkz8GX6oX/AVbFIsopH0bIHBQRU6OZHsuRzwyAieAUbb1QzdNe
1ORu2LqxR2G7Ta7lifQvA26JV/zvoa2Zj+/WC6X4zLXzM3wCSDTPILTVngSHAINx
/KXj4FMawGb63rUqL46sesAVCHmXa8qK1WNileyoY+MAWfmy2mYtQbuYdiOYpmie
s88viJUxSaNgdD+oYSlX3LosFkyp9PrjnRFKI8Kxu//z6Jkb7FI9fjxjCna+6pgL
u9aFg4y5ixGOcDCcOsVfW7vjx/2gMGG59gc78IC04jFCnLaf8cUp0KJQTPDRHUbL
Isqvbz9j7qzJJp2VOmO/ClrdsKhuRDlScDLZTx8jSVNqSJZfJX641RYgzG2nkavt
Hb5UTDDUsMVzqjf9WZxqI15FAgqBguOAyNmpuFwL9/o2DdzkWhNFTn2uXoLJllAC
Az5FcabWYDobhGmHIQMvqTnD8SACuqRrBmzsldvcMQ2Tt6rwXIqqauVLpSfLfLvf
rem0C7E1VLeh3CZfJUCMoPZm6grHNlvwMxWwPz9mYxW+AZ1LYXbHSQ5NnQMelZfT
XuKEV3xJhodwtN8wAl6+jHCRmyXwZEw8actOgSkZS6aLbS7MznXOfX5HcZpcx+YZ
MVUpYIkh91WYWSJ7z9koQLnlat1uB9xzSB5hGY3taI+gybTjH/zHstpleBYYMs6T
OjsD/gfJQD2dUvwPyQ7SwKTgvVSc7Z4iFk0u69753nbTqFDictB5DudaHjxbhLrp
D/uNBLC2DZZ87n78ch7l0tI97khY49hVFb66aszAZouPdVoRJ0bYuJFYLx8q56Lp
uvwTtsDBAAwpua8fUkzSRh3iIYL3FZbDVJBa/8Zk11rO0aOLV+XMmgOuVZXjRQQI
ocDeX/2Ttgp97vL/gpoE4rscma/Qf+hVYa6O/Z6kIZ8E32v9N6Oj3m6WfsW3GLxX
4ziLzcqFuV5YQs7JXmdqV5G0z8pNWGJQ4X9ChFyQflgKbuRLS8Dj1JFXRhDS58SK
65SB+Qrhp6WD1i7Ik/wyEMrFWo9baQ+mjzpQJgCQMB0pkcIyTI+uzyyHNQ6EO/EA
KrJBgv10apJvhLrMzb0g6XCtVqe522JegrWFSTzYymEH02iMdQzJLiPe7Nwg14Um
kZRNboXyps/FitAHkGnDFOIsaLEr2tg2BK5bnu1bLSbPJ2jjGJeyr+42vftA6CLk
69hYbkdoTeQHDPGhxfrSPWtTvkZG9B0lDslgvJc88naB4c0F3aw6QZ9XI4JXGtM1
7F8jjxpB+ac/7S6DPAekl5HTFc25JcE7S/ZQzhqOrqHgndmIMf5dBMsG3/FXBznt
dUuzrTS74pLnhXnMfkcGFejcxuyI9Aa9HjVhgjdn18581m2+723gQ/yK2i8G4PMW
gJ6OT2uKk2mx0CI6dg5A3d1BNjRVvCTTG6wXyhgkd7TO5RcIqIWCYNLi6UZ3tm/R
czv8vn0x9Dpukh6fc4wxJHJfkJAThwexYDUjYjGVTXBZAMslo54srrP5lJYCOi8h
aCoC70EC+2NXifh/CryOxkDzA2/Ku+5uQVl1inL2VE13l053oxuRG2/wEpeaMV1f
oTCOw/zPzZ99z+bbZdx2yqrHnO/J76Ym2oQTFNMcxBUOaG1jMh9+trYm5nWLoGPC
GSuY4Vb5gmSNfDn+JT5WJMvPRfTGMXzjo2UlvN2QrrTtn9a9aNOCVnpOXS04qjjb
4BqR/CoMmhSdRK4Yk0o5NTZqpD9GV5BqlZ5JQsoqHlAYf/TsZX+kLAbGyw9YMUOK
Zidk4BSFFTW78/bFN50Hv2YfYynxC1soVEP7yeP/l0vqwTCTOziE2vTmwvS3O2Vo
cm6lI6M5WG9er/xoee9dhvKlw7nsPoB6v5kyQJtSnFdNwIqZmasOV4gZiZ+vU/zs
UzJ2I4kzbnpyjR14IMt9s8dglb9Rgc/DbiGoSRRbGc3QeMutUQfzmPSIvXHYVaRc
xDCroboP65fYqj/qFR8jhz4axDNPcd/A9sTHAKEZyYzNiy0ru06itEc7fH6UpKjy
KXYRNeP0tzAK8XpvTvVTWoNO0ybLJVAG76TenJb8aexp9Mg4rVP21DvLPq2Th3lt
7VjfPU7F4XWHgrGbvqocK3qRYYOre6N5SSR10H4omFlNZWaQB7PeFWbqeh7cIYFV
6e6ojnE+2AHv2BThEmYnSALb+IPtCK84PaPyYWkpaVyw51XYlT40QOfiKsbqOZWf
4H/hYcEYe2m/E4zqC+t3NyEExifFNOD0aE/CtOd5DL5tbnlwv6fE4T51x2CbBHjj
SQ2+mnvKNaV37hagGPN3hA3xZtCmwUYhWKEDFeDt8QUAaXegg+8PMyJ4BzFN7Dth
iWrcIflJEVua4SROIxRWJSfDhjZKfgYgLAioSv3mPsyvQ85BtrNqL6Q8c6zuc3AL
/AL6AU0V9JMV6GcINWoidOKh2Lp5KLDrAcl2bx1Qj9zBxLYUyonYoQ7PvVEDeCxL
kvjLZxKNbEf0nEgAufst8s/H1Z9icIgytDNJYUGIEOCbdPXmyalO3XRnk38fFx/U
zjSbwsNhaRTQDS3hOExR0XjLejlShHPWg2EMlEun2no7uOpJvUwdAXyRHD1ePR0r
vr4ADaGZrLf9NsQE7pVzofJd0ZCLMox6cVajpF7J74nZX6tdy67+NhdIgFXUvyRY
3XrFxPNdz9xtTqqKg9Im/3A26gxQ4jWIQZ/EV0+QcFouqcd2A1UzMbObFYeskH+A
acmyDeclWPmGiQcD90ooOj+EgbDkVP3vp5AOFZrAF+TMWPrcChMJFiPLsZl/LtXs
1z5lRNPpQxdJL7uNygLsR1WhRaUQ8XSluW/+HAAZXz5jEW1vutAPDZkHNKSRvzQx
j7JwP/NxDCjhuSA50TScCFB+FpDo3Q4h7UJUkCeZQ+qQFlQDRTTf73lILGpsGBSw
+nFeXGn3U7B7PM1mO/dkqe0SgiNzwzo+X5fyjy6E8mh6InIb027L+TUXtG3Av1S8
LADUq7rBZhvi5cxYnu5TfM0wzHl2zK5d+4ZDk8hb3iIf+/q2KjzMPWhiUfGxw6tT
R1fAKZIDzHUFPuooWYinupU77H8EFb+XXbD4n0HVWfv+PKnE4K/9ITiEu1fjSA21
Hln0x720E2DABmCGB3v8Ay7O9GZ5cNo16FvkYrsZyVlqawX+8K9N3E36KlIve0ai
LTVoTwjHc/Qzhs2P4+dtxNqH00zzq4jgeUzc3+pj+dDwhjlCdWt+zBKxT5Vso0Gi
k6a4FVpLM1REUZjhdOEGQF8sNq/LLCN7vt+sJT6URUmqQpKkK1R3XTWoK+8jx1EL
BK3Nv5fduOdmTxfbqDX1gysWuNW9V2nKsrgJewQoQExwx5cS4q6fp0sWa5Mm9+Bk
or+T0nW8n9Zhd2bCb2Q4HO64G5DNRrijTeCTFGXj1lJI6nXXd4CLQEOb75yxTVQG
doKWCs0rKPPigFGFzRDTYNoclu4TXPHMhXYGRThdp6EZN95ofPVsaHC+/pseMzEd
EewxPfSYJZfDmavVVbvVcR4hUHObiK9SqJhQBnbJw+FVrJbhBvx5Qa5PZdPz1mmi
otrlKEpW5jJI/SrnJpYndi0Zdc9qlt2zkJCBPbQA6rZZOT+NmLvJZXJcyg4yjlaF
rW8k/EbBwZwmVU7XtUTwY/YiEiGTN3VfcUyDFXouEfgDEyv2GC3yroRbcp/oFdid
gM/YlfUjR56ZUasko1051skqhlo7caBH3ErsiyLiBH0YGkonwzWQvodhzht4JOb7
N1fMnMfh5+iSpnki5mos31zXIRFFLB/hC/gPHLrGuCG5n3qJIibTxK1ONdIRis4l
hF4SItIodLPtMtQ4XE4IuEJwcmnyFVodFDOUBSl564aThWck8Zp0fAhK2eept7mv
SEv3YYny5t+Mv/qfE8Sz6q9poUwH5tPRnF2mNAcOHbKRQk667BISo5OibE8b/FYN
/iCdYR43pKsTtt4cMvkhfPykrBuzt2cmNY53mu6YLdciM+9D/1q7lK9tLV27eHZr
6I6fcjZ7yqWkEITaS1eLpMhxfymjoxnxXpnf5UxbR23ITsjrBdLHln9C79+q5dYg
WH8spz9LhGpsZc1/LhAQ4bfouqimnxu11nSoOsOZwjjr6ypwL7gPAYYNql8OV5q2
Dy5lQsvxptJSyjXgpaCWxtSO32AJ3m5LqakQrRsPUqrY4iGvA1fl38CS2BoI/D5Q
uSmDSPTTzhTq/yUqFcsaQ6E8CwoergqiUxhUO0ZLc+mbuu/heYPB7i8Xe7sP2xtC
OLwYvET/ku8qTLkkuHA14pQQLk8nfCVQ3Ssa+JTmsQyVTkk1I+7S5KRU5uP1Jbjx
UD7FB1c3yQDA9bjuqPJ/WlFBOkcbxtPUlw0JTI7NCJ+rgVLeGPA2nUk6GldNayyw
CWtELgAoetp6bzNIxP3Uq/55qmNNlvDHiUKdI7JsGbA6F4wSdqTq5ugGweo0ZWNw
LLlsHXGmtgsWEkG4i5CCWyJFGFfkn8gFg2vMpxi+xNRXynFcq418LiHMrRClfamd
DQmGujpyjKKBd9jmVIqS6krQ0Jb0MZzHSf0hDV4iBjFZzGVRogp5KniKUTRn33h+
H/cgdq0RS9P3JrVt/r93Xkk2fjRxABN91DaNa6uQK26/p+HvuHojP/IKX1EHNpdA
Tqt3ALTvVL9kW5WqrwF+oLN071MAC3KeVw5fWmxQPHeQXUZScbKUHWmwUuWr/RF4
eDkDFvMnnUPqR3/dqbz4Y4qYn+ubuMgI2JJeUbi43LLQy9IYCiyBgLijrhHS0E4+
bU+5xJd9AdLekH6SRE19Iid+B440nl+PL87bxfAu+4bGG31OSOvYunGruR7kejmF
+Bgb9pyLp0Vv+P09oZI9Y41nSBqq7dDuErI9QdXKUsPhnJQQYrTHrcLbRgTeTf6e
ZnN5K/DgFASzLdztjtrHuH+i3TUtb9c8z6M5vja+gX5EbBJahZ2TC2ojSPk2c5wA
OjH0OQn7hqYDJuJEms/vCpHkdNpUs7xRv2usnkDcDTxdv7c2YKQMZMzZg2/iAZL3
hY/pv9K45OAk86DzlTUmNvqZIZkiR9JBNpubrhYwb7TlW68fh1r9x4XY0bSNGrlk
e9cFbZ0lfjGftO8pfeKhkVOxgzfNBHfYIbJOZDA51Ugz1hqurTJ9yUviIF4D0C7z
iyP1alpasNVlFThYQpxvFLLthB0vp63oTqSZXZI1e8l+K5WSYPIkSYIiQSHaEL/o
P9ILlQp4WXE/LgZWTbisvKi3QVWWc3VtY5XeVK3ZDpyKFUW6weITxkJbfSnAg/7d
jUY/U0aQkBlT1AeT01Olk6aLiY/OivRiPfIdlnSfRrgrniQvTVmqwBMqjZcbP01R
VzBv+MQh5rwWzaxcVyWyv+PmTaj/B60OYClo8AVzJnxZAIbM1Ws8UCklalG2QQ8v
J3pN7g16HLKKemSx+AZT++17So9d5U+qji9AyYxYfHCx6bb4Qek/t0Uyc84rfoCy
TRViOL//iejD2hyescdG+k4whuTwLnTVKUJLhlaDz7NffIR2C+dBbHBK3wiNphvf
lHx8nGmFkr+mslLEfBqiIayGYK9CJnp735YQByZMSDmr31fVxZvsIURXfhFa9EiQ
WDzpMICDBGscHl1l69S5KUu4JBVpt1FoJ+X0S64gH9psfN+a4ClnB9AtFoU2p2PL
R+73Qn2L6rXB0xmXUKXweDNQW+iym1AHjJqYu+MshDbd2pS/jmQGI/X+Hr58mWOG
fHGbfzCgNifcPXNftjLZ1+MWIp5jHN7TsjAxVPBX70nIcmhg9dxM3xt/5rzJ5ICC
A5bwp2RaS+CMvCWvQLChgwQmTZJTi9Dsh2vuqett3kG75EOwfNw3ah76lvgTl0iw
xvOWnQmDq4ZxAOHEtP8jHkQE4e7o9pfzKPdlIOQkry2SBf9uDAcO/ZokLGs8xQeT
3FdvLvUHZp10wxY/2pbOwd5yt3DTMO67h05dvkM4GVHr1VR9vpUvnIogTeA/C39R
Qvy5GMnyGElitZi1gNUtlPRtkEMTjQcXU++6n5v+ZVwVmFsEJ7eZsBzUVlIa6sp+
Z87fSLsXhkx/iupgvswuf6Scq0dGvlqhlh6KW1QBRMflCFmUfwTDFaCul2MJdzTc
Dqeh9iJf0s1pu0AbS4u623vfja+VyFZqyrdgUfpJdUPRaYEcjUARnDkAmywwPzUu
LKDEacgbd1+OUyrrm2XlKKVMsy4Lx/f68HyQaC1z9A3dannQQ+O8KrzgTwNpJ/PH
bHNj2gxrcT6fbZZ5SzEWuvmrTnDM4c4xKm4/l9mK3YitTAaNABQ6uq6khRLVv+mB
cIW0DzpPwA99tgPEAgydUTqjuvG+L72So/1Pt3CmOLgR/8y7LLoycBjMQdVO+GAn
+ShDJ1YTXqbW5P0vtpmIxaaYQAgTB1xQrpVCqsjmlknJN0wXr4436Ge8gks3W7R3
Kzh2Zu3lwbE43Zau8uEzqCXB+aKk8rrpNKe4+nmoViqthQcdb411pAjBtyRCfk6y
S9SNngwtmlwh/H8si/TnxZymihq/R71pAvyrrGOqYArZ+JHRuZkOnychtmF8EkSA
604nv8Q9nVnQj3rzxEftQwkjfOn8FKoa1/BZSdN2Q88PeHiyijJnt69emGAZCgke
CVIV7pcw8eClJmOJ1FjIdFjnEpKvfxMkgUwdno6Of0LdjCyREbiJ1eZeygOYijuf
za45lWc/YbWs2UbgZ9shfngsWsWBvAgh0bAzqs7urGpeYoLPcrvmiNpGKxfV/r7J
Pr3jj/0KyGVFE/Snss6uW94607C/RMi45Mu4TDuDC+PItG9GIT+Mmwg/kL8XX1sr
S6xfliX881JORRaT//XpIIWf2ShbmqwywIOLvgC6XnAe0XsMoHa8aF1yxHPHAIT6
U1fUefqsJQ0mW+nVsoS9+YZEc+DTRVGa596iHRtOoVYMkYZksOXk5hTEy9+hSXF9
U+ydPbDlu5HEswQ8OsRZ+ZpQ2FFUIQKAlz5VIamqfS872zNTohc9jA2Fb+rZp/vz
yjcKjWxgw58pUGQkZuo7oZ9W64BeQ/H/bXUYkdVjZAslb78YJdtc5kFoS+2NVX+L
bNTHW9AFYtOwYVvpzi0B7MLVBbNin+hfYVqEl8kz3nDjMYiGZXlr4cP0RiJIqAjg
GX/zEymm6AYqKp2Q9xBUK1dSQT5WdvF9qnAv2XMNWRTluXFtyQj+LHdPUj3v7FxU
8jJMz8KT3IP70pkf7QlrCeAoP5BmNYxcMsmI0DwNZ1xJnGAjH6EWWImOfWQK/2SU
qILuJSKHm9dPqpEQjmq+M4KJYXvg+j32mjpqcWQSqndAOfVA1ZXUfC7C3iqVskMN
E6k580PkPOLTfYLg87Nzz5qKa2FHukuAJWmoriHJKHuwPz6A5Bzpor00mj1s0bsj
XwKTylx8zKL9Q8g6lj61EKtvpBHDdfdH+lyvFui39ypKR266/d5+6908aLaihxWK
x6JI2bVqGZ9I/HvReVZXFEljJRxjFB2vSn4/zJjoVlSm9D/dinHUZsA54Exh5d86
r93FETZNTG0wOfJYZRFOiVmsV8ir/MmB+acCQiWXgE95hY7cg0MkouJEuTWy7+hL
pszVfnU2XxAXjxLJCI18fR9YDqCeyKTjcbqGPyg/Mfvdh2gB4lfeOJY+6FiCA0LF
TfdFVbwpzvCUvYIPsEYc7LWTM1T4Fu7SkUFt3OhGNhlcKv6jhI89ZfKlSYsTc5Rd
uN2gjddeqbRJpY2rQMJBL9Rwq84+ajE4AqXrwmZlFdi3ggoPduLJQCWtrnQKyZyt
mUKfVmJaYyfdyPt75zFeyt6knNRd2HwaFuGp5uoQTPMZIU0tlETwC61KuD3+voGL
HjUeweoOtzVOOERca4j6udxO6iJpPwMUVt/6GpF54gzXNugqd/GFjZ2Mr8yL6RKc
Ygt4S3hGeViFw3F62pZNtsoSM0nvVwkXuSIOl70g5XXk/u3yfkFG2nAgHiWQ3CEZ
vBRDmBP4sD1cILAKFVUsdY+v76SzTGG+f2iwaU+8V027J7crEx7Dmw2/kMRLbb6h
Cz3cLk8ozH5W65euOEKcLUozAjLf4/JL0jEwRvp3s969U+h15O5loz+BIWfRL7jb
ljCdThXtbd8Gbkv7hddgCUjUv4bzFVrpRTxqBb7GCtdTb24AqNd2xJqUr4tQMWaE
HTUN7rgh4+X9uYXVXobaWXHBGDGXbv4akXpj2Zlt4sJt5xwCFYGTqLTdF7MTUrk5
idXQegGJSlSzStONVRxIwBGBEnlcyHGUF6Yawm1ApxIjwv2aZDukgkkQfbXYLz4a
uw7EbMM+95tQch6+nFmI1tZkvCVIMZzNmUnMf8JnSFnOZCoUd2AFYUTIXLBCIzzn
wUQSxsXlzouRcNTqDQ1bxly2GNyMaEtkLqnBY35T44t2sfSiNP5sxOIA+XTcfyK9
DeDZJi+t69f0xGXcCzCzf+ytqapN/VgvomOGILzLoj+c0Sj95WVSdO44//PdAKWQ
TmIzQR89uo77PMh3yejQRko5a/eaASGgb14HV7rgRrKlvt7sciiTj4v7FtVORptK
qG+pw42mrOrkAnjX7slRQTlCimH8Cj8OtrdMgAPowtkS15Zf9Rf/ojfE3Nm0fCHL
oGkjiFYKl4RIHwt0u15jaB93DCwg1SUfzZus36pDhkDZ1YtENPUN9hYvEoCQ2kE2
euo4/KtApZ4PGEkxPe02tL1p7OyWaKmwCRro3YdXzwQn5C44TpRmzqZml6AyDsSS
tChZRxiXHG59m7aeMs3dW/QKOCxLIqUcrmEKrDLXpB3euUNBC7JwLVBwpE5gSGhb
Lj0FXccZyeJvW1XWjGqyu8+lh45cIN0wpugZDpx1/EwESOHnk0LUS0assWHWFcXu
KJcbvoiKF+hkawRKqIYn+ydOEfEDjlzYinO2vT4T132Y4PD9E17QLniYaoACXiX4
Z8JiIr50+PCsYAi3vqK++NSXbQZT2VmiVwG65CMhhciICE3l8wXovyXAlKIf4tr6
xSW/A4Hx3f5dVLmeJcXBLDgAgls2qo1GJRtuveRU9IIiiK0FG1qpoOI78/T8Rtzv
ZscGOW9Ntm5muMK9zMCC5YZAYIuXIe14F3xGnpSW/EvfSiE7ui2mUU1O73Z6FCPt
1WymNjEL1H4DcKQBjUlxXQsKEm4INU/TITwQdeIJMERfIw/t+8mk3Vf0kUWwMEot
+bjdJqRWW0KcDYShKwfAaaPJ0I5GqB8SeDLB6NA3anHM1iO8qsu7jYKPypBdUM6o
OVYSq5U9a3JEv+nqRfYS1G74Vf6Csq4NmvHan0GSGaZydyDyT9/0iKHwnK2KDk5q
D7CgcCADeLaJ28cqd2+iI5xdwGBY6AxOT78riPp/dALRBxtoU30mKtQTz8aAD7bm
VrKCKJb9683wIvbMuXDKENOqLBXRTcHU0PIWzYumMlrTF0A8z+nWjSDqOgh/l5bB
9By0Ue9VD63teXzZAirXoN0bM70ddL/4yOkM9mOpVDn7RDalh1gg6QX/yHwuW3RE
Stb5q54f/5dwWv8GGWQ+y5B1v53RgM4ePoaREZvVW7vYe0kwJ1HWQ5ud64afKd1D
14od3IYlJAqtlawNXynEprsy6f2QigVB26C1HVCRjPtRcsSZTHJrsx1WLMySu2TF
INw15uDT9YM6q+e484iLuxX80Aioc7IFg4BXftewxgIKEphuuIsR3IiDIr9CacHn
7oXtdL4FGFI9kRorD7vyt8UDTX/pk98wUBlSSR8/GvrKeuFKb2pXcz0nvdKQL88T
zMI0U9zWLDat6TFnniw76OFHDH8soPAPt1j4P2eCkgrBMYo0oxfwnkWrCG3GRz6U
u5TP6LbTKDLIW1ZroTivRx2ouyD4ewohNz0qJzbGWSQU17HLXtRLkk9uITg1qClr
UzltULfGIA28Dtau7Q/GbWghqh10vjf1R3Z4cdPJqZ7zF4SDaWKq2xfiCAPgUxis
RaEZX10bX/LSPBrJSy/2l+1rn6m7xw2OqgxckWnqgBpWpuDTLa2IvkRRSt5rFSuA
/CKuHTOQkhiKlAb4+TIjEsrgyPvKNnOz3nxnBxDZhdPy8YpOnRIO0jH9s+3ZFZrP
A2h/C/0AS/YJJf3vYAtx1HUY2TEPjLqn9TCPQ9DWdetEvGerqqaxE9Nz+enufBU5
9HB8hdiIFgpMu9w8YKfynYa3CCYALI6HJiGTHW8HcB2h5bQKDZoty/KpMJY9MXqM
N3XfYoxJzKfXX3vNVZBBo3ZeT0xUG3XV4WrTz6wT3VXlPJwwPppR5F6vpkHUgcPO
a48Ngbz7M6n4/H9FlS4rHnfrLN8iU57aMmJNpR/Z2RgyJq0bWyL1yK8LyebDBc6q
kfVuQGzOB/BT4sEOLjXFyAQWZDN/V8mbbswyBljehIqlM7KO64fAUE8o7GQIRUWU
hyEnu6w8xCJFf1Lm7hVPgUHtE7ChI6m3MTtKHUG9UAcxh16fg9lNc3kFtBPdG/kV
pqMia+vKK5sQ8OLBeYQ9AKz9KZ0GLoB6lBxiu9VNReXKLKaz1QzD+cf408zeUXB+
JkyaYF7bwT9ZrR2fPtlMvo7fIDHP1WY6nuSNLvaZwuwsaurj9Qr93tqAAuvta5IA
k+w2R8v90JUoiHM5XDfq0bnnk4hXbbTPv8npXEeOS+1KEqXnBZVA021nTQRDvpma
kcZzz4hQovkxnSjQa7pbSLF2EspuBuoF4Ssjte9XYZxnbvJqcULfb8X6xqXtlutu
1FP6vk6jWJTq60o+ltKg1YAt8SJUE4h05zFPSWZClBhrlB8ktWvUL0g+3v0oNyu6
puXHRxqUXlkOhBbXZ010SoEzRnw42vEwFmMQ/j7xvrwUfSQ/RG1BNzQxyh+iO1VZ
X/zLzWLX4PA12RvHceahz1wskdY7tEs2VsLw7kn9Hzpj1sa0cSW+/5Cc/JGzb8/2
Jm0dg31c8QWXfUc+Rr/eMTtqPpgJTAIm4rA7U1JIdpUVoJX5JBcmOvVBXKqL81N0
e4izGz29Xn5wTAogPgRD0ndZZF4R8vKAYKNnItIKqSMsHWaTdxodqliDynAsiDsQ
hPAkasLgmZy0TCT4/1o0ed+QZOfvav/i4swodmLcDI+3h+ZMCLcmr79cOr0vZQ4U
AJ5FAzFUsyQqTlBoDvCRhYNyv+1xDejSXwK5K2mnYm9rJpPOZnmXse8iE2Zn3RpM
Xqm4se7LcKKPiVBtat4xHidDsOZ0O2L0b2OenqciWyD0ZgsJWxC/9uoZfke23Agj
ODh6SjSV7YLbpMmUynE4qqJoHrwy8AyY2CaNQxOPOSc1AbKRJ4TFgvFrcUJu7NTU
qz7qaomI16GcoRiP1hgowg35Acz8YxlxGYARqs9vWEuY2FnbqJxf/BQAdrHcICK7
XItw4GF1R5yv1k5M5RsNR8CrPAvaNW65Js+j0r9LdY5vi4itvj1aPouJIQL4Nh1d
M/qNv2rcx9/Xl5JMbzC9SEkvP32pLQtU41xe5MHmGKRH6dl0WBegbxNNpdAf43kS
TwSYiJ1D6D87UTB5IF3t1/k44qLurW91sg2+H8g0fHOE+NS0h7QnfDxf9cC48xQN
e2wPyenBEVOrVdQvxAHW9uefWY0tdW0OMBSZKSnzX+hKfJ6TiRSfjDF1z7oTWjRn
KIANrxge3ywIk7/pxpPTpn9uLTtuJo0iJmK+FG81XPlkRD2/ng3uqiRzfajpGI04
Zmy11BJRaBAiETLpbK5zwJ7G0cs3MYuIrvsJUjLupJ5v+9fwlXn++1/dGxa+2fxh
qaFaWsnmEa47/8Zv76iUqMghdm4MkbPGcq8lQCE5cYLuqPpbx1n0cd29J1Vc9nEk
KCGQVB4A7Mcz/wS6VsPT/Ie9Ym6uVtb97dLouRSBu77NGnXRKaucFs/73PDk4PCG
/Rq7Pp5DkGZCNW5jXjYG6wxP7K2pjCkYTBm9/7tNvn9XiBAwyyyaFICVZXfnAG21
wPcwJ9qKPtdpi11Gao45vAi99laT60KCeb04mtqIZNQg0qoIuUvCpPJ0jdtJqP46
qYmg0Kp9V/Ru9PK7QOi26M18fEK+2OxugeRQag3u0oxg1K+95fwzDtOID/4BtoYC
P99GmNqPXdr6g2vMZouRpe6SoHRW/CiCFGgaWuV8hTlyNhbTM3Vcp0+Z/IPU43hI
8WkkRiZXzo4rDTZ/nWG1uWFNgMVha5B13hH9yERxDAYLC18i78E2vCNxXU0whcFK
dDaTfPI6xw7LTL1HDeI+D1uy6n+uu8/G+bQybd/vkvJEsdn0T01n8EpKydpZGVI8
tjOhai8SEGHzBIaax/atlAddEPLUxEOssCtFp+eP4ik94BmJzy+fDEedAVFMP3QL
P3m2kPrygZoYTVPhUI+es0kLtu3t5lOkM7LngT5CN/f4h+F7nQvgR6krc0Zzy/v/
SgBou9FpI6WhcCiGS4OmjmGMlky590NYIGpcrWw1qUg6uPN3luUzK8NzeQcoIPor
V81MamNsMqkknFllD2+CaBxCMNJ0w1v/o1T0KC+4B4cNKM0uCDm7sdSYHdJUBlVK
G/F0vR8idDg4cUrJ1Ps0ofU+guUXIOAJW0lIfWb4Uuo7f9OyLB4EUZHyasC779dW
F5LTNm++6BWtsyofFrPZ6QfV62lZd57Wb0d5ruwqG6uXG5dODn0jmcg/p8GEz04z
3xmcOwtlB3qV9MrMFNOh3uql79MccwxQVMpzOS3VDu1wDc3OWu+3Rc8BOg49exqy
vTwu+6y3sSjBQMcuale9zZKSpqqtL2sXjFpvD0zIbi8m7osx962oR9uhCZLFZHsU
jm8hUSqY8wJ4/igoK/qvCqXgD0fmHRk7+WB1ePOLSgqbXnhK4zDhDrQYQTooDuqe
MnNYH/BR3BJ75xuCSc3QSG8FH0blKfKuHx/5Ev7rJuM5ctSn16aCDadXXaTohBPy
bC/Tr7YJiX+sLPYFa//0po3uFidro9EF7DgTCmkAZifIvPvIphwgdgeFvgOjCaq2
t7FuOCigCS4y5qi4Dw3z4gZHpbB1n93v4Go4OK+R9sDPaSp2Fmzc2PI2FSkD+36Y
8HDZ4gXFcOUvvqLulMXPjdF7ZrX3L3Rs3FqELxsJXjZKDNEEil+2UUQLE4NGzwGG
xZFjCBawHqwR8lda8YoNo5AL9hpxo2lXw2Tup8es5Ls9S73avhOS5SCiQkpPZKDX
enDaA2eo+IfshNqxhNLRsm5raY2qKjfyfI1uASIMFm7cOJJ9ny7XTbWKMogvhJBK
B0FzZ7Qj4Kh47mXFZ2n8iDaA7Wdhu/ctAEWnzqS/RlcrYi3o8g25X+TQD2tcW5iO
tDusL+Z3SClxpNZbNCjfFlM+fX5uvJEcWku6HjeppDH5b/qz5l0vIHDVsFJdETCs
3wfWN6EbIwfCNt6sy683+8qzsqVxdI4cELwLFPq03rBC0zBiF1ptYlFhAKDdXGml
VutBB7+VyLFyEDI2ALp38HOYH09VObRQU0XQwM03hytHRX6PaNBu3DMU30fVJVjB
UpJJhpYrowcCexHHsaVKHwI8LGoQK7uCFiIoCdjtBJZz9HHCUfHuv3E7hdkhcZvm
Gs9FBdouIVfl+EVx69lI0r6Wdr6yhlZ4SAbgNWYs7ku/yk4eZxc7WmvqWt+bdVz7
68DoZeCBr45aZfU+xb4maTop9JtBnGrmjdX1p7E4ToBbmc7s9r8GCm1BBElxEpy5
HcIPF+eXaqJN8YBsnEVEJzPDNKClGorZ0MtzYuOBahhIMicC1b9JebX4BseMMZeQ
rbxWAXXWypWGoObEZI0L8C308mpO87dKgGNsb9jCLXblJsPrfjbQUtfB018e5W2B
4VzPvUqrQoX20tkIdL2xEzM98d9lYe/eNvLoU4CBQS3Ff3ylV8Q9rZhD6Gy5S0eG
wmKgq/H5kLr9CLTT7LaFLLmYxSr8HbyNop/wsNSjd6HOdLGnC0+s/TUvY2GUb/YD
1vZ9garICutzjQ8vJbr+FATEtVnvenawHOkO6LoUjK5Xtvd2Vr9ny8pD3/p17wTC
ZV4Mp8YtD6vaTT38JIjhi/MTgHBusNV4edPhANmPUOHoTlQSlgYicdJIlcNQ1K9L
n+IDhgRNDQFRldsL144foqxoN924Wnob5glu4UEM68G3uaeXWAlv0Wxq8Mlx0o2l
BhiOi39KQZQuPJhGj9gfKO/SxmjtVAOsgXToVnLWbULvtbasboF7ZHfNSCPvb/hT
op/PF2UP0KkFFcU6IxDkEFMo0qUkOMMTv9tNJD0zhPXXtKgilCuUthm3Tu5bVCjK
HcnAeR4zqlh62CDNG+VQTalMTiMhuayHgBi8qqWRKcZ6ef/o1IMMZpRVKZkbFBOi
2j9erzbUWyeBTEcrv8CvWEmGAQDXyWXalbh8pXTjM5YEMLF7PGxmB+Fsc1N1orEo
4iVh1G9/GXI0f32R0/aA3+HPWBqVF+HsLElJXGZz7YlCEvL8I3RfqjyyCnVB+K8G
eBt3RM9Yt/cVG8A1WvnvecIhtjJqUV3ONTaUfOxlAYPwKK/KlGdzELrN792T1SJL
ZZ6Ii1e3S7B8inhZb8UigVg55X+80N8WoKVOQZmjZhqPdbblnhXjW+pgKpYAP2wF
+8H4x+W8zvMTghUFlIVUPCuvT78CX01kykhHBqyFRO6KglMfHrb/J/Xpf1SchHY9
aQeBbNuwz2uPQDb+c5uT689S6zKGVvJyATs5ToFEABGT9lgzsHucMeh926ILuwJ5
anm+jzEFLtd3K05GuIt4cVXhPNi2JrzW+FpRynqnsLzpWiZXzwq5X+IhCCtb900I
tsqhbKsPfMu8o6UD4pAdj7Y6h+rdY2gU6co2N+xcyYOdiamYwMmk6DwkyXB30z2r
USRKXogJYOENMDT+k288h7WiVYOzaTT3RcAy5C+AQUqG11zvg61dUT3TdlP2YWpz
Zswat4/iTC2vX5O/7NZ6H3AKMH5Ri5XzpD/kGxHboGngc3cN/i3mC9OatrsPnmpa
y6/54+bzh2gPjGvWscYMVIy8M2JYJRnlUR9uxX24g7Q37rxy5h+I3rhfePOsZl1m
t8CMpBZrXznQUqe4Nm4d1bvDkm44c30URr/TCcyCdvciuHCRCIRfJvFqg6NCVusC
xkEJlBHW83TP9+OzUV4LLgcdilE72fUhpD4zMc9Y/0tuzoBRJmRYyME8haSJbW9j
Wup0YEkK1fdCSqIRQKf/HgVDiGau09ow1AOAYodYHUAPjHmaAHz+XmLTE7KJNhCd
sJY8AhzqcPe31BQ1duTTNopC1gLK6SrIL69fiv5Tt2BpqA1ae9ir4UIK8vdEyg+9
W76XqP8xokU5EcJm0KY8/L5pstfyJrLYH4rhl6AsTo7ORiO04CUkGFhdLIouEidf
hTgH7PAnKRFyqWW5Ma3IczGHi13Q7P7btXMq8ocRUMYvs6cLxvxzN609DSZPIWqi
ldr9VFrnoqohBDJp/7owud3Suz11QwBxzCZS3tL25w+7KQKJdkyUT3d5p9HpENO1
9WJEYQdE0BOqwdPQEnFJOvCzSr9WHLmOxn404CoPQAutHhPq2pAeBGdUr15rGHul
pkiNfZscYlmSwCs8FX9PuFy3BUmjQTAAyJ7VICE7QyYWgV82k8v06T1zImpwrzPu
pyFuP6bb355rl4XjWUeev9py6BX1gE8n0OvQFkVMm4eRuT9cLol9S5jXBFcE9Z1h
wEsqbyC3LAy4OGO6ur/yJhPjqWvARnXc5XfXPSYsAULfI4phKFSN9L+GyKj8KrMh
IPEY6A1VLK18WywqlZSvFmH1xze42+Xh+mPcjpohdvRMaNz9e9PkQo4ZjgAeC6Sc
egAxcONZ+9xhWemzm/sxfeFzu6Iow9MPg89V63Rf4A0A1EqdA1BztZyNEu1SEQQU
OaWSmDRurMXmSdDup2fgKyoIL9+CZ/+COiUKWWP86UjGhh7XPLtw+3PB2CwVu0YP
CLeP1eDgC//amH3OpVbpi3rPclEWKmQEjQ5hYxNq7hcBX0i6HpgBs047iyD1y1AC
zmBfxwOPL9ye9VrqOmRVnaxdynT+YBmg20I/fC4nnV2q22xrgq4sJPPT+77P26EE
fic0ax6jBw+DEASPJrx51A622fc2YUr0gK6ZDkxRLNF281q+E8tfXVapkoIQZpdL
5lpKfh3k515w/5cq+FZ/muFG9ooDIad/zlUfahdW+WWzybEUlzLnXNnanEEzqOor
AaDL/LaXCKM8IXjvFz28u1L5B5RbbZsNqMt55DTHergVj+4G5mpNGK3dUhc1nlB2
sviKrMYZRX1TLj7BjvKG8naNQr4LkX0Q105a9my3vCwz6292rPxAm8ZfWwFRcRId
AZvcyhGcd69PpP/hRn8dwFzLxErfwVsooR46EXGPLuhxqq6WOFYRtBhXKf82EWR/
ddk1G0ft39W0+SPu7AMAS0moYnNNWrXAHwjhnJaTp/dgrB7cB2jV++1YUea6Rt7p
ZMOsg+ZP+1kb3NivaGtXegfxgun5Jcoivd7YHRwUCbSYpTUQ+UYSWE1WkFPN20ta
g75wfE4mG5CKWvH49a7Kx5sP6zBAhVove3TmdOHYVtPVHUw0K/rzpwnuqPpeUZLO
aq1GPrzysfsI9hJY5bDSNq/TeL94PskDqG+r5+a4HaQBc30mGkpOGToglEyxLKET
RzL2arTegtegbTPm9Mo8js3TfMej3fQncvMTvuR3qJBqvnbjk/hSHZhVGDu67TOA
uRQ4b9qDJvxSeQmNbCJDNjCz+ZMv88pvUNw6f8TZvLJBUqvoXpe9eP9+es5TBepE
s2uJtf4h6sg5wdWeuypOEPZOtBeiUSfTslX5p2td0riX+lYUp0Qo0v1zK3F1Sjg7
cx3+Eg9/RASb7AKqt2GbkND8ytWOEaxiBwH/kiV5W9NQlExe/H6Yo3rrhEDYVTTD
lbqnMw8ydphegsjQiTLTJPkXgosGmyihLnqjPFcguWhwh/W9o345lAX0hZxtAn0E
QvHRFQYDgL3yCt1eeRKQB1wm1zbTqF6ynNw7d/N5DNjKVJD0QAyl3ZBcs/u6AnJB
j/MBsqcHiaATThkpmCZVm91l7fkkAawikiNQk6MKRVa1tZy5vxXc2xYDhArDdVKO
n7/C4moog11WrQkhHUYO6NcnwdolzAP+onEkCk1Rv7WwpVqsnioUtO4oWwCigkl4
shzW2A0Jvf/D252ewKjdEfgc4rawTuZPSL0+CN0bouDv4vVC2CyaY+48ZN1YINmF
LWWHlieElj+45u+TswCCZcJdw7jLQGbY9v3QSE5SejBxnuEjv5qUKaIG7FYmMID0
EdnzwL4HXYoGKf3f410699Sq3m3QfhPLKMH5kEH6pLxj00C1f1Pzwy1B2pjU9kdz
vpJg7bLqTW3rat5g+Lpc/HzqdztVgrAU5HHmtMq6PH3t7910ytuS5tJ8yDRLwmFL
FM+GI6BmgpqE2MAJKEzzQ7PwNKZeBMF9A4Fge9WHkMgIzPNUT43mfVEUi8xy0kEe
rcGFYE5BrDPwJ8cF+vMgrH0ZUUjLm7S3nM/3146C9mysmFRjSyvNgvUTgw7VjRVy
UM+MT+XopkaanbfmUcV0rhOSi7jAP0ivdZggjlXkpJFjNx5BtitOg2TGF+M++PsM
T9Z7xZ8kI/1eHSBjL9Rw2hdIFhN7UNf6B0/wakVE6FBvqdDh5ecVezt5k3TEJAfZ
ktbbvmwkOCZRCtPSa2L4EXKZTo+bZ7cyAe7OWBGpKDQ4Xi79W+UgGA0vtN3k63t7
r90ERMIwogu4Uk41mzrqdOKSi0Cu2FHJJbQzsDjLslJ0QacHzfF/IxEZFBeNferX
c91qdwIJE3dglOvUduaty2H8J+qBcOeU+PFHmZYSmf+7JjPBmFCQtH0galFwdZ9Y
0MuO2aX5h38/bz8quXRnFgACsuEqcrjy4w/hg9N979zYW/fZXWAHbYAA+G3+iWUs
43kOGYnNXw2WGGjyQri/TEJ52kxezvnPygFHDt1G8e95F6v/EalEx3EJdkRYqtW/
Hj4mw+cgFppybGZ1M68kKIbqlsnGKeplCkwdPQvb3YXW/O9p8JEEV8/71ckOzSUf
J/XO40pLcVjiPlhyAUgsMEV1iObSxeeQfXcSz9B95GLwTzppCSNVve9RqT5KUi2U
JZg3gdxvg16SB4tT+NUuOtWwTetgOiqWW9buNiNucgRN0Wd2uPZlPnsq0faAEvuw
7cBPmBXh9mS7js70YjyfMWtr0tF5OFM/H7IdpPH4c2YV9EEErujcR/nyMAGOYkvu
3UTO6Rk9Cs3SUJBU7Yh2y+qX/vQK4WR+6vP2ElFLeh2Z0+wC/KAX2LwFdkmh7L26
33UPr4Gp130GrrBHFkQUZdW4201MR/t61l+3yuoAvMRE/ClULL19IUf71lR++KCD
nHC7goWtz9CJCX6wzs5nNZfS0nWQO+zuf8e87VgsCycJZWl2PYfo9LoU+e87xOB6
weIMsTljDyRh1j1eKACY465POU0ewi37E7oLIpwcWpPUGGhiaESaAACR/N5mtElq
CuxgnjG8N05xhh4GBJC13XHviR5+S0H8HiXfvrbhfz/5TNxwq23uBpV/KPDavHQ5
4c+//SNaOiVLHHJNdaqGygqK2HHLKFqwFcknXfVhef2OF6KWHs82zDp+voYiWEkF
ozxGvt5NSlr7hSewaURzgB3NMWYQ4WFhpsZgv62o5jWl66VTOSA9R2/9GnSBwv9Y
4mfjgibLxGd3m+O9n9N5sPeaC+2xVd11ZOITiN1V85w0XwFPb1gOee4WBLTi/UN1
d9o9SG2uuYGdETa/JFP2xpSXHCEdVXKVMbkv6bMMLmRVYhZQNrXxMM2acHgO8X4U
P6PF7tKLEtRANXFO2J92fvoHmkeUIcP1eQDYjvBeALbOfCWtJTBeQmyzqvlmBvEd
+d5NE40b4ubxtfpBnD7SWe8/frTrqlNODC4ZwnRkrIDxyvw//94WJIeyPd8QgeU2
HcS5yM3bzc5wtsl3+DoFIN1Bva0cyFixqQwgDcLnL2tdX0ojc42iujKrogbgTASr
bW91bkenf9mNh2tfVaAI8OQ/UmtEgP1LDtPJRyJMR7PjJUcYGO2rM3n2LYBgKXwm
etDJKgZieyrdr/DYkUPshi4likSFqu1N1NORfUCchc2NnM8uxIUDg/lmLaEmR/f+
1tPkquWLNhRM4Fsylp6oyHkMDUelwYZKn2VNuONQE1troTZV0kTHWtPN03ASVx1n
FHdUv7vpHj9w2dk1SQVa29Jq+AMGXuZ66ivVXK5wh/jFBJ0Mx5BLFxB4No4JIoXJ
EFAunezFyye31qXXoW42m6kXWG2DzB+GF366AgijTjpHlzLmHG54D7FGwytXbdcy
iq0lAV6fUe/vejyzfhHzYwe+K/2C+1GxnUTDWQ5WRtV+wWP3A0vrnGs5hDVySJaI
VnCjZle4wcWoK8Mgmyr4c1H7OMiGgTSE3myZYz8w9RRzCrs8tqFkI/nNrj9DFLoX
9gPn3iTAzoW7CpiSaNmHqHcSeAZLRW/SfuZj1yRy1Y2AisuXxe6fCqDQox9/Fh7l
6txIA2gPhZzii9UdMR9x2SmWfPoDPWZ6DGz3RIAeVvKm4G+78mU8vwTNw+vcm3Ed
Li4KLfr+DmrW9EtiaklAWbZI3LbmCTtArxfvSt/gwRehFk88j6mUxJd9OjRz6SBE
mWMcDbgUQOcmTno73WBRWhXJZxBQdKt0xZDdg365AR5Prlnaw2m740I+xVPw0ddO
Iwk0nMurQUfy9MyBpP5NVOUPie1gBcd1bwXsi18NtqK62xRdB4Rt0RdLrR/G9Co1
NsYodbNnoOD6dB5yc+dbKxNlMajWYLJMZfcTi3Kg1A9fVtHvoeY3TWdnk5iFWqfc
Ky3oMA3nm5YL6DtXcl6TcYxYG7VmJOSLbQkHzOcD7BzzFcdnrufrLrVRRFAOY7Up
/n8QVwUDZBfXC1LOM/nuSDvFEm7w5DWGwzPnLX8sxZ5AZbWzn5lWh8y7RrL5UpSo
tO0r0kZHrD+mO+4SACE9iaINzc5h/kMMMBX3K9S2Rp6y26kHZIt+J3nCf9+b5wW1
qm2VeBL8undv7vZerair6b+h7an7bke0+Peb5GEsRoBHIFtK44lzaC623n9EP2lb
TlIX5qPAVKO+InE9Bx9o+EShDrIb/x7CwC7JWxsXql/0E/Hspf4K3NplK4ta7t9n
9HlQ0cIKw98GfAJ2IHWIUbDUk2EjaWuy82KSSevC0BJACETN51yswmPdFY2bB6Ko
qMe8bQuSWHa1tlWM6RN3oDSkSH9PLvBNyPu27gpsss2N5qOWO9gGLdogfcGse0PC
NgarPrzKJNSO3SYnRdnQ/088iLp/FOfrCC/0BJuDYhlX61aX/rlYg7hSo6D9Vkk6
u1EFSUq+CkKkzKs/DsXf8BpuPwXqLAcKlVu5Cdz++lPuGzhlJvnoDFeJLHOz+1/W
rMSaq/lBlaoOI+FudKBlPe+1KjqgpGSBAxwjwEewT2GAkuhnq+6HbEqH+0xvcC2Q
K+4vgQP0vqGHZwdgp1ciMpb/eJ5ya6O7xOD9Y6BvsgJzPrJlgpGAdB/1ogUtG4q1
fjvqIdtNgUwkJ0ck2mUn9kY0/ZFY0HfWPaill4AwHihxQqh1RhAxx6S+XFSNXm9n
qaL1FoWQOqvlGoX6v+tC5Jo3FXch0+mO1rTps+Ey9SF6cbgX4I4XhJ++0lPhhcNE
i6l8Xsb76Fzbc8B+JBOsKpG4nM9j6nrlMc6chs42knRU25iEs9i8YxsmhjoZm1cp
B6KMDM9zhdU0tA/N+DumAIH6vX8gfPBUTxYJwaYaSjpi4YIa72eCVV+09a6iXTia
DfdhPxhfXKOvYibSiJ6E3lNgvAciCQoMeOc8ab8fhbyJsWnTBUMqk1d4XEU10Hp9
5TjQ6/bpA8IdE4A5fSy8AtzblZ5IStDL8ukKja+Q+TB00WQdoOf3cjaDw8Yq88J+
oOXJgz40ewLr1931ct7weoBBPiWjB24E3A/uEvrUCTQOWuMJEl9Qdk/mfEEL+KEj
elNTYsIhkid1sGCUFtPVure231r/srCn3of/OuGT1aeub2Jb744cnGJZcFc1xZnr
fbzpLVM9WALo6Qg/TmCiMXhH4HKHCPJtooYS/S5+IU6cEEdBjC9xHLqQqMt5ZPEn
rqjZm+B3Wr57QU6wtxZ8d7ssr4OahGY5+yinKNILHkmVhXLYWJPxoRa16blWa0PF
LozdepkE8SvJwSg7C9ml89+KIZS2uqSInLAhSWXFsIAiFTMm68zMkU2BYNIMYUhG
W1EtKLzJ9OKt3T3XoV2gzbYc+f3NS7M7FbvI9fu0tvnekNpdT38g24ggKNly1H+T
aFQocaSWfxFT+4r2sbYxG1KoMo0nTuvA8axPTTTvihxLQhkO/XU8ATo6eUnGNUSV
rzjJvKAf1Qmzu/Dts9ouYrEfbXTT9/DtDReSpgGINneyeozS51dbjgXrDmdA4bst
8kyP4iW196rsuVjc/htJwjtMkrDN9KW9l5Divp8NblNlVAkTFusufoeSMpS9/9Dt
3nR3rXkF390uIjdd773MxGaLFdk6m+q8zMqHLJZ3QZcT/LuTbiQ35dJn+CN/gxEw
crmao6IVSRBPddRnkMNa3RpT0ZpsmpxMtvrahWwwN9xXmvt93Y5Iud8z2ZKkPxaD
eq7kJa7H0m3GnnsGfBzUYcErCObkAfykO8F4zJAo4n+mzaIwokyZKA4vy5OGYqBc
IrEK7FtK8nCTSuao/51h83/t8ig35e31S3B/rX0Vd1dfYUkEcVsAYMTNJB1bjlB2
1KoKHY/0lthu+Ekh1j0UOC2Vjta4xFe/Imc29Jv3IP7FQYE2nFfwG2ahFArMY7uv
gb48j3QucoLdMBaJvE8KvYfhxhvTkJ3CLp+Cj+i+XypkdTMmNCxYj7qMwlQIXHGH
xPSx+l5Y4FKb0WaAM086Jm/dNrcf0mQk9UlFbaSC77SD5w4kDyTwF/TkfcKHhFp2
mB6vaNCIQyJbZsE3SYWlcaz6gmzD4IrIG1gqU2ID/ntyq3BkAWLvyEZgbtS4tfwr
0dxgkx/a1JrYtbsEqCSP4iyhgx2OjMevjAxUC93m4nF2unNf2GOlI/uaYNwbuHTX
PV5oEjBbDHWLi9fQDhujlsqke+DuTvOPnq9dS3XVcCNA+KTL+d1+5cMQlsmFwxVj
2IktYvA5YBf3XV1wJXrlovqogMTSvLFoQbsKAjIdKixPfvTn/RRPTFbtd7KVVaIc
dEuZQMVkjx/LZ0ltvPpUQj6WG/S7YoaUfXbCC1Fbu5jR2Fi41zj5FSVfUeAusVd5
Z7tRHztnQaFi5aCZne7urudYfRKxu4v8M7J5O8WdOGLRK74p5smWsT6ZEnC9QJ/a
iv3lAieTGGs09ZMc4xAiHvsmNWF1zVUWb+/yWtnmrX4+jPZbhdOFj2FqR7j8L3th
1zHrWdiyBZJSM2seD+I5/cnahINcipyBKxMFAUVREcZgJI0V2u9uFZk9dstrgbLZ
1NkpA7l1n+Uor67KDSqkRJ7YRwgcnv9NdhY4LYvu9sqX7yhI1qu7ZDFHNIoWGMM8
ZqfAvSHcoIlLrWcnsVBxZk3DwiCYkevPNYF5hECNH+UWm167VaRc0+cBXEm6uWrA
83WTiRZjv9OpNUodHpWqjWUczaO5Iya/kZI51uDLPYTKCC4WUtf3j5Yh+ghNoM6s
qNiwO/kUiwLVMIwMpnLk1vxTypReIpAtZ+6iN/3w/z6AJXUzhNi1ZM94k2sP1JF5
j2y6I3HTs9MiN9mjpyTu93KuL5UE3em+GcsGWGDZzGZIoK/Le/UA0jfG3wnz2bZ5
hzavaGoLhyMZDbLgym0Wbkg7hNKQRhNfvVjUtK6e0Y4V7U3+/KZxZdHp/rAt7tsp
zCOZxaw1o37Og2AIbvY+t14DL8J6K52yRcr7Xjs47GojtQO++L0OAfWAZ7hGqGQ7
HF79qVWUq03V79+Vl9qGq4Vqpd2o/iz834KGKNrVIvs0XIZhnWuUd2Gmcyylu2zf
G+3MEgRDKCH7tnHPYjZ2QMb/LU3yagsgqkcg6WrkjhAINEMvOYSPzMQ9mJbAlZMj
ZiKZe4ibC15ewC06w1n4scirS8jm9y1S3E+l+fZ+aADa+hDywDFh130BrqHFhIJB
Twes29PZRoWmZuYMU0lrfTYeIEovyr82jhdN+9ZWQbqonCjja6bUcy/wmlyUu17Z
gqMaXgei3ACuPfcOKuRw5GasdA8mYvR4hBc24ZmMRoaIeL6H9swVi7HJPUFTJbGl
OFC4Bdnin+XOo3FNJHbiEMpHvzHUZGLyTTTGS4qpnoYrnp7q6t6bwl3Xt+kNFdur
Q5/SAzhM9Rp0mLDFCgjebar4EuluAh9DxtZMD6s6QrXJYebRwinmWk4ljy6wBKBg
vqBMe9OderMzT4dUVJSwJ8JRiVRr11IRTd/kj6AGtDlPPFj3L0MFcQPyLer6K2tF
q6NjGZaqclGrX/5LSbknzv/sGA+lWegcDTvtCtoKUKyeuCalftwZNd4zfA0D7/mo
BRbFCxMZN8/9kR8UVUKeuUfIkQ+CoVcaLSL9+qKcq2+uon6raZi9XlizRyf6i0M2
HVjDdOWrMGZTQopmxfBAdn39j7zsmGTQNqKKetRbfZHEYpxRtck8+HabAfi+N2A8
PtN2KT4M5CpkLnxRpmg5RuZtam2MZjzp8NUS6HuPiipzKOLgGdsTntwttb7D8F79
/81NLlMHGSHjc4/O8E8inBd/6vKda92FClOT1Dt0gZRcWwf4Jki+TMFF9Furm75Z
aeNSvgjk8jzycvXM/RH3r2R4rgy3nGKq+Jys2GR4Cu7Hk0JCJ46ZpsqYHeBDRnP4
rf62LaAxpYblin/aJkORKMmxrQmIAoJAKNrbSmk/bpOe5cXKAjWjDTUyJRGsmTjJ
ZubDK/EOzONx+9JWLSP46IRQh6hLuwTJy9YWX/MXvcqylHlYQx+8VABaUhodRykK
2vPeEzRv4iCcy9w5MQDD6YqEr1O4YQCF2RyvpLaxTj0AbLqls4VK+TTmcm9Uj5QY
emdjIq/flCJwBySNRcdUjsq4WiWnRZnlqkCw2gjNaXPfI6O01Q8JPYkmt/VphBRs
ligzheq2XAYKmHpFRGHLBjMFRV8wsPQzy2Kbj39p9Lc1hUt0V1sE5iAIoMtNjwcp
ExeBw3QjBKrxXY0kX0EPGLxiSfYIj5KC0EepkgE0ixlCMMmMvNWdOlGS/5U0qIET
S8/sET452uZLiSfw5uUvNmUQJo8Wkz/PSqUadKzw0OQo7Vu44U/EO4w02wHdEKH8
HgfUGeKvBIvr8pUZ1njwhHhz3H+/K7kQ1xSbh2Hm24BNe9j5T+zUunNxovAeswk2
QLHYrBwYB94t10hT4YLs7tV8Y2RrcKh4NJyw1fwN9Oz3DyAoXrWAYs33JiHeUj/+
E8lxFb2DH9yBwS6oGOSUA4CTdaFB6J+rF7HVw0NcAl5TSe49sLUMNeD55ewu4ZsG
aZ85+6Thhg+aUiXwypmqQD3h5+6sBf5XWHvM+6mTt8orMeT1I7hFDKozWcaQFeml
1jy43f+m0Xi4j4jLbLrFnSIeO9GxItjG4uAKu9Wq985SQXhUiIVoyTz4Bnz5QXY3
VoqT40EVucJjo++0x0OumQgfM9EUlUe44WpBMsggF38e8ZX2NQ75EjC4BRgQWLOf
/rSY3B9e7Mb1tJoB81LAPr9EsqjKK0k/LCpNnT37r22vJ0v0C18h74yw1SICFaGf
aEjUUiksjB9hNKZtpBbNZRVT/zsBjRhS2uKKxfITnlpGHyE5VIertSqsWvoqE5Xf
t3wenVM64xO6cUmBUL5jyYjA4XcQUR4ss5/E5OWIo4qvYuyGyDZ+DlZm7AoN3fJE
YLovJssuJRCmK0IMCdAr8P1eNTFCfv9noZu8uJd4RZ/0uU1Tgh6rtE70aLXovIE9
9UBdkrdlvJ2sSaq/g1nJnvtvCtX5/pVxZs38Hmel3yWi3+cvqRA7QS2Un4mu/o8z
LdQBkXSB/Qg0krCHOoyS5GnMgBEuODmT3FSC4ANTvXFcQAoZ+h9OdP9oK1JRlRGF
+aj6iGNgvMgvmIL5F1/ktiY4hAx4YrXCxjSzkwsLB6A+PLBSF5zEi3xMrODmSxwb
B6tFu6cT6y7JaXK4v3m8V9Tto7YzbKo2LWIxl/eJpnRpkPp7I8QI2l325y8uZV94
eQ17eBQJ4fPNMBLZriTHE4tueYL5iYnoUO3Aw3yXNRxNgG/BBh5j5l3XOnzRquFN
7LtVnLzV3MY4cPb98ybAntT/3SDzNi9cgjJvexZQeBesz2m6otHN1+d9NAmoaN0W
R8yF5DK4cViNQbO3JONTvcX1znioGj8Gt/GoZCxkPxjfZO98rS4DuCKCqvZK/+m4
HRJjHmuvK8F6NKdMQGYrCl1xl58zrMYS2rKFwQ7UKjdQZNISvdbSA5A4I/u8fSzE
ek46H0ma2HNjTKO7BYvf12jppqDxUTqTgmKJ2gERPRh15JOm1h8x0GIhg0u0Ye7n
zTI4KGaEEdHFwd+/BI0np30Yfm+2/SAO7NdMn4TDrBjJ8ex6fNA296sO+TVbplfs
8RktveVvpzRJChfURBmVfsfW1SjMJOTq0wShzfKCg2xsdYh2DQnIuzUSBaDtnU7a
XZBscqXrUpJwjbtJLxRf653APDCBNa6ckwMHLz/q1QBobHWT2rlbGWyf+uXdUse0
m6u+ZQDJi64Bb+odlJmRsv9zo3FjfymzRHgrkWuy1ow8TgZDZc7N54k0eEfurvzV
Wx7gbeG/tW1cO7XVhlyuWvKOvGxgwK+Fqh5gLNX2u6tJcdMTERR+OiIVNMWV1tOO
/2OeL57vRcXL+hnmHKXEZvEF62A5e3ugb1qrHlZIsJtPG1EEHZPOsB+VOicI6sqn
Wpu9u4CbsN+G6qwFOHOykwFFqC6iOSnB4nlCe3FcamjngCLYup8Ep3iAnHELEseS
8JYdgmRtJhYVvZLialO5YPDHMTUpkC+DwltEOykDddxQ5FAmvoDmGRvAxebB1iQ7
Gwf0mM0nMb5HxvDXybDHpF+agcqa2dRHoLNUeDgBwLnNwGW6d2erdhhK/teEBd5l
rJgopmYd7ZB2sKL4zAeSjYObRWRgVM8qzM+Sz2jS3Aw0Zt7dQ0uq0jniEquKkQEN
bjO5Q4wEAOcVAsZY4OlGn+sQfGugLoRwf9P/DdfptcH7u5f7JGqYAHQOmEivOxsv
rx272wmCWHyOcL/7dloM7LTFyyvwWD+5GxXwBvnzamKf2SDd7zpD0UDI6OzsVbyZ
TFcXJBZMmv4Ia+NgR7od3KrN5SpyEy1DiSljXC6yEy0O9MKihOiBrxj6jMEWpPHl
QCndp6bo1A6aXVn8m6Uqo5ubr51AyuzJNHwPugKn47LqJ7Y8BRj8kHcL+7mAcc6F
G0n27+3H72zHpI2vYKd9KtXo60Bp01vpEKBvaTs04v2z9J/LAaXU3TlBm/Uwiux+
JgdzTRzml/bD5EW/sZkPiPdFoiF20BYnAMYPr3deUlnsUCVGAtaAt24+7IQJ3uD7
EpRP5JDCgqgO4zrVgMDRubyu4kzCdX+MUndiLHdxD/BZDXPeLORDYhW8Cny1OZ/I
JzG5qd7zuHoVusiW67PYxNMrvu+AbjvQy0g1UG4ibjt03U3LMWcziaKHFfZuXl/C
Lu69loIYZqBfpI8FGp2zp/X9jWchaBuugXWoka9nwMX8cbxDDd1bUhxQatpNIOC2
WSL1bAduYEzXWPNvzPB/lWvp+deSfnIQ12wflrqEH9Loe1pg3Si3Nu87Ss5gbnQr
MoGpFC1l/2gFggMp4LZPKq/yP33RYZSIM7+U0PYc+4PBRsnJl1A9ZPPJpB5Cf2hP
pR2WwuB1BiTTghuUTG4RlKWFfvCePovl+waysxf2moUPQa19Daq4YZgUJ5RSE/iZ
NKYStaVxKDR2ZYVNqFhhfVk4uhCi3VW4RafSrVmH4/78GhLBPnIF99VIPReIWqdA
McNSobDxhbHcy45GVgi0wa6l1jHY8LczIPbmovLk/foW+ZFEn8RxbAcpxN2jyogc
x1ef0M0MBWyPt6yc8gHLZjBQSV50yehMd3y1RI2j3+WA7PTjjPhNYXZ56VekKc8P
gEv5Hbq/4hMzHGrT0J8KWw1XPwj9IYFShtmG0TvHe24HmbGsg4htnj6qBJGC2N6A
1Y+Wwl8F+I5Eboxx4X3TwAGfze/dc1ebfT2wIUnq7FxNC++Zpf+XVwlW12kMLUHq
qcevPV/jv4KDVx/j7QF9zarVVmza3ChOVIeU2b40m9UBSow1z5vR4RWV6jYflQ9R
WOFpFUeaCOwwp6qcSf8lSCb3JrRD8xEUCNtvEMGS+zxX15GyMhpvVcRoWADlh5Gl
vgn/dau9nWX2hLHTY8O/2WNO7g0VyyXEDKabefZGcwMDb1n7v61fnxy2/Xt1wyyA
kljhOMeVAGvjBzGnl//JVDu/dYTnmSV+/eaDsErel0707YmjHScYFGNUU9JfjOTR
S7PJOMHBxVqikmmIymGY2ROSyGp0PXE4SYLlmRDYagqp9aW2LMG7D5ReXv0fZ0jr
a9jom/I8p+Y+Nh+2CUKfuf8Zv+8QAHdq9dJV7WZItJdkTTb4H7XBcuRdwSwO3m+O
lvfBkRa9mCnvi6iVuJFZE+GsQChCN/2SYLTTWVZwtsLF9XKXDjHpqVlNL6Nlf/ns
7QJqd7m1rtw8tTaPKlbsc3JN8a5qnG7syoiZ5uDydeQL+BLqS7cf5msPxCcTznVN
u2nGccPtK1VZpljG71Oydw0thOz32/zCVn03X2IU3+W6PY0u+ApaglPiPMAUtej+
dp0rEy+1QaKhK0nN4+6wH3YUR9wUoEDUohr/AkOxlMKdRs4gbr0oYvaWmaNDavKj
aOBm7PsxqDOSofh+TGkfWGXNdKsrkotFgQ1oCRmNgoKKCFroCqhDsBUb1RMPPbzN
c79VqgASO4a7bSJIe/pa33FToEuuORGemVZPlJVAlObHEe02LHBquPdz0tzMVcsO
u0lHus087MLTc1q5Qf/YjZg7my7lZHbaxe/SqvEEM2snuSktoy2PVxpTgBGRTjZM
eg6Bg/rBFJR2sFILvrz0GSbi3GoxWCY060YAB/6Z+K0m8res4yfDVG3mz1Hd8XFT
nJO7J9XOXjUl7WlGXouniJRhuw+M0RfOvCsT8XV04+MJUzDOhrecUnMBxYms0rlQ
tQH56odVfFHx9vccOGC05hkp4GVMf+e7bUUAsStc2++KA4TLsw8Fcq21LlT0/d8L
x4fO2EQxokFQehOmKtBdNxT3ze08HNj9b+89S+i8vTt1F6GfuKLMBdERHdhOaPnQ
dx95r5BpIavZ8U2vj4U60uHwtBGiYJpa4HZNsOtluSJOSclyU/JUV6QBgnRLZOC1
qBa6J13M6S21bxkyEQUlUQCW1IF0rCMlFX5JT4y5y7keMHkBl5mRoM3Zy08Nxl0U
uR4jRinsZHCYfHB9iKA8/swRqCBj7gGU/5jF6qXlnQ4f0KzWWNSVABNHX3U7lfEs
p9oqTnRTbQvrKBiAgzHzg48U6qUqNPG8whHdCc7+k9fT84tiOCruxplvoH8ewTSl
NLNuPun+XvBsUFjmgRNq7M93TuNRMmmIvuWmsdvSK+1W/tkBnkJdsWMtXrG3DXex
0scpk6P3Ln2x9jOmABnaS0VB0QKmHir8QCw/jT/Lk8B3/ANbCdwGqUAe7Uos1YkP
w3/YcVQp3mNg2aHMI1ZIUkdu7lTUaAuKZzIGKMw8XEETati8UnZJyKn6eJcQMr6w
iGbbhVdymcJYHhDwASwiTVkCUD9Hw/1uvgHkj1rZ0BC2pNuuPpQsGDFae6r6E4Xh
kVW5tsBMpPaPXcWPZH7T3PCidhpu8/oZ8KheSKiVdiSsUc4sY2gJNgNkXmgpB4RA
Yd+7AF2xhEgyKnhyUeWG/JwW4O0TQVU3Bamov8fhtZRSRE24IEX+u0UWrCwf0J4X
vVgCYQf6O8FkLEXlJcESDqODYVOBclrWjUhxDeKZs88MPZi+teJXQUevlS+nFK35
Dw79LybEZo2QMF8vaOy7HMhpE/wuM8VyeaFOrv9yqHEazb7pS95sEsiQo4Pl0eRa
ItkYn+Z5pHG8I38MIhod0CIxU5Dy52kcMxVXRgrP6qc3D7ZyOkaiJk2IQY1kRlbS
lwYNP5qKk0aZcVAdNA/ddpRJf66jQOaWA7QD4ZUl8p0Wn4sBUOlULLIFRASIv5zY
B5hhOw96wwEs2oGMEzO4U/9pKvY2cb0VR6cVRz5phT0PSX3mCz3tYqxN6OgU2Z/3
qDP5fEXXQGCRiUYN+oW0SpqSk9PaZzM5tw+Ms69FxKKfNkHRDTkw5bfkDR+j81t7
6qXfe9YlDv0BvR9YU0iY4jGTFo2NMPN+OwHsBSiElEVC8q++5Q0yonK9GE8h8VHr
CxDiDzHf69ZZMh42AEECQ7ElVWPiLymRkI8TXH6iq1QFiJPB+92Qv6MGp8SyLHhx
I4cCVYBWu1vsNDB+fA9Q6WgbqKkmlL/JITYCTgMycNhujOK1Xl5Oz39flRlLUhmu
bmiNf8tjZM1o8nFNpMGIHwThdn+8EXd7FtktQv1YY6/YRiKs9ErM9MRoR4v/8aOk
RuvZeZIhtQCWEkgE9JB5aAXZIT78kbcZGi4vLDkyK08JWeZvVZua4AVgZW08OZSM
n5Cix3jIWzIx+mEjyAukEfFlS3/TwHbymTjuaQUNyGDMN0M80wTgs1B/MqJXqvag
Ssd4EtRzyYi3HFi2UqHNtem24Y3A0Qw9hd+UojjWN0gkc7ZF932l5lY9UYKj5Vq3
q4vRtzeuqitw9jvCRwa59aed2QIa6/+IwzLbhhfi7j5cZpUtj0aNthor+e1yyGTE
VPkjpVLr8hV//43lilGQZ8gw4YiDVQeYrfmX/63g8E7cQVlGaylTI6Qs46Iu1xDP
MWjhM1GO8eXDc332VVgh8rqon6QpEt43PC7PERsxfejxZOrPDHa+b7JKwG9sZy1w
ekVxQAgZSSd+gFkxb3pWe/Ye2h9Eyd5MSF7XhZVbbA3rfXxOa4CJQQoFfzoJRH5j
sEjkPtaxjN99ikMRJZ9sdTwRSoya/YvSzqF9xq3fx8arddkRDjMNmCOrqVXRu4ci
0ENkzQoM7a8v+QHAuogMPaRlfxnF38CiKVcqjZp7Z3GhPaT2CJX2/0rleHw+w306
3CBfeS3oyWwq0x+P8Ic3jU5ZMJ3qovhUVXYJGSyvG/WKudEx6Nh13/f1bu12PJxH
h2tl+hyuqD4LK62zDaCw64GowHANjASy1Ask4Bd88EvPaS71Q+TnW/wcpJMEPMJd
f8zn9HwsSwtNADTMyJBBnqtZPtcBrrr4UdAdJH/btf4XbeeCYsUO2OTYDZJZTsRR
nnP5yuls52iaPE+afLmOz0D5DE5hKFtxWnpUNNLGmNbitNkbsY7fztiWdk46Z+L+
lHVosoH7Uw2TxWZ3zEaoxbNqqo36/CA4YuYmbXKj5i0tcWlqh3Y5KYlQ46xamWU6
tsX84lMjc0M4UXMrhOjcUHtMITWZ7GhSkTW32TafZIRAl29Gs0o0Z4wbia3R3yIT
8UL4Fq1/udkWVoiPTtdjkd2evFH8PWqoHo3+QrXQWg+xc4B8CUaqYkPQzcmtQmmR
zyNusIr+mTYoKlcd8RFoJ7Clh9JICLdSeNMvdoygwIQUo4ef+NsNeKTG0odfstxv
WJjipkd2PHA9smKW+W9GpDDEzIWErXxESP45t4nyrzQJM/1M/CXlp0f+PPZJxhAw
FK8SvELNZ33L6riVVd3+itsgW3WVxmf3n06yY+UNcpZExKztTEgU/UFTYEtXfeel
tdwfiE8bIjxLiJpI0OtYgRBqJqlPp76X0TAtReuHXEUA3gee1Dve1TytqF0kVX6s
eK+wv6cltS89kPUp4XvO1jTd7IqLOIYHLAZCK9H5o2AyU4+vo22Iy0yPHCqa+Bjp
77CH686ngwogHogHJt7cnFs0a5FAZgdzWo/aF+PtkfqtJ+4JO87ex0V+kIksu1Df
A2eQpUuGQmneEKECJT33RW2RErd54eiZn3TBlba5qRw1oJubMbFR6jJDfAUM6F6d
KoVAMavMJiPLDv5W60QK2QJudVH3miLPRMHSaU+oodc4xo4JcdoOuFWO6QQtuUsW
Gg5+KC2/+SmOx2NnsDpO/M3+yJxCUEk0XqnxqGJd/vgBG9fGYY+P890XKYRRBEPj
izDV+pq1tykTRsl+SYlnxdvnNysDq4iRpldCuzzr9q8SsnAFlbqB60g4kJM16QTA
+UX+89+5XNLgoxGhW2jvBTXOf2kqbYPE9UOJhpqt5XVSEPI55FJe1gCozAlCtxrO
fwHKmYp7aK5Fu38bLOcVVfd0E3q85wxqYbkm0DgCeYw2VVN1j3saaXM1f2++cXSb
wT5udn9u+HpWixysZSPZ6oDzNQf7nHIPpNzih3B0XapT6IgYvAfUJ9wn88DZ+hh+
p1YpaFYRQCrqzd9tnO8VMcTWGWfvLXRxpUWUSwyvb05St0bibP3IlQBNSaWLKDdA
hDoW3hIYQP+7NSOfOMUgb/zALKmbncEePf/blioxnpVYH8OobpZIXOUGR6aWaqEL
VPY0MszbDNK7M+2I7nylwHv9RI6lzzzOUQjXchPcCx5yPwPMsCfJXRKPf+LiCNCs
bK+sIN8dP3XaciEDxXFlPktDD0mLsqFph30VJnP33RGV2jQaEvzg2RwRmkttfqAJ
81RAAfHzu6MnXt4CiFKCssxe0eF0GTWciyvaFdSO4fN1RWH6ZBHRNKhOUjzVbvbY
UOKGWgm6oC9I2hVxhjvzYeuWNyShpXy36bHPB1uygKd131MussTVYEJ3TxtcNhZV
wiH8ITCOZlA/CfUReLGfXJbnIQ5d4jjdnMGzP9VRsbNqElEgqG2i6UfLYuXxNqIj
rQJrqhCXJBrULgOhLAOuXFpIi9E1WxckMeOtlWp8zVdGwhmZB7FtEXXZnu6oa3/e
fjkvft0Qo9wrpal/lMjP0aBrysFIv/q84FdWKoA35lyIRGhR/mI2fFMl8JnYMOXY
SzJBLpMvEBt9Qv8BlrfZdn87RGVkOmTsiReeKpNUaaPXSJ8bzUJ+ciXtYw5edg/c
W9JW0WwiFW88o7Sy0sEF49hPGasiDTxP6DZhkP2j4tGKVdJ52mIrbx2ibNhmu+j7
wMiYMQu5wtpX05Kuepnzt7G30CgA0iyXh7lQbMTJwYb+nNFjCjFNasmKAD0wCJxk
75HZwnqNj5J9jKRk8OmQzUKtOVFVzy6flCxokzz9CGEHgdTETHnbli3e/CEw5OT9
h+U5Yrxt7cXshLDEqTmFH9c+X0KLmzA19sRE3Fkl9fIhcMWjJNTq980eEak/P2uU
7wxOM2TeJ4xULjPAzV/bq2+MEtYZUYgdjQIs6+EzcQlLwbh9MbFalutSwKEI3nWf
9Tt21Jk68/xLk7HZWE8bz++ubVzCRDrpMR2xy8PniJRNg3onD1rR4e5zYVdzkRel
+SdEQFILPel3QQ2yAVyztt+mZSbxJ15WKQo8yRv+9TIs3uJY+XeJaDJsukROnLkb
zRFN/RdAs/FercVPiLMa9CTruziWyvH0FNw41LVjwGmddoCBY/DQLW4vXPsxIRnh
840I/UywXiTxlAzVkZInTsX8WfX3oxQXe0RQr+k3anp7/yoQ67nGkSYtf/AV8pLB
YtuFo2LGyi6IzVxb5c09qgpfvhyod6F4d4yQGj1NGXyKrqCAr+/HRD80RpMCDXOy
VDt1WGU1uUZ7538FdsNSCnRQDc3SNNf1Gc6IN3HDHsuUKKnumzT97kMpYZYPuWwl
yGrhgo87SUHJbE14dsfS5cZVDgpHCfvljy57pBQbmIWpz50mpDqR5xgEjU0PcXel
FWFsrhrWE/sMy8K78ukSVSBPfwBrDp3l1VK9tf2YYktDv2hL8BhzQiY5tbPZ/wC1
infKphdgEyhh+TcWoiT4C+nEV3CCR/w4s4sYobOW/F4O0iw9VExwelbGS3UBktwa
`pragma protect end_protected
