`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LqEACF85aTdhH7Rb3gacYRTGSe2Wn9eSdy7z1qZ1CvLu6jTouYPc9TavvDJYTGeP
wJEXBTmxcSFFjuSEne9G7egOuODfeEbdK5elfVvqkHYUS6DNr093XuiPLMuRS05d
70hpBbKj9lVUC8UN4kBsoJlxAFyrglUXBeEldn95ekU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
ZME9rPnnQTXeJlKvwQusmIDqXdnPKrDPVIDkNH+mcSLlOS1uE3WqyWtka+k0A/n4
Wt535TDumWJSklE+ogZ4zjUwiBlAO1eXNlaBwGkhAgB/vueoO6yzP7Ykic5R80bB
FcpOdOQQ7CQf/5Uxk9s5ImuWIhsYIxKFWMEWIK4WZdh5BXP8KZlb+1eyPI4QXSZH
D9CXzNmmfr5D2YzSYh+qBw6lGLTtUsGFsbEHM4gQnZibC2VoX5uSafWKfsnzSqvY
6Iswcw38VG606w/3BO9/ZA86dfbmbDdq5AD+F4ZMXGlaONy/1xUnE2SB5EjQyMk+
lC6+srBaxFigSa9Ez/1p9YqxyoxXYaaW9YHg8gcEERaZeoOhkfBHo5qBT9zZz/kg
+mpBdqzoEquTHXjVEr8WWaQ8QOXkCciEtLgfyTKu96oASn85aUhDGmytTVwUHKhd
X/enIAX5huFD/55op3iRtYubU+M44CB5KFqN2OVi/VHJK4kIJtR/2MHqKuU1jv3c
M//M4f6pQA+ji4pq8mGpxXrcAq91W5rlF4e2SRJve5K5vu5w5tuDjBE8rl1Co4vh
gT/T0Y8nEFAIJO/TML18sbOzlOmjy7VTzucBYQjmYfw+wRzc0cSzZlirP4qYndnQ
XGCXb9Op5qs5sLccocyxUp/C7p/2Vh8djLgTl1+B4ARck7tnDjfKFHtrzT0AfPRf
oqfso2mo/bvKCXN3IoOhU7g95ne9tYvhacUpvaWoFboqxU0c9SMXV6NMMPGGybR0
0S3A/9UUcus2J9ozvyoh/sh+mW+hg87RwPCH09hFdHrt+lPWBZEB1w4/xkUqWxZt
3548Xs632D3R+XhmWGcsf4RcVjB9d8ecMV0rWVgGV5d0pVXL6pZuS4JzEb/aYsK9
l3DKb0h3nFRfS1ekLgcfm2XFMUo95BoBIJp1xxN6/rwzWer536/lYIAznrIJBL2A
e6IQ5+lhbAvJKNKFdOBwETKFW218u3J9vz1T8yVGQZa0Lf2+VHBsGdgSMCARu3Tq
SHeDA7G7CUM44vj9WNchOoOoHIhsKtH2rP0MwjV/oXGgoeTz+UYMPrc/D98tW2AH
hyalc0mBR/lhlza70ePVLADtqSV+FoViIGr2QydyUwR6cK3RBBg9NL/xRrKmmgml
p9szbfna8LT7Sh+n4suKo8zN0tTHLojbbFPBAYvM0ACyHoXjTxVLlKJo9DZMQA/S
+oWSjgLwiVyGZI/Zhc1xjsPv53KQiHxYCxITaM/3QpWUgANvC3hI3t37ALNO10Rd
mIH7z4tXTHKHIx4bFgVyA2Ked7v3pgUXL7ag11zkEx0QQD3fDxahy5gpBXRFAoca
ye9gi6z9TzDX/xHXOkg958Tq/ZWC3J631hSzB/E4rUvlpUHm2QCOoRSMfpe9mUVg
e1xtzs0cFZPbzsKMXg5c520Jc8sh0Yt+cGoGHU0e9/HNNqpN9iy6PqxGqwvVPw6U
t+cMmV5SUGW9IQzIfDM8+Furtu3gUcEs1pdcx7lGEIEd5/U7gHyEGRXDPMSVEa3r
HACobZFzBgBnH2b4NVRYsiIs3W4+c8CYxSjQfEtJ/z+3ydsVIYfRsvalQTtEHO8A
lMyyO44E93GLww8iJfexI9NhitWcX+jDWEHV+aGi003fujiXPjlewVE9Xf8Jd5kL
dQCSwR2bTg7lWFffo5+nO4j4iKdRE/cye8rPicPEOMYBYJcPr5MllizwjL93U+Hn
QupbAsR+GYvwWwJCjlTFo8cTzeI8ziDXdZuUG90I2DC2vyXmwjXBjEbddCAppk7X
b2foQMjTixS1iJukIKmNAcpRfx1H5CaMtYB0pDjQet48dwIpNZZLsk+6zFzkJo2j
4xfsetnW+7u6zxj1dFD+Ocgr6ExiIPU9bJvi8b2OL9nJ4xFJnyr/PTYAa30zGxD5
uFglZP5I/5gd3KbOP5Em8/8YNj120zGgexeBxV/lu7R3F7O5jWHxp41UYJs/6qrL
8/qAjvSa/ECd6svh0+1a2KmjQIlDkw4Oek8f608wrplDdmiwadHHYlTSiBG965iV
mrnI1jfoD6yx30ytQi1mBc+rh+GCOHMNPEQkF97mcs6hAdoJhmf6SoagNl6n3Zc+
0qm5s8t7buW2mfi9QP5QE04AO0yZH+Pbbb+rpdi0/AZWdzzOs2Pn0ZUrR03iRatV
IB4NEC2S0+zPEVbL+ywYQ2IitwAsKf9L3bFkY/TyaMf2tpJu+qcBfDDoIbCeV5sR
a8kXwlpoZivfOzvtIa1OMGlQWzSkD+4NTCcwnbb315Y1shULn/t0mwB9nNT84plt
1laRRQam3f8hZdwPHygIujKAfIn4+3IdB5sQvxnYDwad5ItPf3cDDIw5JWrqd0EH
P8a4hz0CkQ6x+EZDm0jAc1vtLmqZcIgqs+Uw8BmQgkcrNE6Y4J/xa7hr0fyRnIJI
BnQh0iF8cT+VAGyQYt1VnQyaJrA7LkkaT1Q3ZBNTeBye0htapq0W+HPZ7Eisw4to
9Dlh+lfctRpQg/lvJe0BYnUXRt2C673D2kp9fygewVZQ4UM7Aj/TjiHWCPR24qVH
/LmvCSevjex5gb9piZJc0v/RcGM/Xs+hFTfojy1eMyQZ3thcmd2NJFmKjYfN5A/E
cf1bpKKRg9JhUIM1EZpRloWOhvkEQise+wRdwcUtfckDcL3tMFHr89XfHhkme3qG
UVAtIOtY/hHMh2IloIzs1X7Q0t4wUd/OUdXU826phHzApu9X5g1xnAddIsKDPxzP
+2JmCS95o6BnoytlotDrZC3gwcRhpFtrKxxSWF5FckadVEVniDUqKkIfn42qZjMG
lEcQvJB3/FTVZfNLBZZ3oEDZiQ/WKRTLJpwRyl/SrnrQ+k/fe93EaNCfek4t8xJB
cqeMsthPzwqucm0zZtY1gHpJgagaWpR8uMFLeee8wrqRF4DDIukW4QUDwA85KuEH
cqegna1Ety75Lys19K1ftUHsq9HmmQwQ4pwlxg5dAWO+rhY/P1MTRffaYb+OizO0
xfVBA+UZ8VnoUe386kOQZLUwkgn85u0OJHXZyfZEF/DX1EHcijw/zgRiMlhh7emP
jl9S1w0AP1XjbtxAs7R/Y/hffng7ur4JNe6NzBDqRbYKPHrQNs1+RsR9fYBROPoF
ckFRr7hScnjyXck5RkQG5cI0JrJCKr8kvgkg7XrV4fDWjxA8uw6Fn8x4u4ergQ3L
Yact0A38Vbg++EtwJfrJDMNj3E3Hu44lwT80h4hDPRVm3leb8rLy9yI/KLx9RkPr
Qkcj3+zbOu3O/eSC7zpEbajmKPZoNylazXFIe43a/g5zX21DvgmwwiuvrpEpxaIz
WUW7pgnpfPf3A/DpaYQgZ/NoytcGZ5YSEz8vNOZ3kxXbKou7ShU/iZhXYf2mJBGx
F2S5w21WHFAFuogM+qNi7G3xLBrKy3XeUZvxXVbVdAHJgk48gBjEQQJWtjmR3Z5Q
6BS03udHA5vX5mTeUEaUf8VQZbW2KvrUDWz5F3Pgci6XHTHjPB8yGcuNwZNQMicV
/Dagna+hInrzaXzhf0sMvnXG7u/b3utu+cFuFtEpLoKq7y+nhkj2gvXtp9dtAcG+
uL/tQCl2y7q8CzVTCwUfQ0JHVZhcGb/yTHF3nVOEfjLTkACsWlOlTI/b/R1aHkXH
HyfSZLW06pTHAKIDxZMVbBx3nnhU3UdBsydK6outNd35pZjPdpdYl/7xXVD1xKVX
IO3FMJNqQc34URPLmb6ySwrV6ATG7neL95KKq2cnwHisD8oRW+YQnW0zMCzWlpMp
n3gDDI2og/yuIC1ud536LnBGpRyBlzCbAMiROUp2xYm5UwHeCXJSgQsW2dzaNu26
lddTmjN+N6oO88EPdJaoL4MHvdgHyxGHNdFSAmE4aCGBkjsWBjao/ULmvfOE2npa
+ZDusrJTwLvvCKUxt9Ly2omzYgzBFV+JaHnZ+JFGVaMMQuuja2F9sCk1zZGvFDLr
OKaw86oVDTiAv8W9FgwzIZlPNCUDzTuuN/yX4YN6BvI0VIGYm6il3R9o2RtTYv3R
bAXdpgPoPzbfvZ/JzriZLg==
`pragma protect end_protected
