`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CEZgb1NDx/NWjKoWppnp0qvUwMk+NsF6XCSNi0CNsz5QEYsSz+Gfw3ntEMlVnFkn
NySYiOjcEu1KuuAWqXVwoevNdXy7Ztjo8UGrXjxhUR6bRlpU2fvRWdXaj2zf5OWJ
T5OizcIDZRNyGl9h7jWjHTJiqN05f3OBXm703tJl3bw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16304)
M6nXYjhK0nxas+zYkod5nySd9lr5HXjmixEwz4i96T6t7YotBVTeYr2m4hNgDeFU
CEITYt7PQT2B11WF1P9mMTFBZYwf4aRGpnNk88jlNmGoPKv6B0nBauWxW6AeRH/W
fgCHmnUEwICErfCJ1RkcrPVd38kNgfGJPEytHQRRm+jNfbPn6/d2T2o0H36/Aw9A
wK3QQpMvnCgm31YahWJgc3/6AqEzoUtSlu5HkcSzBXsYy5EaHC2ZDCww3zhZbv17
fhFGI5aEF3vVfAJXjsKlyTDrjhLmKvuKw8rp5iRGspA+SASNqEyNdrd891IWSASP
XA1iaVVMdwnK9i/11DPsvfsnZKvl2LQ3DLqSdpoeO4ZAw4gOErqxKuIHtbRwipEH
nWJ933zIxxs328AP8ZqfOxvyymOxmWIWlSRq1BDIOjXRO33HKIQDHp+MB3UiVTLn
MAQ2K7ZSBe1c6pFdS0DXquPFSUcc2qrkHgtFTReWyWAYZH5h7OlJqYob5AGA/IaM
HOuSyE7Bj6fw5fUJbXD6H7Ui3BhamLc3vpW+3S77F+986bY8kFb2IoQemFe4P5XS
03wJIC8/dqGN3u49KIeE07mUxGGMa9Kim2qJFmPhc9Nbb5u6pWS5Z9vfRjoBUFqv
ujcetsEkDjVQiVhMTfN7MdE8C2o/5duq7F90xYznJjkCiH38q/Znn4L47JOho1Je
l8u/wCQqSdEbgI8yX5p02j/Bj2trQhWBDJuZvhBlQjopRHfP9S+8O4yoLRi+79pt
4JmrJLOs+ivXMcWJfDdeq3pWTPji4ndYnOfAB9Kn+2tLcUqFB2n1vpf5iYi6B2B0
OEhV0TwwPbKWGzfeVe7lzlDW/4ipXSjJE10D933RSG5QVDDT1cVhiC1hylXcYfKq
76Doge29rQMr+lWBmscLI1ewxDUPffx+CIdrQ5L2aYLbSHs5zCIEhnLs5F1VhXLs
49m7O3zYrosDLJczGIYLjRJkEV1sD/pKFpC42+UqPF9Ax5plN6inQSBnruaDOgnA
RW8Pczj3SJixBEboadTRlPjg3yR9Mrtm1EkUYavw73Eaaib+rAYufP7WBFp+DZ2d
1FGZ5Dw9TOJWGZhd1G882jPsLnegA8ESbddwp8HavPGZx6y71+0cKoGxiSdEZF3W
wXS3DXk0Ct0Uegh6y4xaVF1McPHd4l94TYqHrxOG5JEIIXb5TR+tLk6V0t70yPIp
rDmqBvo1ogu9fcuynuBiXObR6/6sQfzECqrv59sngJoAw+HSmkp3GUCqvsbCYbsJ
rN/UVDpY2YFj3iBS1ELWTKiWjnMxRH5aokjzfGKVjgw/aEfuIj1kL5gID3Qn6aLu
OyeanAO5SeSA/jboiMdTZK8ID/NL7wIFxYVOl/1PB10P0KucKeo0kh+o0zqcoeYQ
vsDDFpE1SEmTB2GV2uOtJapM9SiyGx04bvLgiPQXdDiCtzMewQIbIf+t1Ig5LWMU
i3JU6aApmgq6AVq4NqdrbepVop62ziDp0I/OvDxjMMa3/R/Y5ZAsqmi7jVx6tEbo
wtrhwQ5g5NfzJc0J1tLwI7wmLJilPgzoBGvnR7tey5CCmECiv4TCdqY+r9DHjjFP
q2a6Il2vYUPV34fB4mzEszAYvamR6PFTDvav8FikJCMZtbEprGiDPPwMSz0t8zPK
/sVnlzNnp3fNoorpYZCvgy0roVDpa2kigdhRuwD5DIGBFMU6dAasXGjWx5SDDDvI
W1xX7bIOektj95gxVrI3S1HSE3Q1xpydtPyshEJoUX7fA/FkOHTQSQ9REmdRxFoU
+1U6SodPm0oWc5L+W7Y2F1OG44VkGQtSJqVBfgek3vmSDtAVHS8ZDdMt9oLYkcNC
h0ty8JRGoekmxy7jPEVIlfz/mi7381GtxB6simp/qMpCX23xX7atdlDgKcoL8ukq
Ou63O3v4trDyOaw8n+IwwqyAUXRSvptkxuGIu9KaN60BEn0PbQHpKkF0wQKUdhvb
CjeuRsO+zmmNdrDktJ2GxMDlppHdnvaxtxEAWFtQDdoCygYz+wLZt2r8kT3WCnkj
Ly283O1jfy3dsnwOCNMoFP5Tn5CPfpTwkJ2KKtkZsJj1c1P0vRg6nr2lXZD+aYCN
wM5qMYbG/XXJQY1TQqxFyxmK95W3pBKpy+R2CY26MupnHK+eSSArivBJvoPIomR8
3WbUZS7A8RJ6T4w66eWvUQnSnn0paj2QzAqBXMmAEvvSx3laOygzevGhkjTxahZA
QliG+EuZgwI4SJr3vdhhyjYOjVVmc41FVRWWI8AB7JqT5+sgTlFKlAhBubGZ+4j3
GZ/8dNBll4iSMG6frwstyK/f7IpvjUJ0IConJXd0AJDWSq9e+RlrwPzPjU2eKOIs
KA9QB7fyWxdPVSVvJ/i3imDruUexPMfs1jFi+rcV00wRbOKmKRqK4T2e4jCdj7mH
wg9avp273BufOk0TvuHaznTitJ2dZrRodbOYZn8xvA291mVMwPKzOhj9O/gUxymK
5HQCxpES2VM+QWXIHAdcnr+EUIqD/H9QMZillW7uc1sWt7zv8X5hUWLBDE8RwlX3
0/N/m9+y277pjpywk2AXjdswCpCZFCgkIERGjAcOr0dLkkjeJALMnrzZsSRGubUD
XKkMFwhZ8skmS6ddkqKsSKmj/tkBlNWxdOuwZXd1zBQj5YuIoCxevweV5K0RR1UK
Xh8PB8cOj/fwDVgvzSiKC1DvRy+6/4ZgiE6dpMM1p6ucPQxlkSxwjct+rjacvHjN
5pQRUKpzjxWjbDerAPBrrXsMj0ngva1sw0lDpzUkI7MiCk8UtRYhI4eflE0r4qBV
uV3R6n6jbzXR5SLt/MpI3vEPn0T8u5ssTHklz2BBzFO0odK3NAakrsl7DP+yw8Pc
UhCNPhiDQRTIRDWl1BYOBtLM6AG9V72KmLO1fRCdAG2DnHZe9KmepKpkFagYw6KZ
AZncjtjwDyCuPiPZerDoRrCvlwEGLt+EMXFS4BX5+ahQmjSH8U3QRQH6LpQWltu1
ochrFB22IA2Kb85eK7a2YpMIno5kq8VpjZpvvSqiMmWIwzg+EMuD10OougqRnZWH
MJ+2bM6S4oWRhDyQ+88BxRWwvPEErAtJm7VbcskyVUhvH12mO+Vp1JCvnWoDCm5M
PqeGhJ9NNqj+YcpyML1lU8JleoVf2GgPRMxpLTfUEsIPiqgwYBzEg6YWOxas1mI6
EfV5ZQuMxWT2dXRlCTObIQilRc7STnjsLnf5s4oXPBuQ8EHchjF9yf/xgewts2gS
N1VDwummLfgobFY/JmFiHVMI+ePG8jIOqLgmc5Q5SpE+ez/0B+MuXGnG42B9EtBo
DvK1scbY8zEiIoDyHlLh5qiOe7NgQwJceCRGqDPa82EjjBvMAi/wlay3YI2QzlDt
QPi73exYVYeqKDod3A0pVyBoKxqj15Jve9m/U31b7dFA6C44uTC/NSxdXlfjkiO8
eAQSEML6AD0lmifbfCnwhnar4wDWKgB9+DfScd6u4oHOCEhuwYAJGfkzODMXOoiH
OAEVNE401I4mTBD7M5PFaO+CIbDV53ukZmtK3s7NKLsNssSNVFbl0r5EgDZQKMKA
ahTqccXYKoR2PMUK7CQQo6OyDJWOGTfrAPHsq3UB4Ieh86RhbG3Pmz5BxWIqtlZ3
guAAzy/RwEPeKWAPornO6XBhMfzRakH+jXODln9wedz8DhpfTwtu2GkOmjXJ3vew
kO0h5kuJ3IabGHbHPSvE6H0mfj7ZGBpSwcvxN8L3YCVODEvqJodp2b6Mq5ssRYoC
b+BkEAXyu2Tu1/bXDN9J3u8iiwgxmjILessSyyKnRAk1j3a8r/d6YK1utbguCFqD
OwD4iUvdwObWquT7/RghmRPym0kYx3VyXop6dseguVZ5eU9X5hde4/N6FNwzsffZ
6w6S9+CwnNlDw+CoqJ8rjXxKXwVRt85HiC8PHv7mf2frNRJ/4hBoJCRGhikNrYpb
zqCiKs40pbHwcFiKyLdqHvSdzxsGluWlA+O3cW05FD+4EBNCfse36PaOs0AyV+G3
E14fiCESVPNsnvgMPFPaXHL4fcZ/9j3FSfnxxf4R6hv7PjGOu7hz9/pSXj9x2H25
3wusLgG1cDBYadN1Pwx3qerv3YmUdri06MB8ci2KI7S1igedwouufCrcrAkm+kpg
FvlDaQDcPQUq5H7SAy0J2UTdGyABxxUFIlDESCPsCF9rWIkS8NwDDk2aDggpELXZ
8wQ2bcKqXHYar+ElHx7WwOmHGzTLULXQGmS785NiFLj9suV/0TrEpAK60bV9so1g
dGNmHZJEX4EO7XNikEbbjzUJrAd9mB21YQ4ZvhXwDI3WF1SN+upF/CXcHXkriBcN
xHjcys59XZcqUGp0fACodstfOWWttugBd/IXT/AsohNH5dEjYufUYh99/dqdvzfa
kEZqgKsoYtVIxEvOuEkBmxz1nvHKxP5iltLHrshFnpyDAedE9+R6vADzW0jp2le/
OgBtjObvasIc7PeLvahnzUYUg7O7m9k1sbLdqWtooPMv51oE3spBCTi/5TMtECMI
+ReUBlelyfQOa7xm7UVFI4Z0oai9n/gfAtYle4I14lr+2zE+92jMIM5eBM4Pvmyz
Dj69afqY0lTYCAuMZ0UrKBXYBMmxcV7ZmTV6zbGV4BvQmxCjB/d6TB8uvywAB8OR
HOREZ7SGtJRr3XBnijUNtaJRzjBaIehkL2GgLzVg0qq8+qajtcrTgmOSrcwoq+Ov
7WJBe/5OCSpCs3+TSWLChjkCENpXbNIbxdNF85AaBXNHy0KS1G3Y9X9/321vRsSg
jyAE6iNt+W2L12W4wBq1Z2edJlJcbvPV9yiTHXx+QFAO9mE8BDLRMRYXPb/67kF7
5do5NbaeLfbd0doINQL4G1BdzhT5xP38OYE1dF/QZNak99TJuNvvSOJMgbTW8nir
HBqIzgOWDQJOfarHSUU/GHB6TwiNJYSC8D8VW8Qm/XSb2jxmk29VnQ6MIPjr0xap
i9m/+bin5HexicJ+lQ0lS0oOZRwr1wVgDQlLkAdd7MK5OFcBCMX9KuIGvuvTPdmz
fmv/ch3x6pJETxU4tl/adWXVjUwk0tG36abu1vkGd7ps1vk3ZcWqFgoey87Kv0s0
0iZFTaxy1FB0BCbAkO04GIJg0+ZadTXHam/LWnLz+W28CoJl/XB2x+A3awOMc3gu
v0wl5c2uxFGzJMbliqFQXM9SePVyoTpBQPdgf9EKpmCXtSzHnb5SgybFQcmgvP4t
6NRusNEh74c8fW6h6aw9Yc9jcJ+n6KFD77muquQ9WD2a+kl2vuc4wjLA1krlQKxe
DiG+fpsMfQ5XdPf8jEW5rdBGVOH2HnC5iUHbPtgjY3DxKma7Y78adXhNwdSM2PNG
9HZvwYyTaDbNnNcqJn06auqDNEV9pXaegYTf1+fRQlvMaBnK8aKPtAcyCh1+MBh0
bXLxCf3cFoqnRde9WgoaDBCpf8OBsXsfs2oINtDgezPUDhBd5x68S1oDtlNrm6y6
it0SurRuL9++/XzQq/QGpA5OBOf3d0YLF/pbaQlWdVhJqPd8bKJqP1sGphGzElHL
TESlFF++Eel63HIPRkt0kEcTJLqJUvXUroqihTuSabopAoXZHuuj3EZqPkr61NuF
g+1saykr8tTA0jHpBuDggApGpA42SJr7lkaDrpJzuH+G9kN+lWogBGeseIeAIotm
C8eQS/CS5lTyVyss+5cePI8iYO4nMI9Xfk774+xSsq8cPebQlURUUpcJyK4NKiQT
6CS5EfzfR4xMuTKHHY0SbL9MsduR3OlBRbrg2gVvJmG4ELQQS5WiLgxQiPBVzVfu
4buomVV2zCWXeYn6fEfaUg9y6UT/G+/fzB5h4+Cs6rt/MmbJYo6yIyzpdLCYHYha
Z4r2eHolQ688MTzarzmYKDQ4drHm2XW9tH3/F4WKfrdkUDNJtt24t40pFz0RWAQD
2tz0S8nHvNaiWLB3ouSUr9EP+Adf/I5tU4EZkvkZY+8MjA3GWwrcGaBo1TmhS2An
i8DlxsPFEXY2hBd0EIJq2tZLTxIVamsNEpKibihuiSvFcEoS5Bq+xFrOhZte4l1e
VJL1C9WusAcqeVfNHm4ADrsYTowICdkNWubbJZbSiEtHBSuWqAWfz/ABwyt/YJ8Q
RNCvvfx7nd+mcbm2ovpVrNiA1DiMeZ1GQto4wP+7qQohd8BLr19TN0KM3HDTjhHx
9Iu2hZCbTSBCswef8tQ+xpZkrH3lBbFmI1wbdQvdGzUvfL7Jv30F3LLO/vSJ7tiv
88froWUnidBHNnPUtr07eDpxvuyL8UcIaW9Me73RwaBOiLo6zBkW3aKXaNczgaA/
GZCkbCiNTcTykmb45NJRqa8jszZKxHJS9jAJHfD89Nyr9waokJ/xt+hGQ1k87iQ+
JNVANN0KeiS+5PT5gfWTVmikH1BixFRhA1NxGWloztKCFD65qyKsrryotSQXsiU9
XOgLVIseOlmWGNWyu+H80w7NWmFZ8N2lP8TV5TTHTkUfUr17ZUgNlyjk3eOAbNDL
YThKlulr5Zrs5gGpx9wUvxznyHN3i2DxextEeIkhK4hgiUI4P16Mee8by6t/RhF4
AnXJNmXfhFonbbz7boPW7ehmExT2e2FMzWVxIta9NFGuQdzzQcy56TBbi0hBbGTr
TigfBr8NtOMDe4NYCAOzXAd4R6GNhjNGJz1YbTO5olQS60z7n7kzaxLyr02MSua0
ie/I6r4RaMF1x+JpnFVoYlgJwKCLrtqgt4gn3sxSU8UNJddoEj1BbFiG/hM0ZR7A
/4hZVyTbwjf84IKTnZubxdU9HIHJ6TNkvPaatHtWKXOBPPV9AV7AoKQmlJul059s
VY1JKsxz7nuOfGh8iIzOoaihdKwwV/youitkqnlPg8iDUWmIQK/VriTTJxQWm32m
JG/D5R5HkQ8nkIt7n4/ED48xrdBIjT4mi8F4JXm/C9AvKFO5t9nA7SfbQSfgXDB8
VNl0PBdSI2RSnlCLdNuSvOQIow3rTd1iECKUxotdlh+b3+sK3o370ya65YjwYFZw
/Kx2o/T3UXNxYHSRmfGplneIm2oqFJIo9JeLTnnEuZzx/Lh+S9bo0OC4QBXTwtp+
NHwSC6Oq/WXV2lUTu8BO+MGtvR9YjJ3y5tbiNjQrDLLDyvMMrnlBYec2MWGVYwjV
GFjV1lHABzB41WfeyG5ZO40F2OB9CCiqUofRnDggZN3vP9/zb/0voG66U1SK1+bM
zXj/DJaNrLiOFvezQUDFxPgcjk4X1ohpKWxKYeKoEfshgqp70HES371q9yQMbgSL
gEWL1BiiMOjFoQDzs4nDnAnhkVG508G8PQkd+A87bQYfuauredFogAj8ywZbKoXC
CrCVeXJzQtKs+Na69Bl5+6KzkRs7bCe1GdPFqYIuwk0RRsWxiovnsdchu0NgYvJJ
OKF7pNCsrCryZC7l6B7JuWQSLCCfHNkgA/6o8bpBad7ibh8y+4L37BcX/2bB4TR/
0e1YOY2tdN3vYl6n36bijxkFJpqabfMmaQqbwXlYlEIEBhAS70K40FN+suYz4OIV
nz/Sct4yh5b1q+AnPV2Ue2IuW6gYiNQC18bOy0dm7wlSRgvekssTqGkwFsDYBEmI
lcYOI5oAxeFjiUQabCDMaIpu7UZGkwgrxrbiA9oP5yGUBk0zyfwmzYfJJxjsNArc
S/dhhe4zVpzbAqmGp7pYVTHBQxnhEOnCqqRKWdqBlTNjPyFpux9y3bljSNMXdpBY
BHUQcJ0E3yLgntBLJleeA4WqxjM3Jpg7VDvC8+JplBIpyvOTSRxwhrHiZmItEntT
CMrcQ45kqyLB0U7CN6nw/91UDRA7j5Ajs7s9ozIDmVRm4bm0KvTIWA4QFRG2yWsF
89oPTbWQlJlqDCbqSIATYXXKx1/MrDDXkEmSiEPDAqV4cUXxUsbB5/T+tuw93X8r
RQ6gDzstHgCLXvWM79Kc8LJ6R5rMA3P8nrb44OIKot3L3kDOxDNdUhLyVppwC8Gx
gtqpjtVL4tI4HOkxILRUvZkB53RuGI88PWx2Gmb6eZ6Gw+d4gLHSha0k1mXv0OVE
h8lcbIqSwF7dACg5pAx/OAPP4Ta92rPNOV0tFMgx9AulrJH5aAPmk2+GFhMm3Vw6
Wxy1fFB7uS2dXN2yidFxRA5PGItENrU1PZzriVJrF3Wa3m7PTkKnYPlrlkXLXmq3
hsAhrHRYNo6r+ktv/trrMYI3CjxncwDEPyAW/7GBxD/u3CbliI/gpNWbTEUc9EMy
qJ09UIT8t2ZisMHswgWTEaIVC1iBXT0ZKi1lR1gzgzLQxAbfR16yurEUAUB3HHrq
GV5mu5PzAvn9OWr/vLuUi8BYyOHfBGVStA/BDIerm/sxuVLOPqyujsh7srmGzlz5
XOBaxFBjCM24IgxrZVDeF8DAjqMi8X2ipA6sHP3KDU/FVDsO6vpLCE2jnFX7HUJV
gIQ5bGyk9cd5EI+3FPcQ+VMnFzt28Hrs/SJ/gzviL57+IOiCd1A02PiHCBP68NMu
mjMTX8b13xVm0md67byTxHEzc17alqDPfpxqckB46FkC2Ci6/5xQIH65As/NYrJT
9KM1hXz1cKnsVr/97QA+qKtRCtLzG0CdYfiZktR1mzGAnRDk+WVeFzk7r9ebh53g
X8m+izFOKWk3nxA8fDg/wmGEQ31scE46KpMfc5qCA9CUfSYd7C3tGe7NogC6U1iv
j76VNuGzGA0EpHLC09s0uNoMTZVtCvd3a16pfojxdTfK2fGt8G3zqi2IWabfYL2S
uEWSp8dnXzpBnNSfIddO85yOjiJCYXm1JP4Gdn0mog8/aiGzkBGYJxjKo2DMDZIF
jbyzS1Ft/LBKn3WB8uw4YbjZzG/DGFv4I4ZDTYBqTeo2IJwRRUv43rfG7Bq7CoOb
S9AE1Des51oX38XAkjYfoE0N7KqXFP3Gy3eOa7ywsMnGmKJWURPwgwG7MawmbIHb
eOSr40oT6qzHU745TD1hRE3cT05qt+srkBG3VVhYXQgKHxxTc+ewA5gbSBpAndRo
KZsHQX+pKK6/JANxQL1quIUZSd1XaZ/n+h78TeDK6kiqvOZXYu8qY9GL9BhWONNc
OVY6AowQxCr94bLA2uUDRw5F5uq1O1DLNUVHjBZXq8yDRNaam/fA/JV9yNzfG9+e
YIwDgD1NyCSMWi5J4ieWhEbgSX4CWwZpuCgXqlxSsM6b64kgubgfrYw2vSkQ4jcQ
P6j2LY0gCc/q6VBuL1iIwh2mt7TNypKIGZONJro8qDinMtNNJxjqXVoBGsB6bfxA
auZFqfUfh92QMTN3xxm9h/HEfk7Gb5EYV4NAoRBpu6j2PiR8WJ6DdQCgXKxPzn8H
VgVkIuU/atvTdxJ3y9/rgiXcUaAofjvFCEmnr66NQatB4/e/XWFLKjk8PlVBmw0E
SvlchhGWiU1JJLzzya23rbAwpyhLMAqgGljpBurRPkMfd50z0QnbCS1ma9ot6W5I
oGjhnoXSissdGNF74Gj5WN8UKJi8PulXgIOQvFkdTr39tXQrRWhyASoWjrYDp/RI
A54TrDqo9ZNmN2LbaTVm9L0Z69BzD4nqvf7w/bIC3ehnzOJrkXNfy0JKc6Sqd77t
d9rLAM8AD/yPnY6T38MUtaDPDLof4GD6jJhRu0CWYTyt5WVRzQSvKJTCLcRLOAwj
671G+VF8vDFEaeajW0bHmiKWAURNOuZijsE3dRuf0q6mRBAZ6pocpHUyCr1PBvir
kqsSwBo4VZvcLYpMdzj9af4k2Se3XCSkHViRoP42kTb4fE2wgonYnCd71zt4w1UL
kJAjmg9SOzcjXhRD9yOBjPPAS2SKAC8i17oZ16diTIyEBslA4tMWQkX/auKQODOg
Tu4E6id1zrmN+GaU1gEmuwVkNeFre72hbpOSDb+n56lMbVM0BUafi/Nbi5KrZur1
X8WNLAKTF2Q1uxCSX5fHTJWPRSa6P58fzqUv64wzHmMc7vMaefdH0iLhOxzWWGic
KZMqIkF/pQOiU8+LRJfszbF89F/cXSGAkOZqwqnfwKRI8gbqSdh1w/K3lDSjgWnb
Z7krl3leS8xg/HYJaBKZLzTRszY9PUvufGH/0grf/Q71Y7PrpYhNOKDr6eNc0YO5
lajMiDUKEIpi5CMyZ6/zecqjSPNchivOCa3CXQAZ1R7vttpE0zu1GtTGcEo3OP76
2tyTccrq8H4Lrepb0Fcg8Wcnr8m/w5fiqWQH3KXwlirMeGVdiaSjBJ+khLVvUJc/
qa26TirBdnNhO1mCaFajWbYCAIqbHHSMJPifTGr2Y5bkWA2FsLbrvdzhElJssJ/I
Dr+lA2/2LmBQVCW0P4orlOKX6SBKnIw6hHeRvadBwWHcL2Te0Afko9Tv7+fUpPnk
c9/k0IJifNMBVyrQR2YBD1sS++Ng67pmUxGC2fY48R3WN5x/2e4MTJCGYvV5LndO
uIiG8FMQKU2eJEvFv7lVcdzQVjZBg7UVhZ5QK1BvNZPJaM1b/fGD7GIhRtJImpX6
xbslbhP+0NQlmb7AQ94gO9gVux40aK7F88SE5TKQXaRwvnZqHcsGBYo9Rs/ql0ca
8MO1ew6pSIYWKCAzwhBuCPdL0bRFmxcoTLnGoet/IcPhSl+koqFpN0Xi2x7p+LsN
rh3DaWnmijSvVzsyO3ganGJ4a+fHZtRq8Jfjk3ZFOFBF/mVfKyv21GuK90MmV4uE
fSLiMyVyPUOsoxh9Q+GvlmrwYO3Dz5gtADN/YOHQP+A2K5rLpfeweK2ZiWoOE9pn
mhPhcR2ERvjPE8KeHqB1G7wKTt+uoOrq0v2rXKsWi6mztqlW35T6GAzadHrkxqTK
A33xNdfcqfcNkv/22FqK4cUjYl50sC6RIowu7qBJSqedzsdZgVDfKeb+090UrTmi
kRTLvabJ1kzWb+wkgVZZYXWn1mL4EdM3hwCN3n23yhtSHsrAbY1S5PBCRe00rbh0
c4l+efyl7bmo/pZ4ihBqfx/j0m7qFaW4W3GF4tPIZvF9GGHiQ3w8Oo+/DRRA7peR
DXhTBOxYMu5Hub9pgdQ3kc8X4qkAoDKTyqrA7iuVnw9M6I0OxaoCxVDX0zMRisQ1
Vy32PgNlzBbrOBG3NZZdIB3SNXpoDi5fIZ3s0PlkM29niCT+5jA/Bf8hiIxzwpc4
qZ6nggPgce8CBWiUhy/gl82kC6eSDF4num8rb2fKZrGsNjyhcW6Dz9cX9twpsqHx
UQdsySrQRfbfk1AVHQWOOSOVMg3cyTn8R7v5ToRBA+K0Lwis+aE0QIq+rOR7gOrj
izWVrfineTLHdo0Zp6xUGu854zk/KuiDbjlwT9D5QIbBvars5YzjcgD02UGygObv
0ZeEbFMEQRvSf7HNJIHfnE6/c0v/QyD/kAOBVUL+0G835xGuG4GxoD3uP9jv/NYk
Ym0MU4UcNfnd8n5e3M4GM/SjBVOafPPIHC19eDu8O+ph1ImG4p3d3Fw0WpDbtJJl
OVkXWTXTzDzSsiktiAd+unNLhCxMwFQhv0tyqDretROjXgyEOiRzLmp2ixGAfPOo
E25v3+3ucjj7kyapCaTVXjuTobBUhgQCizH015kB0NNU+KdVcBO2qMX6MqWarJFY
WeRJRDWMFLheWxTDr6sE7DOmL9HIlGFDRQGthy/so5TvDD5ii4rmNh7PwzHwhhfR
0OHdCpn6vHMQ0iwuT2fwv9GYjCisinjpas8/r7VoHpphvBi94M6sdH1SQRwCr2Gn
dijBNmc+cPAwocWHZUxSLaxQ5Cv7xqAhrFd8UumR370gefGSYOAA/DF9ZUrYBL9L
nTjry4ZJfVOrWXRGopJvQpTvw+JNhufEFXDpSc32M1/fdALWP7mw3LsjPQtnUrjr
ljS9pC/rCwMMi+VOMsuk89tmK8a1Q16Xe0mu1nsUJP8E5wf2W2vjw7ju4Q1dkHwY
n8T4GfcSTa66jY7lsc+QK2iaqMFLzJy0K6NZ34rYAGBUTqI+RArrySg5OCa4cXKD
dv1v2rw98CiSvlZ34tIa3N2Oh4Jhq7fWpWP36rREVb4ZlCl4ELDtsXimsTqVoyTM
pf7PrhTZyGeIS8fnacmDPJIi+m8W1EWzfO7su0Ph5DDXRDaujjBiJYwAP4B1+bVn
W8vh9OD7JlNqVH6GN6aoWdfKKSL/wDjjn5hIxl0q1iAjPrmNIw5EwwTee4jUUmCe
7V9f5LIezV86CoCsbrdGJ5o2sSfivRzxLTBnj2ZNH1Iy/8mBpg7POVavx5r8Iz1R
npAW5Vo0cL5tDnUV2jTfbYulHU1yWt2ZReM4hAfltxt/4pqnhQvf6sAXL38ueXZo
ImRQIgdLdpwjYLHu5Wb6CUGrvCCr8O9Y+XWO3hXzHVo2LL18Ui2xbj9MjGc7bfo+
3EdmTTx85l4lzNfllA57qhw6qbRfGllkXDWApPJrRiXZ54iqqsHzKGHG8C0vbSwa
KOdHED20V5EBMqtEou1sMUkF0KByK0Xz5xexF1pcsCwIsNLoZ3F79M9gDwXGPATr
UYWdftbhJl+Wr0M38QiCXHfMAVb2j7Vv7gpG0wHDC3NzhjI58EonKNhIpbfJUkdW
1xJjjzpwVjsNtu7oF7CLr2U7tIQ6kZ2R8k33r702IAdTnF1qAuTYirnQU9+zzJJb
M5sL58uZBYrhlpyJxoqqZ4TCMOpIce7iVkc7qQVSEolYYQEcFDMX2M7ZLB0zxFQ9
GWTFFfTCu26iNxSbf2Bd09/3LFU6EB/OQDW32ajjwP1NkXHqGDUZ1VF4H2NqLQ12
SN1XNIl0RbkBaDAgQK/0ux+GrUre11nB5HEWrzBXJ04NpTAAIEz4NWqRQlXSwCuN
bWvDCkq7MCTNOGuYOiENvHZwoFus+kcrSOsmnnyDmmupqi7LYAr9DWdqd8Po7aV/
bXCsWBEf/amUi/y8Pa/nfn+iANIm9D6RFpGYv5CEsSjSMuppYMFGcz7Sx47/ARhj
e6v/wQr1om2Nh7Df/pffgO9k1aUGTUEJAITRl9ZWkndPhwH07K/TAJdCapzg52De
05M3MkrmoeXuoZWHaF/9xPysiTXIQFLVeJT6blYS3rwQ3W5pJOlgUVrAUeyrsMj0
hg77EgWI7A6kS7JsxFjwG42oIk44V25pP5N43J4x2uX2JtvYD2rlDTewCGQsUShW
klQ6SRyEBhA+vRJWzn7jMi61W+YLGVJFcUD63/vn1LAqp/C6CHpuTCJlcT3OFbpa
HgBNsCS2lDtkynWyQCsnA3BVT9fDz1tm2vng2Icws687yNpyQqdh4wOBpJnb1usK
8uvLTiARQ5Mu3mh63USIFDXKiSQYWUcnYfC7LDZKYNKG7/jE8h0ZOnv3UhtnTb9r
jdkti+q8vGBOGNpxSRhh6Mk02xiapQOo41b3UVQNeShEri870rLyRoWjLLWqcHg1
BC0fJdPiKOJD2WEvpwUJDwJ/f9KD4zyeYWj++/PZkGAa1OFax8vjpVNJKUT8VNG9
ZO33iZUzP0auzBJE6UyxzC3s7R0+z+Oi4mxnbpv6En8bUG+E8bH+u1J0OAKEOVvb
+XldypNDRD6KGmh4vyvkLC0lEON8Bf/lfBfwo3CqnzFfKrkxMcMnMs0SNQ823kz2
UorBXt8FDfbyBOOUMnWWshYCyzQH3YL6LGd2aJScDzkaBUkzrokNev0NO/DB2/Tz
jgkMIkSSKJ74Vp/7s6KHE3s+/uqiscwOKVxO/bQY7onDxiDpKZQALxb/tOsbv68F
5wiXzoedzxSYVxe6nFXacjUn4qBCVs3SnOtvai6ydxSq2plDszl7riNEPkeCBrbY
1fQs6EhoUXcBsjH07QYTzJTaucuBTE+2LPfLL5l3+xtsNLmtz/28Xml9mviJbbLu
lsjIUiE/ULnWt0CHial3eovvBI/EEZHWZWmrBzdJwMnI6j4r2HYN9nsnx0bKbUmD
xb1dF2EfhRVr/dc4VXOwX1aJBfmRX/VyhIfADDvgHuKmvfTPtaM1f9gXyiv9/YwT
H7iIIhe3VD8j1vbqDMNE8k5Fza4tHe4vHxclbTJ+xnLhJLIyKeXDKFj+8HCHo/J1
mwzZtR3Qv3SX5wUTMm+bkBm/IOmvwxQQokXuNQLejrJkkaVQWx2lnS3USTGTxOgX
Jmo9YLvSDz3RwvznMj7dzkNifOMNwIaPJOjxqx+cg28OvVd4/tHUXpNLMj6lSLp4
brrZuNXbkOXX3XByH6gVWbWIRX1u6DUDQt/hkiCioenfbVUL1V5wFRl6g/6jVqgj
SZnHRpKcR1lg09qlx1bGkL2/36r9PpPYmAiykVmmVurr76czDuHPf23jWNnRBdpY
8Wg+p5tG2lc+e6ltS2TeiVuYXk7bLdEaDGDVmDbVjWfewO79JmuusBglVGFCqXo1
7LsBBvCRkeslsQ9KMaQX885Se2h5VKiUwAWwFFe2vRzYJCMxMxNGHIw8eARZa5QI
IUvXe3VhbqdNSSQMcEtoq/1p7b4eDxmhBY7cEfs5f7ZXvkGEfEWo5UpXilUZ0r/d
gxdGFJLm3WqYM5YYrzUoLYvOB8nmUXwv9aMj3hATaGinT2hovqI+6CFDq2CqbRHa
hfEHHIkL8wvM1XVt2LLqVxolSmm+L2O+RCSJkf1aDMOgP0+E/Sn7XhGzJZowh3zS
7Rd5D5EIe62FdU3qef+tHBqAoqjLDLA4TpBT4GoPL8z5DqFWSnv3ejas3O/zX4rw
l1oG4F9gDrCre1jgEuENwdfupNVcWVe40eppsVrmBtMchkQQQHL5F5TB10T95nKB
IXpQK4X8c0aj4yE9av95DPOmEQ7qMsFttgkzPCngUkubsF8GceZvhgqGPzIKhumo
hvPC7IS/aygtuMPdP2PyIosdVe3XOrMH3jcUz1gg5iEAXK4FDPJX6DHkkdvA25/l
IFUS/aDWSiH64ry/rFDTYMFezhFt1fWcEs+JO9wTTHNCUQhKi9EUpSjsQMvrckJn
uSWqF3gM47WrhSXWaRQnIT7Agq3BVNe63I9w0kpnPY6eR3XNnhbAAWt95z7Znign
oSI4Tu5uazDGYac15A7CvGi3wuFJnfmTd5jsRis0ysE2RUCwG1bUI0B0ufdZKzw+
p+4wpU4v2mQcE6wSJ+hbNvj95fzYaUvwNOgpahAUdCftfv+lJtaOAQEQrLS3aJS3
DeV31LmCjbN78yDp2sUOKvv+k06mKttCZvaqKZZidorOoPVNncV/o04DhSIbjcH0
PhBxN6V8rJSQjNR5CPXgOUfWjPP5kbNuc2weZIF/KnAK8Oe6/wm3yFGhxevOYLEW
+9OxBVI5osDDCpilsohZ3LSIEjgGcbxWnD8uRAWDQo14LXgZD6fblCijFqGLxX7R
rZQSllyh+7LsUwnk24uRGk0uZoWihzIkvzQ/tSgiD343sG9YdcLrMmM3wvNQw3we
DoE92UQooEQmmNEH4ffHBumEJTd9FyzpY14rx/BB9o2d8BkZg9tw99asckHuvySM
5j3B0dp9+c31LvdYpxv3yKVEhGxslNuaNg2IYjcMz70wSLA51BG3gnMdLw0BpUZT
qD1NNTodddPDwIhe1M2LQVfM8gaH08SuzfzBXpmdYDmffQyLiwnb6r1I9rlBZ71q
xmoZvbZCGbN4BPNMp0uQLTdKOwBP5hvYnzYT4u6asyghyeMCsVzte+EqSMHOSiAF
GOKmJZjCl9vSaiVWIZsDhXitQBOUW9vw7aRRrNsPemExYUYmwX9BDUb6R/11K/RY
gJbV8r/c+4q96FUeUZLb/ooE82DcEG6f5zQB1N0vn44Hf2fdlyvhYWgORDnYHgkL
2jFAHRobSfhXMhBsVjdfPUWG3dSHdc+6Q2Aa9p9EJ+luFIVQlQjc64/BD8WwsYQz
EWloEshaUsM8jXYtBgiNvYLI0VfyRa+19Z2SQQ1i7o2jRKn9x8w77RWsLqFdh5t8
uwATJFA93OPKHoKTwbAM/puFHVefovzxlyPfoDlHgatktdaqgtDV8V49OWGS7xV3
QKtiWm/B96vpdlaDniIcVyVF870CdMCqAEbxgVBFz6awm89SCPlpvxwXHghLrQSe
R535XISO42ZDgk4P/J9J4T+XoMo3nY/DFkZO5zTW8nxCUmcX4YnFAK+86WQtC34Z
WXHED/tn3WbD8c1X+mNSiXmhtPZvyRGZezzJHBjQBWW/PequS9F9IdTa5cSsb6+2
MxKpkTqmBFbZ8t5drkYB04Z+Bm812ISzmu33e3aDoiFYnpzlwuw9NK844+wWhhQh
KeZBozbsgDd+VljKOpNN0keXDhAwdEcFz33OTPYqYwaA1vsTyAXuepEd97/YxdqF
3SAjBuFu4vmfnbQkxUG7ECY9iuyMztb7Zm98U/tCjsGDO4GB7esrAL7nDLBCVw4d
5kFo6YztRFK3rx7NlMoeHjugq856t0tiZ02d5E2mogPIwVSs2a+UZJYiIhSHHZFI
VWvyW5lEMdJLiOOZnHSV/3WchwV88Udx0ZYoh+6ub3ey5GzlSxJtAugtCfSF5Vnn
1zd/dQBOwW/TjmDdCfxiGcXdR+9rdnsowcD1F02dhiZPJOREBPhAime6OVzWytHf
sriA3PSr4yQcK2LWP269zSUiupLOb2TFm/LfcKcQp7sMjKuCe62cO2wd23Ij4kRx
2IPbLhgg9rPf2kNwi1dhL2vUafgJfSenfXVZitEQ4G95vpSauYl/NGT4Rs/PP2oe
znu11Frq1KNsOA9PEbtl05KtrliogWGLN/zW3dPmY4wTFlpEgrlBxM+pVB0kNEua
HVYQHDVjydJMUwqYSCSHEIT06FklMN4BwokQNndhO520uQBaiq8NTRLNnrRAtfkC
zXoLV5QJzDned0EyjQvi+KW0VNpuzo7Im1Pnpf9EpMbPXxRW6Ouzn2p2WRMPTXI+
5h7hrvb5mIds2fJXXv7e5Gx0/d0248ZfH5d4cDc6sJpfpVXeqtK/nHchziTmlbLc
yCQtsrm9VivwiBckA8d21uR4BXe7m+UBTpPrio47QJLdlyCyPbStQ/3iTBLj3nFI
M2ruCkH9MV+mkIqSngFbtvnKcR7tyCCK2MuSspamZ/RSvaXdHf/mJ561ktO687B5
LMFktddiDzLQQ1RhBz5HQfwmIGTgNh6dvEV1fw6OL+0P5tIcF8b7BGJ/tLQ0/ca2
yJyXL1BKV5nxbbEZgjZRPqP4C1zoG8QgMswGmsgRDQ4DRdqwJVWmsedHStiEuJqP
KjV50FBPh1d2UTu+1tCTBzqUsxr5HpARMBYfWtEZX9WYosSdz+QoCoDdZhTsihVD
wPvVd7lQmzXNAE+8BfS0fb8ntzxtpZdJhtrKbXbM/TVrgzWlb4c0G+4dXc/uUHB/
WNFe4uEsWEreswk1uzUROPchJ8MzYbAIwvzTKW+FrJxD0NyFLwqkOW6QEZHjWApW
3lVKTUfaw1mKXHdl9Kv6SH8zWcvmQY7Fh6zSTVoWPV+dhnKxwTO9GJCmGEgGDzQm
8PYjbdnxiJWg5RPWDuBM4fNjCoroDmC6tXIPVi3f1ENoKrCWLG9WfljA+mo/3wxF
BE73N0Ml/GMhTSQ3p65Wdhb4FQFJv3ody+xuv2QhRdfF1dDBmrY/REz5HUJprhwh
JPzQtZ0b7CCPH6d04gskU3dWKdmJlTM/YhIdTHD2DWF3lJWwquDfmJQwL2R+kSI+
pir4VKqYvnshYz7w8a8frDgBNwIDMHm9RkxLr/tjvC28H3TdvErnw78JFspweC/N
tlP5riD6ujchCRNf1RXkWLNrjKFRhgX2PLBf7KzIqJrVIvAcBFJ+Xehe1jC/7NJR
aoCN61x9nIYQ+dgd+pwxm7bcEoEZ5JeSFPPx08JGuOERUY/Fh3hIdMxPwD269753
IJ+tX97EDprXkF8fZX6Q91NgaobWtzJMHU853doJJlDV1jvY+sxREkVcjFTZ5062
x9vFPujaLXgJSUBpS3JfAsy2TOYQ+Da+oVXCZqlQlRywriD3fc5ddfbgzHgB8DCG
BwqxTuLjNFJmPwKQFg6ijeC9GOVkXF3L7CMEF+8hFUXzd6ZKgHVZXIrdEgS9Jr1o
ysUtHYe3TzR9agj7XZEaDO6830wUFiEoULKAYOln5NGY7tSnfnddzy83/klwwZlM
rgU4w/1vrQUR0+FLwfGCIKWBFV0hWIlay7Q+bxUUOEb1v6/buGOIJs2X6be8D9vn
tzhbDNbyz+Ut9vWxnfHQ+01T3XS9bL3wwF0pYmv5zqirflMrR3z3Gq7LYyAhctRy
i+phi88CRuB3dwu0RtQ0C84CmRvCKnhlesgJHDqDiL/8C7T7eNMqGmbL/wGCUCpZ
7aN8HGO7QtZ957WIuttokD2U5DJ8aOovSVhf42WJVW6DHj9GQlDeaPDwXAFlqMln
pppEU4q0ZO0O+WvhCqPZM7PPQ57qFX9IQnfR+8uDhw3ZT283Ag0tfVczcbCY/xOX
Z40zeXG4Hr09KTKJlTCIckRREbBfLyBM6+NDuRga68KgoDmRYT2C+wrXPdK/xd2X
Yl4v/6Wu935FpyFW35QLzm+/28u/K9Tos6fc5gUAc2lO7JHtVxPqw6p22atV47j2
z86DKCueERXkwvjC9PJIxy+B72qvNGuDvCV0JF2bpuviiykG/jKw3Y+TI+vUht5Y
/S8rbnpbqbNflwaHDUNm6yTsmK56NpWZ2JN3eoLGtVKo4BOx8xBKlHAmurUJP54j
hIzPJimH4qOZh7K9TwQWqwMHFV27HedWTNQBuYb4rkIgFgwg6f92khszQS7VnOCN
yexSaSOC6eQaIgykxfBDUB0DbfL6wjLyrYOddcMblB17gtK34aHYqZWrgRDZwP2V
zIp/oIJ3e5W6zXgaf/xxuDwKC8AlOwJMVMenTfET+LpxVQ4PNVwVBiDbucYBDu57
pWs50H8eOUUvTDzngg/rSIxz0St5B0L39Mfe4Bo1XzWPapJikd/Ur1E2zD1nR3YU
Ls6NeSKYtgsVCeq9F04GbUw/Et5KHWaA8XubdbpRr01cHW3nz34D3S6DT6n6/0kH
xRCmcLtmiAKSR98nwxFqebHc3cLv/aPUZiEg0+FiU8aM9EiGn4PlGeBlaCjqgm9A
F+ibF0t3cOe6l2HsRwFJhDVkmJbnYPI3a8cv4tQro9KLJ1NCmbxlzUBLMoVtezjd
2R1+3WA9ZjEw6WvbgWuYfgqML5IM8iCq+Ufw4c07eQtLJ+6TAW7RXF0HBQPKZJGG
aQJswkeidPOyscuTpZVi8nfNlhEvTjiBaPYxMxr2wwAxdrEy6uS2rl6Lb2UCtmS6
qXsspPFI9nISPzQMU7lhOtAJlcvVSHQauJOHsmwTbZDSLJp5xS1XbF5bNRos2ZJS
eREsxrW/059WfDVNk+sPu2LSVk3I4CpN8uVbcVBTPP6m7M3RO4h29FYby6z9irxp
qHtVlaxZhs43Fz4Of8rQfrGvtLvnoHN9R9YSR+AYVd/4yV0NUpHCly1cT26+Muaf
YXJrsu1LTjpul7Prpl4JtihCJkPfkYKmOJQKUxpZ7SQzv7pOck4iiF2s3Q7x9aWN
sD+sYT79FkJl+YOWX0CerNWDgCFFRoOzHRVopU8Chj54+6eR65w/tD/GaEyNDpky
7cHzGiJceAtssaysrAfd45UMCwFlDU7eCVBCPoL0qQxCH9qzGh7aQ4SrNQJbUr2y
RI5MpPiKjUDTf2EeUto+EoaIY1db1n2OZDbdozn2DprdlwLninRfOEdSOA+rxro5
DG1MVLiwjZ5sIYlneklC0+IbZZaOU36uQ9YAv8va1rQM/9PuQmiNjippU42iAF0U
V2pfUFDwU+iNIdHBEsZ7CRv8/FVtf5KeZwidntTApp5ma4vaPwPQXhjojNYr/LkM
sTzw911Rt+ZQ2mZbAMCTGaP9QI2ydKYg8SMkYhfzBkkXtxwIvx86DUCJm+zYWAAG
hxWeaJLnAGSLGAwHRsZD0UTDiaaHMd62ta6kEDzbhSpspLKebWGPy8p8CZggvSeI
UXerX9yqBKWz/qEKpNvephVM+XalPgI7HUnFFCLGGp3QYO3Svm8ab0oPmwWpSrGj
FASvPTsZtDg7Hqga2JHZr0EA2e4wGtZQn2IDixgCzKDTsvm2iQyc8tLt1q2zsXJr
OLJxvbtD9dB3NTzEISwyp1Lxsk1N0fIn0rWyjJ219DF6uw46P9Aaj3m5GM2vbPt/
+ANMN2JwyPUrRRD5nX68kwfa/XQuzsxn3vCKvPejR44xuWAbvdah14rg7L57v7RQ
tWVhfMVYE+EBqSTDjNptdFjcdHyzMUR/F/73RCRXXwLzkYQ3y04ucOhUQERAc65n
D51ehd3zPi02/PZl6u6SlRYyAnSGBC8RE49QJALUMhruR3qAvAzxue566VXC90ws
b9L7rBe9sI/t63ag3XAKsNcvRKwx4OpCMjW8wD2v1JyXm/boFWdHkvJSalwAsajE
edusb6Puzu0yrZ8c8Op/C/p0xye49i47AW0FCTH5Oxj6BBwG5efBK6Tpf38WTQtd
VyjJGDnIOevHs6DKDTkW5vbXe01JIHEpm213sxv1H393bwIO9QUgJXsInIVBcutB
pwe7uJEjWOF8YEkA2ioe6rmfJUPj9l0CJ3+bDjY8WIhqSiuhqZnY6aP5ziIWo2Ah
zY43R7SG7Yed7r7ZHJD4xlHv12eOQlW32+miIm8nGiP2kEcm+8jzrRUZUPclB4Ia
10EkzvW45COIfqfVWYqK+Vo3iek7jzy6Rwzlzl55ioG0npid3DEKgCrlsxvez3Eu
ga3ypsTOF+G1zU7gTB0V9VZfTd3rLXd2uQcht648ht5LtJUw4emzZpCrS2erLB5N
Zm22RCDZF+VI5UL7hmxnSBPXWu81FrJDt47kBHdgiEbAvdvP6jngWLd6joM/+yrb
y7QNuLlsjdmG1K+hnD3WoGBZ3ELkzkbLAqg4eY/7GaAC0Dm9C/jQ4L5HYvFX+ce3
pjMXrhLI4N2bOlEdfqa5DTKviu9sESJJAWojsFul/10byjAW4xA6QHug97bEZuMW
D6W1p/Z57vVekqaz1I0SHNqLXAWdNgP07+kJ53KgA5YAqjS6kjFt0PGNiAaiUOJ9
ZtWsPpn77wvSrKQmq6Ih78gqu0WyOl7wEjkcFyenpH3XG2NmSHcodCFz2oiToGYF
RIbGvt/LpVfNScQpsdkPfmTuAP6A+WrKRQIETemqBmSKQYUFMb9CJAMgg9vt/NWP
B9Py5Wg0n1CH7cJpeJqYcVPY9Q97RZu8vd4d3iTzVVUmfa9GpMHpQIBWszPCs6Uf
eXdAyYbbQar3/YyVFMy4NsU+7kfbhB/3ITWbTmuvEeTsP+D/oLzInHgtOWc9QVmw
j+nvSAhG6H29u3mFtU/vMikZ+uQfPpddoHPFVtj9QrXsMV+Kocy5Bv45FS7pFqWC
YpQLPcK8SlqByzZEFTM5DwoHyTB2yJxkfY4bzB5xk9fKtsQntm1lHlUbw8Q91BY5
o6GV5+vGodo6kGCCmUloF3+itWsiUL2+a7Ufkjb8W5zVBYSCkbB9GOlVlKW6al3Z
17seertZMYdNV7KqiMsYpxNwCmedSLLBA3H6BWhNhsoKFZNQjtHAwdXSfIsQaBFm
WQfqXk7g703NGow2zXmCAIc6/VkREEDCoqA0btUrZgwZKTxAGzNqeXK/Ip51PfVw
AMR9a3Ai7rrJENIKanw/u0T6Fyvz/da9CKGJdFxHLSINZJQZnMvKWlSN91+bOcvk
aNwpEKQsCP3LjfN+nwz4qF9yLV3aSbPDUlCMXdVW5Zz4TU3vhVeo+LzYmi/4FpLN
2igbR8DtNBHd5BDu+Cyr7XIXTWKA79vrq4UmF6Zs/k4=
`pragma protect end_protected
