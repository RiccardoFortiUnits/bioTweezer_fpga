// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Fc/W5iv+Dt0Kw43mpNFJtqfkjGxIBq0163LG9YnD7oA1qYGHkuXJ3yvPjoI1xf8niZozboBVjIv6
NR66HVNjZfKfPHKCWBFGnBRpDx2CpDxY/HWoFOhBIZ4JWgudeRq20Ydk/Z/p8HZovuUzBYiFR5rM
1B/0VMaibViOBAIC3jlpoUomlIhTjjFMR31eJmORbCLjfaqcmHFoRn0BAZ3zsy9ZD4OksUbPa8pU
RtxZPQh6Q25uUW8U5Hep6mp+oaSFLNGsBf5AHRMDniCSD/CYTrdRNRfbL2CXYz/gaFsbtWfJwcsL
Lonqvu1VjotpnJRXATlJGZPqvf/+STtr0zGqjg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22832)
pTNRxBGP/ngdAwqkjNQZyZEM9AmgHTl1x1JzENXfhRqDvKdv6WOWh2sPK4YPWkqxMQ2gW5/GPE0D
7MYzIbBNYZFcwDZ8DOum2ihQby8cqmOUfs4MT53rc7nSaVFaq8WJniG6QS0kAOCgEJ3WJ4qnTrdJ
RREYY7Z10Fpa6DzE3EMF8SLzxpbSQlqnD5l7yNbOAN/Vb2vgFryYOkMUpdgTmql4G5/20hI8G6Ss
o1iOgMgQLW2nlLwuxTTgvUNxdg0DxKy9HqT7o+cR3wb5Ki2YPLXAfQDykDqB+fCpIJZreOUMHMDB
GfzK2HkiZ3zGK9wfGynnQNdSXo6PBDnxw8CyQZRGmavlh9w65bqZy4nRMjaog/zKtxqIYUt+a2u+
nAGwevmuTiqPwuesppnbOUzWcJBj6fuyOPiZ3e922fkQimfgRx3H+bBBJnq6Q4o0uqazGGpaktYY
AgswcyObY8So0XOQuizjOXWPxjhENXwtKYxZSOWLKWGcIX4hxWkJDrldbhjHzHiX6HJY34i2fhmS
iV4HM7KtQR6oyYFrEtj9/UbM+Hex4MK4J0NEPHtP0jNVmK6M0zakZZUCQp5KL988fvl4G6/z8b46
LSgRP4wdhnmrYUJOiDby5jJBOM7PxXSBNwow3Nwng8SGO6l87P6QeB4vKaqPL+8kxzeCc+JD0DzA
PrMkWcpCcSrEngPxBkT1TNGvGGDaWgR6gB/5GRTt7f//mNUbs0N5OAcK5cjScDccCch7Dv+BsYwL
Sm89VjerA9HsfG9sjDmeo5dXVOiu19yDap2qV9oTUbDWQFr4XVdn/U9TTo4zNGlUd+RLZRr56v1I
3paGl+fdkTOHNzHy5EFHJ7C94tbUMBhmZr1nhszOudLarpfrRfo5D5qrApAUiXJfZyOMrck0nusl
gK34v/8WXY+9tdkp/e9pEOMd+Tqi65spsNemiC3MUabY8O8TWLY4rt9ewjN4XSoGhxY9wBDG9CHZ
dJURTsueDdjoI9R2b8PFj0qsgvCb1OdkZjT9tSqFsivLWgUebJkUPG/59hxIP4LXb0KcxD8kZZzx
STSrBRC2VcAKidsy0kVc2RvtiZU8U17e+uf4wVQkk9PFXIzChcUU8HUqHVF25vnMYnh8LZO1w6Rz
e2Bcs3p5Fg1jNdMnGiPBglBnpfycyPhDFihipJJxiPh001skYu6JOlqmZxtLj/K2wdsaiHNiXPFE
yLoB2SBziLu4Dog5Rfcxo/XfK70SMv1vfLIRtMyycBMvweeNIyBzb/puDqqyTxhHNx+pvFbhtDIH
iXmsPIFLs9lz9GKaldVsoFBA/aN43BZ/SWXDh2o2UA3/93kqobaJhxTPqIiZiY0J6Yvxx3aQNiRc
v7pcmZtj20EJxANeHCPwpPgTI+3wwrFdQ8c6pXSAYRzjFfZT11fbO309EwqPKHZxENyudmv1o0E4
/TFNp0fXeS9E97yfh/cpF4xBmmfXscD6NvZbWRnWz2AdJa0Pbtx0Jh4JP05rt5NHSvtNDIDZd8wO
Zx91uU4Bb1Q4DQs6Dk/EAIDxaK/jXRaTCubIrzy94DeM8UE+oTJVoHymjJyTUygbNdn/TcCGridK
CEcz/xqLgprVkL50nMgSzr+ZRLVBKSnPWKOIiup0/AV8eei/LlPluC9YoYm8BwQlN+LXCln2z02a
9BAsWeNwa6svW2dW2DOTgfDMd3NY+nvhTHuOPRvnXk/NHgPadJt+e7aLPLovLeqfvFoY6XVP6I2L
DMwW6PB6DDMcP2hicQUwICjelGImF5X/Em3A5pfHu49QnwHdoqEglWteJLKykytyGfaGZikd8KVX
69jHNUW2krBy0kEJPL6uheyUrTnvYK8S0PLsfcbxB4IkmXrikrVdc2+M+wHk+5k0+4Wm+EeqIIw4
5fwSk+6yvbEFTPm2fkTh2fYmPkd5jG4+oY98JLDEVk1EtoTXBjXusrlnBWAyhHh5BFxJLRJog2Zl
0v0FlqvlkZUQh/VzSjAKt0ph5SllvDAdt9SMaTtA64hyQznRaoDeShkjCQ6Xi8AMKAubvws8VTYJ
HbGGrskPOqutogDIf1nNh4+QKwTjvBpO5ysVheeZe6ZJ6KC5OjQx2XzEPArTpjjvSs5cnTucG8NF
ODViCVZ3P1/rEXZu25FGMFpdPHLz+n1/ZSC6+uXJv2z05RRhcH9fLxu5NU+JimWtmHXXk7I6pasP
igR7ILHwOa8e2auWlaCqwV/FhW35D/7eXOMELM1a9lPd9A0VU0hsKzY+yYUHOeucazBYJo6lhHx+
z129u68Ycx3N305EWE0PcrUobFCwKHBW8l8rvsxNu3uohfn0UahQf8LoX+5otZY4SjaZVv8AUNX/
vTyvRZU5/iFlhYJFaBi3kip2s8IenkiaOiAsKinxXnbFKFIugCtvf0B/np+JIng/R5hHq9PqlBZq
kY16rogCs/JR89boOO2tgMgIwrJkETcInlCHtG5gYVow8A1k1xD+Mr3M1XyTiR12utESlozxxfnt
kMGZd3oG0QtJPxY6sKxH6ZGoYr0B1vk+/95KZ6IXw8pHQVWCPG0sWwRRAivj6uQcXL+xJXjl1UQN
2Edp8aVKerEq38w1Yxg7rgjEof7OTBrKYbViNp6akJOuf78EVtk9hvrOoTKv5G2dGxXmy5HX7cQ1
kd3fIbrB69/3UVV/VQVPetOQ6awybLlSJush2ecGGi8AOe/VSxqf4ZvGkC8VNf7XJ/iBIWjUkfd9
StxVxV6Vc14xVZSxEcrfoIJRmp9hJSPJVjBgJvW4UX5TRXvHprtlwLkJ9JlK6nNaQOWHCmy8qVRu
FBZov6Oss2YFu40CjHGznm/XITGGcy2P5o3xQ6/RZGnejHx+jSuqRNQ0/UdUY1ebOdgY1tRNNPEI
leCYPL9D6ZP3BTVWtBU0f7MKGMkPEzG10XUi7lSq9ibXv1pPV8K6YSNSBQgD4g+pq1IXejYM8i3M
Z5cWlGtNulWdMB6UfcNBJnxQn616fy4a0G70QBc3FlUusxASHTXn1qmRqDLEy8AtN/eJbFhaaMEZ
RTPUORdYilMdjhfYbMQ0SZpI3yibBQlfospvNmzuqKrgEWPoYzcfE8V9HVOQnuGjermwdf6yJMHU
CbOQMy8j3s0S5/TbVCA8yL0n8LAAkReio7E21CuKZ7phXkYxZrpqIz+lnd9j2E4UIJPIQMgR/NBe
Gn/y9xt5KDFz38UFe9HSx1b8DlPykUURIGNtfTjdpIykLvKAlli6Ie44G9uVo5t1arRY/JqQ48O7
vPITagta6XV6xuGnkmPvOEtuf91rozLJy1okfuPzHfFeitX/V6yrYQNPW9853O3MAJCqWLtcnOLU
jfGdv4Mn/8p7jq59NQbELpw0xhHal6Jg1zBTPx3zBpXmEYyUyvE/gNwCYv98LxHp3YDiDqcTE8Tw
D7kvRVWUx1H0GTzoJo/Hyu5erzMvAhn6DHZzJ0N+uN50yYE61QStQ6imvyLixaggiuPYOAY5kV0z
gkXH0QZdR18VeJRhTv2YCQ4aJfM4ghahsoULLOBbh6mA8dF7B9Z80Ibni5tsQu9prmO7tlFNexSX
Na2g1DStQl47ZlddE8RBI0CaussSXijMJwFyHeG1f3rF8THzd/BpZf+L1aMqnFrHbo6DeOdo4rug
zsDaaOQyn92UOmGeEj+e89fPnnMwB+8/cc7KADql4hjzLUon0larS2Rp9PptRDT1WHDVj7oAxukV
7iXhqz108yutvE4drayN4Bi59e7K7enu/FPkI/tWU4OcmkewNaptmDO34Tgf8j4TgXVZubwVNdhW
7QkA+2uVd798QMn7fYCezTuS9xX8zQuaqJWzdWmQXX9sSIAAJjd+iyCxVCsQU1QHyGIwU8QxTpnR
+nfXDR/mRJsOss3dsSLF3SFGdxIevuX+5auVzsdQtseu8lu4kHjc7xE13fbG4E8xHZShqK7MkyVZ
tQUTIP4zQ4LatYDpHpKOgu9OcWCrnxed56Lc17SRMplHfK5dnn8uhiOS3xySumiK8MIhsHK26f0a
LlWwcggjFTTMZryx1hDqLBxN8PCQtZjwLbtPr+76nieuNJIMeajtQx39EX2KFcOd1CtnzkRb2frf
ZqF/4LT/zlqp3HnXafA6pf8QhhQE8O1W2+cnuwDBBZxZMX7L0U3pn3s3sDALq676McwEP/iE2gGk
jpQ8sclNYdjE3uK6W+iGxNmkN2qA5+ZG6umpb+oLiQyH4pY23UcQLlQQZtPcQSoiN6x1cLSoCf/n
jL0j2+kLoyvh4ghswgvJsLer8qWGhJo6VLLL5MGOoVqs7TTaMZXJoMwJMFc6k7IxJbWPCauMQGxr
xfvawE7XgUkr5ezlYTchcE7ai7VB0Ucy7DuDHnBBd6Tzyt8hN8fTWobq3yR/jDHVPpwKunlvPofQ
GKDMdx1Oczc54OOeVfN9V0+lwkuyqBB1nh/gdTXmG0DuLgPmlPj2tv0UvxauK13MDsc+Fss1slcP
YrL56EnL8CPmflHjGcwD3KKZBsWFNoC3UxQQ5YKEcr8HZAbZ4L5aY52m44qlaISBjs6GN4dzotm5
6O+kOne3MkQaJUaLUlW0qM1chUPYW6WWAaJR/YhvAfEVu03RnTntytmSKT0QSyNVN4MHpmbi4Atr
NzTZPB4jcv41SI4bvSjooYMI3oaLxiP4pPvoi/lTciLO5X0r1a0/5y86OvFLPjUpMgvhtkOLne1L
cWAJAuh075sqeU0Q1bGfY41ABLTv9FL9AG1v8x0vgokvvmE0PkWQwq1ATRRrymw0L4sQmX7zuOvI
6JpOsGPJkhw6SWC5mMd24nKQOo388FJdAAU6SN19x+FUX/6QYh39Dz1N+mW5BQv43wihZW1ZhdRu
ZeStrZTAe8he6EYyblTcrXS9mYif4vFudMpQW4JFbxB9lmGY5RtbR+wvg6SsLu0p/MciitCBmvzw
ohvjPqmgCLino4ccZiTAZBYn5jTXNmH81nzQBOfc4OQ/1TXQLSGj22//CJ4pzLZTcN8kNYqeFE5W
Ky2aUOfQh90tzaC2touGoSISUsWekCu3z9VlXspcJbZA1gQ1Fy2zth90qtJrGbJXnl1AmLp4+NGh
t2KVHyYHJfb/R9flEzECmzRfoBB9RT7NY/Wrb67ZAbskgg+JoDU1iZlZosaAemPwUvT4aZwR31MS
wzH2YasMO5uy3B1x61UxUYTvH+iG3LVJqcxtRXS46pXAgH3Tw5tQbWWRsMmpXAqAODjJvph68nI0
QhreXfE3EyOjJkAVMWoJlLZaGTn+XmVySgqA9THvR+XvNc1Uy+SFPgjljp1WLwAoNCHyg0NtAdmp
ZBKu7pAiKAkSkm+erD5B5QZDH5pZsEajcSLFVaQlr5C/j6xEjCmEuMn5r3pgAOusRIAZDOxZTx/q
iarNTQliF3z96LEaV7bPAC6+bMDKMGOtKuKtC1QgSofHDggGxqsNZkIw+xgG1E0XdS0WKJylLApk
rZlyycY88fbuKdeYHX3baqCbx0vNdQNxFDxZ3jho9+AMQkrS1u8tMmORMgUg5hws6RtfhgE6uTGy
Mj2yJLfhHtMB9T+0Efl0YFeccETRWwdx3q7KzGsZPixkJ3rBEko3XbTx2Tb4yuLKko9gDk/WsSEt
E5gMQNa7d9RdDgVsldcfQEm78fB71q2aLjAdHNQOjVDsh6IIVL/UgBf7Gw0zUb+ODdL/fEnGY/zO
7f0E3HsBPUPV3QzDikRe8QTzV+SouesyM/tDfgyrQZSdnbYI5b1S1XNNkv+KaW9ZcjZgnNNJkuZx
Q8z/sFHBAVLa2ThO9xoOFIeK6oNythF4nAWzRRCsIz/nhAqseUu9LO2bYRGxUdJ6kcgO4bA7CIfP
/iIqcSS4wQDd3vwdJhbnaFpOMdLc+jfCtrOU2SJSKtM4qZroPuRWhMfsrfPtHp5pczFbEvGbHfdI
AxdA9BvzJYr4IkpDttrk2wUdy4HZZkDHsbqQQRqwy7cDpzAIimg97/hFaiVsZ3yToy9TsfMFWLMV
Z7KETxACEQTh+luzOzdBi5FnRsGhi0GlEn6Gwu0VmeP3Nn1MoVjzdjSoowV3uV52t/YDiyIDfySu
YcIhSjUZptQHocdtxRu012738PPcfJznxl/YsPI6ayBf4B3k0WL/AMyEoU3W/m9zqlJ2hZW4KmI5
Dh+RipKJGIeEQOHGXl0qK/Tu9HmSvOW3O0mx/RPl5lDe8HMIcgw8f+5cy+NIqjnGkQINgkz9aNNp
KSOFq5iSKvre4h3Ya490bXrpRqcCmNGdssTiaNpL7NTt0i1jC+ywZcAGURPgK4iwC9ArU6/lPjin
/gwVIFaIoX960ybXHfgQKcp/kn9wPaEBcrtiXXEi68OtZPV33CbbmPWguHKjNR1MXoayAkQiq9dp
Db8qCXJj+k11wz4Vak8dtj1M3j1XSOGkjxbX653y+Ys5OkZLVxViJhunBLx4PNHCzGr0mHzV+suF
yNZapf81M/Hhr/x5+kUgunJ7P4xaGuONiY+dlWivGNmG4Y+/RZ40x5lmYSjxKc+eF88ygHSfI4iV
9cQJl/RtNiWtlhMLI2Nk+AcRlRrbEkGedFpOXQ+mLYYBEAy6Do8DcLz888Y1lowM71iytP9y5+sb
YU9orzB/+1QITl1a3wF3XA5Xa7QMLB+/8Lyxs8CfBqNklwQVJ1AiDAeKvz5/dloA1FplzC5MVvy/
cBU0dk9pkpMkYOj74BSBV4wpx+XHepM95fkTWceqBfwMgd+B/fkhNQ50rclt8lE6JR1uiwxVI3up
aApLv5WbTSoWJ32uTaUsH/L2XoOsqjHZsgCwI58nKN4rKgsRWzTqUsN2NItGJncKRqnwP9A2bb+l
utQdNC1kt+/plSdfE4ug8RGH3s/Zt4WyQUisWAjHbk6rezJqKlig/vBs4iOaeTwNCQV7G0UXAWEo
iNjBRFs9SL4HToH4F62A2YZm30J9Q09DGyVURbA0u0vlYdLZBX/HOfRjUwd+nT/WVdRnUWvjIptB
q/t+dz0KkM7qIRdgV+cz8viFDZv69oYRvbVJB7UxnfOaPwtLCM9M6pce8U8Q5gYMVupEd4+/a309
HpIj56dabeHauqyxpclJir5WmAdgVg5Jgu9pEqZQIXgLGcOt+I4AOi0w9kD9YpvLA8lbqCJuSkap
8O0z4/iYApBhbUQfN/jS2yDpkgiubP/M8qugb4jPDiwI8DIFxqJnSopN/S+Ql7lU7n20jtSt4FSB
ksjUwsfTI1nQlY2vyQvfS+GBLoi+YAddJAiULa3yiJlFe9RC3PEeDpbTCqx84UFcG4/TqR1E8Xy7
xuWkv8k4cxWJ3cVeoa/cn+osvmN3lZB+A5Z07TWmC6L6GZaArWmdDXQE99Q02XBi7ch0RMFQsbN0
O6O/yuLTl9NQPlFSa7ZfK3wkirH6aWRNDwGOhW3wvgy+SL2tTOojz9/mZS+XVAfMmSSvxXwIh9Ol
5z+dMZjf8G6BkcuPK/Yc2/CT7GI3Nyur6YIG26pmRhr3vgBGEsmQz/IFl3pXrSiULG7hLbrcNy63
jLvAAFTasqxcAdDOyo90raJ6PsxZLLTKLfy6F7Gk+iodFTFtIO5xUtCtl9WSf8XnE9+tvSBiXacC
CjTZkB2Q/lR6hb/UcqlvrMMYL1y0Mi1tVW7+7G1r+S5+rr/Zmw47hxf5E/4bIYZG6zV+WlSX+Ahx
VzOKUoMfmM913mSkB4P+L2eQdNsoJJx4/DzslBOgOq51PwcC8rGBDiYG4k2YUFjrzGXOcuCpvDkD
78tyaR1Omc+x21mN0eHpPpunBoQK/Xd7GKleZhEYC80XJj6aXpWJMnwFPDZCXYZlQjmd1JqE9/sE
8GbJgM8WAkkr089h0ic0aG5SkY352TRaXJBNM8Dt0Q1lxu+MqB9CYR2ROsku4amBV5dGnk9Jrfgb
l/jRaz5VrAPYU5Pgtr4YaHF9khrGQSu+LClYULyaK4Icj3rubwFRNFjfMXLDz1bjEdepMqCebWsa
qNu5kkJnA0h/4nyjdI8lF9n2pv+FAQjrHPYie1ZlHHbHuR3R6ovzrTyx4/kg/fPy5HPvWHQs6U3I
CegTqwiNnq+TAmkS+wZ/I6AJTv+GAMz4598vIiX9N8PAeXGjSuXutjaMEBpk/YJpgSRlV450kAPl
ng7cHXPQFLQHug7K6WXv0txnjtd+JIKdcoWp/tWLtDaX6QmO8gQkxe7JbqQU53MPjbD50nvMtJOz
+pCMyomXKBLNdO43AKIwwW/7NwhtQfLfiVcgsMfxmTJXiRTc88yu9fNjF2FVTlFvAOeyhfR7ivRH
ySeultrh6mVQ8nMezFh7KCZ02pyu1d2TSJsSwmOEgZc8ZqKa7kBaVqV8x+9RHvD5wMFOoQdGGbMW
0Fg3tyo27H3dLykfXy/8zfCqXeNzbK0jRjApWmsbfPDtAXIe4S3SEYGhgd8Yx+7EdJ35IsAVN2dd
kEZf8vP16yu7FWDApYe1sxmz+DiX1WE/9r4wUPyZ2bFvRoUq6gJPpPchkPvtJPHbBu24ed+NkRO6
2gfIC7zJWDRPYO0wSJh3OnVLDAHqj5cw5YcX+Kp8erd0b86iJEINxDadWx9gkJ4rT0BY5IijqSCI
KjnJMLKzDTYZHNGGZpzL8GOFvx2NozMM6pqDyX+4CZ0OoUeRK5wuowWOHVGYyTV124l7yOU2ehI8
cyJHhZEH05wMncZRjljapTP2OMS0xySkHpgqRTbmxBbBkOFezEYfK+FNPpCkkvrDSCcf0cA3aTKp
FavenmdpzDwfG0A4O1FLofISNdr4BVIpuZCHkz/TH9VWSNIq9jso5lKK38rucGuwFP+QWQrQPeA7
aenUGSEOEARmZFfQUHtVlh6WQ2pZhykl8Ke+yR7Ap1O7tXB4FaIZrdLn+dWV86znXnHTWrK01Zwb
T7PgxBLVf/39hL4tbPo2LtK/xVIqHCEmx6tGj9niIRy6VY6HPNmkNq6EbilsfrdtPlWYKcHcOr+9
RES188hoV6iTc2Bi2FVE3iFnxvuaM8D/SNP0fvqKad6QwQTPttlIHFiCilbT3P6Eoz7cP+gmaL+H
vpmLeI0MkCDz1lh7inVidq9G3eQJquNJRJdgm8FE73Ch/SnaVjyfTMFW8yQ00TDUtOFYEY/Ev65D
OzNc9nwVbgcoeKxJxDbJGZfUgs6EXKXFcLz6OiF/23JKL8w1F+fD0ZWMMbvjcpr2b8EQHFuKC8G1
wbaHODgLRdbrkyr+gBy0LHfzQC6bAUT79HCN84MzAyOUHmts4kdB3Bcsertq0t9Na0/0lxRfFerB
/ecpWIDzQpLFzRl3sejlavR1IDcKjmrrZdMPHfSB6hUb1b3LEfM7vEeKOPcYd6PV+GuvE04Jg5Fx
zQCK3BqeAAZZ/7T2LEJP15Enq9XYnAtzXIjO6s4y1EvN/fxTumyW9yDgPP5fmedXJpapE9xlHwkl
M8NlvKsf53r+A3cFJmwFBJS4/YgEU0LT/bWeSYzJ9Ivce4vbvrJDfUHIrI3ithU2bXwKpVLpYYFQ
zBiLmRayK3Biltkl7TrI8HdFITlLCLq3dVK7xN06BaEQxURmww8i14TXVrs2ArhT1eLS2CQODRwI
LokA1GJz4Ue3X9IfNcRRQOYMbj7GFNk6dFcKKDd5nxoieu68UWgi4fSm++exL3VjT87ZTvKcLMGK
aGjcpTdFScLg/4a43ovs7lESFzUjLgZVtJkisBBUcR8gzrvVYOQ9LqX36qM9IT17PNS1F4Cj06nh
EGJHnSh2Ht1ApgpavW/bDyyePegIcAPCFNEMq5oVc5DE6qATPJrUmK4+tKTdaJy5PDoqve3gXHns
s5B4B+684E+bfd4aXLDp5QYVgbJZjVHVB0RZTl7vTc+ZMT5sVE/OFsMaZCgm2zvUrOc/Ofx+74a3
JKhzMBF8+17TJesLhG1H+nTX7iFJeR6V43VdkU1XzGCYFuSNgyXYfr+QTlSY1B+TX6OUeZjsbazI
ViIk3h2xv3mJvNsrPSLulQOMXCyuts5GcSERYH2WwSqDWKdfQmpLkNPDvTouLATgrM8agyDm7YF4
hCrt1pP8lQghBgZNVf3boKIaee9sYM1EDQeLIBKchmqW3O3JVgC979K7pMO3s3ER7+bnYEx4fk+9
UG5cnPExaIjCiGDAMGJxrbkbOIcjafK5uNEE9T/OjZWlCalT6GxJ1isyFCq1QB1s4eeRm1LwpOUa
PnDRxMv66fEkXVivqHewhI/UXgDhTld1RXK560uwbryC+Zlm3gaVnlPagKTMiFsIK55J5MY6vM2F
o5pswxKbPF8F7hRbZ6OLvI7erXwOiUu9Ecyu5JWxpkM8flh/vUhQnopAhx1XflhzpPbTGsVDrNO4
yYD6zW2ZM0rEM8hP5YIV+8G1rHqzJMgdftGjLcOSpe+oeVYlxroh+8WbdflGGUNaZ4BaOT3mRLW0
UwRVKFCufN0DefwMYwnDAUhLT6zR8feaIgNV6mIrNf8kuCY4joiaGQQ4AkcE16iaVDBDBr9qUe64
KbUbsIsCqyRraVtCYMayeAJQ02LJ4bJ3X7fG7HvZJ5I3UHRTwCsDjc3C5cMbmS2op6xYubgHw+vz
4KWLnOn/KW7JxX/DHuIl7fwl9kjjrdOHuaUQrZaQwCzh0Ed1aOxc5eybf2f35OyspDKgmB40CSZe
K8CfP2OOIN1k91zQCTez3motRfGk6Lri3E4zwC0WgzT//36vKuIhd7DS+0hszyglGrA8wtsp23FV
Ptl70e0nKFPbcJRjCuPVM/HoyU0Y0+firyrfCKkDLzB3Co4wLYhoKs/u7s+BGLGCbTYikCRGdX3E
W0qqK7JGUBRazBNPzD3sRxtLJODDR8WubbKyfMlw8Faz7rSvF3l3VKbAP88EPevaD91x/mgL3Nqd
KLOg71SAMR36P2QExkaYHGeegAzwh1mJzZcqsmvJSOlhx1jFgsYaltg9JoAsPHbAa3BDky16NZXH
m+VMovhI1EqH5iJabHZyLrBaT2cFQJMimXU2dp8qcXG1C69BbmoQRheSaqrFUsuYr+y4C8wZJxm8
A9sMLVo5u5IqOAFBQw/9B2lzAh3P83OvT33zvlCn7TrU47uqYAHmOSh43aYEjekyOPBHwhEis8AV
GnPx7yO9ka3UmDarmvJZpn+t8/xU0WutSnj03p061UUkeYbL9H2Z/U1vtJDxisLUVQ78tqZihm51
1lbzGVq5j3EzI6CGoLlkqXNdSVboVhMGwmgD78IBiYr5qgpbRDQ2/AfOeRrUSRkzf46wR6w+o9Ub
2T4XM+Ez1UecXNEUPBNpUoSOgut+hmLODzzuuyZAgUzRu44gfhFqSfdrro3S6tjgmDsTAOvy3Zkw
k8aR34UW1Bs6g7Ol/MQzUyNxlTzIH2Y+6lNQvjY71gO8ffsHJBYVxj+KiWrJhxXisVo5pZUjmEIg
7FuJzcaAuc39q009I3b2SiNEyFnni/n5LXNKAOhHHSqfySpSsyvZl4TRxsTc8hXPvaTcAydwtrqZ
azFrgC9mGy/Xc5/8wsfjtG1kopN7e9HMhJsG3QC4mIYAMl23dv/URN8/TXSdzLY1iuuSrrj0s/NY
HLzeQQt+8bEhNdQw1NTTurUzUAis8zoGbCfy49lW3qkLAx2FS7+9PQb0rxNVTnBt2gYrKaHFxzv6
9wEMOEeyk4v+yQxFXHtkbR6R9DGN2VR0xnilsEYaOmQnfGaRokopwW2PgiGMHehvxNBzUPLpxw4/
HPtF+TtFoZbk3/BXg0FBfphl+kNVjM7zIFuO3CIfZPrCqEj6WAWUzwguNh2Ffs5E87V72faGXI6L
2/vaopY+DLhQ+YgIJRbzGZ7Lpp4C2J9dcfGZ2N5eu/i9fQPW0bQb+zODshW75Al3Nce0/esk/Dw3
OHeRSZQlO/XRkN2kTyaCnQYy9SrayYS8xvSfK2T+K7UfzZrr6UNmb6mHGsioGAKbZazgHWUV0RcL
YxNGB49WNeivcAiAY5ylUmW0IC1Fbl2g9a1gPw/Q8ccHA0kjlrOdEHDUELb5ITpPSE8/w24T/IYu
ReKHRmyGKzc3J0jKN1yP0XPUDl4L2aULe6gJjvmbW3/C8drkwQ92TWMl2uYyJ6oU6/VfegdAEF4i
/i5WmGzPKM+PHVxSXCYrFunx89xXdLjveHDQU9+ezPhdCrnzQCyVJkeeiu7VGKLr3RX7s5QJjjn5
L/rppCjC6hmSCvl+6XuojWgg2sC7PRnGe54q7zC4bOlDvqLJyYXAT86ioevWjkuAV7iVmS2p++oX
vOE3aaUHm5UXj7vPX9cIbpBi9T1BirxA7GZKdg7eOY6i2xxbgFMyeIj0wFd6IKnwyjADTOpbC7Ll
y85VNw4qjc3nydHsA+zlPg/JeB6py10F80e4bypOW8KFcSdVqbcCzMse0sslpmBS73+FBzgTXN2f
hVGfg47cesDlYxu7/z2E/bzr+Qj6GAGYJn3FkVJWvGdOaMYmiyq7TwpHd1ReVCW2et5wAdJ6uzO4
ikS/rMxM/q940OB2Q6np4PvQs0UE1xcjOoywOy459rFPjdxd5JnqGsH5RpfHqr9BtkA+Md4qrvQi
nINlaXOeMj3gkHk4IqYMHnEETyOOcFrffAKWrKdlG9dey+CG0Nnx1pX+UWbo6azoAPjaA/+KH04m
wzDVcAhwrztM+sBlMEYK89Rz5xXFnDpXHA7sjfDWrcxCnyBxI9DkhvcbqN7s3f/MzZdsUo0EBeWN
7eIcr/W9ouRJ6xpHQN7ZKJbUQt3Ic2hTQwVlPss9hWReH0Tv2qY2rP1oz6yqXKtusPFE1PpTnRtf
YvL1jq00CNqtQZDgdKr25pRGYqIMcrCHcl3lE8Wn1SlkMSgM7YoCTvwE7iaCqs/MvKvuH+aqwZ7P
uEt1qW4vRdAjCE56Ccpmd9erDgSWzPK4AcYQJvhNAr7vgIn4qDIduU4vMpl+7GUH9xFQb28NSLf4
TBAA1Wrs5ETZNsV4T36RKE0fuwKJLE39JIt80mgkg0d5Ngo6kCQS24JHQ382AeLXwfOwxwBMX3EB
pW79kObmoZvddaFploQNwwQZyHG9PeeTf9vh1EzDT7x8dAHYap9+mcvAR4brptp5EmDOnvFmb1Wh
tOsRNjQnuNmjrrSuQM1vPFqkR1ExZoslxI+k+zDGDtuwL5l4Z4chPv6KazDCI38qd8AFfv81Gy4r
bJ2y6mGldOJalfC7hY8gHdpOQLhFqEBlyBoQKLItEFtXNfrrg0rbJ4mKtLuMCkVhAZMzTpnVJShF
z2QCx/JgLFRkzWVAiOT9L/43gpNTkbSb9XRcr8IHkzrmCQDdorDRq9amThWqCH1rwZQ92uN09qrQ
NliiTp6KJwmhK7MNMBbpkFsYYpCrdeoMdV1jzrj55jEq74R6iTPKAoVOVnWscRbuyMhK4KxEuX9U
q/gHN0Eqz5RBWy8AYUIsFkW0ukbUXi5CHHNSAW3cgjknbhJj14j7KaNdapaP1yL54VkSQGnXImvc
XMW/KvunGhTplPtR1SOBf4G1KVSFtqvsLPnF/pWYE0IIaxUEHMHcEgpAOcM4imU3nqezf3h82v1W
CykhTRpBE2P4tsiYDo4VPnaz4DemuzZlNPJhjKliJQvNOFE4VIvOBTj5+8Uk3EMwwjA6nwTIA9Yf
g3HlMnVq9Y7ERlBmkcruOqs0DXROnpAPPQ3dQ5zeFMJGZFocjilGIjN+fQrlBiUyP9vZ5CjCIWtd
15EgTOsNmGByUwxqnB7mvK29W7oLIzPdjSJShNpNgsxLYi2v6tyJiQrgJ3jcxN0gEfM0iBISKqOo
r2rxZA8hf1sOLZ1YbiNjjwmGTyIHqVpgiVKPAqgsORgbzSBW5ICWM3083bF4QQO/BdmmomIx14oD
fatVjZRGgrmLyoWOfjQsubjBTpZnnRXBOvs7/8Wo3VSgQBXT5hoC2/C/Jkis4xPLGETmKYh0Y2RQ
eHfb4nj7C4xA9BNadoUMIwhSsrN9hT+SAh0AYp5GEBA88vYXc8DRDsYMUtum+zLtHQU2xToR/k6L
nFD6vejOD5FA3jmxXl7y2r3V4MUTT/zAche5gmYLnssyn6dLeViEk8skAYj53MfrZ9V2DNUqY11N
FLRlIgChKXg8KOVsyMjqTSWPAdZUJx+sq0qFrOaROF5pg5rYnl6c5ziODBnvGwjupX2wxDAl3S0v
CfWL4UnnAnwdsJw74nfZ0azxjR5sf/38eo+ky0MaN2TW9MgbCsutwvWgAMk+aO/ynFgJBy1Y2Ro4
49clEZ7rl1ZTNJhwLOK5DnJrnFLMX5wlmyzDf5cM5Rsdy6TI88pccBcmI8Iz9LyVfv8M/LkDCutq
A2vwYZEOs0LsdT96ZfpYbqwt1SbK/6xgN5fPonMH2aQB+YmLhaCPqJ6+RXmBo+V1VFUt+8p9iIK9
xzxqU8CWLI0gXy+RrkgbkOTXTvFB/joeqhW0JtM69SQwop1YiaBpH0JHPUoMGxgdh15KP0jnVKfm
9IJJrD36BAYRjRK2mEpfAa+Tcy/qRVRO7yPR0VxiVAygazHPbZxxSp4G1GhQ1ltt/Y+b/1iMJjus
qLFJ4tFyMKd94JeT5WkpIie+zvj2WbQz9N+Omm2+dbyUowCL5lT77GB8h8osnbH//DRgnEbVA2XG
jWT+ZY+s0A4be8iH6wemXzU2e0rf7Wmx8ziLstUFzj+CpBxZcM4XJQeT+f+hpcpPqHXGHWtbKc+b
1SIw0Kk8mhuCfJwVCzYQx06x0kgzNwV779vT906R8fDWlAht2YxLfz7R4y1FuY8C++ICRR6W6nCj
LXP4nzxrT5z/P2NapOVY9Rk+JFJuq7dQjYSZmCFAV03jjE6reWMClU5lII/tLjMGyVpSEee4g+FS
3PldxjFpy672lPulaME2Jooko4m8rmNbqDQkMK1KSUQHT2exn8nMyFV4l+GPlZQS55ovDtA9AK3O
KMPdSUcsLP5M656MbYMKkSB7QBsYAxZKDOez6EU+vC7TCNVZQl6DbtXPkFwEHCYYU+QpIBjHgcJA
uIzwBE5Om5MSPE+PWWUKf7z621UegTykvxwxXTMdbXU2sDi1CXEXrfbE5V6FTIVSicngxKtzTZcS
F2Ycfs355FvSITRKefmA2klrPqXwI21yVIrSiVBL6rbyAQhZXoLhC/H5ocujdDSThBbhHLlMQg08
F/G85pjYSw87NJOkNlqQzm+7+IxgRVd/oVywl8LLdcJvQpHk0TLy2rMRvYmcZIqToONy/aqGijA0
mQ7xnVlJNYHp1JDpct7ro5n/+0eMri8+6Q9Ubmz3KcLvpCKnq8s7x6m9QkxyMNgxfyQ7BJyAAJM5
NSjUsN6Ag/UDEedeF5bT+3zqH4t5o7RWsxFsOSD/Za/PjUH35HhXAbyYbS88SvYb6cAXnEgkURwL
yOdH7E6HmDLPy4tIEYaBab29y//xtkl+WZ7uni5mU5MPea5ecTdwBZSV/9e4NinbrnLkGUcxubtB
dDEg1scDACWB1wmUu4Mf8YkytkZOLJ2azwhawdozaSfRliCUEJbrvzbdCxGKM3wHp5DaeWymRAZP
2eKU19KxdFHELuk3WI2ETyF5RbVohmEYNgrR0rt+eyhfWokQzPyBYkZ9dkgVRqwG7mv/axy4UFwT
uyhHu8ffQVSrXL0Gv37A63Wge37TvWf822R66MhwqJjIPy0IRQICi3L/Bw7J8xCTEvkrmieYcDH1
1iVW4CkS6MLRuwuS+U1sLfzYDtLN//xg3SrtoBUE/Ueek8eTpPkqKpNRedotEfjU68Rag8/BAnf4
50cbA5EbfR5X+1RqK3qYWm7/InKSRtL2SDA2yJIJ9arsaeEHDd3Wa+Bdos5AC3qK3fnL4rPoPFpt
WwI2lEPLFobezqUr2IuC9H8WGhDPKg2Ha6XqegU8QIIxp9mt8OqT395116Hjt3BU5oCkYVVNf8SZ
R+L6rvs/N3POvWqBU7n8xJ9i7LEwJ2Y9W5ZdVU1T3tSXQXKxBgUKwuexMtb64VEE3gdHWGaNTJsk
B53n74Mn+hha8w16rUHm9lE8JCvegbH2PXflFjkmQDUii7vkkDIVE070EnBRkmZLvdSpfmXvh6xl
4CMgPm5JRH4OzB7tVCderdPaPxh2aF/1MXMAANlZrNC3GgzflQvI2BS2VK8PRfXFkXLlBO0qMZ7d
sYB310sHcekIBKrrRATwvGvFxaLgTya04T+/8lAAyeyNUm3L/zNoXmPH4dUkpJ4/IzaTf95jj8hY
f5DSEHZu5cqeMs+SuOVeywszV2GoJKwPKaYsQgBYu1TAnA6ZhNGY1B7BzivZLW0h7X9y0Hw/qhro
f3rYWP5sHbBy9cnD3hpQFTnzHGS1b9abfTxdJavZQ4raVVd+rO9ixZJtctIhgGIuRVJWWzQLA6Tx
hcnypgpRvhEHPxqNL2IhokrQguYM05bh7218oVoNP/bcaWTU07rykImY6hdZbNfVUONuM9cLF+fh
4UhORk3PC8byJisZp1xlXkxoCByp30Qqav7mfRs8IQ4bViZVxp9jlx55zhIBLKGyW2lxxBlcWysx
q54QdsjeaCsmPZL7wlzUekI7ZFuP92UrD6wmjRTTOxcI27RlbRSxKL5XjvXi/4xFLVtSbUtOLrQx
mJZQhJbXwfvZSboVpsOTHlEysJAeYgzHmVGR/3zuLf5WLOaZKt9YPXHzjPOUq2Pq3n8goY9RFdjV
UgWUEIabLBRLBZZsERXHHW3DbOR/g0jZzdM36N5o+aVW73lzjq9h0T0B1hgnsri20cYOeDti9Aw3
Ne9zo10tl/49zW0ZQzqx0Uy3++lB7/LLO5gHXF7wbmRHeN9LECDHQ4JEuA21CbKlt1vsIrmoQhFW
l8tScQ/4CybN/HntEjAiV3Dbtoe8+cCYLPTDuKpj7sL1LLb+g8WsuLC4N0q++5ZAD3IAnYzpE2qF
7SlwJdR3npQ7xwWm/vZdN7MbTrgi82wEwtjtTUeMYFiRi/Oyma17mxJjvQBu5IrSWs1vJStMw8IF
PbQl5tNVsEH6cFIlf4IdT2YGb24HfKIrO6sVDaStF18yv9/4zN8uvBwIDZ6ysE21QVqMPsWf9+DE
HNv176vDkcqJ75VrOV9rAE8740VfqFUecp0+gqlHoUj9fyPc/AR8LooT9beGHP70Qx/QD4Efm/MH
KhExI1NB6zSmTiNUzG/uo7nqE66fiSBXjc0oL+c4pcfpGaJGkAhH/pNfvusc8k/BeBVx1Ww6Sy3O
4pVm1TYfKUQmgzFeCsF0oD0AoAm4OKDjvcEKD6ruyaursHwmZn2xoH3JdeBb5JHVfY0DcXtkhANw
xexAjMGU7leIhTSZwYqjysJccHP7IvRDP7FFBdPaxcxHzWJRAGpHpB4Aqmy7u7fFsBGwXw2eQjiT
SBAcBEcKjBgQDmFqMlK++/oJfdnjRSBTEgk2JBgJZpLvjXDUv/xt8WlCMMtiCO4Q7dXkJN/hF7CQ
KEPNfS6uxkaVEWYd4SKc0Wgv/cyYKTR+TypV7MJAFjYcTU6FAfcLQ1qHIUUHDWDhqMM4+ZcfHCxM
22XOXLiRXaxAT+uIohjyAP6s5CrmI5n56JYtu4Lnrcv8FYKEk/j2vfWLgbgE6q6UDGVZdQ5gqL5A
GAHkJBJsXRfl8bDgkn5aGPOe7QCXTGf69rXWifxnD2RZ4Wb+Z2VdeqaDDhxyDsJ1xkBNYql/MSsg
pqbh8DFYrdny0HtT4R2HYbSwDiBG96U90Eq+KikjziBjHCJGxCLH6k1Xog+qpLEh78fi6108v5xC
MR7QgVHbhYJ4TgWI1OKzKJvfCXJmZ1zwpJYtN4WxWBShLwfwapsZDjaEwEmriq73K8ccY4cytYJ3
VN/8UvYzV6q/OVTJgo6VZkA17eQYdAAtAtZcA8n9N72Qj4TJmWiVz+ueO2kZdjE6NWwGG7//u4Jt
dkhU1hs8DtPz068x8Ak6vRd8OCWmWRVH7fKjZ/P0cXT2ey31+ENtsUwaXLZ5lPCdYlKw6Aro0HPx
BSLY3Rs/csHIgzf8014VXxi8xFILE+AJXwadZWo42X1WfcVrewaDCKbl70Nd+p127YZ7a6NwYrZS
1U4c+0K/fW8ZGOVj1H+np7kvkacLBTZBPTzHF8gzLXQDCq/IfkH0pzN3B+0faZsrEq0gohiZMe6H
yEv1yKQqKPSoPttA/PyE+9nLpwjl/oRhIAUMLjH8hCmhwucCJ9Yono4dS1ph9p/SaeDItJGCO2R7
/AaD9cQtzS3lWounxEZ71Kd45MtS6BiChecJWm74b+BtN+enzwTnPcvYd2Yq17cxYrQveFqZl6ya
StfixcxqbvMbX7uBA0cmBswfx6ABIUlqsXMRA57pexheISbCGSYNrpk9kUO9VnM7GU5NkRy/0kZf
NZgO7hoRoMT7tAx2J3aK45M6bVQcjczQYQ//wOtvl+Pva5i9u5SelovNfA0tXzc9ic+h0FNNLxgq
TH2PWOmVP0pwq2V4N+Kuk10C3In5G92YFdfUAqGdU4ApA5/QdH9Pnv2UWE4JztKOP0jGS9iV6nYL
oa2gx4L6V5I5c3FMgiIwtf0/CVgTTQ6xIxZzF6obGFfZ/9qBWv01NxV8oF5UJ0BUcq6bePwwn6bJ
X3J0QfkFXxwVcubsnQMg5WL2E9m7WJ6aEbiDG9ZMmLCBK+xugq2AmdCF8yVUNJ6u5ksDOyF5Hn27
fFrq5FmnISBAbNuQ6mXEHTV5tgKsvxigwkTpRnlPAl14o5/WLI1ViVohCeCOYpr5/35aoShnuxNx
FKJFSoFreBzbJsmUk1jOuf1c4S/ed658mlVhjPUcsV0lGMJsVexj7p40DL1uaUcE7S21vpY9/HAh
ghgl/XsSMW9x2oguP5iGJilOiNsuenwEIKFeijVzhFHIL9SEfMKjeMODX8Hbt/l1XNvSb3ap0e6M
BJSDGdWGdSaUBvDusG/Q9ibNUsZWTEDVjDGk4wh4w6M9lV/Wlmu7e1R4A/N6eT1UwSYwlRoakYdQ
JvDctkXnYp76zGGWhCc6J/r8misu7tKOkrCz5uffAyfop4KP15aREwGQyjOlbxCRHK+g6n4CMw81
Vv7WbLIMqnSDqjnVmv9KeWY9xcYLXcf8L2DSYaN2j1viD8MuJNlmyHdq2NW0/Swt9cjLWAAxH7/B
GNUcC0XgpHqcm3BBrF5SFnPJ2nV4hqQF7AZM1s2ui1kUND13McKph402PUNWcdS+gdQIyP3ewt4/
TDciaz8lbiKNe2cUDipHmN+Thrmp9WnhihHpS8mXS3SwapmqRw7JU7kS7xB2jNY6PFolHqKHNh7X
Yn56/PouWevSyp5mLhXD4GUpqzhwsbHbT01LgfhcJjlVuWt3e5dKJzv4pKso8J2m3cWjPdf9TlN2
IctG2M4vYjGXAV2ost0dLlh6/8YZeqOtmphg8xymkeyHCYWElyD2wHQl/Uzu5qSolJQKPY6zJ1u1
9B9BS5T8UoO13zJOdhmb5TbCm1Gjm0Lo5dbIx12ZY5ckKi8UymPJXwhWMErDU0Vfn3hxkQVUFu3m
H1q9e1+0Xwd/yot4st1MDuVW8DgReFKybEnzuqBiU0O6zjqQNYoPanFNpS/UgGr+sEK488Itj+6i
lx56Hfj5mv8aRB9Aug0sTD/3gi1esxHD4XEtn2Z+8oI6l3rnURK6DvyaQ4Xmi2fFpmT7n3Znr1FB
mO75m6nyrHnYsuLl2pl14jXhoi5lQqFtBMgaPqphsW3yDwjRF3ClZj3fLyZzz2ZjWudFzy3bX4Uv
GGMTzwb4KcpAHJorNoCotsxV0d31sJlzw8GPwinMJvcMnog8022j8v9HA5C/ZFuIUj59cSyprZrM
OMG+KCJk7VkobmJE+y74RB53Crntn7D+2bfnyJKSbrBdFweWrCiLF2kRcc5VepP5A9cBSo8SDgro
2bevjCXlcSAfvGHArjaX27U8VQ5nNzjzGjwOf1NlcAcw9Byke1HZtWyF8OuEWQEHRdER9gYPeTs4
RpqMw3y3wJrq7WsUllqYZUQk3mk3zNjUdlzssb74t0jXgzHATPjizkxuo9uZweeZVpGZzzyACwUM
FMpTgGNKSpoKYXxAoxTFmNng9ngMfoR1Rn79N34x1Ghp24+ctJ7QO08HV3jnrsL7R4BMDpGvR5JQ
QVbi7w0n+kPG+vhXFbd3RKrEUgV9nsxqWzwEbiamrbid07wxqmoQb+EMh1hDpCVeNkbhUzOkOU7m
RgUMnTIPH2UhlKdOaeqVKsRZJdtEyA6DHvd6z9SPuUGk0f1BNb2s7o/H0Ycy0j5KkZfoCrv+SJ2t
3iXAcCfJ2eS3zmxfyRQ5mpEoRxlnfVHmw48psE63PTevQWCeKoLaqFTcQNIlV/t0tnIZNLi2dSAD
xHG1mWOqIp9N9F/5hBwfOO45uyDM7VbUaiBbFodiqI8g1Va1W0GcEm31aBROVeOs1h84iXxUEz8z
7DTMgOjMNatkmv8wKatZar1itY6uG+W35SnGeWUUqZtwNYNXSpQ5RwAlzu8q9FSFyMMurK0JaomC
ClX/QAv2+Bhrz6f9HWtK+gdJ1gYK8Lf/EIwgkG9uZ5cPCicJTejTviTs2WgSUq1bZQOYRn4Cj3cU
ARl+FaQxJ2UEf8aCxMHPV57f1ovNjwp3rXvpvwnrC2wF3mE+9mQ5XdXYk2cfMp2VBj6vU1ZbCnOH
j26inCOOoqn6bPbaygP0Ym9L/ZDDl3/l0xt2udTtpVCOrYSN0Tt39rR1VGb+1XBSOfxVIisHaVgZ
JbhM09cLXh3I+Hz7MBy1giYpdICtzzfkHft+zpykiFW6QmG0w7HTLCZ+XDEW2maGO3W/fq+LeZpS
7qw1JerwIIaTmBqbTSaNBcnA3yUkD+/G1CX4ep3NFyNKuY5E2Mi06E8wl20B0vW3pu684uJi0tlR
4r7jeZ91NG9o00vJHcTQuo97ajDz0i+l9Skr0x/UYoKckPPrx/InaUHlD2MslAqH4zyMkLk+SmMw
msxbv6TSTqvvacLIjQsCH4oA9qLs5MyxBcTpL3lLX2fFYjFr1kgUO5WiMDCR0r00Ir38GwL0g9hV
5QCa2eSM0gsUSrMYhr5zSO4rbKo/GlQrls4y0UdvISbp6RVzgP8hl8r3e6ywFLckLzSOLGgr6Yt8
lqAI7JbXIAsDzNgFB8WDnhsQDZkCwrpXY4rDFTNlccDRb7R4nXAwglkS0qelnwPeM2CPYFO1o7O9
W3j0OtSgEOP9hRsIS2uesWYT+K0Sr9vsba5ieYywXl15XJGKHg3LeQ7zyQv4DQ0rmMoJTUyZv8fJ
9PAJkr/KU8wio/cYinUvdtVne2HPA2D7v4+1gk8EobYKGDI4Bk9O3M8s5SuYR66o/PTKSjK7erjK
npVOU5sMgmW32OuDRXwlNUIGPQK+OnexLj9kQnxVAm/ogY/s3SWfjEBLeUfd7HYZFV/tkupOIh63
woEItMV5xiVquCUOB3EkpJspQqRloQBGC8prgDmhCsyzQlWLPEWN2zuD6w4WOURja+oq05hq60UE
4pkjgCE5tgeoox4/Kd6BhJyf+teVmHi9vfwp/SQD4rISf4ISXtMdC+7SumKX6JMurNK+alBp8cWs
4noNJx7NJo/sOZoSLebLWpIqHybvIXf1VcGaimywFlN4DUePGBOCdESj9VUEqSdi9G+fK/X5W9fz
P8aepngObxQVol/NNy13eYdpTCSgvJrhJEyG0idtqU1MM+Bodgd4uhwYweGCbf35fQck4mwA770o
ISfs0NHh6TMUAwKok7y2GfSuH+klyEfj4UP7TTRHVrQ82/qZ0z6E7Xlwr9NE/kCawGyZ3o4TOUGQ
VkyXJCZ78NMBdKfX0BYmHid5VrqSJ9u95FXtkEGpZCt/9zJ9RCXMRkGJTMvakl4rY73UlUX6hBeB
khTRpuPcVTSWpF+9zcXXIriu0JHZyRjOYw2u+2sBPyB0zLU2rG5hPeWw8DHU+r4JVwSP205zSC+J
s6Gey9Neh41FFLYw5qXfOgEPyh+p4GtbAhpWcIP4RhXPxlrZRub7rJr0YquwWwRsXuszbfAqviah
ySTZK48OV4evwJ90tAI6G4e/u+NZ2XdgZxHffjX2LH7iJ3TiluD9GPbZbbVIcVQsPTYHFj8oKDX7
5JbILjFc/jGqkmgdy1vM3gvcs/izT3ZgHNuf65fWmeob0mg/HoYUw3t+fXr72AkXeTp+w63j3nyT
V+bVu+krfcDOUhrQDBXfhwg/oOzq2QNg7VicNjWwqwh2ikgRIZeSDf9+LbBinR6Ls7QpRQ1JQxvB
u7bD3VviAVqD3UNOCIs3uKezogcbJneNfb09YAjXJMKYdfrYtDUS/5yt1fob4dqcYE3nLbHWwkIe
/blXDrBwGuFsdih5kIZL6HF/oqUuYdKD3G+vLsRmzivbttp7xPWQlTk1zehzriS7wRQ9mX0KxaHO
XunCO3w4X/Gxsiwyr8YgiyqJwgwurVUFQJr3oRrose/3CEM8cu4ZYrKyc8HO6ClIGKjuvlh355XA
0wL1AsAxMSF7chwrJ/3LEkezDQCnmSFEqzzY3IqpOQ4csTfIVmSnBdYBvB3Ft2IxSH2yNbA5xApS
V9fkPSrBjUbTwbLqOe3IjhK5+zsbNmukebu0659XWMM0hi2kExvQPc7gdGGL++OhI7PtV+HdoYA3
42TXB+qD4xzGpdk8B6HOkBDfYmYOLP9WzixDVhFIiTA0SHRZNOhEURrDzM9hUnPwc/UVOqpgGrbX
QFZk+d/S+ieH+TCeDczldP2dVuOso2cFEautWYUq6uW5L2Ohdx/TkXk97OdwxDHgL5kq2ujt34Gf
E+AxvqVn85/eyzVapBB8D3+RagozUMYcGrPMzlwFue+RH9S7HKhbPciUQOa5086O0jj/mLvM40QZ
tuasHP21obR4efDtbZGqTl/VqBrxOj/xUdqZESgBD8cQbTNvRZBH+xp9fCmT/UOKCKLrBqr+8iT9
RIZz7FCy9dLn0ZEztwAoC04Nu5Nrv1hWMtwfDDAg5JrcpT8LEe2TNwG9hBnsgQmx1N4fPNy+aS/f
sZwcAa1FrsO8wY2ZGn4Ez4X0mvWK970Kla/2av0eHyxhqslf5EC+1osG8Gcga0x/95OkzfTbDa2r
CXLX5c0xnXe0QZmvD0VDNQfqKWd3Ub5UPX8jIwKCZB4T/QTGa3DNup8n+JidlvrW9hqju7+R/PNc
9aVs5E92KzAarp/gNHXsrzUplB06FJdgq5fJB2RApEWfd5scif+FpkDMd65I2fwfOVHOgJMPJCzk
yPpoOUJW9onH6NdyKtJ1UFR8yDlaWNYRkoWzED/ckb9LOpP9Dg1gHqmbUqXrkFgyZRDV+z1Bb9KW
Hxb9Wg3mgpFD9y5/CTpw42lwjmfc1gGEXh/guOJpBHs7SHNKt5ei4P/Jasv6gepd8fLaetxifAdP
D0vfRJNOtLaUGYUC3pqz+HQJTR71vlaFkCZ7g5ZQKbNvWv6h0PUfH3SdI/MprmK9n3okYgRAWFrk
TP2iPv7VSERvMl10h5tK5YAvYtwL2zE0t+rddT2bQh3VAWrKNFBehJiTFo1MF+QeLTNd/ThUeoJc
fZBOTbePOPdo9FfccPBmHcUPLdW9MjMRmMctHu+TCBzxf36gK9pYY9av2QVaHhVWmdm3uOzOhoI6
OFaijArs8QQbcrIRuHvXLtSW760l90G82GVBlRGFWOxjm0Cp9kXrHBBPFwE50WK5C7qvumSAngWZ
UE6Z0bALBh3bCrz9638ApFRegM+4GmxLilzP3kNcD7GR6qCqZ1NnjywIp7f7LBJ5kkgTkovL1cSH
ysnEMP6NPYVrK0G9wYBcTsLJUIsokyFehCzej1wlStwtyXEDDGZj4T9S5+N+Uhqe59CC8Dc81Njb
aiHBeltJM4Wd4dyAuGdXhuWJ9Az7ehMgSpDPsCf1jFAdju2VhsVYEMGhIsZR5UHKv6yEvQkQOPCm
V9AfQy3siqp/knbGAzcRvZk29YzkuFrKR6itH0AkKcGCHZ1sd/AyoDnjNhU1SdE/7cNeLrvVplzn
0RTpcUviiDsPvm0Glvty+dr8nE18uCmiAqCwsOK0uOmaPWAJvk0bQ763HkzdYQa9dtZvVHKiudYA
iHMtRKVzHzGWSy/tjeslE4wlbhQ1CaqH7pFraptkk/yvSIjwV0XANee7uhKgbzVnnmbhdxsnZXzz
w6BM/Rjm+h14+ueeWFfpUYlJyhDhoQrzr1enSD9v19+WiwtFYEHp2MpgBLI/7T2pHQOFGDZ0RkIA
aqRaXDjxd0Rt9XxQB9IG9Tarx7t6YBODzk0sHKfSOoF9DYRihmiq8I1QW/bddwg3MT4mUXhiDf19
EEcose7er1bVfA+msUWdaP4Wy/vqDtyX9VXcB7YfYoYUkpN42zA/Z9tgNT/Hccuo7iO8XBqKseG1
mIbzKJsuDbJb0U3JNfmsELTHZ3wMcqLM4YOMi+DFYLMYFxlAfVTr76V8IMRY2yE/hi3K83Ql+SNW
WDMOQ+zBjltxhN9Y8zpf8KGoPPZlGV0BxP+RjjrBolkz18MgSWoKsUKXl7MWBLt73vlwkuEcp+nV
lLMhMsh5vkg4mowoo9iHo/Bru+iKkA9Ws4beRGpgWHg8lc1g7ebtVCVMnWWDgKigYpA8Nj1w9tTL
qvq6TEdGhFL3cs4VaDlU16JwtPk5aaNOLrZbIzdZCS9Qf5jWx9Aemqj1986CcQefAhMZY4qLqhrv
zHYxw3kGAVm5455Moi30UoPWYddTOyRshPMBh9fzuSYd/mpZMYlhiXGK/IWTziZ7nhOwuYbNV0z8
xNsEssuedkUjuLgga6WdrNu4WRz0aC8SkGaY3FvwHQR0f4a0q1ViV4e0wMCl+OeXfOoH9ezgqrXR
DMJE78om/CAuMnFE2O5NJwWDx+pKJbwqNkzfNb8eUX5scyT/zkD6+9d5hFz3I6aqp/yEiFHU7lnW
c7pkdu07feJbJHg7B4RTIorKkthA++CGnTGmJqfWiCHwLDvNoETfbu3AWXHQfPW+dGQAHXakNUah
evKqBXDWcyJVOTUnDv/coP2LeA2diU2S0FeE98p/FlIVF62d7xxl+cCuLql3Hj8pPjrsisZ4Fcjb
OyRHCBfaKn5+p0mGMHo976+UC/XWGCR44mQCaPSOFU4bBHzA3wSoiHXewT20QKbFsCeuaFKHFAq1
5ADS32EBi43IzpTMty+sFzTn8r7tvA3oT+tLcSfr07OFZhxWA+mrS9a+SAz7Fpz0Na5SPgnp83kP
n4bKBS//VbZEQtjQU0kAbv17HmSEDzPPcfH1foJsBp7u7HaBYTwSgfaQdUNXEVNUzik6lMdrtlB6
YzEQVqBXChjAxcxjVYpWWzDSk2Wl3hZgQVTepdKuA0b/MnkQ70kPoW2PLR0k9zj1L1xxJdX+/ASm
zk3bPphIYJ1MigpGHdF5ZDbZq38Zcl9ON3/aJZpyke5wpqt5j9HXudPGAxocEBjWJVoS3NryJjKC
0/kCpZhckWGSd94auwX8WReBw6W9lX/I3+Zf91HFjU7DTCAJvux0gAUhNgvfZh7rDM805p2etZvN
HlLOzYQAsl6trkT5WbwPd3x02NyJ1vW1wdAS9687R4N8yweDVVRv9IjMm+YyHqEED34g8E0UQaPg
sJNITQq+ZBR4aJCRIdnfRM5fPr4YEC2zzJ3hvShv04sQW6L6x8ybq1EPTBX0IH1pLwc0vdtg+9tH
4aS/2UQbeHgU08z8fXyzUooGJTrB8zO4PhPafRiJ6pAWJ+spVs2eIe55ouB/FkE3GuazHhQzVKl6
OlX5BChXPUSsgQ4wL7YdijU5MDCChYcAAt0h6KgkE2jWCU89ddqXdmBWL5xyHafjMqIitZ54OlRY
ZMm+URVZv3QUkS9hJ1/JzwK8SlhEr80mXsRmeWl629tG1C+KOJYe1n+rGcmC4qLlgCyAhaRA5jjR
wgdXgUwsAoe+amkIEk+xJD4saEolmNfkA7LOP5iSOC5PayY5QiiTkjpwY5rpIDktoREDgRGpsWce
/z7crTad//e+IC2aG4A47PjKwk7EEPirRd3dRRirzwue0jG+6xqO8Vt69jgfco/iigbyFNUgqwoa
+1A4z8X+VFwLQTp0bi4EnBnxzYnrbs8u0qoYBOJ+gLMGbnW/lbsbPMLrdmFo+fAA1ZqFyJwUVbtn
Q0fgoiJAefHx4xZlPihJcVEHz5JMnkRLSh7beeP481VM+sifiq18AFOu4z8UpbCZrb90ZLYLetvy
T/DsRDsfw+DLMR2WzsPmvubekiAns49IENjMUhfD8P3BmRv9JJ2Are0Pskgv95wE1zvcUNxpqmFD
WEkTgcyFxpXNd8juDovir1IS6iv5IeKl4Xu2tpVQGoylHt6IUmCBKqHYkiHMG9SxICKLvBC5exIW
DwtnGWUyHhVWDsWtUNAtPmgdqIGZFpofL/29bt1kmVJ93RdAPCDDu3iO8R/xeeAg+i//sfAgVr/H
UKQml9bLZexA81lL+BRtwXnZ/YhpEK7t7PQfOLT+hOO/6Gk2UjWt56H4awZTRGUrfC4kmzUZB6kz
tC4upud16xz3W0elVIuyJSo8/5eGlK0VwI4yTFNQDQkVtc3YNnGPPT7q51HUmj3Llc5lJf+DOsBC
8Kva5Oz3RToNO+RSsIeV3CFIXohtXTxIA3VoDD4BR5QG66VpqqwyzokjXieXtZ0g8QOSMuDR7FR0
Ztac3o8YGK/ng0wNL/UWlxIoQMbpUanV/RuwFzjVVFpXY+i7lL0Ne08YGbW7x3TD452VQ09XcmWr
ZevHw5wcYDqCLbMQkgFBhhV52Ga4typ9eRTBQAeZg9RSua6FNQZHnxD8VP6RJNTgV4X4wChTOGoa
PgfYHnbpvMOwyrKJmZQZdOoogV55N+3qnb2Q6Pr2Q605wKt7lZvbkFGHrp5VjZZozTX9ztF4a9cf
wIHuFOACqevcvIkDkLH5g9jpb7Pn9Z0vYKc/qC/gvShMmq2WrLUchS9VRpErBfjovA89UsCmjTBp
MIONK9o/C9VzrOWLqiAE0fSN7Tt9spqWx7JkRaAV4WzMnIht2G3dqkW1kcWz1ytmCCpJs4aWhw/b
XiSDU9V058ACEMX/U1AJXA2qTvbAk43gM/ybzdc/MNoP4E2TTER8pptDmkb1OSWf04dB6HsbQJ7v
Vkp90h5pTm0ysoC6m+zDB4E25brGA2RScGbjCE4vihq/Xna1txdiEqlVnmMEOSVRoMdX8gTRpH5y
IYfN5QUvLUlkSs084Zu554grH2v4VmE6Pocykk/d1cA3JEt9VLtPogcgUfwLN/AHke5p+cdmdYpU
8dj60nMBbpkyGAAksjLhUpNetK0zuNvKPjQ7mbE+QZCsqQXWMare7AzUBAAJYJYxQnEf+0i/61gy
IkK6pAmenkjBYPPZUIgqLVg+mFA6XZsBMEa/dzRvQLo2E2wh5yb3ixzNlasrAmiwYKE0XztCkjUu
LqMr1cdvLZ1KlUJH3y4+ohX7A3tI2i/2sSrVSRREYbCnkrQl7cPzr4Cj+lWfzHmugNA3gVccpRm4
XtpGZ5cENpikBjUh+8PUCx21Mn1Nl8k7RbGagbNp6vKIKVeIGrlRp+15AciQqvLvfI5bXLhRfmlv
xif03tIQBf4C5niY9r7/EqIrgL2xOavXwZ/ZZ6QiDBbeo/0cWkxE3ixA9TjLqustI3JBJ4GJiyJA
GwrJs92gZBy4X3PSGiJ8z7PJggPfqUp3sDa3pqIlR7OV8aW5x3oeEufXS9i9srBZSPvfhnhmvxFM
7U4UqInvhPGjCJe+qI2qkqOi5ZzHZnF50HRKBUy1dbQKFdYV1C+db9AievNSryWUK4mSbf+F4ZMn
ae6VHTOrgOLNJ8nbUUQhjYxkoeP8sqpp3oyKPpkDe5gXyp6qQ4phEU//AsBmVijUvKVkxkaMes0b
8QHDFdvuD2wglu7S+h6bgcSN8SCQtMUkQXrScqWA6dUyCjUYWIn0uVF7nn3IH/u0rLXbvNe+14uz
CMMA54C6tRpvDDFck2yH79W8mpENFhJLPOEH/LFeqoFxiSpOyUoq9vxWvQJSFjZvvAmFSplKo0B8
WSUqNsFyHvow1wPMZeamzRNhi23IYHKeDUgaoad3LH0N8Tlr0nYA3dmSDK1pPludrZn9oRcfGzun
Y5HNj6nMsX5B8iWjMxpf5xyhFaHp46P3mjohwb5bPM6nlSAPUBa/7v1e1uXY4fSjC14lUaCAZoUR
mQlTTHH9nYxfhJec8+mKY2VscBUq7DWc081CLyJZf6TFnMGlcJHKK++6xGyxXGP6fJMtQywKKiTJ
4kRgzwHPbjxCQiavXMG7awUUoTIxGgbMG5YcRxM/ImKAf/MyZMyE4K0+g6ZakGR4FpaZskeV9K0v
NTELjPy5UDS9N9TtpSumKrLCQgpAT49PtqJTUcIxvpt7yMDjPuZC2DauNCPpRdTgxnPvANgsHeas
39vtZuFRXok/0T3wahHI9wBGweqBfTl7UHiOE3nHZfMmBeLu51fn62zgAgacM61etL4O5av4ddLL
ulUXEILhOkdDNgPUtV2bnq3jga4fsjduGhtANmr/dCRj//bqAqhYkkja/N3eBiObgYb0n08sOwxA
4zBxgAbc+H3PDezrIrH6TpSWO/S/70JSRvgIcXhESrgnOkuk9mflGMidtzKujlfpgd6U/0CH8q4j
xz9bebGLYqCuYOQv7cqz8DPFne6M3nnrys19rsVGeW0vhFEIhXJtodiMF5XgUUrWHKdWhhN+u5S0
yJdKcueKN4L0Z4ZUqCgmJrnyy/ysYEQ3YQYb4PawcD2aJJsqyhP5T8CoM9K0PB0XSli8FxlBY1Nf
JOOGHYpuP4SNxRowWjhWgzdY/ABu0QOPNO/oCn42/vHcOmDnTPHoW+mKDapMJlmJzr3xKraPjx6a
70IlOr8y77cnYuwR7Dx2omF7ynRci5R0qJ7btSLKW0naAfzIm+W8HWOqDirfCT5jdOfK0BobDOz4
SENbBAN9PT46aIJVDsK0p7gnJaA90GJExT1WyPX9vC+Od08scnH2Zz87O7slC1p6sPXtneX1kRVi
zmvXylcaHwXzErSvqm8gC8DOyOHY9LWpErpUgSecLsE/P7srCnvEEjpbrGhKuNtyz6dcmDx8ZHqb
V/X2j1mCYDs8wyKrJ6uQkjtgwgNw1Kglfph/vczaqqngYakm8Qa5agQJofh21wr1UoJk35Inzbhv
tITWOCtrCPp7a23d6FH4D8Yf+c3SrIIvaCEBfBXfXKG1kCoWO4aTWz4wPhn0d32yRbtWd7pwyMnQ
8FfNQ+33Ept43RuWK7Q0sysb4ecs5NbJPYl98vWlEyzEVeFj7Ay1oXpfhIHGTHn6wCz9TDTsIMkI
GeGrnJv3uwyhT7juckt05pxtTm0e+bIawqx0ZUj5e/DWeV7n47wLjyjWqYoxd8LHA0fzTVV1Df2c
L2r27kUiP8hRLHVBqlltoFE8SlvqzxPUY/FRMnmXxiHClJ6eR/djEXvXbtHJopT98Fq39jhSlqRz
nwvw+kZpIG6uS0gF6Xe9EJQX4RqBUU70Ny6TQ7WKmXjDzDasMBD4rDIJ9OT9SGFyCNUVtMe2oBv7
Drf9DLbnqkiwVYngIW+7RpegxFH5NtpVKKILfbvndkJLrJl5O14pLoTDS3KkG72bg+G2SM5Awooj
TN8qqJ/ZqAR94Rp2Z2aMZqmP8sAPoNuaeAbmmpjHT9Q4zvScGdK25j7wQ3jt9PNv71uHOOqJu3Ob
d/tIGLeilq9aKX8DRdGWpn+WczLe65OpWOB+eMSbUg2UtTNYj4xeDJay9TavfD6+v4NZ7pNNyeK8
RZkNNCLKj9USOCYJvOSgmcOweJfVFQ3OeZngVWziuS9qApHAj3IBiRWva/cJ8eYFqyP+KBJgXM3u
8c4PXbrN1rFXQP6f/AF+0cqyursT8evBt9Q5dTp8TZvc4Q+FNkRJjwod/mGsekLQcVUl9oaAX0ys
En1A3ysPzrggiV3HpId6jxv/pBAnfe/Y/o13BGMf9tb33o4uRvO6YXdnmnr02gleNK3cH2/zNNHW
V/lJXNQDfwh61hiBQa8Qng01HbuvdcrTJsRRNyaijJtTxkrhcNFaMtl/wIEz7rRenzsFBaYhVf8m
eJALHg9Uwx9FU3+9mE9/hbi/WT6ErUTmyqpiiQmPe+jzzjvSAwoGGEfWZfNzMo430+SHB5e72C2d
j8lu37SnO3kSXSjXsCzO4okS0vmN4iWs0CfzUIIByR4RKSd+VBGqWgGgEymR3H3WqW2tay+hfuGp
Wgvf3NJnSXAql3wfb+yFN1Z4EF10TBOA/A8NrkrRviV/7uB4dlD4tZxLyC8mKBgShcrZony9xrxY
Wcrlcc2p++2/JyXSQ/wrB0Xo35g82x481S5v/ZKefQK1v39hO2eULAbu8GMawavJ2Tr12lplUPDI
OLFhD3/XmTLVshDGf6yjZ2g3SleiVJGBRrrLvvwm9hSu+935SIb/bDHlmzM+o2fhCt2lrpUcZCbx
5CSaPnQyHSKHnvCtNlAxl1SalOAkKjZXsgJlL9sSlvs=
`pragma protect end_protected
